VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cic_block
  CLASS BLOCK ;
  FOREIGN cic_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 280.000 ;
  PIN io_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 -4.000 30.730 4.000 ;
    END
  END io_adr_i[0]
  PIN io_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 -4.000 37.630 4.000 ;
    END
  END io_adr_i[1]
  PIN io_cs_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 -4.000 16.930 4.000 ;
    END
  END io_cs_i
  PIN io_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 -4.000 44.070 4.000 ;
    END
  END io_dat_i[0]
  PIN io_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 -4.000 112.610 4.000 ;
    END
  END io_dat_i[10]
  PIN io_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 -4.000 119.050 4.000 ;
    END
  END io_dat_i[11]
  PIN io_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 -4.000 125.950 4.000 ;
    END
  END io_dat_i[12]
  PIN io_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 -4.000 132.850 4.000 ;
    END
  END io_dat_i[13]
  PIN io_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 -4.000 139.750 4.000 ;
    END
  END io_dat_i[14]
  PIN io_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 -4.000 146.650 4.000 ;
    END
  END io_dat_i[15]
  PIN io_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 -4.000 50.970 4.000 ;
    END
  END io_dat_i[1]
  PIN io_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 -4.000 57.870 4.000 ;
    END
  END io_dat_i[2]
  PIN io_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 -4.000 64.770 4.000 ;
    END
  END io_dat_i[3]
  PIN io_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 -4.000 71.670 4.000 ;
    END
  END io_dat_i[4]
  PIN io_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 -4.000 78.570 4.000 ;
    END
  END io_dat_i[5]
  PIN io_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 -4.000 85.010 4.000 ;
    END
  END io_dat_i[6]
  PIN io_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 -4.000 91.910 4.000 ;
    END
  END io_dat_i[7]
  PIN io_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 -4.000 98.810 4.000 ;
    END
  END io_dat_i[8]
  PIN io_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 -4.000 105.710 4.000 ;
    END
  END io_dat_i[9]
  PIN io_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 276.000 4.510 284.000 ;
    END
  END io_dat_o[0]
  PIN io_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 276.000 92.370 284.000 ;
    END
  END io_dat_o[10]
  PIN io_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 276.000 101.110 284.000 ;
    END
  END io_dat_o[11]
  PIN io_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 276.000 110.310 284.000 ;
    END
  END io_dat_o[12]
  PIN io_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 276.000 119.050 284.000 ;
    END
  END io_dat_o[13]
  PIN io_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 276.000 127.790 284.000 ;
    END
  END io_dat_o[14]
  PIN io_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 276.000 136.530 284.000 ;
    END
  END io_dat_o[15]
  PIN io_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 276.000 13.250 284.000 ;
    END
  END io_dat_o[1]
  PIN io_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 276.000 21.990 284.000 ;
    END
  END io_dat_o[2]
  PIN io_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 276.000 30.730 284.000 ;
    END
  END io_dat_o[3]
  PIN io_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 276.000 39.470 284.000 ;
    END
  END io_dat_o[4]
  PIN io_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 276.000 48.210 284.000 ;
    END
  END io_dat_o[5]
  PIN io_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 276.000 57.410 284.000 ;
    END
  END io_dat_o[6]
  PIN io_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 276.000 66.150 284.000 ;
    END
  END io_dat_o[7]
  PIN io_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 276.000 74.890 284.000 ;
    END
  END io_dat_o[8]
  PIN io_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 276.000 83.630 284.000 ;
    END
  END io_dat_o[9]
  PIN io_eo[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 147.600 154.000 148.200 ;
    END
  END io_eo[0]
  PIN io_eo[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 168.000 154.000 168.600 ;
    END
  END io_eo[10]
  PIN io_eo[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 170.040 154.000 170.640 ;
    END
  END io_eo[11]
  PIN io_eo[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 172.080 154.000 172.680 ;
    END
  END io_eo[12]
  PIN io_eo[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 174.120 154.000 174.720 ;
    END
  END io_eo[13]
  PIN io_eo[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 176.160 154.000 176.760 ;
    END
  END io_eo[14]
  PIN io_eo[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 178.200 154.000 178.800 ;
    END
  END io_eo[15]
  PIN io_eo[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 180.240 154.000 180.840 ;
    END
  END io_eo[16]
  PIN io_eo[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 182.280 154.000 182.880 ;
    END
  END io_eo[17]
  PIN io_eo[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 184.320 154.000 184.920 ;
    END
  END io_eo[18]
  PIN io_eo[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 186.360 154.000 186.960 ;
    END
  END io_eo[19]
  PIN io_eo[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 149.640 154.000 150.240 ;
    END
  END io_eo[1]
  PIN io_eo[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 188.400 154.000 189.000 ;
    END
  END io_eo[20]
  PIN io_eo[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 190.440 154.000 191.040 ;
    END
  END io_eo[21]
  PIN io_eo[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 192.480 154.000 193.080 ;
    END
  END io_eo[22]
  PIN io_eo[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 194.520 154.000 195.120 ;
    END
  END io_eo[23]
  PIN io_eo[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 196.560 154.000 197.160 ;
    END
  END io_eo[24]
  PIN io_eo[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 198.600 154.000 199.200 ;
    END
  END io_eo[25]
  PIN io_eo[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 200.640 154.000 201.240 ;
    END
  END io_eo[26]
  PIN io_eo[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 202.680 154.000 203.280 ;
    END
  END io_eo[27]
  PIN io_eo[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 204.720 154.000 205.320 ;
    END
  END io_eo[28]
  PIN io_eo[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 206.760 154.000 207.360 ;
    END
  END io_eo[29]
  PIN io_eo[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 151.680 154.000 152.280 ;
    END
  END io_eo[2]
  PIN io_eo[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 208.800 154.000 209.400 ;
    END
  END io_eo[30]
  PIN io_eo[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 210.840 154.000 211.440 ;
    END
  END io_eo[31]
  PIN io_eo[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 212.880 154.000 213.480 ;
    END
  END io_eo[32]
  PIN io_eo[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 214.920 154.000 215.520 ;
    END
  END io_eo[33]
  PIN io_eo[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 216.960 154.000 217.560 ;
    END
  END io_eo[34]
  PIN io_eo[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 219.000 154.000 219.600 ;
    END
  END io_eo[35]
  PIN io_eo[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 221.040 154.000 221.640 ;
    END
  END io_eo[36]
  PIN io_eo[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 223.080 154.000 223.680 ;
    END
  END io_eo[37]
  PIN io_eo[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 225.120 154.000 225.720 ;
    END
  END io_eo[38]
  PIN io_eo[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 227.160 154.000 227.760 ;
    END
  END io_eo[39]
  PIN io_eo[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 153.720 154.000 154.320 ;
    END
  END io_eo[3]
  PIN io_eo[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 229.200 154.000 229.800 ;
    END
  END io_eo[40]
  PIN io_eo[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 231.240 154.000 231.840 ;
    END
  END io_eo[41]
  PIN io_eo[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 233.280 154.000 233.880 ;
    END
  END io_eo[42]
  PIN io_eo[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 235.320 154.000 235.920 ;
    END
  END io_eo[43]
  PIN io_eo[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 237.360 154.000 237.960 ;
    END
  END io_eo[44]
  PIN io_eo[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 239.400 154.000 240.000 ;
    END
  END io_eo[45]
  PIN io_eo[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 241.440 154.000 242.040 ;
    END
  END io_eo[46]
  PIN io_eo[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 243.480 154.000 244.080 ;
    END
  END io_eo[47]
  PIN io_eo[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 245.520 154.000 246.120 ;
    END
  END io_eo[48]
  PIN io_eo[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 247.560 154.000 248.160 ;
    END
  END io_eo[49]
  PIN io_eo[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 155.760 154.000 156.360 ;
    END
  END io_eo[4]
  PIN io_eo[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 249.600 154.000 250.200 ;
    END
  END io_eo[50]
  PIN io_eo[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 251.640 154.000 252.240 ;
    END
  END io_eo[51]
  PIN io_eo[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 253.680 154.000 254.280 ;
    END
  END io_eo[52]
  PIN io_eo[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 255.720 154.000 256.320 ;
    END
  END io_eo[53]
  PIN io_eo[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 257.760 154.000 258.360 ;
    END
  END io_eo[54]
  PIN io_eo[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 259.800 154.000 260.400 ;
    END
  END io_eo[55]
  PIN io_eo[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 261.840 154.000 262.440 ;
    END
  END io_eo[56]
  PIN io_eo[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 263.880 154.000 264.480 ;
    END
  END io_eo[57]
  PIN io_eo[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 265.920 154.000 266.520 ;
    END
  END io_eo[58]
  PIN io_eo[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 267.960 154.000 268.560 ;
    END
  END io_eo[59]
  PIN io_eo[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 157.800 154.000 158.400 ;
    END
  END io_eo[5]
  PIN io_eo[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 270.000 154.000 270.600 ;
    END
  END io_eo[60]
  PIN io_eo[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 272.040 154.000 272.640 ;
    END
  END io_eo[61]
  PIN io_eo[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 274.080 154.000 274.680 ;
    END
  END io_eo[62]
  PIN io_eo[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 276.120 154.000 276.720 ;
    END
  END io_eo[63]
  PIN io_eo[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 159.840 154.000 160.440 ;
    END
  END io_eo[6]
  PIN io_eo[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 161.880 154.000 162.480 ;
    END
  END io_eo[7]
  PIN io_eo[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 163.920 154.000 164.520 ;
    END
  END io_eo[8]
  PIN io_eo[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 165.960 154.000 166.560 ;
    END
  END io_eo[9]
  PIN io_i_0_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 0.720 4.000 1.320 ;
    END
  END io_i_0_ci
  PIN io_i_0_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 17.040 4.000 17.640 ;
    END
  END io_i_0_in1[0]
  PIN io_i_0_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 33.360 4.000 33.960 ;
    END
  END io_i_0_in1[1]
  PIN io_i_0_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 49.680 4.000 50.280 ;
    END
  END io_i_0_in1[2]
  PIN io_i_0_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 66.000 4.000 66.600 ;
    END
  END io_i_0_in1[3]
  PIN io_i_0_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 82.320 4.000 82.920 ;
    END
  END io_i_0_in1[4]
  PIN io_i_0_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 98.640 4.000 99.240 ;
    END
  END io_i_0_in1[5]
  PIN io_i_0_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 114.960 4.000 115.560 ;
    END
  END io_i_0_in1[6]
  PIN io_i_0_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 131.280 4.000 131.880 ;
    END
  END io_i_0_in1[7]
  PIN io_i_1_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2.760 4.000 3.360 ;
    END
  END io_i_1_ci
  PIN io_i_1_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 19.080 4.000 19.680 ;
    END
  END io_i_1_in1[0]
  PIN io_i_1_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 35.400 4.000 36.000 ;
    END
  END io_i_1_in1[1]
  PIN io_i_1_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 51.720 4.000 52.320 ;
    END
  END io_i_1_in1[2]
  PIN io_i_1_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 68.040 4.000 68.640 ;
    END
  END io_i_1_in1[3]
  PIN io_i_1_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 84.360 4.000 84.960 ;
    END
  END io_i_1_in1[4]
  PIN io_i_1_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 100.680 4.000 101.280 ;
    END
  END io_i_1_in1[5]
  PIN io_i_1_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 117.000 4.000 117.600 ;
    END
  END io_i_1_in1[6]
  PIN io_i_1_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 133.320 4.000 133.920 ;
    END
  END io_i_1_in1[7]
  PIN io_i_2_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 4.800 4.000 5.400 ;
    END
  END io_i_2_ci
  PIN io_i_2_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 21.120 4.000 21.720 ;
    END
  END io_i_2_in1[0]
  PIN io_i_2_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 37.440 4.000 38.040 ;
    END
  END io_i_2_in1[1]
  PIN io_i_2_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 53.760 4.000 54.360 ;
    END
  END io_i_2_in1[2]
  PIN io_i_2_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 70.080 4.000 70.680 ;
    END
  END io_i_2_in1[3]
  PIN io_i_2_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 86.400 4.000 87.000 ;
    END
  END io_i_2_in1[4]
  PIN io_i_2_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 102.720 4.000 103.320 ;
    END
  END io_i_2_in1[5]
  PIN io_i_2_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 119.040 4.000 119.640 ;
    END
  END io_i_2_in1[6]
  PIN io_i_2_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 135.360 4.000 135.960 ;
    END
  END io_i_2_in1[7]
  PIN io_i_3_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 6.840 4.000 7.440 ;
    END
  END io_i_3_ci
  PIN io_i_3_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 23.160 4.000 23.760 ;
    END
  END io_i_3_in1[0]
  PIN io_i_3_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 39.480 4.000 40.080 ;
    END
  END io_i_3_in1[1]
  PIN io_i_3_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 55.800 4.000 56.400 ;
    END
  END io_i_3_in1[2]
  PIN io_i_3_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 72.120 4.000 72.720 ;
    END
  END io_i_3_in1[3]
  PIN io_i_3_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 88.440 4.000 89.040 ;
    END
  END io_i_3_in1[4]
  PIN io_i_3_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 104.760 4.000 105.360 ;
    END
  END io_i_3_in1[5]
  PIN io_i_3_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 121.080 4.000 121.680 ;
    END
  END io_i_3_in1[6]
  PIN io_i_3_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 137.400 4.000 138.000 ;
    END
  END io_i_3_in1[7]
  PIN io_i_4_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 8.880 4.000 9.480 ;
    END
  END io_i_4_ci
  PIN io_i_4_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 25.200 4.000 25.800 ;
    END
  END io_i_4_in1[0]
  PIN io_i_4_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 41.520 4.000 42.120 ;
    END
  END io_i_4_in1[1]
  PIN io_i_4_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 57.840 4.000 58.440 ;
    END
  END io_i_4_in1[2]
  PIN io_i_4_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 74.160 4.000 74.760 ;
    END
  END io_i_4_in1[3]
  PIN io_i_4_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 90.480 4.000 91.080 ;
    END
  END io_i_4_in1[4]
  PIN io_i_4_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 106.800 4.000 107.400 ;
    END
  END io_i_4_in1[5]
  PIN io_i_4_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 123.120 4.000 123.720 ;
    END
  END io_i_4_in1[6]
  PIN io_i_4_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 139.440 4.000 140.040 ;
    END
  END io_i_4_in1[7]
  PIN io_i_5_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 10.920 4.000 11.520 ;
    END
  END io_i_5_ci
  PIN io_i_5_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 27.240 4.000 27.840 ;
    END
  END io_i_5_in1[0]
  PIN io_i_5_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 43.560 4.000 44.160 ;
    END
  END io_i_5_in1[1]
  PIN io_i_5_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 59.880 4.000 60.480 ;
    END
  END io_i_5_in1[2]
  PIN io_i_5_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 76.200 4.000 76.800 ;
    END
  END io_i_5_in1[3]
  PIN io_i_5_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 92.520 4.000 93.120 ;
    END
  END io_i_5_in1[4]
  PIN io_i_5_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 108.840 4.000 109.440 ;
    END
  END io_i_5_in1[5]
  PIN io_i_5_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 125.160 4.000 125.760 ;
    END
  END io_i_5_in1[6]
  PIN io_i_5_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 141.480 4.000 142.080 ;
    END
  END io_i_5_in1[7]
  PIN io_i_6_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 12.960 4.000 13.560 ;
    END
  END io_i_6_ci
  PIN io_i_6_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 29.280 4.000 29.880 ;
    END
  END io_i_6_in1[0]
  PIN io_i_6_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 45.600 4.000 46.200 ;
    END
  END io_i_6_in1[1]
  PIN io_i_6_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 61.920 4.000 62.520 ;
    END
  END io_i_6_in1[2]
  PIN io_i_6_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 78.240 4.000 78.840 ;
    END
  END io_i_6_in1[3]
  PIN io_i_6_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 94.560 4.000 95.160 ;
    END
  END io_i_6_in1[4]
  PIN io_i_6_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 110.880 4.000 111.480 ;
    END
  END io_i_6_in1[5]
  PIN io_i_6_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 127.200 4.000 127.800 ;
    END
  END io_i_6_in1[6]
  PIN io_i_6_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 143.520 4.000 144.120 ;
    END
  END io_i_6_in1[7]
  PIN io_i_7_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 15.000 4.000 15.600 ;
    END
  END io_i_7_ci
  PIN io_i_7_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 31.320 4.000 31.920 ;
    END
  END io_i_7_in1[0]
  PIN io_i_7_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 47.640 4.000 48.240 ;
    END
  END io_i_7_in1[1]
  PIN io_i_7_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 63.960 4.000 64.560 ;
    END
  END io_i_7_in1[2]
  PIN io_i_7_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 80.280 4.000 80.880 ;
    END
  END io_i_7_in1[3]
  PIN io_i_7_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 96.600 4.000 97.200 ;
    END
  END io_i_7_in1[4]
  PIN io_i_7_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 112.920 4.000 113.520 ;
    END
  END io_i_7_in1[5]
  PIN io_i_7_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 129.240 4.000 129.840 ;
    END
  END io_i_7_in1[6]
  PIN io_i_7_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 145.560 4.000 146.160 ;
    END
  END io_i_7_in1[7]
  PIN io_o_0_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 0.720 154.000 1.320 ;
    END
  END io_o_0_co
  PIN io_o_0_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 17.040 154.000 17.640 ;
    END
  END io_o_0_out[0]
  PIN io_o_0_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 33.360 154.000 33.960 ;
    END
  END io_o_0_out[1]
  PIN io_o_0_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 49.680 154.000 50.280 ;
    END
  END io_o_0_out[2]
  PIN io_o_0_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 66.000 154.000 66.600 ;
    END
  END io_o_0_out[3]
  PIN io_o_0_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 82.320 154.000 82.920 ;
    END
  END io_o_0_out[4]
  PIN io_o_0_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 98.640 154.000 99.240 ;
    END
  END io_o_0_out[5]
  PIN io_o_0_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 114.960 154.000 115.560 ;
    END
  END io_o_0_out[6]
  PIN io_o_0_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 131.280 154.000 131.880 ;
    END
  END io_o_0_out[7]
  PIN io_o_1_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 2.760 154.000 3.360 ;
    END
  END io_o_1_co
  PIN io_o_1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 19.080 154.000 19.680 ;
    END
  END io_o_1_out[0]
  PIN io_o_1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 35.400 154.000 36.000 ;
    END
  END io_o_1_out[1]
  PIN io_o_1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 51.720 154.000 52.320 ;
    END
  END io_o_1_out[2]
  PIN io_o_1_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 68.040 154.000 68.640 ;
    END
  END io_o_1_out[3]
  PIN io_o_1_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 84.360 154.000 84.960 ;
    END
  END io_o_1_out[4]
  PIN io_o_1_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 100.680 154.000 101.280 ;
    END
  END io_o_1_out[5]
  PIN io_o_1_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 117.000 154.000 117.600 ;
    END
  END io_o_1_out[6]
  PIN io_o_1_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 133.320 154.000 133.920 ;
    END
  END io_o_1_out[7]
  PIN io_o_2_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 4.800 154.000 5.400 ;
    END
  END io_o_2_co
  PIN io_o_2_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 21.120 154.000 21.720 ;
    END
  END io_o_2_out[0]
  PIN io_o_2_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 37.440 154.000 38.040 ;
    END
  END io_o_2_out[1]
  PIN io_o_2_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 53.760 154.000 54.360 ;
    END
  END io_o_2_out[2]
  PIN io_o_2_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 70.080 154.000 70.680 ;
    END
  END io_o_2_out[3]
  PIN io_o_2_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 86.400 154.000 87.000 ;
    END
  END io_o_2_out[4]
  PIN io_o_2_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 102.720 154.000 103.320 ;
    END
  END io_o_2_out[5]
  PIN io_o_2_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 119.040 154.000 119.640 ;
    END
  END io_o_2_out[6]
  PIN io_o_2_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 135.360 154.000 135.960 ;
    END
  END io_o_2_out[7]
  PIN io_o_3_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 6.840 154.000 7.440 ;
    END
  END io_o_3_co
  PIN io_o_3_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 23.160 154.000 23.760 ;
    END
  END io_o_3_out[0]
  PIN io_o_3_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 39.480 154.000 40.080 ;
    END
  END io_o_3_out[1]
  PIN io_o_3_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 55.800 154.000 56.400 ;
    END
  END io_o_3_out[2]
  PIN io_o_3_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 72.120 154.000 72.720 ;
    END
  END io_o_3_out[3]
  PIN io_o_3_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 88.440 154.000 89.040 ;
    END
  END io_o_3_out[4]
  PIN io_o_3_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 104.760 154.000 105.360 ;
    END
  END io_o_3_out[5]
  PIN io_o_3_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 121.080 154.000 121.680 ;
    END
  END io_o_3_out[6]
  PIN io_o_3_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 137.400 154.000 138.000 ;
    END
  END io_o_3_out[7]
  PIN io_o_4_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 8.880 154.000 9.480 ;
    END
  END io_o_4_co
  PIN io_o_4_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 25.200 154.000 25.800 ;
    END
  END io_o_4_out[0]
  PIN io_o_4_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 41.520 154.000 42.120 ;
    END
  END io_o_4_out[1]
  PIN io_o_4_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 57.840 154.000 58.440 ;
    END
  END io_o_4_out[2]
  PIN io_o_4_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 74.160 154.000 74.760 ;
    END
  END io_o_4_out[3]
  PIN io_o_4_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 90.480 154.000 91.080 ;
    END
  END io_o_4_out[4]
  PIN io_o_4_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 106.800 154.000 107.400 ;
    END
  END io_o_4_out[5]
  PIN io_o_4_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 123.120 154.000 123.720 ;
    END
  END io_o_4_out[6]
  PIN io_o_4_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 139.440 154.000 140.040 ;
    END
  END io_o_4_out[7]
  PIN io_o_5_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 10.920 154.000 11.520 ;
    END
  END io_o_5_co
  PIN io_o_5_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 27.240 154.000 27.840 ;
    END
  END io_o_5_out[0]
  PIN io_o_5_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 43.560 154.000 44.160 ;
    END
  END io_o_5_out[1]
  PIN io_o_5_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 59.880 154.000 60.480 ;
    END
  END io_o_5_out[2]
  PIN io_o_5_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 76.200 154.000 76.800 ;
    END
  END io_o_5_out[3]
  PIN io_o_5_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 92.520 154.000 93.120 ;
    END
  END io_o_5_out[4]
  PIN io_o_5_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 108.840 154.000 109.440 ;
    END
  END io_o_5_out[5]
  PIN io_o_5_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 125.160 154.000 125.760 ;
    END
  END io_o_5_out[6]
  PIN io_o_5_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 141.480 154.000 142.080 ;
    END
  END io_o_5_out[7]
  PIN io_o_6_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 12.960 154.000 13.560 ;
    END
  END io_o_6_co
  PIN io_o_6_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 29.280 154.000 29.880 ;
    END
  END io_o_6_out[0]
  PIN io_o_6_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 45.600 154.000 46.200 ;
    END
  END io_o_6_out[1]
  PIN io_o_6_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 61.920 154.000 62.520 ;
    END
  END io_o_6_out[2]
  PIN io_o_6_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 78.240 154.000 78.840 ;
    END
  END io_o_6_out[3]
  PIN io_o_6_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 94.560 154.000 95.160 ;
    END
  END io_o_6_out[4]
  PIN io_o_6_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 110.880 154.000 111.480 ;
    END
  END io_o_6_out[5]
  PIN io_o_6_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 127.200 154.000 127.800 ;
    END
  END io_o_6_out[6]
  PIN io_o_6_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 143.520 154.000 144.120 ;
    END
  END io_o_6_out[7]
  PIN io_o_7_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 15.000 154.000 15.600 ;
    END
  END io_o_7_co
  PIN io_o_7_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 31.320 154.000 31.920 ;
    END
  END io_o_7_out[0]
  PIN io_o_7_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 47.640 154.000 48.240 ;
    END
  END io_o_7_out[1]
  PIN io_o_7_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 63.960 154.000 64.560 ;
    END
  END io_o_7_out[2]
  PIN io_o_7_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 80.280 154.000 80.880 ;
    END
  END io_o_7_out[3]
  PIN io_o_7_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 96.600 154.000 97.200 ;
    END
  END io_o_7_out[4]
  PIN io_o_7_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 112.920 154.000 113.520 ;
    END
  END io_o_7_out[5]
  PIN io_o_7_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 129.240 154.000 129.840 ;
    END
  END io_o_7_out[6]
  PIN io_o_7_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 145.560 154.000 146.160 ;
    END
  END io_o_7_out[7]
  PIN io_vci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 -4.000 3.590 4.000 ;
    END
  END io_vci
  PIN io_vco
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 -4.000 10.030 4.000 ;
    END
  END io_vco
  PIN io_vi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 276.000 145.270 284.000 ;
    END
  END io_vi
  PIN io_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 -4.000 23.830 4.000 ;
    END
  END io_we_i
  PIN io_wo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 147.600 4.000 148.200 ;
    END
  END io_wo[0]
  PIN io_wo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 168.000 4.000 168.600 ;
    END
  END io_wo[10]
  PIN io_wo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 170.040 4.000 170.640 ;
    END
  END io_wo[11]
  PIN io_wo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 172.080 4.000 172.680 ;
    END
  END io_wo[12]
  PIN io_wo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 174.120 4.000 174.720 ;
    END
  END io_wo[13]
  PIN io_wo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 176.160 4.000 176.760 ;
    END
  END io_wo[14]
  PIN io_wo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 178.200 4.000 178.800 ;
    END
  END io_wo[15]
  PIN io_wo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 180.240 4.000 180.840 ;
    END
  END io_wo[16]
  PIN io_wo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 182.280 4.000 182.880 ;
    END
  END io_wo[17]
  PIN io_wo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 184.320 4.000 184.920 ;
    END
  END io_wo[18]
  PIN io_wo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 186.360 4.000 186.960 ;
    END
  END io_wo[19]
  PIN io_wo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 149.640 4.000 150.240 ;
    END
  END io_wo[1]
  PIN io_wo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 188.400 4.000 189.000 ;
    END
  END io_wo[20]
  PIN io_wo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 190.440 4.000 191.040 ;
    END
  END io_wo[21]
  PIN io_wo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 192.480 4.000 193.080 ;
    END
  END io_wo[22]
  PIN io_wo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 194.520 4.000 195.120 ;
    END
  END io_wo[23]
  PIN io_wo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 196.560 4.000 197.160 ;
    END
  END io_wo[24]
  PIN io_wo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 198.600 4.000 199.200 ;
    END
  END io_wo[25]
  PIN io_wo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 200.640 4.000 201.240 ;
    END
  END io_wo[26]
  PIN io_wo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 202.680 4.000 203.280 ;
    END
  END io_wo[27]
  PIN io_wo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 204.720 4.000 205.320 ;
    END
  END io_wo[28]
  PIN io_wo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 206.760 4.000 207.360 ;
    END
  END io_wo[29]
  PIN io_wo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 151.680 4.000 152.280 ;
    END
  END io_wo[2]
  PIN io_wo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 208.800 4.000 209.400 ;
    END
  END io_wo[30]
  PIN io_wo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 210.840 4.000 211.440 ;
    END
  END io_wo[31]
  PIN io_wo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 212.880 4.000 213.480 ;
    END
  END io_wo[32]
  PIN io_wo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 214.920 4.000 215.520 ;
    END
  END io_wo[33]
  PIN io_wo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 216.960 4.000 217.560 ;
    END
  END io_wo[34]
  PIN io_wo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 219.000 4.000 219.600 ;
    END
  END io_wo[35]
  PIN io_wo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 221.040 4.000 221.640 ;
    END
  END io_wo[36]
  PIN io_wo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 223.080 4.000 223.680 ;
    END
  END io_wo[37]
  PIN io_wo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 225.120 4.000 225.720 ;
    END
  END io_wo[38]
  PIN io_wo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 227.160 4.000 227.760 ;
    END
  END io_wo[39]
  PIN io_wo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 153.720 4.000 154.320 ;
    END
  END io_wo[3]
  PIN io_wo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 229.200 4.000 229.800 ;
    END
  END io_wo[40]
  PIN io_wo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 231.240 4.000 231.840 ;
    END
  END io_wo[41]
  PIN io_wo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 233.280 4.000 233.880 ;
    END
  END io_wo[42]
  PIN io_wo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 235.320 4.000 235.920 ;
    END
  END io_wo[43]
  PIN io_wo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 237.360 4.000 237.960 ;
    END
  END io_wo[44]
  PIN io_wo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 239.400 4.000 240.000 ;
    END
  END io_wo[45]
  PIN io_wo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 241.440 4.000 242.040 ;
    END
  END io_wo[46]
  PIN io_wo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 243.480 4.000 244.080 ;
    END
  END io_wo[47]
  PIN io_wo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 245.520 4.000 246.120 ;
    END
  END io_wo[48]
  PIN io_wo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 247.560 4.000 248.160 ;
    END
  END io_wo[49]
  PIN io_wo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 155.760 4.000 156.360 ;
    END
  END io_wo[4]
  PIN io_wo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 249.600 4.000 250.200 ;
    END
  END io_wo[50]
  PIN io_wo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 251.640 4.000 252.240 ;
    END
  END io_wo[51]
  PIN io_wo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 253.680 4.000 254.280 ;
    END
  END io_wo[52]
  PIN io_wo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 255.720 4.000 256.320 ;
    END
  END io_wo[53]
  PIN io_wo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 257.760 4.000 258.360 ;
    END
  END io_wo[54]
  PIN io_wo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 259.800 4.000 260.400 ;
    END
  END io_wo[55]
  PIN io_wo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 261.840 4.000 262.440 ;
    END
  END io_wo[56]
  PIN io_wo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 263.880 4.000 264.480 ;
    END
  END io_wo[57]
  PIN io_wo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 265.920 4.000 266.520 ;
    END
  END io_wo[58]
  PIN io_wo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 267.960 4.000 268.560 ;
    END
  END io_wo[59]
  PIN io_wo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 157.800 4.000 158.400 ;
    END
  END io_wo[5]
  PIN io_wo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 270.000 4.000 270.600 ;
    END
  END io_wo[60]
  PIN io_wo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 272.040 4.000 272.640 ;
    END
  END io_wo[61]
  PIN io_wo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 274.080 4.000 274.680 ;
    END
  END io_wo[62]
  PIN io_wo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 276.120 4.000 276.720 ;
    END
  END io_wo[63]
  PIN io_wo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 159.840 4.000 160.440 ;
    END
  END io_wo[6]
  PIN io_wo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 161.880 4.000 162.480 ;
    END
  END io_wo[7]
  PIN io_wo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 163.920 4.000 164.520 ;
    END
  END io_wo[8]
  PIN io_wo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 165.960 4.000 166.560 ;
    END
  END io_wo[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 278.160 154.000 278.760 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 278.160 4.000 278.760 ;
    END
  END wb_rst_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 120.520 10.640 122.120 266.800 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 74.200 10.640 75.800 266.800 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.880 10.640 29.480 266.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.360 10.640 98.960 266.800 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 266.800 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 145.215 266.645 ;
      LAYER met1 ;
        RECT 3.290 5.140 146.670 270.260 ;
      LAYER met2 ;
        RECT 3.320 275.720 3.950 278.645 ;
        RECT 4.790 275.720 12.690 278.645 ;
        RECT 13.530 275.720 21.430 278.645 ;
        RECT 22.270 275.720 30.170 278.645 ;
        RECT 31.010 275.720 38.910 278.645 ;
        RECT 39.750 275.720 47.650 278.645 ;
        RECT 48.490 275.720 56.850 278.645 ;
        RECT 57.690 275.720 65.590 278.645 ;
        RECT 66.430 275.720 74.330 278.645 ;
        RECT 75.170 275.720 83.070 278.645 ;
        RECT 83.910 275.720 91.810 278.645 ;
        RECT 92.650 275.720 100.550 278.645 ;
        RECT 101.390 275.720 109.750 278.645 ;
        RECT 110.590 275.720 118.490 278.645 ;
        RECT 119.330 275.720 127.230 278.645 ;
        RECT 128.070 275.720 135.970 278.645 ;
        RECT 136.810 275.720 144.710 278.645 ;
        RECT 145.550 275.720 146.640 278.645 ;
        RECT 3.320 4.280 146.640 275.720 ;
        RECT 3.870 0.835 9.470 4.280 ;
        RECT 10.310 0.835 16.370 4.280 ;
        RECT 17.210 0.835 23.270 4.280 ;
        RECT 24.110 0.835 30.170 4.280 ;
        RECT 31.010 0.835 37.070 4.280 ;
        RECT 37.910 0.835 43.510 4.280 ;
        RECT 44.350 0.835 50.410 4.280 ;
        RECT 51.250 0.835 57.310 4.280 ;
        RECT 58.150 0.835 64.210 4.280 ;
        RECT 65.050 0.835 71.110 4.280 ;
        RECT 71.950 0.835 78.010 4.280 ;
        RECT 78.850 0.835 84.450 4.280 ;
        RECT 85.290 0.835 91.350 4.280 ;
        RECT 92.190 0.835 98.250 4.280 ;
        RECT 99.090 0.835 105.150 4.280 ;
        RECT 105.990 0.835 112.050 4.280 ;
        RECT 112.890 0.835 118.490 4.280 ;
        RECT 119.330 0.835 125.390 4.280 ;
        RECT 126.230 0.835 132.290 4.280 ;
        RECT 133.130 0.835 139.190 4.280 ;
        RECT 140.030 0.835 146.090 4.280 ;
      LAYER met3 ;
        RECT 4.400 277.760 145.600 278.625 ;
        RECT 4.000 277.120 146.000 277.760 ;
        RECT 4.400 275.720 145.600 277.120 ;
        RECT 4.000 275.080 146.000 275.720 ;
        RECT 4.400 273.680 145.600 275.080 ;
        RECT 4.000 273.040 146.000 273.680 ;
        RECT 4.400 271.640 145.600 273.040 ;
        RECT 4.000 271.000 146.000 271.640 ;
        RECT 4.400 269.600 145.600 271.000 ;
        RECT 4.000 268.960 146.000 269.600 ;
        RECT 4.400 267.560 145.600 268.960 ;
        RECT 4.000 266.920 146.000 267.560 ;
        RECT 4.400 265.520 145.600 266.920 ;
        RECT 4.000 264.880 146.000 265.520 ;
        RECT 4.400 263.480 145.600 264.880 ;
        RECT 4.000 262.840 146.000 263.480 ;
        RECT 4.400 261.440 145.600 262.840 ;
        RECT 4.000 260.800 146.000 261.440 ;
        RECT 4.400 259.400 145.600 260.800 ;
        RECT 4.000 258.760 146.000 259.400 ;
        RECT 4.400 257.360 145.600 258.760 ;
        RECT 4.000 256.720 146.000 257.360 ;
        RECT 4.400 255.320 145.600 256.720 ;
        RECT 4.000 254.680 146.000 255.320 ;
        RECT 4.400 253.280 145.600 254.680 ;
        RECT 4.000 252.640 146.000 253.280 ;
        RECT 4.400 251.240 145.600 252.640 ;
        RECT 4.000 250.600 146.000 251.240 ;
        RECT 4.400 249.200 145.600 250.600 ;
        RECT 4.000 248.560 146.000 249.200 ;
        RECT 4.400 247.160 145.600 248.560 ;
        RECT 4.000 246.520 146.000 247.160 ;
        RECT 4.400 245.120 145.600 246.520 ;
        RECT 4.000 244.480 146.000 245.120 ;
        RECT 4.400 243.080 145.600 244.480 ;
        RECT 4.000 242.440 146.000 243.080 ;
        RECT 4.400 241.040 145.600 242.440 ;
        RECT 4.000 240.400 146.000 241.040 ;
        RECT 4.400 239.000 145.600 240.400 ;
        RECT 4.000 238.360 146.000 239.000 ;
        RECT 4.400 236.960 145.600 238.360 ;
        RECT 4.000 236.320 146.000 236.960 ;
        RECT 4.400 234.920 145.600 236.320 ;
        RECT 4.000 234.280 146.000 234.920 ;
        RECT 4.400 232.880 145.600 234.280 ;
        RECT 4.000 232.240 146.000 232.880 ;
        RECT 4.400 230.840 145.600 232.240 ;
        RECT 4.000 230.200 146.000 230.840 ;
        RECT 4.400 228.800 145.600 230.200 ;
        RECT 4.000 228.160 146.000 228.800 ;
        RECT 4.400 226.760 145.600 228.160 ;
        RECT 4.000 226.120 146.000 226.760 ;
        RECT 4.400 224.720 145.600 226.120 ;
        RECT 4.000 224.080 146.000 224.720 ;
        RECT 4.400 222.680 145.600 224.080 ;
        RECT 4.000 222.040 146.000 222.680 ;
        RECT 4.400 220.640 145.600 222.040 ;
        RECT 4.000 220.000 146.000 220.640 ;
        RECT 4.400 218.600 145.600 220.000 ;
        RECT 4.000 217.960 146.000 218.600 ;
        RECT 4.400 216.560 145.600 217.960 ;
        RECT 4.000 215.920 146.000 216.560 ;
        RECT 4.400 214.520 145.600 215.920 ;
        RECT 4.000 213.880 146.000 214.520 ;
        RECT 4.400 212.480 145.600 213.880 ;
        RECT 4.000 211.840 146.000 212.480 ;
        RECT 4.400 210.440 145.600 211.840 ;
        RECT 4.000 209.800 146.000 210.440 ;
        RECT 4.400 208.400 145.600 209.800 ;
        RECT 4.000 207.760 146.000 208.400 ;
        RECT 4.400 206.360 145.600 207.760 ;
        RECT 4.000 205.720 146.000 206.360 ;
        RECT 4.400 204.320 145.600 205.720 ;
        RECT 4.000 203.680 146.000 204.320 ;
        RECT 4.400 202.280 145.600 203.680 ;
        RECT 4.000 201.640 146.000 202.280 ;
        RECT 4.400 200.240 145.600 201.640 ;
        RECT 4.000 199.600 146.000 200.240 ;
        RECT 4.400 198.200 145.600 199.600 ;
        RECT 4.000 197.560 146.000 198.200 ;
        RECT 4.400 196.160 145.600 197.560 ;
        RECT 4.000 195.520 146.000 196.160 ;
        RECT 4.400 194.120 145.600 195.520 ;
        RECT 4.000 193.480 146.000 194.120 ;
        RECT 4.400 192.080 145.600 193.480 ;
        RECT 4.000 191.440 146.000 192.080 ;
        RECT 4.400 190.040 145.600 191.440 ;
        RECT 4.000 189.400 146.000 190.040 ;
        RECT 4.400 188.000 145.600 189.400 ;
        RECT 4.000 187.360 146.000 188.000 ;
        RECT 4.400 185.960 145.600 187.360 ;
        RECT 4.000 185.320 146.000 185.960 ;
        RECT 4.400 183.920 145.600 185.320 ;
        RECT 4.000 183.280 146.000 183.920 ;
        RECT 4.400 181.880 145.600 183.280 ;
        RECT 4.000 181.240 146.000 181.880 ;
        RECT 4.400 179.840 145.600 181.240 ;
        RECT 4.000 179.200 146.000 179.840 ;
        RECT 4.400 177.800 145.600 179.200 ;
        RECT 4.000 177.160 146.000 177.800 ;
        RECT 4.400 175.760 145.600 177.160 ;
        RECT 4.000 175.120 146.000 175.760 ;
        RECT 4.400 173.720 145.600 175.120 ;
        RECT 4.000 173.080 146.000 173.720 ;
        RECT 4.400 171.680 145.600 173.080 ;
        RECT 4.000 171.040 146.000 171.680 ;
        RECT 4.400 169.640 145.600 171.040 ;
        RECT 4.000 169.000 146.000 169.640 ;
        RECT 4.400 167.600 145.600 169.000 ;
        RECT 4.000 166.960 146.000 167.600 ;
        RECT 4.400 165.560 145.600 166.960 ;
        RECT 4.000 164.920 146.000 165.560 ;
        RECT 4.400 163.520 145.600 164.920 ;
        RECT 4.000 162.880 146.000 163.520 ;
        RECT 4.400 161.480 145.600 162.880 ;
        RECT 4.000 160.840 146.000 161.480 ;
        RECT 4.400 159.440 145.600 160.840 ;
        RECT 4.000 158.800 146.000 159.440 ;
        RECT 4.400 157.400 145.600 158.800 ;
        RECT 4.000 156.760 146.000 157.400 ;
        RECT 4.400 155.360 145.600 156.760 ;
        RECT 4.000 154.720 146.000 155.360 ;
        RECT 4.400 153.320 145.600 154.720 ;
        RECT 4.000 152.680 146.000 153.320 ;
        RECT 4.400 151.280 145.600 152.680 ;
        RECT 4.000 150.640 146.000 151.280 ;
        RECT 4.400 149.240 145.600 150.640 ;
        RECT 4.000 148.600 146.000 149.240 ;
        RECT 4.400 147.200 145.600 148.600 ;
        RECT 4.000 146.560 146.000 147.200 ;
        RECT 4.400 145.160 145.600 146.560 ;
        RECT 4.000 144.520 146.000 145.160 ;
        RECT 4.400 143.120 145.600 144.520 ;
        RECT 4.000 142.480 146.000 143.120 ;
        RECT 4.400 141.080 145.600 142.480 ;
        RECT 4.000 140.440 146.000 141.080 ;
        RECT 4.400 139.040 145.600 140.440 ;
        RECT 4.000 138.400 146.000 139.040 ;
        RECT 4.400 137.000 145.600 138.400 ;
        RECT 4.000 136.360 146.000 137.000 ;
        RECT 4.400 134.960 145.600 136.360 ;
        RECT 4.000 134.320 146.000 134.960 ;
        RECT 4.400 132.920 145.600 134.320 ;
        RECT 4.000 132.280 146.000 132.920 ;
        RECT 4.400 130.880 145.600 132.280 ;
        RECT 4.000 130.240 146.000 130.880 ;
        RECT 4.400 128.840 145.600 130.240 ;
        RECT 4.000 128.200 146.000 128.840 ;
        RECT 4.400 126.800 145.600 128.200 ;
        RECT 4.000 126.160 146.000 126.800 ;
        RECT 4.400 124.760 145.600 126.160 ;
        RECT 4.000 124.120 146.000 124.760 ;
        RECT 4.400 122.720 145.600 124.120 ;
        RECT 4.000 122.080 146.000 122.720 ;
        RECT 4.400 120.680 145.600 122.080 ;
        RECT 4.000 120.040 146.000 120.680 ;
        RECT 4.400 118.640 145.600 120.040 ;
        RECT 4.000 118.000 146.000 118.640 ;
        RECT 4.400 116.600 145.600 118.000 ;
        RECT 4.000 115.960 146.000 116.600 ;
        RECT 4.400 114.560 145.600 115.960 ;
        RECT 4.000 113.920 146.000 114.560 ;
        RECT 4.400 112.520 145.600 113.920 ;
        RECT 4.000 111.880 146.000 112.520 ;
        RECT 4.400 110.480 145.600 111.880 ;
        RECT 4.000 109.840 146.000 110.480 ;
        RECT 4.400 108.440 145.600 109.840 ;
        RECT 4.000 107.800 146.000 108.440 ;
        RECT 4.400 106.400 145.600 107.800 ;
        RECT 4.000 105.760 146.000 106.400 ;
        RECT 4.400 104.360 145.600 105.760 ;
        RECT 4.000 103.720 146.000 104.360 ;
        RECT 4.400 102.320 145.600 103.720 ;
        RECT 4.000 101.680 146.000 102.320 ;
        RECT 4.400 100.280 145.600 101.680 ;
        RECT 4.000 99.640 146.000 100.280 ;
        RECT 4.400 98.240 145.600 99.640 ;
        RECT 4.000 97.600 146.000 98.240 ;
        RECT 4.400 96.200 145.600 97.600 ;
        RECT 4.000 95.560 146.000 96.200 ;
        RECT 4.400 94.160 145.600 95.560 ;
        RECT 4.000 93.520 146.000 94.160 ;
        RECT 4.400 92.120 145.600 93.520 ;
        RECT 4.000 91.480 146.000 92.120 ;
        RECT 4.400 90.080 145.600 91.480 ;
        RECT 4.000 89.440 146.000 90.080 ;
        RECT 4.400 88.040 145.600 89.440 ;
        RECT 4.000 87.400 146.000 88.040 ;
        RECT 4.400 86.000 145.600 87.400 ;
        RECT 4.000 85.360 146.000 86.000 ;
        RECT 4.400 83.960 145.600 85.360 ;
        RECT 4.000 83.320 146.000 83.960 ;
        RECT 4.400 81.920 145.600 83.320 ;
        RECT 4.000 81.280 146.000 81.920 ;
        RECT 4.400 79.880 145.600 81.280 ;
        RECT 4.000 79.240 146.000 79.880 ;
        RECT 4.400 77.840 145.600 79.240 ;
        RECT 4.000 77.200 146.000 77.840 ;
        RECT 4.400 75.800 145.600 77.200 ;
        RECT 4.000 75.160 146.000 75.800 ;
        RECT 4.400 73.760 145.600 75.160 ;
        RECT 4.000 73.120 146.000 73.760 ;
        RECT 4.400 71.720 145.600 73.120 ;
        RECT 4.000 71.080 146.000 71.720 ;
        RECT 4.400 69.680 145.600 71.080 ;
        RECT 4.000 69.040 146.000 69.680 ;
        RECT 4.400 67.640 145.600 69.040 ;
        RECT 4.000 67.000 146.000 67.640 ;
        RECT 4.400 65.600 145.600 67.000 ;
        RECT 4.000 64.960 146.000 65.600 ;
        RECT 4.400 63.560 145.600 64.960 ;
        RECT 4.000 62.920 146.000 63.560 ;
        RECT 4.400 61.520 145.600 62.920 ;
        RECT 4.000 60.880 146.000 61.520 ;
        RECT 4.400 59.480 145.600 60.880 ;
        RECT 4.000 58.840 146.000 59.480 ;
        RECT 4.400 57.440 145.600 58.840 ;
        RECT 4.000 56.800 146.000 57.440 ;
        RECT 4.400 55.400 145.600 56.800 ;
        RECT 4.000 54.760 146.000 55.400 ;
        RECT 4.400 53.360 145.600 54.760 ;
        RECT 4.000 52.720 146.000 53.360 ;
        RECT 4.400 51.320 145.600 52.720 ;
        RECT 4.000 50.680 146.000 51.320 ;
        RECT 4.400 49.280 145.600 50.680 ;
        RECT 4.000 48.640 146.000 49.280 ;
        RECT 4.400 47.240 145.600 48.640 ;
        RECT 4.000 46.600 146.000 47.240 ;
        RECT 4.400 45.200 145.600 46.600 ;
        RECT 4.000 44.560 146.000 45.200 ;
        RECT 4.400 43.160 145.600 44.560 ;
        RECT 4.000 42.520 146.000 43.160 ;
        RECT 4.400 41.120 145.600 42.520 ;
        RECT 4.000 40.480 146.000 41.120 ;
        RECT 4.400 39.080 145.600 40.480 ;
        RECT 4.000 38.440 146.000 39.080 ;
        RECT 4.400 37.040 145.600 38.440 ;
        RECT 4.000 36.400 146.000 37.040 ;
        RECT 4.400 35.000 145.600 36.400 ;
        RECT 4.000 34.360 146.000 35.000 ;
        RECT 4.400 32.960 145.600 34.360 ;
        RECT 4.000 32.320 146.000 32.960 ;
        RECT 4.400 30.920 145.600 32.320 ;
        RECT 4.000 30.280 146.000 30.920 ;
        RECT 4.400 28.880 145.600 30.280 ;
        RECT 4.000 28.240 146.000 28.880 ;
        RECT 4.400 26.840 145.600 28.240 ;
        RECT 4.000 26.200 146.000 26.840 ;
        RECT 4.400 24.800 145.600 26.200 ;
        RECT 4.000 24.160 146.000 24.800 ;
        RECT 4.400 22.760 145.600 24.160 ;
        RECT 4.000 22.120 146.000 22.760 ;
        RECT 4.400 20.720 145.600 22.120 ;
        RECT 4.000 20.080 146.000 20.720 ;
        RECT 4.400 18.680 145.600 20.080 ;
        RECT 4.000 18.040 146.000 18.680 ;
        RECT 4.400 16.640 145.600 18.040 ;
        RECT 4.000 16.000 146.000 16.640 ;
        RECT 4.400 14.600 145.600 16.000 ;
        RECT 4.000 13.960 146.000 14.600 ;
        RECT 4.400 12.560 145.600 13.960 ;
        RECT 4.000 11.920 146.000 12.560 ;
        RECT 4.400 10.520 145.600 11.920 ;
        RECT 4.000 9.880 146.000 10.520 ;
        RECT 4.400 8.480 145.600 9.880 ;
        RECT 4.000 7.840 146.000 8.480 ;
        RECT 4.400 6.440 145.600 7.840 ;
        RECT 4.000 5.800 146.000 6.440 ;
        RECT 4.400 4.400 145.600 5.800 ;
        RECT 4.000 3.760 146.000 4.400 ;
        RECT 4.400 2.360 145.600 3.760 ;
        RECT 4.000 1.720 146.000 2.360 ;
        RECT 4.400 0.855 145.600 1.720 ;
  END
END cic_block
END LIBRARY

