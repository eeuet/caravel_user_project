magic
tech sky130A
magscale 1 2
timestamp 1623880151
<< locali >>
rect 8033 51255 8067 51357
rect 15945 49147 15979 49385
rect 21925 43639 21959 43809
rect 25237 41123 25271 41225
rect 19533 38335 19567 38505
rect 4629 36091 4663 36193
rect 7297 33983 7331 34153
rect 14197 31671 14231 31773
rect 22753 31671 22787 31977
rect 19441 27931 19475 28169
rect 11529 27319 11563 27421
rect 13185 24599 13219 24905
rect 17325 19703 17359 20009
rect 8953 19159 8987 19261
rect 19441 16031 19475 16201
rect 22017 12155 22051 12257
rect 8309 11543 8343 11849
rect 14197 11543 14231 11645
rect 29009 11067 29043 12121
rect 4169 8823 4203 8925
rect 14197 7395 14231 7497
rect 15853 7259 15887 7497
rect 25605 5015 25639 5253
rect 22293 3927 22327 4029
rect 19533 3383 19567 3621
rect 13553 2975 13587 3145
<< viali >>
rect 5181 53193 5215 53227
rect 7113 53193 7147 53227
rect 8033 53193 8067 53227
rect 9781 53193 9815 53227
rect 12449 53193 12483 53227
rect 13369 53193 13403 53227
rect 18613 53193 18647 53227
rect 19165 53193 19199 53227
rect 20453 53193 20487 53227
rect 21189 53193 21223 53227
rect 23213 53193 23247 53227
rect 23949 53193 23983 53227
rect 4537 53125 4571 53159
rect 15209 53125 15243 53159
rect 16681 53125 16715 53159
rect 22017 53125 22051 53159
rect 25605 53125 25639 53159
rect 6009 53057 6043 53091
rect 1869 52989 1903 53023
rect 4353 52989 4387 53023
rect 19349 52989 19383 53023
rect 24685 52989 24719 53023
rect 25789 52989 25823 53023
rect 27077 52989 27111 53023
rect 2789 52921 2823 52955
rect 5089 52921 5123 52955
rect 5825 52921 5859 52955
rect 7021 52921 7055 52955
rect 7941 52921 7975 52955
rect 9689 52921 9723 52955
rect 12357 52921 12391 52955
rect 13277 52921 13311 52955
rect 15025 52921 15059 52955
rect 16497 52921 16531 52955
rect 18521 52921 18555 52955
rect 20361 52921 20395 52955
rect 21097 52921 21131 52955
rect 21833 52921 21867 52955
rect 23121 52921 23155 52955
rect 23857 52921 23891 52955
rect 26341 52921 26375 52955
rect 1961 52853 1995 52887
rect 2881 52853 2915 52887
rect 24501 52853 24535 52887
rect 26433 52853 26467 52887
rect 27169 52853 27203 52887
rect 20085 52649 20119 52683
rect 22661 52649 22695 52683
rect 23305 52649 23339 52683
rect 23949 52649 23983 52683
rect 27905 52581 27939 52615
rect 1869 52513 1903 52547
rect 2605 52513 2639 52547
rect 4068 52513 4102 52547
rect 5641 52513 5675 52547
rect 7389 52513 7423 52547
rect 8217 52513 8251 52547
rect 12541 52513 12575 52547
rect 18236 52513 18270 52547
rect 20269 52513 20303 52547
rect 20913 52513 20947 52547
rect 21373 52513 21407 52547
rect 22845 52513 22879 52547
rect 23489 52513 23523 52547
rect 24133 52513 24167 52547
rect 24777 52513 24811 52547
rect 25421 52513 25455 52547
rect 25973 52513 26007 52547
rect 26709 52513 26743 52547
rect 2789 52445 2823 52479
rect 3801 52445 3835 52479
rect 7481 52445 7515 52479
rect 12817 52445 12851 52479
rect 13921 52445 13955 52479
rect 17969 52445 18003 52479
rect 21465 52445 21499 52479
rect 28089 52445 28123 52479
rect 24593 52377 24627 52411
rect 25237 52377 25271 52411
rect 26893 52377 26927 52411
rect 1961 52309 1995 52343
rect 5181 52309 5215 52343
rect 5733 52309 5767 52343
rect 7757 52309 7791 52343
rect 8309 52309 8343 52343
rect 19349 52309 19383 52343
rect 20729 52309 20763 52343
rect 26065 52309 26099 52343
rect 26617 52105 26651 52139
rect 4537 52037 4571 52071
rect 23213 52037 23247 52071
rect 2789 51969 2823 52003
rect 8447 51969 8481 52003
rect 11621 51969 11655 52003
rect 15301 51969 15335 52003
rect 16129 51969 16163 52003
rect 27445 51969 27479 52003
rect 2605 51901 2639 51935
rect 6009 51901 6043 51935
rect 6377 51901 6411 51935
rect 8217 51901 8251 51935
rect 9505 51901 9539 51935
rect 9781 51901 9815 51935
rect 11877 51901 11911 51935
rect 19993 51901 20027 51935
rect 21833 51901 21867 51935
rect 23673 51901 23707 51935
rect 25789 51901 25823 51935
rect 26525 51901 26559 51935
rect 27261 51901 27295 51935
rect 27997 51901 28031 51935
rect 1869 51833 1903 51867
rect 4353 51833 4387 51867
rect 11161 51833 11195 51867
rect 15209 51833 15243 51867
rect 16396 51833 16430 51867
rect 20260 51833 20294 51867
rect 22100 51833 22134 51867
rect 1961 51765 1995 51799
rect 7849 51765 7883 51799
rect 8309 51765 8343 51799
rect 13001 51765 13035 51799
rect 14749 51765 14783 51799
rect 15117 51765 15151 51799
rect 17509 51765 17543 51799
rect 21373 51765 21407 51799
rect 23765 51765 23799 51799
rect 25881 51765 25915 51799
rect 28089 51765 28123 51799
rect 3433 51561 3467 51595
rect 4353 51561 4387 51595
rect 4721 51561 4755 51595
rect 5733 51561 5767 51595
rect 7205 51561 7239 51595
rect 7297 51561 7331 51595
rect 10425 51561 10459 51595
rect 10793 51561 10827 51595
rect 12449 51561 12483 51595
rect 12817 51561 12851 51595
rect 15761 51561 15795 51595
rect 18337 51561 18371 51595
rect 20453 51561 20487 51595
rect 20821 51561 20855 51595
rect 22569 51561 22603 51595
rect 22937 51561 22971 51595
rect 5641 51493 5675 51527
rect 14648 51493 14682 51527
rect 28181 51493 28215 51527
rect 1869 51425 1903 51459
rect 2605 51425 2639 51459
rect 3341 51425 3375 51459
rect 4813 51425 4847 51459
rect 8125 51425 8159 51459
rect 8401 51425 8435 51459
rect 10885 51425 10919 51459
rect 13645 51425 13679 51459
rect 16221 51425 16255 51459
rect 18705 51425 18739 51459
rect 19533 51425 19567 51459
rect 24389 51425 24423 51459
rect 26709 51425 26743 51459
rect 27997 51425 28031 51459
rect 4997 51357 5031 51391
rect 7481 51357 7515 51391
rect 8033 51357 8067 51391
rect 10977 51357 11011 51391
rect 12909 51357 12943 51391
rect 13093 51357 13127 51391
rect 14381 51357 14415 51391
rect 18797 51357 18831 51391
rect 18889 51357 18923 51391
rect 20913 51357 20947 51391
rect 21097 51357 21131 51391
rect 23029 51357 23063 51391
rect 23121 51357 23155 51391
rect 24133 51357 24167 51391
rect 2789 51289 2823 51323
rect 1961 51221 1995 51255
rect 6837 51221 6871 51255
rect 8033 51221 8067 51255
rect 9689 51221 9723 51255
rect 13737 51221 13771 51255
rect 16313 51221 16347 51255
rect 19625 51221 19659 51255
rect 25513 51221 25547 51255
rect 26801 51221 26835 51255
rect 4445 51017 4479 51051
rect 27353 51017 27387 51051
rect 2789 50949 2823 50983
rect 8125 50949 8159 50983
rect 10149 50949 10183 50983
rect 16589 50949 16623 50983
rect 7389 50881 7423 50915
rect 7665 50881 7699 50915
rect 9781 50881 9815 50915
rect 12357 50881 12391 50915
rect 15393 50881 15427 50915
rect 17141 50881 17175 50915
rect 20545 50881 20579 50915
rect 21741 50881 21775 50915
rect 23673 50881 23707 50915
rect 1869 50813 1903 50847
rect 4353 50813 4387 50847
rect 5825 50813 5859 50847
rect 5917 50813 5951 50847
rect 6101 50813 6135 50847
rect 7297 50813 7331 50847
rect 8401 50813 8435 50847
rect 12173 50813 12207 50847
rect 13001 50813 13035 50847
rect 13645 50813 13679 50847
rect 13829 50813 13863 50847
rect 15209 50813 15243 50847
rect 16957 50813 16991 50847
rect 17785 50813 17819 50847
rect 20361 50813 20395 50847
rect 21557 50813 21591 50847
rect 22569 50813 22603 50847
rect 23397 50813 23431 50847
rect 25237 50813 25271 50847
rect 26065 50813 26099 50847
rect 26709 50813 26743 50847
rect 2605 50745 2639 50779
rect 6561 50745 6595 50779
rect 8125 50745 8159 50779
rect 27261 50745 27295 50779
rect 27997 50745 28031 50779
rect 1961 50677 1995 50711
rect 8309 50677 8343 50711
rect 10241 50677 10275 50711
rect 11805 50677 11839 50711
rect 12265 50677 12299 50711
rect 13093 50677 13127 50711
rect 13829 50677 13863 50711
rect 14841 50677 14875 50711
rect 15301 50677 15335 50711
rect 17049 50677 17083 50711
rect 17877 50677 17911 50711
rect 19993 50677 20027 50711
rect 20453 50677 20487 50711
rect 21189 50677 21223 50711
rect 21649 50677 21683 50711
rect 22385 50677 22419 50711
rect 23029 50677 23063 50711
rect 23489 50677 23523 50711
rect 25329 50677 25363 50711
rect 25881 50677 25915 50711
rect 26525 50677 26559 50711
rect 28089 50677 28123 50711
rect 3433 50473 3467 50507
rect 5641 50473 5675 50507
rect 9413 50473 9447 50507
rect 12633 50473 12667 50507
rect 14197 50473 14231 50507
rect 14289 50473 14323 50507
rect 18245 50473 18279 50507
rect 21281 50473 21315 50507
rect 23305 50473 23339 50507
rect 24225 50473 24259 50507
rect 24777 50473 24811 50507
rect 3341 50405 3375 50439
rect 27997 50405 28031 50439
rect 1869 50337 1903 50371
rect 2605 50337 2639 50371
rect 5549 50337 5583 50371
rect 5733 50337 5767 50371
rect 7113 50337 7147 50371
rect 7573 50337 7607 50371
rect 8033 50337 8067 50371
rect 9229 50337 9263 50371
rect 9505 50337 9539 50371
rect 9689 50337 9723 50371
rect 16221 50337 16255 50371
rect 16405 50337 16439 50371
rect 18337 50337 18371 50371
rect 19441 50337 19475 50371
rect 19625 50337 19659 50371
rect 21373 50337 21407 50371
rect 22661 50337 22695 50371
rect 23489 50337 23523 50371
rect 23949 50337 23983 50371
rect 24041 50337 24075 50371
rect 24961 50337 24995 50371
rect 25605 50337 25639 50371
rect 26249 50337 26283 50371
rect 26893 50337 26927 50371
rect 7665 50269 7699 50303
rect 12541 50269 12575 50303
rect 12725 50269 12759 50303
rect 14381 50269 14415 50303
rect 18429 50269 18463 50303
rect 19349 50269 19383 50303
rect 20085 50269 20119 50303
rect 21189 50269 21223 50303
rect 24225 50269 24259 50303
rect 28181 50269 28215 50303
rect 2789 50201 2823 50235
rect 26065 50201 26099 50235
rect 1961 50133 1995 50167
rect 12173 50133 12207 50167
rect 13829 50133 13863 50167
rect 16313 50133 16347 50167
rect 17877 50133 17911 50167
rect 20821 50133 20855 50167
rect 22845 50133 22879 50167
rect 25421 50133 25455 50167
rect 26709 50133 26743 50167
rect 11989 49929 12023 49963
rect 18521 49929 18555 49963
rect 20085 49929 20119 49963
rect 21189 49929 21223 49963
rect 21833 49929 21867 49963
rect 27997 49929 28031 49963
rect 2053 49793 2087 49827
rect 15117 49793 15151 49827
rect 17693 49793 17727 49827
rect 17877 49793 17911 49827
rect 2605 49725 2639 49759
rect 2789 49725 2823 49759
rect 7849 49725 7883 49759
rect 7941 49725 7975 49759
rect 11897 49725 11931 49759
rect 12081 49725 12115 49759
rect 12817 49725 12851 49759
rect 13001 49725 13035 49759
rect 13461 49725 13495 49759
rect 13645 49725 13679 49759
rect 15393 49725 15427 49759
rect 16773 49725 16807 49759
rect 18429 49725 18463 49759
rect 18613 49725 18647 49759
rect 19993 49725 20027 49759
rect 21097 49725 21131 49759
rect 21281 49725 21315 49759
rect 21741 49725 21775 49759
rect 22569 49725 22603 49759
rect 22753 49725 22787 49759
rect 23949 49725 23983 49759
rect 24133 49725 24167 49759
rect 25513 49725 25547 49759
rect 25789 49725 25823 49759
rect 27905 49725 27939 49759
rect 1869 49657 1903 49691
rect 17601 49657 17635 49691
rect 12909 49589 12943 49623
rect 13829 49589 13863 49623
rect 17233 49589 17267 49623
rect 22753 49589 22787 49623
rect 24041 49589 24075 49623
rect 26893 49589 26927 49623
rect 5917 49385 5951 49419
rect 15945 49385 15979 49419
rect 23029 49385 23063 49419
rect 23121 49385 23155 49419
rect 25421 49385 25455 49419
rect 27997 49385 28031 49419
rect 1869 49249 1903 49283
rect 2605 49249 2639 49283
rect 4160 49249 4194 49283
rect 5733 49249 5767 49283
rect 5917 49249 5951 49283
rect 7665 49249 7699 49283
rect 7932 49249 7966 49283
rect 10149 49249 10183 49283
rect 10241 49249 10275 49283
rect 10425 49249 10459 49283
rect 10517 49249 10551 49283
rect 10977 49249 11011 49283
rect 11161 49249 11195 49283
rect 12265 49249 12299 49283
rect 13553 49249 13587 49283
rect 13737 49249 13771 49283
rect 14289 49249 14323 49283
rect 14749 49249 14783 49283
rect 3893 49181 3927 49215
rect 12357 49181 12391 49215
rect 12633 49181 12667 49215
rect 13829 49181 13863 49215
rect 17417 49317 17451 49351
rect 27905 49317 27939 49351
rect 16037 49249 16071 49283
rect 20085 49249 20119 49283
rect 20269 49249 20303 49283
rect 24501 49249 24535 49283
rect 24593 49249 24627 49283
rect 24685 49249 24719 49283
rect 24869 49249 24903 49283
rect 25789 49249 25823 49283
rect 26893 49249 26927 49283
rect 21373 49181 21407 49215
rect 23213 49181 23247 49215
rect 25881 49181 25915 49215
rect 26065 49181 26099 49215
rect 2789 49113 2823 49147
rect 14427 49113 14461 49147
rect 15945 49113 15979 49147
rect 1961 49045 1995 49079
rect 5273 49045 5307 49079
rect 9045 49045 9079 49079
rect 9965 49045 9999 49079
rect 10977 49045 11011 49079
rect 13369 49045 13403 49079
rect 14565 49045 14599 49079
rect 14657 49045 14691 49079
rect 16129 49045 16163 49079
rect 17509 49045 17543 49079
rect 22661 49045 22695 49079
rect 24225 49045 24259 49079
rect 26709 49045 26743 49079
rect 7849 48841 7883 48875
rect 14933 48841 14967 48875
rect 21741 48841 21775 48875
rect 28089 48841 28123 48875
rect 3249 48773 3283 48807
rect 6285 48773 6319 48807
rect 9781 48773 9815 48807
rect 14749 48773 14783 48807
rect 25513 48773 25547 48807
rect 4905 48705 4939 48739
rect 8401 48705 8435 48739
rect 11897 48705 11931 48739
rect 13093 48705 13127 48739
rect 14933 48705 14967 48739
rect 15025 48705 15059 48739
rect 21281 48705 21315 48739
rect 23857 48705 23891 48739
rect 27445 48705 27479 48739
rect 1869 48637 1903 48671
rect 5549 48637 5583 48671
rect 5641 48637 5675 48671
rect 9965 48637 9999 48671
rect 10333 48637 10367 48671
rect 10885 48637 10919 48671
rect 12909 48637 12943 48671
rect 13277 48637 13311 48671
rect 13645 48637 13679 48671
rect 15117 48637 15151 48671
rect 17325 48637 17359 48671
rect 17509 48637 17543 48671
rect 21373 48637 21407 48671
rect 23029 48637 23063 48671
rect 23213 48637 23247 48671
rect 24317 48637 24351 48671
rect 25237 48637 25271 48671
rect 25513 48637 25547 48671
rect 25697 48637 25731 48671
rect 26709 48637 26743 48671
rect 27261 48637 27295 48671
rect 27997 48637 28031 48671
rect 2136 48569 2170 48603
rect 4721 48569 4755 48603
rect 6561 48569 6595 48603
rect 6837 48569 6871 48603
rect 8217 48569 8251 48603
rect 22385 48569 22419 48603
rect 22569 48569 22603 48603
rect 23397 48569 23431 48603
rect 4261 48501 4295 48535
rect 4629 48501 4663 48535
rect 6745 48501 6779 48535
rect 8309 48501 8343 48535
rect 10057 48501 10091 48535
rect 10149 48501 10183 48535
rect 17693 48501 17727 48535
rect 24133 48501 24167 48535
rect 24225 48501 24259 48535
rect 26525 48501 26559 48535
rect 4353 48297 4387 48331
rect 4813 48297 4847 48331
rect 5181 48297 5215 48331
rect 7113 48297 7147 48331
rect 10057 48297 10091 48331
rect 11069 48297 11103 48331
rect 24409 48297 24443 48331
rect 3240 48229 3274 48263
rect 8493 48229 8527 48263
rect 10885 48229 10919 48263
rect 20177 48229 20211 48263
rect 20729 48229 20763 48263
rect 27997 48229 28031 48263
rect 1869 48161 1903 48195
rect 7113 48161 7147 48195
rect 7297 48161 7331 48195
rect 8401 48161 8435 48195
rect 9781 48161 9815 48195
rect 9873 48161 9907 48195
rect 11161 48161 11195 48195
rect 17325 48161 17359 48195
rect 17509 48161 17543 48195
rect 18153 48161 18187 48195
rect 18337 48161 18371 48195
rect 19257 48161 19291 48195
rect 20085 48161 20119 48195
rect 20269 48161 20303 48195
rect 20913 48161 20947 48195
rect 21005 48161 21039 48195
rect 23213 48161 23247 48195
rect 24225 48161 24259 48195
rect 24363 48161 24397 48195
rect 24593 48161 24627 48195
rect 25605 48161 25639 48195
rect 26249 48161 26283 48195
rect 26893 48161 26927 48195
rect 2973 48093 3007 48127
rect 5273 48093 5307 48127
rect 5457 48093 5491 48127
rect 8585 48093 8619 48127
rect 10057 48093 10091 48127
rect 18429 48093 18463 48127
rect 19073 48093 19107 48127
rect 23029 48093 23063 48127
rect 2053 48025 2087 48059
rect 8033 48025 8067 48059
rect 17325 48025 17359 48059
rect 17969 48025 18003 48059
rect 18889 48025 18923 48059
rect 24041 48025 24075 48059
rect 28181 48025 28215 48059
rect 10885 47957 10919 47991
rect 19073 47957 19107 47991
rect 19165 47957 19199 47991
rect 20729 47957 20763 47991
rect 23397 47957 23431 47991
rect 25421 47957 25455 47991
rect 26065 47957 26099 47991
rect 26709 47957 26743 47991
rect 2605 47753 2639 47787
rect 24225 47753 24259 47787
rect 6653 47685 6687 47719
rect 18521 47685 18555 47719
rect 20085 47685 20119 47719
rect 3249 47617 3283 47651
rect 15669 47617 15703 47651
rect 20269 47617 20303 47651
rect 21281 47617 21315 47651
rect 27997 47617 28031 47651
rect 4537 47549 4571 47583
rect 5825 47549 5859 47583
rect 5917 47549 5951 47583
rect 6469 47549 6503 47583
rect 7113 47549 7147 47583
rect 7573 47549 7607 47583
rect 9505 47549 9539 47583
rect 9689 47549 9723 47583
rect 10333 47549 10367 47583
rect 10517 47549 10551 47583
rect 10977 47549 11011 47583
rect 18061 47549 18095 47583
rect 18429 47549 18463 47583
rect 18705 47549 18739 47583
rect 19993 47549 20027 47583
rect 21373 47549 21407 47583
rect 24133 47549 24167 47583
rect 25605 47549 25639 47583
rect 25881 47549 25915 47583
rect 27813 47549 27847 47583
rect 1869 47481 1903 47515
rect 2973 47481 3007 47515
rect 8401 47481 8435 47515
rect 15936 47481 15970 47515
rect 1961 47413 1995 47447
rect 3065 47413 3099 47447
rect 4629 47413 4663 47447
rect 7205 47413 7239 47447
rect 8493 47413 8527 47447
rect 9873 47413 9907 47447
rect 10425 47413 10459 47447
rect 11069 47413 11103 47447
rect 17049 47413 17083 47447
rect 20269 47413 20303 47447
rect 21741 47413 21775 47447
rect 26985 47413 27019 47447
rect 4905 47209 4939 47243
rect 5917 47209 5951 47243
rect 18337 47209 18371 47243
rect 19809 47209 19843 47243
rect 20821 47209 20855 47243
rect 24317 47209 24351 47243
rect 25421 47209 25455 47243
rect 2053 47141 2087 47175
rect 4813 47141 4847 47175
rect 9597 47141 9631 47175
rect 10609 47141 10643 47175
rect 25789 47141 25823 47175
rect 26709 47141 26743 47175
rect 27905 47141 27939 47175
rect 1869 47073 1903 47107
rect 2605 47073 2639 47107
rect 3341 47073 3375 47107
rect 4077 47073 4111 47107
rect 5733 47073 5767 47107
rect 7113 47073 7147 47107
rect 7297 47073 7331 47107
rect 8401 47073 8435 47107
rect 9413 47073 9447 47107
rect 10241 47073 10275 47107
rect 10425 47073 10459 47107
rect 12633 47073 12667 47107
rect 13645 47073 13679 47107
rect 13829 47073 13863 47107
rect 14381 47073 14415 47107
rect 14648 47073 14682 47107
rect 17877 47073 17911 47107
rect 18337 47073 18371 47107
rect 19165 47073 19199 47107
rect 19349 47073 19383 47107
rect 19993 47073 20027 47107
rect 20085 47073 20119 47107
rect 20269 47073 20303 47107
rect 20361 47073 20395 47107
rect 21005 47073 21039 47107
rect 21097 47073 21131 47107
rect 21281 47073 21315 47107
rect 22937 47073 22971 47107
rect 24225 47073 24259 47107
rect 26893 47073 26927 47107
rect 5549 47005 5583 47039
rect 7573 47005 7607 47039
rect 9689 47005 9723 47039
rect 12817 47005 12851 47039
rect 19257 47005 19291 47039
rect 21189 47005 21223 47039
rect 25881 47005 25915 47039
rect 26065 47005 26099 47039
rect 2789 46937 2823 46971
rect 9137 46937 9171 46971
rect 18015 46937 18049 46971
rect 18153 46937 18187 46971
rect 28089 46937 28123 46971
rect 3433 46869 3467 46903
rect 4169 46869 4203 46903
rect 8585 46869 8619 46903
rect 13737 46869 13771 46903
rect 15761 46869 15795 46903
rect 23029 46869 23063 46903
rect 6101 46665 6135 46699
rect 8493 46665 8527 46699
rect 9597 46665 9631 46699
rect 27997 46665 28031 46699
rect 13185 46597 13219 46631
rect 14749 46597 14783 46631
rect 16221 46597 16255 46631
rect 20821 46597 20855 46631
rect 22753 46597 22787 46631
rect 25789 46597 25823 46631
rect 10149 46529 10183 46563
rect 11805 46529 11839 46563
rect 13645 46529 13679 46563
rect 15301 46529 15335 46563
rect 16865 46529 16899 46563
rect 23305 46529 23339 46563
rect 27353 46529 27387 46563
rect 1409 46461 1443 46495
rect 4261 46461 4295 46495
rect 4445 46461 4479 46495
rect 4905 46461 4939 46495
rect 6009 46461 6043 46495
rect 6193 46461 6227 46495
rect 8401 46461 8435 46495
rect 8585 46461 8619 46495
rect 9965 46461 9999 46495
rect 16589 46461 16623 46495
rect 17417 46461 17451 46495
rect 19993 46461 20027 46495
rect 20177 46461 20211 46495
rect 20361 46461 20395 46495
rect 20821 46461 20855 46495
rect 21005 46461 21039 46495
rect 23949 46461 23983 46495
rect 24133 46461 24167 46495
rect 25973 46461 26007 46495
rect 26433 46461 26467 46495
rect 27905 46461 27939 46495
rect 1654 46393 1688 46427
rect 13737 46393 13771 46427
rect 15117 46393 15151 46427
rect 27169 46393 27203 46427
rect 2789 46325 2823 46359
rect 4353 46325 4387 46359
rect 4997 46325 5031 46359
rect 10057 46325 10091 46359
rect 11253 46325 11287 46359
rect 11621 46325 11655 46359
rect 11713 46325 11747 46359
rect 13645 46325 13679 46359
rect 15209 46325 15243 46359
rect 16681 46325 16715 46359
rect 17509 46325 17543 46359
rect 23121 46325 23155 46359
rect 23213 46325 23247 46359
rect 24317 46325 24351 46359
rect 26525 46325 26559 46359
rect 4905 46121 4939 46155
rect 4997 46121 5031 46155
rect 10057 46121 10091 46155
rect 11161 46121 11195 46155
rect 23029 46121 23063 46155
rect 23397 46121 23431 46155
rect 25421 46121 25455 46155
rect 3433 46053 3467 46087
rect 19993 46053 20027 46087
rect 24317 46053 24351 46087
rect 27905 46053 27939 46087
rect 1869 45985 1903 46019
rect 5733 45985 5767 46019
rect 9965 45985 9999 46019
rect 10793 45985 10827 46019
rect 12265 45985 12299 46019
rect 13093 45985 13127 46019
rect 13645 45985 13679 46019
rect 14473 45985 14507 46019
rect 14933 45985 14967 46019
rect 15669 45985 15703 46019
rect 17325 45985 17359 46019
rect 17509 45985 17543 46019
rect 17693 45985 17727 46019
rect 18153 45985 18187 46019
rect 19809 45985 19843 46019
rect 24225 45985 24259 46019
rect 24593 45985 24627 46019
rect 24777 45985 24811 46019
rect 25605 45985 25639 46019
rect 26249 45985 26283 46019
rect 26893 45985 26927 46019
rect 3525 45917 3559 45951
rect 3617 45917 3651 45951
rect 5089 45917 5123 45951
rect 10885 45917 10919 45951
rect 13737 45917 13771 45951
rect 15025 45917 15059 45951
rect 23489 45917 23523 45951
rect 23581 45917 23615 45951
rect 28089 45917 28123 45951
rect 2053 45849 2087 45883
rect 5825 45849 5859 45883
rect 13001 45849 13035 45883
rect 26065 45849 26099 45883
rect 3065 45781 3099 45815
rect 4537 45781 4571 45815
rect 12357 45781 12391 45815
rect 15761 45781 15795 45815
rect 18245 45781 18279 45815
rect 26709 45781 26743 45815
rect 1593 45577 1627 45611
rect 8125 45577 8159 45611
rect 23029 45577 23063 45611
rect 4261 45509 4295 45543
rect 9689 45509 9723 45543
rect 14841 45509 14875 45543
rect 16313 45509 16347 45543
rect 17877 45509 17911 45543
rect 22569 45509 22603 45543
rect 25329 45509 25363 45543
rect 2237 45441 2271 45475
rect 4813 45441 4847 45475
rect 6469 45441 6503 45475
rect 11161 45441 11195 45475
rect 11437 45441 11471 45475
rect 15393 45441 15427 45475
rect 23581 45441 23615 45475
rect 1961 45373 1995 45407
rect 3157 45373 3191 45407
rect 4629 45373 4663 45407
rect 9505 45373 9539 45407
rect 13461 45373 13495 45407
rect 13645 45373 13679 45407
rect 13737 45373 13771 45407
rect 15209 45373 15243 45407
rect 16865 45373 16899 45407
rect 17785 45373 17819 45407
rect 18153 45373 18187 45407
rect 18429 45373 18463 45407
rect 21189 45373 21223 45407
rect 23397 45373 23431 45407
rect 25237 45373 25271 45407
rect 25881 45373 25915 45407
rect 26065 45373 26099 45407
rect 27077 45373 27111 45407
rect 27629 45373 27663 45407
rect 2053 45305 2087 45339
rect 7941 45305 7975 45339
rect 13277 45305 13311 45339
rect 16589 45305 16623 45339
rect 21456 45305 21490 45339
rect 27813 45305 27847 45339
rect 3249 45237 3283 45271
rect 4721 45237 4755 45271
rect 5825 45237 5859 45271
rect 6193 45237 6227 45271
rect 6285 45237 6319 45271
rect 8146 45237 8180 45271
rect 8309 45237 8343 45271
rect 12541 45237 12575 45271
rect 15301 45237 15335 45271
rect 16773 45237 16807 45271
rect 23489 45237 23523 45271
rect 25973 45237 26007 45271
rect 26893 45237 26927 45271
rect 2881 45033 2915 45067
rect 4353 45033 4387 45067
rect 4445 45033 4479 45067
rect 22845 45033 22879 45067
rect 23397 45033 23431 45067
rect 24409 45033 24443 45067
rect 16037 44965 16071 44999
rect 19870 44965 19904 44999
rect 24041 44965 24075 44999
rect 24257 44965 24291 44999
rect 27905 44965 27939 44999
rect 1869 44897 1903 44931
rect 2973 44897 3007 44931
rect 5733 44897 5767 44931
rect 6837 44897 6871 44931
rect 7021 44897 7055 44931
rect 7573 44897 7607 44931
rect 7941 44897 7975 44931
rect 8309 44897 8343 44931
rect 9505 44897 9539 44931
rect 9689 44897 9723 44931
rect 13185 44897 13219 44931
rect 13461 44897 13495 44931
rect 14289 44897 14323 44931
rect 14933 44897 14967 44931
rect 17693 44897 17727 44931
rect 18153 44897 18187 44931
rect 18429 44897 18463 44931
rect 18981 44897 19015 44931
rect 19625 44897 19659 44931
rect 22661 44897 22695 44931
rect 22845 44897 22879 44931
rect 23305 44897 23339 44931
rect 23489 44897 23523 44931
rect 25145 44897 25179 44931
rect 25329 44897 25363 44931
rect 26249 44897 26283 44931
rect 26893 44897 26927 44931
rect 3157 44829 3191 44863
rect 4537 44829 4571 44863
rect 8769 44829 8803 44863
rect 12909 44829 12943 44863
rect 13093 44829 13127 44863
rect 13645 44829 13679 44863
rect 14105 44829 14139 44863
rect 14841 44829 14875 44863
rect 16129 44829 16163 44863
rect 16313 44829 16347 44863
rect 6837 44761 6871 44795
rect 14657 44761 14691 44795
rect 15669 44761 15703 44795
rect 28089 44761 28123 44795
rect 1961 44693 1995 44727
rect 2513 44693 2547 44727
rect 3985 44693 4019 44727
rect 5825 44693 5859 44727
rect 9229 44693 9263 44727
rect 9505 44693 9539 44727
rect 19165 44693 19199 44727
rect 21005 44693 21039 44727
rect 24225 44693 24259 44727
rect 24869 44693 24903 44727
rect 25145 44693 25179 44727
rect 26065 44693 26099 44727
rect 26709 44693 26743 44727
rect 3157 44489 3191 44523
rect 6469 44489 6503 44523
rect 24041 44489 24075 44523
rect 1961 44421 1995 44455
rect 7757 44421 7791 44455
rect 11161 44421 11195 44455
rect 16129 44421 16163 44455
rect 18245 44421 18279 44455
rect 19993 44421 20027 44455
rect 22017 44421 22051 44455
rect 23489 44421 23523 44455
rect 2421 44353 2455 44387
rect 5457 44353 5491 44387
rect 7113 44353 7147 44387
rect 9597 44353 9631 44387
rect 9781 44353 9815 44387
rect 13553 44353 13587 44387
rect 17417 44353 17451 44387
rect 18337 44353 18371 44387
rect 25513 44353 25547 44387
rect 2513 44285 2547 44319
rect 3065 44285 3099 44319
rect 6837 44285 6871 44319
rect 6929 44285 6963 44319
rect 8033 44285 8067 44319
rect 9505 44285 9539 44319
rect 10241 44285 10275 44319
rect 11345 44285 11379 44319
rect 13277 44285 13311 44319
rect 13461 44285 13495 44319
rect 16037 44285 16071 44319
rect 16221 44285 16255 44319
rect 16957 44285 16991 44319
rect 17141 44285 17175 44319
rect 18061 44285 18095 44319
rect 18797 44285 18831 44319
rect 20177 44285 20211 44319
rect 21281 44285 21315 44319
rect 22201 44285 22235 44319
rect 23397 44285 23431 44319
rect 24041 44285 24075 44319
rect 24317 44285 24351 44319
rect 27997 44285 28031 44319
rect 2421 44217 2455 44251
rect 5181 44217 5215 44251
rect 7757 44217 7791 44251
rect 10333 44217 10367 44251
rect 17877 44217 17911 44251
rect 25758 44217 25792 44251
rect 4813 44149 4847 44183
rect 5273 44149 5307 44183
rect 7941 44149 7975 44183
rect 9781 44149 9815 44183
rect 18981 44149 19015 44183
rect 21465 44149 21499 44183
rect 24225 44149 24259 44183
rect 26893 44149 26927 44183
rect 28089 44149 28123 44183
rect 3433 43945 3467 43979
rect 5641 43945 5675 43979
rect 7757 43945 7791 43979
rect 8401 43945 8435 43979
rect 10977 43945 11011 43979
rect 24685 43945 24719 43979
rect 1869 43877 1903 43911
rect 4528 43877 4562 43911
rect 9842 43877 9876 43911
rect 13369 43877 13403 43911
rect 15025 43877 15059 43911
rect 17693 43877 17727 43911
rect 20729 43877 20763 43911
rect 25329 43877 25363 43911
rect 26709 43877 26743 43911
rect 2605 43809 2639 43843
rect 3157 43809 3191 43843
rect 3341 43809 3375 43843
rect 7021 43809 7055 43843
rect 7665 43809 7699 43843
rect 8309 43809 8343 43843
rect 8493 43809 8527 43843
rect 9137 43809 9171 43843
rect 13277 43809 13311 43843
rect 14841 43809 14875 43843
rect 17601 43809 17635 43843
rect 18797 43809 18831 43843
rect 19441 43809 19475 43843
rect 20821 43809 20855 43843
rect 21925 43809 21959 43843
rect 23581 43809 23615 43843
rect 24409 43809 24443 43843
rect 25513 43809 25547 43843
rect 26157 43809 26191 43843
rect 27997 43809 28031 43843
rect 4261 43741 4295 43775
rect 6837 43741 6871 43775
rect 7205 43741 7239 43775
rect 9597 43741 9631 43775
rect 18889 43741 18923 43775
rect 19349 43741 19383 43775
rect 21005 43741 21039 43775
rect 2789 43673 2823 43707
rect 18797 43673 18831 43707
rect 24501 43741 24535 43775
rect 24685 43741 24719 43775
rect 25973 43673 26007 43707
rect 1961 43605 1995 43639
rect 8953 43605 8987 43639
rect 20361 43605 20395 43639
rect 21925 43605 21959 43639
rect 23765 43605 23799 43639
rect 26801 43605 26835 43639
rect 28089 43605 28123 43639
rect 2697 43401 2731 43435
rect 4353 43401 4387 43435
rect 4997 43401 5031 43435
rect 5825 43401 5859 43435
rect 10149 43401 10183 43435
rect 21373 43401 21407 43435
rect 25329 43401 25363 43435
rect 28089 43401 28123 43435
rect 26525 43333 26559 43367
rect 22385 43265 22419 43299
rect 27445 43265 27479 43299
rect 2605 43197 2639 43231
rect 4261 43197 4295 43231
rect 4905 43197 4939 43231
rect 5733 43197 5767 43231
rect 5917 43197 5951 43231
rect 9505 43197 9539 43231
rect 10333 43197 10367 43231
rect 10885 43197 10919 43231
rect 15025 43197 15059 43231
rect 17601 43197 17635 43231
rect 18797 43197 18831 43231
rect 19993 43197 20027 43231
rect 20260 43197 20294 43231
rect 23029 43197 23063 43231
rect 24317 43197 24351 43231
rect 25237 43197 25271 43231
rect 26065 43197 26099 43231
rect 26709 43197 26743 43231
rect 1869 43129 1903 43163
rect 11152 43129 11186 43163
rect 15292 43129 15326 43163
rect 18613 43129 18647 43163
rect 18981 43129 19015 43163
rect 22201 43129 22235 43163
rect 23121 43129 23155 43163
rect 27261 43129 27295 43163
rect 27997 43129 28031 43163
rect 1961 43061 1995 43095
rect 9597 43061 9631 43095
rect 12265 43061 12299 43095
rect 16405 43061 16439 43095
rect 17417 43061 17451 43095
rect 21833 43061 21867 43095
rect 22293 43061 22327 43095
rect 24133 43061 24167 43095
rect 25881 43061 25915 43095
rect 11161 42789 11195 42823
rect 12449 42789 12483 42823
rect 12541 42789 12575 42823
rect 18696 42789 18730 42823
rect 23121 42789 23155 42823
rect 25145 42789 25179 42823
rect 1869 42721 1903 42755
rect 2605 42721 2639 42755
rect 3709 42721 3743 42755
rect 4537 42721 4571 42755
rect 4721 42721 4755 42755
rect 7665 42721 7699 42755
rect 8861 42721 8895 42755
rect 9873 42721 9907 42755
rect 10793 42721 10827 42755
rect 10977 42721 11011 42755
rect 18429 42721 18463 42755
rect 21465 42721 21499 42755
rect 21557 42721 21591 42755
rect 23857 42721 23891 42755
rect 24041 42721 24075 42755
rect 26709 42721 26743 42755
rect 27997 42721 28031 42755
rect 3617 42653 3651 42687
rect 10057 42653 10091 42687
rect 12725 42653 12759 42687
rect 13737 42653 13771 42687
rect 14013 42653 14047 42687
rect 15117 42653 15151 42687
rect 23029 42653 23063 42687
rect 23213 42653 23247 42687
rect 24133 42653 24167 42687
rect 2789 42585 2823 42619
rect 9045 42585 9079 42619
rect 25421 42585 25455 42619
rect 1961 42517 1995 42551
rect 3985 42517 4019 42551
rect 4629 42517 4663 42551
rect 7757 42517 7791 42551
rect 12081 42517 12115 42551
rect 19809 42517 19843 42551
rect 22661 42517 22695 42551
rect 25605 42517 25639 42551
rect 26801 42517 26835 42551
rect 28089 42517 28123 42551
rect 22201 42313 22235 42347
rect 24317 42313 24351 42347
rect 2789 42245 2823 42279
rect 13645 42245 13679 42279
rect 15301 42245 15335 42279
rect 17325 42245 17359 42279
rect 25513 42245 25547 42279
rect 4353 42177 4387 42211
rect 9597 42177 9631 42211
rect 9781 42177 9815 42211
rect 12265 42177 12299 42211
rect 16681 42177 16715 42211
rect 18705 42177 18739 42211
rect 23489 42177 23523 42211
rect 26065 42177 26099 42211
rect 1409 42109 1443 42143
rect 4261 42109 4295 42143
rect 4445 42109 4479 42143
rect 4905 42109 4939 42143
rect 9505 42109 9539 42143
rect 15117 42109 15151 42143
rect 22109 42109 22143 42143
rect 22293 42109 22327 42143
rect 23121 42109 23155 42143
rect 23305 42109 23339 42143
rect 23949 42109 23983 42143
rect 24133 42109 24167 42143
rect 25237 42109 25271 42143
rect 25421 42109 25455 42143
rect 28181 42109 28215 42143
rect 1654 42041 1688 42075
rect 12510 42041 12544 42075
rect 14933 42041 14967 42075
rect 17601 42041 17635 42075
rect 17877 42041 17911 42075
rect 18521 42041 18555 42075
rect 26332 42041 26366 42075
rect 4997 41973 5031 42007
rect 9781 41973 9815 42007
rect 16037 41973 16071 42007
rect 16405 41973 16439 42007
rect 16497 41973 16531 42007
rect 17785 41973 17819 42007
rect 27445 41973 27479 42007
rect 27997 41973 28031 42007
rect 1501 41769 1535 41803
rect 1869 41769 1903 41803
rect 7665 41769 7699 41803
rect 8769 41769 8803 41803
rect 9505 41769 9539 41803
rect 10333 41769 10367 41803
rect 17509 41769 17543 41803
rect 19533 41769 19567 41803
rect 19625 41769 19659 41803
rect 26341 41769 26375 41803
rect 13185 41701 13219 41735
rect 28181 41701 28215 41735
rect 2881 41633 2915 41667
rect 3709 41633 3743 41667
rect 7573 41633 7607 41667
rect 8861 41633 8895 41667
rect 9321 41633 9355 41667
rect 9597 41633 9631 41667
rect 9781 41633 9815 41667
rect 10241 41633 10275 41667
rect 13829 41633 13863 41667
rect 14013 41633 14047 41667
rect 17325 41633 17359 41667
rect 17509 41633 17543 41667
rect 21465 41633 21499 41667
rect 24041 41633 24075 41667
rect 24225 41633 24259 41667
rect 24501 41633 24535 41667
rect 25329 41633 25363 41667
rect 26433 41633 26467 41667
rect 26617 41633 26651 41667
rect 27997 41633 28031 41667
rect 1961 41565 1995 41599
rect 2145 41565 2179 41599
rect 2973 41565 3007 41599
rect 4629 41565 4663 41599
rect 7757 41565 7791 41599
rect 8401 41565 8435 41599
rect 8585 41565 8619 41599
rect 13185 41565 13219 41599
rect 13277 41565 13311 41599
rect 19717 41565 19751 41599
rect 25237 41565 25271 41599
rect 25697 41565 25731 41599
rect 26157 41565 26191 41599
rect 3249 41497 3283 41531
rect 3985 41497 4019 41531
rect 4905 41497 4939 41531
rect 13921 41497 13955 41531
rect 24133 41497 24167 41531
rect 4169 41429 4203 41463
rect 5089 41429 5123 41463
rect 7205 41429 7239 41463
rect 12725 41429 12759 41463
rect 19165 41429 19199 41463
rect 21557 41429 21591 41463
rect 8125 41225 8159 41259
rect 25237 41225 25271 41259
rect 25329 41225 25363 41259
rect 1869 41157 1903 41191
rect 6377 41157 6411 41191
rect 6837 41157 6871 41191
rect 24133 41157 24167 41191
rect 27537 41157 27571 41191
rect 7389 41089 7423 41123
rect 9505 41089 9539 41123
rect 15761 41089 15795 41123
rect 21097 41089 21131 41123
rect 23305 41089 23339 41123
rect 25237 41089 25271 41123
rect 4261 41021 4295 41055
rect 4997 41021 5031 41055
rect 7205 41021 7239 41055
rect 8033 41021 8067 41055
rect 9772 41021 9806 41055
rect 12909 41021 12943 41055
rect 13057 41021 13091 41055
rect 13415 41021 13449 41055
rect 15485 41021 15519 41055
rect 17601 41021 17635 41055
rect 22017 41021 22051 41055
rect 22201 41021 22235 41055
rect 23121 41021 23155 41055
rect 23857 41021 23891 41055
rect 25513 41021 25547 41055
rect 26157 41021 26191 41055
rect 26801 41021 26835 41055
rect 28181 41021 28215 41055
rect 2145 40953 2179 40987
rect 2421 40953 2455 40987
rect 3065 40953 3099 40987
rect 5264 40953 5298 40987
rect 13185 40953 13219 40987
rect 13277 40953 13311 40987
rect 17846 40953 17880 40987
rect 21005 40953 21039 40987
rect 27353 40953 27387 40987
rect 2329 40885 2363 40919
rect 3157 40885 3191 40919
rect 4353 40885 4387 40919
rect 7297 40885 7331 40919
rect 10885 40885 10919 40919
rect 13553 40885 13587 40919
rect 17049 40885 17083 40919
rect 18981 40885 19015 40919
rect 20545 40885 20579 40919
rect 20913 40885 20947 40919
rect 22201 40885 22235 40919
rect 25973 40885 26007 40919
rect 26617 40885 26651 40919
rect 27997 40885 28031 40919
rect 2513 40681 2547 40715
rect 5733 40681 5767 40715
rect 7389 40681 7423 40715
rect 15393 40681 15427 40715
rect 21373 40681 21407 40715
rect 2881 40613 2915 40647
rect 4721 40613 4755 40647
rect 7481 40613 7515 40647
rect 20260 40613 20294 40647
rect 27905 40613 27939 40647
rect 1869 40545 1903 40579
rect 3709 40545 3743 40579
rect 5641 40545 5675 40579
rect 5825 40545 5859 40579
rect 7205 40545 7239 40579
rect 11161 40545 11195 40579
rect 12725 40545 12759 40579
rect 12817 40545 12851 40579
rect 12909 40545 12943 40579
rect 13093 40545 13127 40579
rect 14013 40545 14047 40579
rect 17877 40545 17911 40579
rect 18061 40545 18095 40579
rect 18889 40545 18923 40579
rect 19073 40545 19107 40579
rect 19993 40545 20027 40579
rect 23397 40545 23431 40579
rect 23857 40545 23891 40579
rect 25973 40545 26007 40579
rect 2973 40477 3007 40511
rect 3157 40477 3191 40511
rect 14289 40477 14323 40511
rect 17969 40477 18003 40511
rect 18797 40477 18831 40511
rect 19533 40477 19567 40511
rect 26065 40477 26099 40511
rect 26157 40477 26191 40511
rect 4997 40409 5031 40443
rect 1961 40341 1995 40375
rect 3801 40341 3835 40375
rect 4169 40341 4203 40375
rect 5181 40341 5215 40375
rect 6929 40341 6963 40375
rect 10977 40341 11011 40375
rect 12449 40341 12483 40375
rect 25605 40341 25639 40375
rect 27997 40341 28031 40375
rect 5549 40001 5583 40035
rect 6469 40001 6503 40035
rect 7941 40001 7975 40035
rect 13185 40001 13219 40035
rect 16221 40001 16255 40035
rect 20269 40001 20303 40035
rect 21281 40001 21315 40035
rect 22201 40001 22235 40035
rect 22937 40001 22971 40035
rect 24113 40001 24147 40035
rect 25881 40001 25915 40035
rect 4445 39933 4479 39967
rect 5089 39933 5123 39967
rect 5181 39933 5215 39967
rect 6377 39933 6411 39967
rect 6561 39933 6595 39967
rect 8171 39933 8205 39967
rect 8309 39933 8343 39967
rect 8401 39933 8435 39967
rect 8585 39933 8619 39967
rect 10701 39933 10735 39967
rect 13461 39933 13495 39967
rect 13553 39933 13587 39967
rect 13645 39933 13679 39967
rect 13829 39933 13863 39967
rect 15209 39933 15243 39967
rect 15301 39933 15335 39967
rect 15393 39933 15427 39967
rect 15577 39933 15611 39967
rect 16497 39933 16531 39967
rect 16589 39933 16623 39967
rect 16681 39933 16715 39967
rect 16865 39933 16899 39967
rect 18429 39933 18463 39967
rect 21097 39933 21131 39967
rect 22293 39933 22327 39967
rect 22477 39933 22511 39967
rect 23397 39933 23431 39967
rect 23581 39933 23615 39967
rect 24317 39933 24351 39967
rect 25421 39933 25455 39967
rect 26137 39933 26171 39967
rect 27905 39933 27939 39967
rect 1869 39865 1903 39899
rect 2605 39865 2639 39899
rect 2789 39865 2823 39899
rect 5825 39865 5859 39899
rect 10968 39865 11002 39899
rect 18245 39865 18279 39899
rect 18613 39865 18647 39899
rect 20085 39865 20119 39899
rect 23489 39865 23523 39899
rect 24041 39865 24075 39899
rect 1961 39797 1995 39831
rect 12081 39797 12115 39831
rect 14933 39797 14967 39831
rect 20729 39797 20763 39831
rect 21189 39797 21223 39831
rect 24225 39797 24259 39831
rect 25237 39797 25271 39831
rect 27261 39797 27295 39831
rect 27997 39797 28031 39831
rect 4629 39593 4663 39627
rect 12081 39593 12115 39627
rect 13921 39593 13955 39627
rect 18061 39593 18095 39627
rect 22661 39593 22695 39627
rect 3709 39525 3743 39559
rect 4537 39525 4571 39559
rect 5273 39525 5307 39559
rect 10701 39525 10735 39559
rect 27997 39525 28031 39559
rect 1869 39457 1903 39491
rect 2605 39457 2639 39491
rect 3893 39457 3927 39491
rect 3985 39457 4019 39491
rect 7021 39457 7055 39491
rect 8033 39457 8067 39491
rect 8401 39457 8435 39491
rect 8677 39457 8711 39491
rect 9689 39457 9723 39491
rect 9873 39457 9907 39491
rect 10333 39457 10367 39491
rect 10481 39457 10515 39491
rect 10609 39457 10643 39491
rect 10839 39457 10873 39491
rect 12311 39457 12345 39491
rect 12449 39457 12483 39491
rect 12541 39457 12575 39491
rect 12725 39457 12759 39491
rect 14151 39457 14185 39491
rect 14289 39457 14323 39491
rect 14386 39457 14420 39491
rect 14565 39457 14599 39491
rect 15025 39457 15059 39491
rect 15118 39457 15152 39491
rect 15301 39457 15335 39491
rect 15393 39457 15427 39491
rect 15531 39457 15565 39491
rect 18245 39457 18279 39491
rect 18961 39457 18995 39491
rect 22569 39457 22603 39491
rect 24501 39457 24535 39491
rect 26893 39457 26927 39491
rect 5457 39389 5491 39423
rect 6837 39389 6871 39423
rect 8861 39389 8895 39423
rect 18705 39389 18739 39423
rect 24409 39389 24443 39423
rect 24869 39389 24903 39423
rect 2789 39321 2823 39355
rect 3985 39321 4019 39355
rect 9137 39321 9171 39355
rect 1961 39253 1995 39287
rect 7205 39253 7239 39287
rect 9781 39253 9815 39287
rect 10977 39253 11011 39287
rect 15669 39253 15703 39287
rect 20085 39253 20119 39287
rect 26709 39253 26743 39287
rect 28089 39253 28123 39287
rect 3249 39049 3283 39083
rect 5917 39049 5951 39083
rect 7757 39049 7791 39083
rect 8493 39049 8527 39083
rect 1869 38981 1903 39015
rect 11621 38981 11655 39015
rect 18981 38981 19015 39015
rect 25881 38981 25915 39015
rect 26525 38981 26559 39015
rect 28181 38981 28215 39015
rect 1501 38913 1535 38947
rect 7297 38913 7331 38947
rect 9781 38913 9815 38947
rect 10517 38913 10551 38947
rect 3249 38845 3283 38879
rect 4353 38845 4387 38879
rect 4445 38845 4479 38879
rect 4537 38845 4571 38879
rect 4721 38845 4755 38879
rect 5181 38845 5215 38879
rect 5365 38845 5399 38879
rect 5825 38845 5859 38879
rect 6837 38845 6871 38879
rect 7021 38845 7055 38879
rect 7757 38845 7791 38879
rect 7953 38845 7987 38879
rect 8401 38845 8435 38879
rect 9873 38845 9907 38879
rect 10057 38845 10091 38879
rect 10977 38845 11011 38879
rect 11125 38845 11159 38879
rect 11483 38845 11517 38879
rect 14933 38845 14967 38879
rect 16635 38845 16669 38879
rect 16773 38845 16807 38879
rect 16865 38845 16899 38879
rect 17049 38845 17083 38879
rect 17601 38845 17635 38879
rect 22569 38845 22603 38879
rect 22753 38845 22787 38879
rect 26065 38845 26099 38879
rect 26709 38845 26743 38879
rect 27261 38845 27295 38879
rect 27997 38845 28031 38879
rect 2973 38777 3007 38811
rect 3157 38777 3191 38811
rect 11253 38777 11287 38811
rect 11345 38777 11379 38811
rect 17846 38777 17880 38811
rect 27445 38777 27479 38811
rect 1961 38709 1995 38743
rect 5273 38709 5307 38743
rect 14749 38709 14783 38743
rect 16405 38709 16439 38743
rect 22753 38709 22787 38743
rect 19533 38505 19567 38539
rect 20085 38505 20119 38539
rect 1685 38437 1719 38471
rect 2697 38437 2731 38471
rect 4537 38437 4571 38471
rect 5733 38437 5767 38471
rect 10701 38437 10735 38471
rect 17570 38437 17604 38471
rect 3617 38369 3651 38403
rect 3985 38369 4019 38403
rect 4353 38369 4387 38403
rect 4997 38369 5031 38403
rect 5641 38369 5675 38403
rect 8953 38369 8987 38403
rect 10425 38369 10459 38403
rect 10518 38369 10552 38403
rect 10793 38369 10827 38403
rect 10890 38369 10924 38403
rect 13441 38369 13475 38403
rect 15117 38369 15151 38403
rect 27905 38437 27939 38471
rect 19993 38369 20027 38403
rect 20821 38369 20855 38403
rect 21005 38369 21039 38403
rect 22937 38369 22971 38403
rect 24492 38369 24526 38403
rect 26249 38369 26283 38403
rect 26893 38369 26927 38403
rect 9045 38301 9079 38335
rect 9229 38301 9263 38335
rect 13185 38301 13219 38335
rect 17325 38301 17359 38335
rect 19533 38301 19567 38335
rect 20269 38301 20303 38335
rect 23029 38301 23063 38335
rect 23121 38301 23155 38335
rect 24225 38301 24259 38335
rect 1961 38233 1995 38267
rect 5089 38233 5123 38267
rect 8585 38233 8619 38267
rect 2145 38165 2179 38199
rect 2789 38165 2823 38199
rect 11069 38165 11103 38199
rect 14565 38165 14599 38199
rect 15209 38165 15243 38199
rect 18705 38165 18739 38199
rect 19625 38165 19659 38199
rect 21189 38165 21223 38199
rect 22569 38165 22603 38199
rect 25605 38165 25639 38199
rect 26065 38165 26099 38199
rect 26709 38165 26743 38199
rect 27997 38165 28031 38199
rect 4353 37961 4387 37995
rect 22201 37961 22235 37995
rect 27261 37961 27295 37995
rect 2513 37893 2547 37927
rect 16129 37893 16163 37927
rect 16865 37893 16899 37927
rect 20821 37825 20855 37859
rect 23029 37825 23063 37859
rect 25881 37825 25915 37859
rect 25973 37825 26007 37859
rect 2421 37757 2455 37791
rect 2789 37757 2823 37791
rect 3157 37757 3191 37791
rect 4261 37757 4295 37791
rect 4445 37757 4479 37791
rect 5089 37757 5123 37791
rect 10149 37757 10183 37791
rect 11989 37757 12023 37791
rect 15485 37757 15519 37791
rect 15633 37757 15667 37791
rect 15853 37757 15887 37791
rect 15950 37757 15984 37791
rect 20085 37757 20119 37791
rect 20269 37757 20303 37791
rect 21088 37757 21122 37791
rect 23121 37757 23155 37791
rect 23305 37757 23339 37791
rect 27169 37757 27203 37791
rect 27905 37757 27939 37791
rect 1593 37689 1627 37723
rect 5356 37689 5390 37723
rect 10416 37689 10450 37723
rect 12234 37689 12268 37723
rect 14841 37689 14875 37723
rect 15761 37689 15795 37723
rect 16681 37689 16715 37723
rect 23765 37689 23799 37723
rect 25789 37689 25823 37723
rect 1685 37621 1719 37655
rect 6469 37621 6503 37655
rect 11529 37621 11563 37655
rect 13369 37621 13403 37655
rect 14933 37621 14967 37655
rect 20269 37621 20303 37655
rect 25421 37621 25455 37655
rect 27997 37621 28031 37655
rect 28089 37417 28123 37451
rect 2053 37349 2087 37383
rect 4721 37349 4755 37383
rect 5365 37349 5399 37383
rect 9229 37349 9263 37383
rect 9965 37349 9999 37383
rect 12081 37349 12115 37383
rect 13185 37349 13219 37383
rect 14565 37349 14599 37383
rect 14657 37349 14691 37383
rect 15945 37349 15979 37383
rect 20361 37349 20395 37383
rect 20453 37349 20487 37383
rect 21281 37349 21315 37383
rect 25053 37349 25087 37383
rect 27997 37349 28031 37383
rect 1869 37281 1903 37315
rect 2605 37281 2639 37315
rect 3525 37281 3559 37315
rect 4629 37281 4663 37315
rect 4813 37281 4847 37315
rect 5273 37281 5307 37315
rect 5457 37281 5491 37315
rect 9045 37281 9079 37315
rect 9873 37281 9907 37315
rect 10057 37281 10091 37315
rect 12311 37281 12345 37315
rect 12430 37281 12464 37315
rect 12530 37281 12564 37315
rect 12725 37281 12759 37315
rect 13461 37281 13495 37315
rect 13550 37281 13584 37315
rect 13645 37281 13679 37315
rect 13829 37281 13863 37315
rect 14381 37281 14415 37315
rect 14749 37281 14783 37315
rect 15761 37281 15795 37315
rect 18317 37281 18351 37315
rect 23101 37281 23135 37315
rect 24685 37281 24719 37315
rect 24869 37281 24903 37315
rect 25881 37281 25915 37315
rect 26065 37281 26099 37315
rect 26525 37281 26559 37315
rect 3617 37213 3651 37247
rect 9321 37213 9355 37247
rect 18061 37213 18095 37247
rect 20545 37213 20579 37247
rect 22845 37213 22879 37247
rect 25789 37213 25823 37247
rect 2789 37145 2823 37179
rect 3893 37145 3927 37179
rect 8769 37145 8803 37179
rect 14933 37077 14967 37111
rect 19441 37077 19475 37111
rect 19993 37077 20027 37111
rect 21373 37077 21407 37111
rect 24225 37077 24259 37111
rect 25973 36873 26007 36907
rect 28089 36873 28123 36907
rect 4353 36805 4387 36839
rect 7205 36805 7239 36839
rect 11713 36805 11747 36839
rect 15209 36805 15243 36839
rect 18061 36805 18095 36839
rect 26617 36805 26651 36839
rect 13829 36737 13863 36771
rect 17049 36737 17083 36771
rect 4261 36669 4295 36703
rect 4445 36669 4479 36703
rect 5181 36669 5215 36703
rect 5825 36669 5859 36703
rect 9689 36669 9723 36703
rect 11989 36669 12023 36703
rect 12081 36669 12115 36703
rect 12173 36669 12207 36703
rect 12357 36669 12391 36703
rect 13645 36669 13679 36703
rect 15669 36669 15703 36703
rect 15945 36669 15979 36703
rect 18705 36669 18739 36703
rect 20729 36669 20763 36703
rect 21465 36669 21499 36703
rect 25421 36669 25455 36703
rect 25881 36669 25915 36703
rect 26065 36669 26099 36703
rect 26801 36669 26835 36703
rect 27445 36669 27479 36703
rect 1869 36601 1903 36635
rect 2605 36601 2639 36635
rect 2789 36601 2823 36635
rect 4997 36601 5031 36635
rect 5365 36601 5399 36635
rect 6070 36601 6104 36635
rect 15025 36601 15059 36635
rect 17877 36601 17911 36635
rect 27997 36601 28031 36635
rect 1961 36533 1995 36567
rect 9505 36533 9539 36567
rect 18521 36533 18555 36567
rect 20545 36533 20579 36567
rect 21557 36533 21591 36567
rect 25237 36533 25271 36567
rect 27261 36533 27295 36567
rect 3065 36329 3099 36363
rect 4905 36329 4939 36363
rect 5549 36329 5583 36363
rect 8309 36329 8343 36363
rect 9229 36329 9263 36363
rect 14105 36329 14139 36363
rect 15209 36329 15243 36363
rect 22753 36329 22787 36363
rect 25421 36329 25455 36363
rect 27997 36261 28031 36295
rect 1685 36193 1719 36227
rect 2973 36193 3007 36227
rect 3157 36193 3191 36227
rect 3801 36193 3835 36227
rect 4629 36193 4663 36227
rect 4721 36193 4755 36227
rect 4913 36193 4947 36227
rect 5457 36193 5491 36227
rect 7196 36193 7230 36227
rect 9137 36193 9171 36227
rect 10747 36193 10781 36227
rect 10885 36193 10919 36227
rect 10977 36193 11011 36227
rect 11161 36193 11195 36227
rect 12265 36193 12299 36227
rect 13921 36193 13955 36227
rect 14105 36193 14139 36227
rect 15485 36193 15519 36227
rect 15577 36193 15611 36227
rect 15669 36193 15703 36227
rect 15853 36193 15887 36227
rect 17647 36193 17681 36227
rect 17766 36193 17800 36227
rect 17866 36193 17900 36227
rect 18061 36193 18095 36227
rect 18705 36193 18739 36227
rect 18972 36193 19006 36227
rect 22983 36193 23017 36227
rect 23121 36193 23155 36227
rect 23213 36193 23247 36227
rect 23397 36193 23431 36227
rect 25605 36193 25639 36227
rect 26249 36193 26283 36227
rect 26893 36193 26927 36227
rect 1777 36125 1811 36159
rect 2421 36125 2455 36159
rect 6929 36125 6963 36159
rect 9413 36125 9447 36159
rect 17417 36125 17451 36159
rect 4629 36057 4663 36091
rect 8769 36057 8803 36091
rect 28181 36057 28215 36091
rect 3893 35989 3927 36023
rect 10517 35989 10551 36023
rect 12081 35989 12115 36023
rect 20085 35989 20119 36023
rect 26065 35989 26099 36023
rect 26709 35989 26743 36023
rect 7389 35785 7423 35819
rect 11069 35785 11103 35819
rect 12081 35785 12115 35819
rect 13645 35785 13679 35819
rect 28089 35785 28123 35819
rect 1869 35717 1903 35751
rect 2053 35717 2087 35751
rect 18245 35717 18279 35751
rect 22569 35717 22603 35751
rect 23029 35717 23063 35751
rect 9781 35649 9815 35683
rect 25237 35649 25271 35683
rect 3065 35581 3099 35615
rect 3341 35581 3375 35615
rect 4261 35581 4295 35615
rect 7205 35581 7239 35615
rect 9505 35581 9539 35615
rect 11713 35581 11747 35615
rect 11805 35581 11839 35615
rect 11897 35581 11931 35615
rect 13277 35581 13311 35615
rect 13369 35581 13403 35615
rect 13461 35581 13495 35615
rect 14749 35581 14783 35615
rect 15945 35581 15979 35615
rect 16773 35581 16807 35615
rect 18521 35581 18555 35615
rect 18613 35581 18647 35615
rect 18705 35581 18739 35615
rect 18901 35581 18935 35615
rect 21189 35581 21223 35615
rect 23213 35581 23247 35615
rect 23903 35581 23937 35615
rect 24041 35581 24075 35615
rect 24133 35581 24167 35615
rect 24317 35581 24351 35615
rect 27261 35581 27295 35615
rect 27997 35581 28031 35615
rect 1593 35513 1627 35547
rect 7021 35513 7055 35547
rect 16957 35513 16991 35547
rect 21434 35513 21468 35547
rect 23673 35513 23707 35547
rect 25482 35513 25516 35547
rect 27445 35513 27479 35547
rect 2881 35445 2915 35479
rect 3249 35445 3283 35479
rect 4445 35445 4479 35479
rect 14841 35445 14875 35479
rect 16037 35445 16071 35479
rect 26617 35445 26651 35479
rect 2421 35241 2455 35275
rect 3617 35241 3651 35275
rect 9965 35241 9999 35275
rect 12817 35241 12851 35275
rect 13461 35241 13495 35275
rect 14749 35241 14783 35275
rect 16129 35241 16163 35275
rect 17693 35241 17727 35275
rect 23489 35241 23523 35275
rect 26433 35241 26467 35275
rect 1593 35173 1627 35207
rect 19165 35173 19199 35207
rect 20913 35173 20947 35207
rect 23949 35173 23983 35207
rect 25298 35173 25332 35207
rect 27997 35173 28031 35207
rect 2513 35105 2547 35139
rect 2697 35105 2731 35139
rect 3249 35105 3283 35139
rect 3341 35105 3375 35139
rect 3433 35105 3467 35139
rect 4445 35105 4479 35139
rect 4712 35105 4746 35139
rect 7941 35105 7975 35139
rect 9781 35105 9815 35139
rect 9965 35105 9999 35139
rect 10701 35105 10735 35139
rect 10793 35105 10827 35139
rect 10885 35105 10919 35139
rect 11069 35105 11103 35139
rect 12413 35105 12447 35139
rect 12541 35105 12575 35139
rect 12633 35105 12667 35139
rect 13277 35105 13311 35139
rect 13461 35105 13495 35139
rect 14565 35105 14599 35139
rect 14749 35105 14783 35139
rect 15301 35105 15335 35139
rect 15945 35105 15979 35139
rect 17923 35105 17957 35139
rect 18061 35105 18095 35139
rect 18153 35105 18187 35139
rect 18337 35105 18371 35139
rect 18981 35105 19015 35139
rect 19855 35105 19889 35139
rect 19993 35105 20027 35139
rect 20085 35105 20119 35139
rect 20269 35105 20303 35139
rect 21169 35105 21203 35139
rect 21281 35105 21315 35139
rect 21373 35105 21407 35139
rect 21557 35105 21591 35139
rect 23085 35105 23119 35139
rect 23203 35105 23237 35139
rect 23305 35105 23339 35139
rect 24225 35105 24259 35139
rect 24317 35105 24351 35139
rect 24409 35105 24443 35139
rect 24593 35105 24627 35139
rect 25053 35105 25087 35139
rect 1685 34901 1719 34935
rect 2237 34901 2271 34935
rect 5825 34901 5859 34935
rect 7757 34901 7791 34935
rect 10425 34901 10459 34935
rect 15393 34901 15427 34935
rect 19625 34901 19659 34935
rect 28089 34901 28123 34935
rect 1685 34697 1719 34731
rect 4997 34697 5031 34731
rect 16221 34697 16255 34731
rect 17325 34697 17359 34731
rect 18245 34697 18279 34731
rect 22845 34697 22879 34731
rect 23857 34697 23891 34731
rect 25237 34697 25271 34731
rect 27353 34697 27387 34731
rect 12173 34629 12207 34663
rect 13553 34629 13587 34663
rect 28181 34629 28215 34663
rect 5917 34561 5951 34595
rect 7297 34561 7331 34595
rect 9781 34561 9815 34595
rect 1869 34493 1903 34527
rect 2053 34493 2087 34527
rect 2789 34493 2823 34527
rect 4537 34493 4571 34527
rect 5181 34493 5215 34527
rect 5273 34493 5307 34527
rect 6193 34493 6227 34527
rect 9505 34493 9539 34527
rect 11805 34493 11839 34527
rect 11897 34493 11931 34527
rect 11989 34493 12023 34527
rect 15853 34493 15887 34527
rect 15945 34493 15979 34527
rect 16037 34493 16071 34527
rect 16957 34493 16991 34527
rect 17049 34493 17083 34527
rect 17141 34493 17175 34527
rect 17877 34493 17911 34527
rect 17969 34493 18003 34527
rect 18061 34493 18095 34527
rect 19993 34493 20027 34527
rect 20249 34493 20283 34527
rect 22477 34493 22511 34527
rect 22569 34493 22603 34527
rect 22673 34493 22707 34527
rect 23489 34493 23523 34527
rect 23581 34493 23615 34527
rect 23673 34493 23707 34527
rect 25421 34493 25455 34527
rect 26065 34493 26099 34527
rect 26709 34493 26743 34527
rect 2605 34425 2639 34459
rect 4353 34425 4387 34459
rect 4997 34425 5031 34459
rect 13369 34425 13403 34459
rect 27261 34425 27295 34459
rect 27997 34425 28031 34459
rect 10885 34357 10919 34391
rect 21373 34357 21407 34391
rect 25881 34357 25915 34391
rect 26525 34357 26559 34391
rect 3893 34153 3927 34187
rect 5273 34153 5307 34187
rect 7297 34153 7331 34187
rect 11069 34153 11103 34187
rect 24685 34153 24719 34187
rect 25973 34153 26007 34187
rect 4537 34085 4571 34119
rect 1869 34017 1903 34051
rect 2053 34017 2087 34051
rect 2605 34017 2639 34051
rect 3801 34017 3835 34051
rect 5181 34017 5215 34051
rect 5365 34017 5399 34051
rect 12817 34085 12851 34119
rect 15117 34085 15151 34119
rect 16405 34085 16439 34119
rect 18061 34085 18095 34119
rect 19257 34085 19291 34119
rect 21281 34085 21315 34119
rect 26709 34085 26743 34119
rect 27905 34085 27939 34119
rect 7656 34017 7690 34051
rect 10977 34017 11011 34051
rect 11161 34017 11195 34051
rect 12633 34017 12667 34051
rect 13369 34017 13403 34051
rect 14013 34017 14047 34051
rect 14749 34017 14783 34051
rect 14841 34017 14875 34051
rect 14933 34017 14967 34051
rect 16037 34017 16071 34051
rect 16129 34017 16163 34051
rect 16221 34017 16255 34051
rect 17693 34017 17727 34051
rect 17785 34017 17819 34051
rect 17877 34017 17911 34051
rect 18889 34017 18923 34051
rect 18981 34017 19015 34051
rect 19073 34017 19107 34051
rect 20877 34017 20911 34051
rect 21005 34017 21039 34051
rect 21097 34017 21131 34051
rect 24869 34017 24903 34051
rect 25513 34017 25547 34051
rect 26157 34017 26191 34051
rect 28089 34017 28123 34051
rect 7297 33949 7331 33983
rect 7389 33949 7423 33983
rect 13553 33949 13587 33983
rect 2789 33881 2823 33915
rect 4629 33813 4663 33847
rect 8769 33813 8803 33847
rect 14197 33813 14231 33847
rect 25329 33813 25363 33847
rect 26801 33813 26835 33847
rect 1593 33609 1627 33643
rect 5089 33609 5123 33643
rect 7849 33609 7883 33643
rect 27261 33609 27295 33643
rect 27997 33609 28031 33643
rect 5733 33541 5767 33575
rect 8493 33473 8527 33507
rect 12817 33473 12851 33507
rect 13737 33473 13771 33507
rect 25605 33473 25639 33507
rect 25973 33473 26007 33507
rect 1501 33405 1535 33439
rect 2421 33405 2455 33439
rect 2697 33405 2731 33439
rect 3157 33405 3191 33439
rect 3341 33405 3375 33439
rect 4997 33405 5031 33439
rect 5641 33405 5675 33439
rect 9689 33405 9723 33439
rect 12725 33405 12759 33439
rect 12909 33405 12943 33439
rect 13369 33405 13403 33439
rect 13553 33405 13587 33439
rect 15025 33405 15059 33439
rect 16037 33405 16071 33439
rect 16773 33405 16807 33439
rect 18153 33405 18187 33439
rect 21465 33405 21499 33439
rect 21741 33405 21775 33439
rect 21833 33405 21867 33439
rect 23673 33405 23707 33439
rect 24041 33405 24075 33439
rect 25789 33405 25823 33439
rect 25881 33405 25915 33439
rect 26065 33405 26099 33439
rect 27169 33405 27203 33439
rect 27905 33405 27939 33439
rect 4353 33337 4387 33371
rect 8217 33337 8251 33371
rect 20085 33337 20119 33371
rect 20269 33337 20303 33371
rect 21649 33337 21683 33371
rect 23857 33337 23891 33371
rect 23949 33337 23983 33371
rect 4445 33269 4479 33303
rect 8309 33269 8343 33303
rect 9873 33269 9907 33303
rect 15209 33269 15243 33303
rect 16221 33269 16255 33303
rect 16957 33269 16991 33303
rect 18337 33269 18371 33303
rect 22017 33269 22051 33303
rect 24225 33269 24259 33303
rect 27997 33065 28031 33099
rect 4905 32997 4939 33031
rect 13093 32997 13127 33031
rect 14473 32997 14507 33031
rect 18153 32997 18187 33031
rect 18981 32997 19015 33031
rect 19073 32997 19107 33031
rect 27905 32997 27939 33031
rect 1501 32929 1535 32963
rect 1869 32929 1903 32963
rect 4169 32929 4203 32963
rect 4813 32929 4847 32963
rect 8677 32929 8711 32963
rect 9505 32929 9539 32963
rect 10701 32929 10735 32963
rect 10885 32929 10919 32963
rect 12173 32929 12207 32963
rect 12265 32929 12299 32963
rect 12357 32929 12391 32963
rect 13001 32929 13035 32963
rect 13185 32929 13219 32963
rect 14105 32929 14139 32963
rect 14289 32929 14323 32963
rect 14381 32929 14415 32963
rect 14565 32929 14599 32963
rect 14749 32929 14783 32963
rect 18797 32929 18831 32963
rect 19165 32929 19199 32963
rect 20637 32929 20671 32963
rect 25053 32929 25087 32963
rect 25237 32929 25271 32963
rect 25329 32929 25363 32963
rect 25421 32929 25455 32963
rect 26433 32929 26467 32963
rect 3985 32861 4019 32895
rect 4077 32861 4111 32895
rect 4261 32861 4295 32895
rect 8769 32861 8803 32895
rect 8861 32861 8895 32895
rect 20269 32861 20303 32895
rect 20453 32861 20487 32895
rect 20545 32861 20579 32895
rect 20729 32861 20763 32895
rect 22569 32861 22603 32895
rect 22845 32861 22879 32895
rect 26249 32861 26283 32895
rect 26341 32861 26375 32895
rect 26525 32861 26559 32895
rect 2697 32793 2731 32827
rect 25605 32793 25639 32827
rect 3801 32725 3835 32759
rect 8309 32725 8343 32759
rect 9597 32725 9631 32759
rect 10793 32725 10827 32759
rect 12541 32725 12575 32759
rect 18245 32725 18279 32759
rect 19349 32725 19383 32759
rect 23949 32725 23983 32759
rect 26065 32725 26099 32759
rect 1501 32521 1535 32555
rect 8401 32521 8435 32555
rect 18521 32521 18555 32555
rect 20821 32521 20855 32555
rect 21281 32521 21315 32555
rect 23029 32521 23063 32555
rect 23673 32521 23707 32555
rect 25789 32521 25823 32555
rect 4813 32453 4847 32487
rect 7205 32453 7239 32487
rect 13645 32453 13679 32487
rect 13829 32453 13863 32487
rect 16129 32453 16163 32487
rect 6469 32385 6503 32419
rect 7757 32385 7791 32419
rect 10057 32385 10091 32419
rect 13369 32385 13403 32419
rect 18705 32385 18739 32419
rect 18981 32385 19015 32419
rect 21557 32385 21591 32419
rect 21741 32385 21775 32419
rect 23857 32385 23891 32419
rect 23949 32385 23983 32419
rect 24041 32385 24075 32419
rect 1777 32317 1811 32351
rect 2053 32317 2087 32351
rect 2513 32317 2547 32351
rect 2881 32317 2915 32351
rect 3065 32317 3099 32351
rect 5089 32317 5123 32351
rect 6285 32317 6319 32351
rect 8309 32317 8343 32351
rect 9873 32317 9907 32351
rect 10977 32317 11011 32351
rect 11069 32317 11103 32351
rect 11161 32317 11195 32351
rect 11345 32317 11379 32351
rect 12081 32317 12115 32351
rect 12173 32317 12207 32351
rect 12265 32317 12299 32351
rect 12449 32317 12483 32351
rect 15945 32317 15979 32351
rect 17417 32317 17451 32351
rect 17785 32317 17819 32351
rect 18797 32317 18831 32351
rect 18889 32317 18923 32351
rect 20269 32317 20303 32351
rect 20453 32317 20487 32351
rect 20637 32317 20671 32351
rect 21465 32317 21499 32351
rect 21640 32317 21674 32351
rect 23213 32317 23247 32351
rect 24133 32317 24167 32351
rect 25237 32317 25271 32351
rect 25605 32317 25639 32351
rect 26801 32317 26835 32351
rect 5365 32249 5399 32283
rect 7481 32249 7515 32283
rect 17601 32249 17635 32283
rect 17693 32249 17727 32283
rect 20545 32249 20579 32283
rect 25421 32249 25455 32283
rect 25513 32249 25547 32283
rect 27068 32249 27102 32283
rect 5273 32181 5307 32215
rect 5917 32181 5951 32215
rect 6377 32181 6411 32215
rect 7665 32181 7699 32215
rect 9505 32181 9539 32215
rect 9965 32181 9999 32215
rect 10701 32181 10735 32215
rect 11805 32181 11839 32215
rect 17969 32181 18003 32215
rect 28181 32181 28215 32215
rect 2053 31977 2087 32011
rect 2421 31977 2455 32011
rect 4905 31977 4939 32011
rect 5273 31977 5307 32011
rect 8861 31977 8895 32011
rect 10701 31977 10735 32011
rect 14565 31977 14599 32011
rect 18337 31977 18371 32011
rect 22753 31977 22787 32011
rect 24133 31977 24167 32011
rect 24961 31977 24995 32011
rect 25973 31977 26007 32011
rect 3240 31909 3274 31943
rect 7849 31909 7883 31943
rect 12909 31909 12943 31943
rect 1409 31841 1443 31875
rect 2237 31841 2271 31875
rect 2513 31841 2547 31875
rect 2973 31841 3007 31875
rect 5365 31841 5399 31875
rect 7067 31841 7101 31875
rect 8769 31841 8803 31875
rect 8953 31841 8987 31875
rect 10517 31841 10551 31875
rect 10701 31841 10735 31875
rect 12173 31841 12207 31875
rect 13553 31841 13587 31875
rect 14289 31841 14323 31875
rect 14565 31841 14599 31875
rect 15117 31841 15151 31875
rect 15807 31841 15841 31875
rect 15945 31841 15979 31875
rect 16037 31841 16071 31875
rect 16221 31841 16255 31875
rect 17325 31841 17359 31875
rect 17509 31841 17543 31875
rect 17601 31841 17635 31875
rect 17693 31841 17727 31875
rect 18521 31841 18555 31875
rect 21245 31841 21279 31875
rect 21373 31841 21407 31875
rect 21465 31841 21499 31875
rect 1501 31773 1535 31807
rect 5549 31773 5583 31807
rect 6929 31773 6963 31807
rect 13093 31773 13127 31807
rect 13645 31773 13679 31807
rect 14197 31773 14231 31807
rect 18613 31773 18647 31807
rect 18705 31773 18739 31807
rect 18797 31773 18831 31807
rect 8125 31705 8159 31739
rect 27905 31909 27939 31943
rect 22937 31841 22971 31875
rect 23029 31841 23063 31875
rect 23121 31841 23155 31875
rect 24317 31841 24351 31875
rect 24869 31841 24903 31875
rect 26157 31841 26191 31875
rect 26709 31841 26743 31875
rect 4353 31637 4387 31671
rect 7297 31637 7331 31671
rect 8309 31637 8343 31671
rect 12357 31637 12391 31671
rect 14197 31637 14231 31671
rect 15577 31637 15611 31671
rect 17877 31637 17911 31671
rect 21649 31637 21683 31671
rect 22753 31637 22787 31671
rect 23305 31637 23339 31671
rect 26801 31637 26835 31671
rect 27997 31637 28031 31671
rect 2605 31433 2639 31467
rect 4721 31433 4755 31467
rect 6377 31433 6411 31467
rect 22201 31433 22235 31467
rect 27537 31433 27571 31467
rect 2513 31365 2547 31399
rect 4629 31365 4663 31399
rect 7297 31365 7331 31399
rect 11161 31365 11195 31399
rect 16773 31365 16807 31399
rect 5733 31297 5767 31331
rect 7389 31297 7423 31331
rect 10057 31297 10091 31331
rect 19993 31297 20027 31331
rect 21373 31297 21407 31331
rect 23673 31297 23707 31331
rect 25513 31297 25547 31331
rect 1501 31229 1535 31263
rect 3157 31229 3191 31263
rect 4261 31229 4295 31263
rect 5641 31229 5675 31263
rect 6285 31229 6319 31263
rect 7849 31229 7883 31263
rect 9781 31229 9815 31263
rect 11897 31229 11931 31263
rect 12265 31229 12299 31263
rect 12541 31229 12575 31263
rect 13001 31229 13035 31263
rect 15393 31229 15427 31263
rect 15649 31229 15683 31263
rect 17325 31229 17359 31263
rect 17601 31229 17635 31263
rect 18889 31229 18923 31263
rect 20269 31229 20303 31263
rect 22477 31229 22511 31263
rect 22569 31229 22603 31263
rect 22661 31229 22695 31263
rect 22845 31229 22879 31263
rect 23949 31229 23983 31263
rect 24041 31229 24075 31263
rect 24133 31229 24167 31263
rect 24317 31229 24351 31263
rect 25237 31229 25271 31263
rect 2145 31161 2179 31195
rect 6929 31161 6963 31195
rect 11989 31161 12023 31195
rect 27445 31161 27479 31195
rect 1593 31093 1627 31127
rect 3249 31093 3283 31127
rect 7941 31093 7975 31127
rect 13185 31093 13219 31127
rect 18981 31093 19015 31127
rect 26617 31093 26651 31127
rect 4721 30889 4755 30923
rect 5365 30821 5399 30855
rect 15577 30821 15611 30855
rect 18521 30821 18555 30855
rect 19165 30821 19199 30855
rect 22845 30821 22879 30855
rect 26709 30821 26743 30855
rect 1869 30753 1903 30787
rect 2605 30753 2639 30787
rect 3801 30753 3835 30787
rect 4629 30753 4663 30787
rect 7573 30753 7607 30787
rect 7941 30753 7975 30787
rect 8033 30753 8067 30787
rect 8401 30753 8435 30787
rect 12173 30753 12207 30787
rect 12357 30753 12391 30787
rect 12449 30753 12483 30787
rect 13737 30753 13771 30787
rect 13921 30753 13955 30787
rect 14289 30753 14323 30787
rect 14565 30753 14599 30787
rect 15209 30753 15243 30787
rect 15301 30753 15335 30787
rect 15393 30753 15427 30787
rect 16129 30753 16163 30787
rect 17509 30753 17543 30787
rect 17785 30753 17819 30787
rect 19441 30753 19475 30787
rect 19533 30753 19567 30787
rect 19625 30753 19659 30787
rect 19809 30753 19843 30787
rect 20821 30753 20855 30787
rect 20913 30753 20947 30787
rect 21005 30753 21039 30787
rect 23121 30753 23155 30787
rect 23213 30753 23247 30787
rect 23305 30753 23339 30787
rect 23489 30753 23523 30787
rect 24225 30753 24259 30787
rect 28181 30753 28215 30787
rect 5549 30685 5583 30719
rect 17325 30685 17359 30719
rect 17601 30685 17635 30719
rect 17693 30685 17727 30719
rect 18705 30685 18739 30719
rect 23949 30685 23983 30719
rect 2789 30617 2823 30651
rect 8677 30617 8711 30651
rect 26893 30617 26927 30651
rect 1961 30549 1995 30583
rect 3985 30549 4019 30583
rect 12449 30549 12483 30583
rect 16221 30549 16255 30583
rect 21189 30549 21223 30583
rect 25329 30549 25363 30583
rect 27997 30549 28031 30583
rect 17693 30345 17727 30379
rect 24041 30345 24075 30379
rect 6101 30277 6135 30311
rect 6745 30277 6779 30311
rect 14841 30277 14875 30311
rect 16589 30277 16623 30311
rect 18981 30277 19015 30311
rect 26157 30277 26191 30311
rect 3341 30209 3375 30243
rect 21465 30209 21499 30243
rect 3065 30141 3099 30175
rect 3157 30141 3191 30175
rect 4813 30141 4847 30175
rect 4905 30141 4939 30175
rect 5089 30141 5123 30175
rect 5549 30141 5583 30175
rect 6009 30141 6043 30175
rect 6653 30141 6687 30175
rect 9597 30141 9631 30175
rect 11989 30141 12023 30175
rect 12357 30141 12391 30175
rect 12817 30141 12851 30175
rect 13277 30141 13311 30175
rect 13461 30141 13495 30175
rect 14749 30141 14783 30175
rect 14933 30141 14967 30175
rect 15669 30141 15703 30175
rect 17509 30141 17543 30175
rect 18613 30141 18647 30175
rect 18705 30141 18739 30175
rect 18797 30141 18831 30175
rect 20637 30141 20671 30175
rect 20729 30141 20763 30175
rect 20821 30141 20855 30175
rect 21005 30141 21039 30175
rect 21741 30141 21775 30175
rect 23673 30141 23707 30175
rect 23765 30141 23799 30175
rect 23857 30141 23891 30175
rect 25697 30141 25731 30175
rect 26341 30141 26375 30175
rect 27997 30141 28031 30175
rect 1869 30073 1903 30107
rect 11897 30073 11931 30107
rect 15853 30073 15887 30107
rect 16405 30073 16439 30107
rect 20361 30073 20395 30107
rect 26893 30073 26927 30107
rect 1961 30005 1995 30039
rect 3341 30005 3375 30039
rect 9689 30005 9723 30039
rect 22845 30005 22879 30039
rect 25513 30005 25547 30039
rect 26985 30005 27019 30039
rect 28089 30005 28123 30039
rect 14381 29801 14415 29835
rect 16037 29801 16071 29835
rect 25973 29801 26007 29835
rect 3402 29733 3436 29767
rect 5641 29733 5675 29767
rect 10425 29733 10459 29767
rect 27997 29733 28031 29767
rect 2145 29665 2179 29699
rect 5549 29665 5583 29699
rect 8484 29665 8518 29699
rect 13737 29665 13771 29699
rect 14289 29665 14323 29699
rect 14473 29665 14507 29699
rect 15117 29665 15151 29699
rect 15209 29665 15243 29699
rect 15301 29665 15335 29699
rect 15485 29665 15519 29699
rect 15945 29665 15979 29699
rect 16129 29665 16163 29699
rect 26157 29665 26191 29699
rect 26709 29665 26743 29699
rect 2237 29597 2271 29631
rect 2329 29597 2363 29631
rect 3157 29597 3191 29631
rect 5733 29597 5767 29631
rect 8217 29597 8251 29631
rect 10517 29597 10551 29631
rect 10609 29597 10643 29631
rect 28181 29597 28215 29631
rect 5181 29529 5215 29563
rect 9597 29529 9631 29563
rect 10057 29529 10091 29563
rect 26893 29529 26927 29563
rect 1777 29461 1811 29495
rect 4537 29461 4571 29495
rect 27997 29257 28031 29291
rect 4261 29189 4295 29223
rect 6837 29189 6871 29223
rect 8033 29189 8067 29223
rect 1409 29121 1443 29155
rect 4813 29121 4847 29155
rect 5457 29121 5491 29155
rect 10701 29121 10735 29155
rect 25697 29121 25731 29155
rect 1676 29053 1710 29087
rect 4629 29053 4663 29087
rect 7941 29053 7975 29087
rect 8217 29053 8251 29087
rect 9781 29053 9815 29087
rect 10793 29053 10827 29087
rect 10977 29053 11011 29087
rect 11437 29053 11471 29087
rect 11897 29053 11931 29087
rect 15025 29053 15059 29087
rect 15301 29053 15335 29087
rect 25513 29053 25547 29087
rect 26985 29053 27019 29087
rect 27629 29053 27663 29087
rect 27997 29053 28031 29087
rect 28181 29053 28215 29087
rect 4721 28985 4755 29019
rect 5724 28985 5758 29019
rect 11989 28985 12023 29019
rect 15209 28985 15243 29019
rect 26249 28985 26283 29019
rect 26433 28985 26467 29019
rect 27169 28985 27203 29019
rect 2789 28917 2823 28951
rect 9873 28917 9907 28951
rect 15301 28917 15335 28951
rect 27721 28917 27755 28951
rect 2605 28713 2639 28747
rect 4445 28713 4479 28747
rect 5089 28713 5123 28747
rect 5825 28713 5859 28747
rect 7941 28713 7975 28747
rect 8401 28713 8435 28747
rect 9137 28713 9171 28747
rect 9505 28713 9539 28747
rect 10793 28713 10827 28747
rect 12173 28713 12207 28747
rect 26801 28713 26835 28747
rect 1869 28645 1903 28679
rect 10701 28645 10735 28679
rect 13829 28645 13863 28679
rect 15485 28645 15519 28679
rect 25666 28645 25700 28679
rect 2513 28577 2547 28611
rect 3157 28577 3191 28611
rect 3341 28577 3375 28611
rect 4353 28577 4387 28611
rect 4997 28577 5031 28611
rect 5733 28577 5767 28611
rect 5917 28577 5951 28611
rect 7113 28577 7147 28611
rect 7205 28577 7239 28611
rect 7297 28577 7331 28611
rect 8309 28577 8343 28611
rect 12081 28577 12115 28611
rect 13737 28577 13771 28611
rect 14013 28577 14047 28611
rect 14197 28577 14231 28611
rect 15209 28577 15243 28611
rect 18981 28577 19015 28611
rect 20260 28577 20294 28611
rect 24777 28577 24811 28611
rect 24961 28577 24995 28611
rect 27997 28577 28031 28611
rect 8585 28509 8619 28543
rect 9597 28509 9631 28543
rect 9781 28509 9815 28543
rect 10977 28509 11011 28543
rect 15485 28509 15519 28543
rect 19993 28509 20027 28543
rect 25421 28509 25455 28543
rect 2053 28441 2087 28475
rect 10333 28441 10367 28475
rect 15301 28441 15335 28475
rect 19165 28441 19199 28475
rect 28181 28441 28215 28475
rect 3249 28373 3283 28407
rect 7481 28373 7515 28407
rect 21373 28373 21407 28407
rect 24869 28373 24903 28407
rect 2697 28169 2731 28203
rect 5089 28169 5123 28203
rect 6193 28169 6227 28203
rect 7941 28169 7975 28203
rect 10149 28169 10183 28203
rect 17233 28169 17267 28203
rect 19441 28169 19475 28203
rect 24225 28169 24259 28203
rect 27997 28169 28031 28203
rect 1777 28101 1811 28135
rect 12265 28101 12299 28135
rect 3157 28033 3191 28067
rect 10793 28033 10827 28067
rect 12081 28033 12115 28067
rect 16681 28033 16715 28067
rect 1961 27965 1995 27999
rect 4261 27965 4295 27999
rect 4905 27965 4939 27999
rect 6101 27965 6135 27999
rect 6285 27965 6319 27999
rect 6929 27965 6963 27999
rect 7113 27965 7147 27999
rect 7205 27965 7239 27999
rect 7665 27965 7699 27999
rect 9505 27965 9539 27999
rect 10517 27965 10551 27999
rect 11989 27965 12023 27999
rect 13093 27965 13127 27999
rect 15301 27965 15335 27999
rect 15577 27965 15611 27999
rect 17877 27965 17911 27999
rect 20913 27965 20947 27999
rect 23857 27965 23891 27999
rect 23995 27965 24029 27999
rect 24133 27965 24167 27999
rect 24317 27965 24351 27999
rect 26341 27965 26375 27999
rect 27721 27965 27755 27999
rect 3249 27897 3283 27931
rect 10609 27897 10643 27931
rect 17969 27897 18003 27931
rect 18337 27897 18371 27931
rect 19441 27897 19475 27931
rect 20177 27897 20211 27931
rect 20453 27897 20487 27931
rect 20545 27897 20579 27931
rect 21281 27897 21315 27931
rect 25881 27897 25915 27931
rect 25973 27897 26007 27931
rect 27445 27897 27479 27931
rect 27813 27897 27847 27931
rect 3157 27829 3191 27863
rect 4353 27829 4387 27863
rect 6745 27829 6779 27863
rect 8125 27829 8159 27863
rect 9597 27829 9631 27863
rect 11621 27829 11655 27863
rect 13185 27829 13219 27863
rect 17601 27829 17635 27863
rect 18705 27829 18739 27863
rect 18889 27829 18923 27863
rect 21465 27829 21499 27863
rect 25605 27829 25639 27863
rect 26709 27829 26743 27863
rect 26893 27829 26927 27863
rect 27629 27829 27663 27863
rect 1593 27625 1627 27659
rect 3433 27625 3467 27659
rect 7205 27625 7239 27659
rect 9137 27625 9171 27659
rect 20177 27625 20211 27659
rect 20361 27625 20395 27659
rect 23857 27625 23891 27659
rect 24777 27625 24811 27659
rect 24869 27625 24903 27659
rect 28018 27625 28052 27659
rect 2697 27557 2731 27591
rect 3801 27557 3835 27591
rect 6929 27557 6963 27591
rect 7113 27557 7147 27591
rect 8493 27557 8527 27591
rect 12081 27557 12115 27591
rect 12725 27557 12759 27591
rect 16221 27557 16255 27591
rect 22753 27557 22787 27591
rect 23121 27557 23155 27591
rect 23535 27557 23569 27591
rect 24593 27557 24627 27591
rect 25697 27557 25731 27591
rect 26709 27557 26743 27591
rect 27813 27557 27847 27591
rect 1869 27489 1903 27523
rect 1961 27489 1995 27523
rect 2329 27489 2363 27523
rect 7205 27489 7239 27523
rect 7665 27489 7699 27523
rect 8401 27489 8435 27523
rect 9045 27489 9079 27523
rect 9229 27489 9263 27523
rect 12449 27489 12483 27523
rect 13277 27489 13311 27523
rect 13369 27489 13403 27523
rect 13473 27489 13507 27523
rect 14657 27489 14691 27523
rect 17693 27489 17727 27523
rect 18337 27489 18371 27523
rect 18521 27489 18555 27523
rect 18981 27489 19015 27523
rect 20085 27489 20119 27523
rect 20637 27489 20671 27523
rect 23029 27489 23063 27523
rect 24961 27489 24995 27523
rect 25605 27489 25639 27523
rect 25831 27489 25865 27523
rect 25973 27489 26007 27523
rect 3893 27421 3927 27455
rect 3985 27421 4019 27455
rect 11529 27421 11563 27455
rect 12541 27421 12575 27455
rect 13645 27421 13679 27455
rect 17785 27421 17819 27455
rect 19625 27421 19659 27455
rect 24041 27353 24075 27387
rect 25145 27353 25179 27387
rect 25973 27353 26007 27387
rect 2881 27285 2915 27319
rect 7849 27285 7883 27319
rect 11529 27285 11563 27319
rect 20545 27285 20579 27319
rect 26801 27285 26835 27319
rect 27997 27285 28031 27319
rect 28181 27285 28215 27319
rect 2421 27081 2455 27115
rect 6009 27081 6043 27115
rect 12357 27081 12391 27115
rect 13001 27081 13035 27115
rect 13645 27081 13679 27115
rect 17509 27081 17543 27115
rect 18797 27081 18831 27115
rect 27537 27081 27571 27115
rect 3249 27013 3283 27047
rect 14841 27013 14875 27047
rect 18521 27013 18555 27047
rect 23581 27013 23615 27047
rect 27261 27013 27295 27047
rect 13093 26945 13127 26979
rect 13829 26945 13863 26979
rect 1961 26877 1995 26911
rect 2605 26877 2639 26911
rect 3065 26877 3099 26911
rect 10885 26877 10919 26911
rect 11989 26877 12023 26911
rect 12081 26877 12115 26911
rect 12173 26877 12207 26911
rect 12817 26877 12851 26911
rect 12909 26877 12943 26911
rect 13553 26877 13587 26911
rect 15025 26877 15059 26911
rect 16497 26877 16531 26911
rect 16589 26877 16623 26911
rect 18797 26877 18831 26911
rect 18981 26877 19015 26911
rect 25329 26877 25363 26911
rect 27537 26877 27571 26911
rect 27721 26877 27755 26911
rect 4997 26809 5031 26843
rect 5089 26809 5123 26843
rect 5457 26809 5491 26843
rect 13829 26809 13863 26843
rect 14749 26809 14783 26843
rect 14933 26809 14967 26843
rect 16221 26809 16255 26843
rect 16957 26809 16991 26843
rect 22569 26809 22603 26843
rect 22661 26809 22695 26843
rect 23029 26809 23063 26843
rect 23397 26809 23431 26843
rect 25513 26809 25547 26843
rect 26617 26809 26651 26843
rect 1777 26741 1811 26775
rect 4721 26741 4755 26775
rect 5825 26741 5859 26775
rect 10977 26741 11011 26775
rect 17325 26741 17359 26775
rect 22293 26741 22327 26775
rect 26709 26741 26743 26775
rect 1777 26537 1811 26571
rect 2513 26537 2547 26571
rect 3249 26537 3283 26571
rect 4537 26537 4571 26571
rect 9873 26537 9907 26571
rect 13001 26537 13035 26571
rect 15209 26537 15243 26571
rect 15945 26537 15979 26571
rect 18521 26537 18555 26571
rect 10977 26469 11011 26503
rect 11069 26469 11103 26503
rect 15301 26469 15335 26503
rect 16037 26469 16071 26503
rect 25973 26469 26007 26503
rect 26893 26469 26927 26503
rect 27997 26469 28031 26503
rect 1961 26401 1995 26435
rect 2421 26401 2455 26435
rect 3065 26401 3099 26435
rect 5365 26401 5399 26435
rect 8033 26401 8067 26435
rect 9045 26401 9079 26435
rect 9229 26401 9263 26435
rect 9321 26401 9355 26435
rect 9781 26401 9815 26435
rect 10793 26401 10827 26435
rect 12817 26401 12851 26435
rect 14473 26401 14507 26435
rect 15117 26401 15151 26435
rect 15393 26401 15427 26435
rect 15853 26401 15887 26435
rect 16129 26401 16163 26435
rect 18429 26401 18463 26435
rect 18613 26401 18647 26435
rect 25237 26401 25271 26435
rect 26709 26401 26743 26435
rect 4629 26333 4663 26367
rect 4813 26333 4847 26367
rect 8125 26333 8159 26367
rect 8401 26333 8435 26367
rect 4169 26265 4203 26299
rect 5549 26265 5583 26299
rect 10517 26265 10551 26299
rect 25421 26265 25455 26299
rect 26157 26265 26191 26299
rect 28181 26265 28215 26299
rect 9045 26197 9079 26231
rect 14565 26197 14599 26231
rect 6745 25993 6779 26027
rect 7481 25993 7515 26027
rect 11437 25993 11471 26027
rect 13277 25993 13311 26027
rect 26341 25993 26375 26027
rect 17693 25925 17727 25959
rect 4445 25857 4479 25891
rect 11897 25857 11931 25891
rect 11989 25857 12023 25891
rect 16313 25857 16347 25891
rect 18705 25857 18739 25891
rect 18981 25857 19015 25891
rect 24317 25857 24351 25891
rect 26065 25857 26099 25891
rect 1869 25789 1903 25823
rect 2973 25789 3007 25823
rect 6929 25789 6963 25823
rect 7389 25789 7423 25823
rect 7757 25789 7791 25823
rect 8309 25789 8343 25823
rect 9505 25789 9539 25823
rect 9761 25789 9795 25823
rect 11805 25789 11839 25823
rect 14749 25789 14783 25823
rect 16589 25789 16623 25823
rect 18613 25789 18647 25823
rect 21189 25789 21223 25823
rect 25973 25789 26007 25823
rect 26801 25789 26835 25823
rect 2053 25721 2087 25755
rect 6653 25721 6687 25755
rect 6837 25721 6871 25755
rect 13185 25721 13219 25755
rect 15669 25721 15703 25755
rect 15853 25721 15887 25755
rect 21434 25721 21468 25755
rect 24133 25721 24167 25755
rect 27068 25721 27102 25755
rect 3157 25653 3191 25687
rect 5457 25653 5491 25687
rect 10885 25653 10919 25687
rect 14933 25653 14967 25687
rect 22569 25653 22603 25687
rect 28181 25653 28215 25687
rect 4813 25449 4847 25483
rect 7941 25449 7975 25483
rect 8493 25449 8527 25483
rect 9321 25449 9355 25483
rect 10701 25449 10735 25483
rect 13185 25449 13219 25483
rect 15393 25449 15427 25483
rect 18337 25449 18371 25483
rect 18705 25449 18739 25483
rect 26617 25449 26651 25483
rect 26801 25449 26835 25483
rect 1777 25381 1811 25415
rect 19778 25381 19812 25415
rect 21465 25381 21499 25415
rect 25513 25381 25547 25415
rect 25881 25381 25915 25415
rect 26249 25381 26283 25415
rect 2513 25313 2547 25347
rect 2789 25313 2823 25347
rect 3985 25313 4019 25347
rect 4721 25313 4755 25347
rect 7757 25313 7791 25347
rect 7941 25313 7975 25347
rect 8401 25313 8435 25347
rect 8585 25313 8619 25347
rect 9229 25313 9263 25347
rect 9413 25313 9447 25347
rect 10609 25313 10643 25347
rect 13093 25313 13127 25347
rect 13993 25313 14027 25347
rect 14086 25313 14120 25347
rect 14202 25313 14236 25347
rect 14381 25313 14415 25347
rect 15669 25313 15703 25347
rect 15761 25313 15795 25347
rect 15853 25313 15887 25347
rect 16037 25313 16071 25347
rect 22569 25313 22603 25347
rect 22661 25313 22695 25347
rect 23121 25313 23155 25347
rect 24501 25313 24535 25347
rect 25789 25313 25823 25347
rect 27997 25313 28031 25347
rect 3433 25245 3467 25279
rect 18797 25245 18831 25279
rect 18981 25245 19015 25279
rect 19533 25245 19567 25279
rect 24593 25245 24627 25279
rect 24777 25245 24811 25279
rect 1961 25177 1995 25211
rect 21649 25177 21683 25211
rect 4169 25109 4203 25143
rect 13737 25109 13771 25143
rect 20913 25109 20947 25143
rect 22937 25109 22971 25143
rect 23029 25109 23063 25143
rect 24133 25109 24167 25143
rect 28089 25109 28123 25143
rect 10241 24905 10275 24939
rect 13185 24905 13219 24939
rect 13737 24905 13771 24939
rect 15577 24905 15611 24939
rect 16129 24905 16163 24939
rect 24133 24905 24167 24939
rect 26617 24905 26651 24939
rect 27445 24905 27479 24939
rect 10701 24769 10735 24803
rect 10793 24769 10827 24803
rect 1869 24701 1903 24735
rect 5089 24701 5123 24735
rect 11989 24701 12023 24735
rect 12081 24701 12115 24735
rect 12173 24701 12207 24735
rect 12357 24701 12391 24735
rect 1593 24633 1627 24667
rect 1961 24633 1995 24667
rect 2329 24633 2363 24667
rect 4721 24633 4755 24667
rect 4997 24633 5031 24667
rect 5457 24633 5491 24667
rect 22293 24837 22327 24871
rect 17785 24769 17819 24803
rect 27997 24769 28031 24803
rect 13369 24701 13403 24735
rect 13461 24701 13495 24735
rect 13553 24701 13587 24735
rect 15173 24701 15207 24735
rect 15301 24701 15335 24735
rect 15393 24701 15427 24735
rect 16405 24701 16439 24735
rect 16497 24701 16531 24735
rect 16589 24701 16623 24735
rect 16773 24701 16807 24735
rect 17601 24701 17635 24735
rect 20453 24701 20487 24735
rect 20913 24701 20947 24735
rect 22109 24701 22143 24735
rect 22753 24701 22787 24735
rect 25237 24701 25271 24735
rect 27813 24701 27847 24735
rect 27905 24701 27939 24735
rect 20177 24633 20211 24667
rect 20545 24633 20579 24667
rect 22998 24633 23032 24667
rect 25482 24633 25516 24667
rect 2697 24565 2731 24599
rect 2881 24565 2915 24599
rect 5825 24565 5859 24599
rect 6009 24565 6043 24599
rect 10609 24565 10643 24599
rect 13185 24565 13219 24599
rect 21281 24565 21315 24599
rect 21465 24565 21499 24599
rect 1777 24361 1811 24395
rect 6929 24361 6963 24395
rect 13277 24361 13311 24395
rect 15209 24361 15243 24395
rect 16405 24361 16439 24395
rect 21373 24361 21407 24395
rect 5181 24293 5215 24327
rect 5273 24293 5307 24327
rect 19717 24293 19751 24327
rect 25973 24293 26007 24327
rect 26157 24293 26191 24327
rect 26709 24293 26743 24327
rect 27997 24293 28031 24327
rect 1961 24225 1995 24259
rect 3148 24225 3182 24259
rect 6837 24225 6871 24259
rect 7389 24225 7423 24259
rect 12357 24225 12391 24259
rect 12449 24225 12483 24259
rect 12541 24225 12575 24259
rect 12725 24225 12759 24259
rect 13185 24225 13219 24259
rect 13369 24225 13403 24259
rect 14105 24225 14139 24259
rect 16001 24225 16035 24259
rect 16129 24225 16163 24259
rect 16221 24225 16255 24259
rect 18061 24225 18095 24259
rect 21465 24225 21499 24259
rect 21649 24225 21683 24259
rect 22569 24225 22603 24259
rect 22753 24225 22787 24259
rect 24133 24225 24167 24259
rect 2881 24157 2915 24191
rect 5365 24157 5399 24191
rect 7665 24157 7699 24191
rect 13829 24157 13863 24191
rect 18337 24157 18371 24191
rect 24225 24157 24259 24191
rect 24501 24157 24535 24191
rect 21189 24089 21223 24123
rect 28181 24089 28215 24123
rect 4261 24021 4295 24055
rect 4813 24021 4847 24055
rect 12081 24021 12115 24055
rect 22661 24021 22695 24055
rect 26801 24021 26835 24055
rect 2513 23817 2547 23851
rect 3157 23817 3191 23851
rect 7113 23817 7147 23851
rect 17785 23817 17819 23851
rect 21281 23817 21315 23851
rect 27997 23817 28031 23851
rect 6469 23749 6503 23783
rect 7941 23749 7975 23783
rect 6561 23681 6595 23715
rect 8401 23681 8435 23715
rect 11713 23681 11747 23715
rect 12817 23681 12851 23715
rect 17325 23681 17359 23715
rect 26249 23681 26283 23715
rect 2697 23613 2731 23647
rect 3341 23613 3375 23647
rect 4261 23613 4295 23647
rect 7021 23613 7055 23647
rect 11437 23613 11471 23647
rect 13645 23613 13679 23647
rect 15485 23613 15519 23647
rect 16957 23613 16991 23647
rect 17049 23613 17083 23647
rect 17141 23613 17175 23647
rect 18061 23613 18095 23647
rect 18153 23613 18187 23647
rect 18245 23613 18279 23647
rect 18429 23613 18463 23647
rect 20913 23613 20947 23647
rect 21051 23613 21085 23647
rect 21189 23613 21223 23647
rect 21373 23613 21407 23647
rect 26709 23613 26743 23647
rect 26893 23613 26927 23647
rect 27353 23613 27387 23647
rect 1869 23545 1903 23579
rect 2053 23545 2087 23579
rect 6101 23545 6135 23579
rect 8493 23545 8527 23579
rect 15669 23545 15703 23579
rect 26065 23545 26099 23579
rect 4445 23477 4479 23511
rect 8401 23477 8435 23511
rect 13737 23477 13771 23511
rect 2513 23273 2547 23307
rect 3249 23273 3283 23307
rect 3617 23273 3651 23307
rect 4813 23273 4847 23307
rect 7297 23273 7331 23307
rect 9689 23273 9723 23307
rect 13645 23273 13679 23307
rect 14381 23273 14415 23307
rect 2053 23205 2087 23239
rect 17693 23205 17727 23239
rect 17877 23205 17911 23239
rect 24961 23205 24995 23239
rect 27997 23205 28031 23239
rect 1869 23137 1903 23171
rect 2697 23137 2731 23171
rect 3709 23137 3743 23171
rect 4721 23137 4755 23171
rect 6837 23137 6871 23171
rect 8116 23137 8150 23171
rect 10057 23137 10091 23171
rect 10149 23137 10183 23171
rect 10885 23137 10919 23171
rect 13553 23137 13587 23171
rect 14289 23137 14323 23171
rect 15025 23137 15059 23171
rect 15669 23137 15703 23171
rect 25697 23137 25731 23171
rect 26525 23137 26559 23171
rect 3893 23069 3927 23103
rect 7849 23069 7883 23103
rect 10241 23069 10275 23103
rect 26617 23069 26651 23103
rect 7113 23001 7147 23035
rect 15209 23001 15243 23035
rect 15853 23001 15887 23035
rect 25145 23001 25179 23035
rect 25881 23001 25915 23035
rect 28181 23001 28215 23035
rect 9229 22933 9263 22967
rect 10977 22933 11011 22967
rect 26893 22933 26927 22967
rect 8493 22729 8527 22763
rect 9597 22729 9631 22763
rect 25513 22729 25547 22763
rect 28181 22729 28215 22763
rect 17785 22661 17819 22695
rect 20177 22661 20211 22695
rect 22753 22661 22787 22695
rect 24225 22661 24259 22695
rect 25375 22661 25409 22695
rect 6745 22593 6779 22627
rect 11621 22593 11655 22627
rect 12541 22593 12575 22627
rect 12725 22593 12759 22627
rect 24041 22593 24075 22627
rect 26801 22593 26835 22627
rect 1409 22525 1443 22559
rect 4261 22525 4295 22559
rect 6653 22525 6687 22559
rect 8401 22525 8435 22559
rect 8585 22525 8619 22559
rect 9505 22525 9539 22559
rect 10885 22525 10919 22559
rect 10977 22525 11011 22559
rect 11161 22525 11195 22559
rect 12449 22525 12483 22559
rect 15577 22525 15611 22559
rect 15669 22525 15703 22559
rect 15761 22525 15795 22559
rect 16405 22525 16439 22559
rect 16681 22525 16715 22559
rect 20361 22525 20395 22559
rect 21649 22525 21683 22559
rect 23857 22525 23891 22559
rect 24225 22525 24259 22559
rect 25237 22525 25271 22559
rect 25697 22525 25731 22559
rect 26157 22525 26191 22559
rect 26341 22525 26375 22559
rect 1676 22457 1710 22491
rect 21373 22457 21407 22491
rect 21557 22457 21591 22491
rect 21925 22457 21959 22491
rect 22569 22457 22603 22491
rect 26249 22457 26283 22491
rect 27068 22457 27102 22491
rect 2789 22389 2823 22423
rect 4353 22389 4387 22423
rect 7481 22389 7515 22423
rect 12081 22389 12115 22423
rect 15945 22389 15979 22423
rect 21741 22389 21775 22423
rect 23949 22389 23983 22423
rect 25605 22389 25639 22423
rect 2053 22185 2087 22219
rect 2421 22185 2455 22219
rect 5733 22185 5767 22219
rect 8125 22185 8159 22219
rect 8585 22185 8619 22219
rect 10241 22185 10275 22219
rect 10885 22185 10919 22219
rect 14657 22185 14691 22219
rect 15761 22185 15795 22219
rect 23857 22185 23891 22219
rect 24041 22185 24075 22219
rect 25329 22185 25363 22219
rect 27905 22185 27939 22219
rect 4445 22117 4479 22151
rect 4721 22117 4755 22151
rect 4813 22117 4847 22151
rect 5549 22117 5583 22151
rect 8493 22117 8527 22151
rect 22753 22117 22787 22151
rect 23121 22117 23155 22151
rect 23489 22117 23523 22151
rect 26065 22117 26099 22151
rect 26433 22117 26467 22151
rect 1593 22049 1627 22083
rect 3249 22049 3283 22083
rect 5181 22049 5215 22083
rect 7021 22049 7055 22083
rect 7113 22049 7147 22083
rect 10149 22049 10183 22083
rect 10793 22049 10827 22083
rect 12137 22049 12171 22083
rect 12265 22049 12299 22083
rect 12357 22049 12391 22083
rect 13277 22049 13311 22083
rect 16017 22049 16051 22083
rect 16110 22049 16144 22083
rect 16221 22049 16255 22083
rect 16405 22049 16439 22083
rect 18337 22049 18371 22083
rect 18604 22049 18638 22083
rect 20729 22049 20763 22083
rect 20913 22049 20947 22083
rect 21097 22049 21131 22083
rect 21373 22049 21407 22083
rect 21649 22049 21683 22083
rect 23029 22049 23063 22083
rect 25605 22049 25639 22083
rect 25697 22049 25731 22083
rect 27813 22049 27847 22083
rect 27997 22049 28031 22083
rect 2513 21981 2547 22015
rect 2605 21981 2639 22015
rect 8769 21981 8803 22015
rect 13553 21981 13587 22015
rect 20545 21981 20579 22015
rect 1409 21913 1443 21947
rect 26617 21913 26651 21947
rect 3341 21845 3375 21879
rect 12541 21845 12575 21879
rect 19717 21845 19751 21879
rect 4721 21641 4755 21675
rect 6929 21641 6963 21675
rect 7021 21641 7055 21675
rect 10241 21641 10275 21675
rect 12541 21641 12575 21675
rect 13001 21641 13035 21675
rect 19073 21641 19107 21675
rect 21465 21641 21499 21675
rect 23765 21641 23799 21675
rect 26617 21641 26651 21675
rect 27445 21641 27479 21675
rect 2881 21573 2915 21607
rect 5365 21505 5399 21539
rect 6745 21505 6779 21539
rect 6929 21505 6963 21539
rect 10885 21505 10919 21539
rect 18797 21505 18831 21539
rect 27997 21505 28031 21539
rect 5181 21437 5215 21471
rect 7113 21437 7147 21471
rect 10609 21437 10643 21471
rect 10701 21437 10735 21471
rect 12137 21437 12171 21471
rect 12265 21437 12299 21471
rect 12357 21437 12391 21471
rect 13231 21437 13265 21471
rect 13369 21437 13403 21471
rect 13461 21437 13495 21471
rect 13639 21437 13673 21471
rect 15577 21437 15611 21471
rect 15669 21437 15703 21471
rect 15761 21437 15795 21471
rect 15945 21437 15979 21471
rect 18889 21437 18923 21471
rect 22385 21437 22419 21471
rect 25237 21437 25271 21471
rect 25504 21437 25538 21471
rect 27813 21437 27847 21471
rect 27905 21437 27939 21471
rect 1593 21369 1627 21403
rect 1869 21369 1903 21403
rect 1961 21369 1995 21403
rect 2329 21369 2363 21403
rect 20453 21369 20487 21403
rect 20545 21369 20579 21403
rect 20913 21369 20947 21403
rect 22630 21369 22664 21403
rect 2697 21301 2731 21335
rect 5089 21301 5123 21335
rect 15301 21301 15335 21335
rect 18429 21301 18463 21335
rect 20177 21301 20211 21335
rect 21281 21301 21315 21335
rect 1501 21097 1535 21131
rect 2697 21097 2731 21131
rect 3341 21097 3375 21131
rect 3709 21097 3743 21131
rect 3801 21097 3835 21131
rect 7021 21097 7055 21131
rect 15393 21097 15427 21131
rect 18245 21097 18279 21131
rect 21097 21097 21131 21131
rect 21465 21097 21499 21131
rect 22569 21097 22603 21131
rect 23029 21097 23063 21131
rect 24317 21097 24351 21131
rect 24501 21097 24535 21131
rect 17969 21029 18003 21063
rect 18153 21029 18187 21063
rect 21306 21029 21340 21063
rect 24225 21029 24259 21063
rect 25605 21029 25639 21063
rect 26709 21029 26743 21063
rect 1685 20961 1719 20995
rect 2789 20961 2823 20995
rect 6837 20961 6871 20995
rect 7113 20961 7147 20995
rect 7297 20961 7331 20995
rect 9229 20961 9263 20995
rect 9689 20961 9723 20995
rect 10793 20961 10827 20995
rect 10885 20961 10919 20995
rect 10977 20961 11011 20995
rect 12357 20961 12391 20995
rect 12449 20961 12483 20995
rect 12546 20961 12580 20995
rect 12725 20961 12759 20995
rect 13553 20961 13587 20995
rect 13645 20961 13679 20995
rect 13737 20961 13771 20995
rect 15025 20961 15059 20995
rect 15117 20961 15151 20995
rect 15209 20961 15243 20995
rect 15853 20961 15887 20995
rect 18245 20961 18279 20995
rect 21189 20961 21223 20995
rect 22937 20961 22971 20995
rect 24133 20961 24167 20995
rect 25421 20961 25455 20995
rect 26893 20961 26927 20995
rect 27997 20961 28031 20995
rect 2697 20893 2731 20927
rect 3893 20893 3927 20927
rect 9965 20893 9999 20927
rect 20821 20893 20855 20927
rect 23121 20893 23155 20927
rect 16037 20825 16071 20859
rect 23949 20825 23983 20859
rect 2237 20757 2271 20791
rect 9045 20757 9079 20791
rect 9781 20757 9815 20791
rect 9873 20757 9907 20791
rect 11161 20757 11195 20791
rect 12081 20757 12115 20791
rect 13921 20757 13955 20791
rect 28089 20757 28123 20791
rect 1777 20553 1811 20587
rect 2973 20553 3007 20587
rect 4537 20553 4571 20587
rect 11345 20553 11379 20587
rect 13277 20553 13311 20587
rect 20821 20553 20855 20587
rect 22017 20553 22051 20587
rect 27353 20553 27387 20587
rect 22477 20485 22511 20519
rect 7665 20417 7699 20451
rect 8125 20417 8159 20451
rect 21557 20417 21591 20451
rect 1961 20349 1995 20383
rect 2881 20349 2915 20383
rect 3065 20349 3099 20383
rect 4445 20349 4479 20383
rect 6101 20349 6135 20383
rect 6377 20349 6411 20383
rect 7757 20349 7791 20383
rect 9965 20349 9999 20383
rect 10221 20349 10255 20383
rect 12403 20349 12437 20383
rect 12522 20349 12556 20383
rect 12633 20349 12667 20383
rect 12817 20349 12851 20383
rect 13461 20349 13495 20383
rect 15025 20349 15059 20383
rect 15117 20349 15151 20383
rect 15209 20349 15243 20383
rect 15393 20349 15427 20383
rect 16681 20349 16715 20383
rect 17049 20349 17083 20383
rect 21005 20349 21039 20383
rect 21649 20349 21683 20383
rect 22661 20349 22695 20383
rect 27261 20349 27295 20383
rect 16589 20281 16623 20315
rect 25789 20281 25823 20315
rect 25973 20281 26007 20315
rect 26525 20281 26559 20315
rect 26709 20281 26743 20315
rect 27997 20281 28031 20315
rect 28181 20281 28215 20315
rect 6745 20213 6779 20247
rect 12173 20213 12207 20247
rect 14749 20213 14783 20247
rect 16313 20213 16347 20247
rect 17417 20213 17451 20247
rect 17601 20213 17635 20247
rect 2513 20009 2547 20043
rect 4537 20009 4571 20043
rect 10057 20009 10091 20043
rect 17325 20009 17359 20043
rect 4629 19941 4663 19975
rect 8217 19941 8251 19975
rect 9321 19941 9355 19975
rect 1869 19873 1903 19907
rect 2697 19873 2731 19907
rect 3157 19873 3191 19907
rect 7297 19873 7331 19907
rect 7481 19873 7515 19907
rect 8125 19873 8159 19907
rect 9137 19873 9171 19907
rect 9413 19873 9447 19907
rect 9965 19873 9999 19907
rect 10149 19873 10183 19907
rect 4721 19805 4755 19839
rect 2053 19737 2087 19771
rect 3341 19737 3375 19771
rect 8861 19737 8895 19771
rect 27997 19941 28031 19975
rect 17601 19873 17635 19907
rect 18869 19873 18903 19907
rect 24961 19873 24995 19907
rect 25697 19873 25731 19907
rect 26525 19873 26559 19907
rect 17693 19805 17727 19839
rect 18613 19805 18647 19839
rect 26617 19805 26651 19839
rect 25881 19737 25915 19771
rect 28181 19737 28215 19771
rect 4169 19669 4203 19703
rect 17325 19669 17359 19703
rect 17969 19669 18003 19703
rect 19993 19669 20027 19703
rect 25053 19669 25087 19703
rect 26893 19669 26927 19703
rect 7205 19465 7239 19499
rect 9505 19465 9539 19499
rect 11897 19465 11931 19499
rect 16129 19465 16163 19499
rect 18245 19465 18279 19499
rect 21465 19465 21499 19499
rect 28181 19465 28215 19499
rect 6285 19397 6319 19431
rect 4721 19329 4755 19363
rect 4813 19329 4847 19363
rect 6009 19329 6043 19363
rect 10149 19329 10183 19363
rect 15025 19329 15059 19363
rect 21306 19329 21340 19363
rect 23857 19329 23891 19363
rect 24317 19329 24351 19363
rect 25789 19329 25823 19363
rect 2513 19261 2547 19295
rect 3157 19261 3191 19295
rect 3341 19261 3375 19295
rect 6929 19261 6963 19295
rect 7205 19261 7239 19295
rect 7389 19261 7423 19295
rect 7849 19261 7883 19295
rect 8953 19261 8987 19295
rect 11253 19261 11287 19295
rect 12081 19261 12115 19295
rect 14749 19261 14783 19295
rect 16865 19261 16899 19295
rect 17141 19261 17175 19295
rect 20821 19261 20855 19295
rect 22109 19261 22143 19295
rect 22201 19261 22235 19295
rect 23949 19261 23983 19295
rect 25605 19261 25639 19295
rect 26801 19261 26835 19295
rect 1869 19193 1903 19227
rect 2053 19193 2087 19227
rect 3249 19193 3283 19227
rect 4629 19193 4663 19227
rect 7941 19193 7975 19227
rect 21925 19193 21959 19227
rect 27068 19193 27102 19227
rect 2697 19125 2731 19159
rect 4261 19125 4295 19159
rect 6469 19125 6503 19159
rect 8953 19125 8987 19159
rect 9873 19125 9907 19159
rect 9965 19125 9999 19159
rect 11345 19125 11379 19159
rect 21097 19125 21131 19159
rect 21189 19125 21223 19159
rect 22023 19125 22057 19159
rect 25237 19125 25271 19159
rect 25697 19125 25731 19159
rect 1593 18921 1627 18955
rect 2881 18921 2915 18955
rect 3617 18921 3651 18955
rect 5457 18921 5491 18955
rect 5641 18921 5675 18955
rect 6929 18921 6963 18955
rect 8125 18921 8159 18955
rect 9873 18921 9907 18955
rect 10885 18921 10919 18955
rect 13645 18921 13679 18955
rect 26525 18921 26559 18955
rect 2697 18853 2731 18887
rect 4353 18853 4387 18887
rect 4629 18853 4663 18887
rect 5089 18853 5123 18887
rect 9045 18853 9079 18887
rect 10793 18853 10827 18887
rect 14933 18853 14967 18887
rect 18521 18853 18555 18887
rect 19257 18853 19291 18887
rect 20361 18853 20395 18887
rect 22753 18853 22787 18887
rect 23857 18853 23891 18887
rect 24685 18853 24719 18887
rect 25421 18853 25455 18887
rect 25697 18853 25731 18887
rect 25789 18853 25823 18887
rect 1869 18785 1903 18819
rect 1961 18785 1995 18819
rect 2329 18785 2363 18819
rect 3433 18785 3467 18819
rect 4721 18785 4755 18819
rect 6837 18785 6871 18819
rect 7941 18785 7975 18819
rect 8125 18785 8159 18819
rect 8953 18785 8987 18819
rect 9781 18785 9815 18819
rect 12541 18785 12575 18819
rect 14749 18785 14783 18819
rect 16313 18785 16347 18819
rect 17509 18785 17543 18819
rect 17785 18785 17819 18819
rect 18153 18785 18187 18819
rect 19533 18785 19567 18819
rect 19625 18785 19659 18819
rect 19993 18785 20027 18819
rect 21189 18785 21223 18819
rect 21327 18785 21361 18819
rect 21649 18785 21683 18819
rect 23029 18785 23063 18819
rect 23121 18785 23155 18819
rect 23489 18785 23523 18819
rect 24593 18785 24627 18819
rect 26157 18785 26191 18819
rect 27997 18785 28031 18819
rect 9229 18717 9263 18751
rect 10977 18717 11011 18751
rect 12265 18717 12299 18751
rect 15025 18717 15059 18751
rect 21465 18717 21499 18751
rect 14473 18649 14507 18683
rect 20545 18649 20579 18683
rect 24041 18649 24075 18683
rect 28181 18649 28215 18683
rect 8585 18581 8619 18615
rect 10425 18581 10459 18615
rect 16129 18581 16163 18615
rect 21557 18581 21591 18615
rect 26709 18581 26743 18615
rect 4353 18377 4387 18411
rect 5457 18377 5491 18411
rect 17141 18377 17175 18411
rect 18337 18377 18371 18411
rect 20821 18377 20855 18411
rect 24133 18377 24167 18411
rect 26617 18377 26651 18411
rect 27445 18377 27479 18411
rect 9689 18309 9723 18343
rect 14841 18309 14875 18343
rect 23673 18309 23707 18343
rect 2421 18241 2455 18275
rect 4905 18241 4939 18275
rect 6009 18241 6043 18275
rect 10977 18241 11011 18275
rect 18797 18241 18831 18275
rect 18981 18241 19015 18275
rect 22293 18241 22327 18275
rect 25237 18241 25271 18275
rect 27905 18241 27939 18275
rect 28089 18241 28123 18275
rect 3065 18173 3099 18207
rect 3249 18173 3283 18207
rect 9505 18173 9539 18207
rect 10241 18173 10275 18207
rect 11621 18173 11655 18207
rect 14749 18173 14783 18207
rect 16221 18173 16255 18207
rect 16589 18173 16623 18207
rect 16971 18173 17005 18207
rect 18705 18173 18739 18207
rect 20729 18173 20763 18207
rect 20913 18173 20947 18207
rect 21189 18173 21223 18207
rect 22549 18173 22583 18207
rect 24133 18173 24167 18207
rect 24317 18173 24351 18207
rect 25493 18173 25527 18207
rect 27813 18173 27847 18207
rect 2237 18105 2271 18139
rect 3157 18105 3191 18139
rect 4629 18105 4663 18139
rect 5825 18105 5859 18139
rect 16129 18105 16163 18139
rect 1869 18037 1903 18071
rect 2329 18037 2363 18071
rect 4813 18037 4847 18071
rect 5917 18037 5951 18071
rect 10333 18037 10367 18071
rect 11989 18037 12023 18071
rect 15853 18037 15887 18071
rect 2789 17833 2823 17867
rect 3249 17833 3283 17867
rect 5263 17833 5297 17867
rect 9689 17833 9723 17867
rect 10241 17833 10275 17867
rect 10701 17833 10735 17867
rect 14197 17833 14231 17867
rect 17509 17833 17543 17867
rect 22661 17833 22695 17867
rect 26065 17833 26099 17867
rect 1676 17765 1710 17799
rect 4537 17765 4571 17799
rect 5733 17765 5767 17799
rect 5825 17765 5859 17799
rect 8576 17765 8610 17799
rect 14657 17765 14691 17799
rect 27997 17765 28031 17799
rect 1409 17697 1443 17731
rect 3617 17697 3651 17731
rect 3709 17697 3743 17731
rect 4445 17697 4479 17731
rect 7021 17697 7055 17731
rect 10609 17697 10643 17731
rect 12081 17697 12115 17731
rect 14565 17697 14599 17731
rect 17785 17697 17819 17731
rect 17969 17697 18003 17731
rect 22569 17697 22603 17731
rect 22753 17697 22787 17731
rect 25973 17697 26007 17731
rect 26709 17697 26743 17731
rect 26893 17697 26927 17731
rect 3893 17629 3927 17663
rect 5733 17629 5767 17663
rect 7113 17629 7147 17663
rect 8309 17629 8343 17663
rect 10885 17629 10919 17663
rect 12357 17629 12391 17663
rect 14749 17629 14783 17663
rect 17693 17629 17727 17663
rect 17877 17629 17911 17663
rect 28181 17561 28215 17595
rect 7389 17493 7423 17527
rect 13461 17493 13495 17527
rect 3065 17289 3099 17323
rect 5181 17289 5215 17323
rect 9689 17289 9723 17323
rect 26893 17289 26927 17323
rect 1777 17221 1811 17255
rect 19993 17221 20027 17255
rect 21649 17221 21683 17255
rect 5825 17153 5859 17187
rect 7573 17153 7607 17187
rect 18981 17153 19015 17187
rect 21281 17153 21315 17187
rect 28089 17153 28123 17187
rect 1961 17085 1995 17119
rect 2973 17085 3007 17119
rect 5549 17085 5583 17119
rect 7297 17085 7331 17119
rect 9597 17085 9631 17119
rect 10977 17085 11011 17119
rect 20177 17085 20211 17119
rect 26065 17085 26099 17119
rect 18797 17017 18831 17051
rect 26249 17017 26283 17051
rect 26801 17017 26835 17051
rect 5641 16949 5675 16983
rect 6929 16949 6963 16983
rect 7389 16949 7423 16983
rect 11161 16949 11195 16983
rect 18337 16949 18371 16983
rect 18705 16949 18739 16983
rect 21741 16949 21775 16983
rect 27445 16949 27479 16983
rect 27813 16949 27847 16983
rect 27905 16949 27939 16983
rect 1777 16745 1811 16779
rect 3065 16745 3099 16779
rect 3893 16745 3927 16779
rect 5089 16745 5123 16779
rect 5733 16745 5767 16779
rect 8309 16745 8343 16779
rect 10517 16745 10551 16779
rect 16221 16745 16255 16779
rect 7174 16677 7208 16711
rect 15086 16677 15120 16711
rect 18766 16677 18800 16711
rect 26709 16677 26743 16711
rect 27997 16677 28031 16711
rect 1961 16609 1995 16643
rect 2605 16609 2639 16643
rect 3249 16609 3283 16643
rect 3709 16609 3743 16643
rect 4997 16609 5031 16643
rect 5641 16609 5675 16643
rect 10333 16609 10367 16643
rect 14841 16609 14875 16643
rect 17601 16609 17635 16643
rect 18521 16609 18555 16643
rect 21005 16609 21039 16643
rect 23857 16609 23891 16643
rect 24952 16609 24986 16643
rect 26893 16609 26927 16643
rect 28181 16609 28215 16643
rect 6929 16541 6963 16575
rect 17693 16541 17727 16575
rect 17969 16541 18003 16575
rect 20913 16541 20947 16575
rect 21097 16541 21131 16575
rect 21189 16541 21223 16575
rect 23949 16541 23983 16575
rect 24225 16541 24259 16575
rect 24685 16541 24719 16575
rect 2421 16473 2455 16507
rect 19901 16405 19935 16439
rect 20729 16405 20763 16439
rect 26065 16405 26099 16439
rect 4997 16201 5031 16235
rect 16957 16201 16991 16235
rect 19441 16201 19475 16235
rect 21649 16201 21683 16235
rect 23581 16201 23615 16235
rect 25237 16201 25271 16235
rect 26893 16201 26927 16235
rect 3157 16133 3191 16167
rect 25789 16065 25823 16099
rect 1869 15997 1903 16031
rect 4905 15997 4939 16031
rect 10793 15997 10827 16031
rect 13461 15997 13495 16031
rect 17509 15997 17543 16031
rect 17601 15997 17635 16031
rect 19441 15997 19475 16031
rect 20269 15997 20303 16031
rect 22661 15997 22695 16031
rect 23029 15997 23063 16031
rect 25605 15997 25639 16031
rect 25697 15997 25731 16031
rect 26709 15997 26743 16031
rect 27261 15997 27295 16031
rect 27537 15997 27571 16031
rect 2789 15929 2823 15963
rect 15945 15929 15979 15963
rect 16037 15929 16071 15963
rect 16405 15929 16439 15963
rect 20536 15929 20570 15963
rect 22569 15929 22603 15963
rect 1961 15861 1995 15895
rect 3249 15861 3283 15895
rect 10885 15861 10919 15895
rect 13277 15861 13311 15895
rect 15669 15861 15703 15895
rect 16773 15861 16807 15895
rect 22293 15861 22327 15895
rect 23397 15861 23431 15895
rect 4997 15657 5031 15691
rect 20085 15657 20119 15691
rect 26249 15657 26283 15691
rect 26433 15657 26467 15691
rect 1869 15589 1903 15623
rect 2053 15589 2087 15623
rect 4077 15589 4111 15623
rect 10977 15589 11011 15623
rect 11069 15589 11103 15623
rect 18981 15589 19015 15623
rect 19236 15589 19270 15623
rect 19337 15589 19371 15623
rect 25145 15589 25179 15623
rect 25421 15589 25455 15623
rect 25513 15589 25547 15623
rect 25881 15589 25915 15623
rect 2973 15521 3007 15555
rect 3985 15521 4019 15555
rect 4353 15521 4387 15555
rect 4813 15521 4847 15555
rect 8576 15521 8610 15555
rect 12081 15521 12115 15555
rect 12337 15521 12371 15555
rect 14177 15521 14211 15555
rect 16037 15521 16071 15555
rect 19717 15521 19751 15555
rect 27997 15521 28031 15555
rect 3433 15453 3467 15487
rect 4169 15453 4203 15487
rect 8309 15453 8343 15487
rect 10977 15453 11011 15487
rect 13921 15453 13955 15487
rect 10517 15385 10551 15419
rect 16221 15385 16255 15419
rect 20269 15385 20303 15419
rect 3249 15317 3283 15351
rect 4353 15317 4387 15351
rect 9689 15317 9723 15351
rect 13461 15317 13495 15351
rect 15301 15317 15335 15351
rect 28089 15317 28123 15351
rect 2881 15113 2915 15147
rect 7021 15113 7055 15147
rect 9505 15113 9539 15147
rect 10701 15113 10735 15147
rect 12081 15113 12115 15147
rect 13185 15113 13219 15147
rect 17693 15113 17727 15147
rect 21925 15113 21959 15147
rect 26341 15113 26375 15147
rect 28181 15113 28215 15147
rect 7573 14977 7607 15011
rect 10057 14977 10091 15011
rect 11161 14977 11195 15011
rect 11345 14977 11379 15011
rect 26065 14977 26099 15011
rect 1869 14909 1903 14943
rect 2329 14909 2363 14943
rect 4261 14909 4295 14943
rect 5457 14909 5491 14943
rect 5917 14909 5951 14943
rect 9873 14909 9907 14943
rect 12357 14909 12391 14943
rect 12449 14909 12483 14943
rect 12541 14909 12575 14943
rect 12725 14909 12759 14943
rect 13415 14909 13449 14943
rect 13553 14909 13587 14943
rect 13645 14909 13679 14943
rect 13829 14909 13863 14943
rect 17325 14909 17359 14943
rect 17417 14909 17451 14943
rect 21649 14909 21683 14943
rect 21787 14909 21821 14943
rect 22109 14909 22143 14943
rect 25973 14909 26007 14943
rect 26801 14909 26835 14943
rect 27068 14909 27102 14943
rect 1593 14841 1627 14875
rect 1949 14841 1983 14875
rect 5549 14841 5583 14875
rect 7481 14841 7515 14875
rect 17141 14841 17175 14875
rect 2697 14773 2731 14807
rect 4353 14773 4387 14807
rect 5181 14773 5215 14807
rect 6285 14773 6319 14807
rect 6469 14773 6503 14807
rect 7389 14773 7423 14807
rect 9965 14773 9999 14807
rect 11069 14773 11103 14807
rect 17509 14773 17543 14807
rect 22109 14773 22143 14807
rect 1777 14569 1811 14603
rect 2421 14569 2455 14603
rect 5273 14569 5307 14603
rect 10149 14569 10183 14603
rect 10977 14569 11011 14603
rect 13553 14569 13587 14603
rect 17693 14569 17727 14603
rect 17877 14569 17911 14603
rect 21097 14569 21131 14603
rect 21373 14569 21407 14603
rect 22661 14569 22695 14603
rect 26893 14569 26927 14603
rect 12449 14501 12483 14535
rect 12633 14501 12667 14535
rect 25789 14501 25823 14535
rect 25973 14501 26007 14535
rect 27997 14501 28031 14535
rect 1961 14433 1995 14467
rect 2605 14433 2639 14467
rect 3525 14433 3559 14467
rect 3709 14433 3743 14467
rect 4261 14433 4295 14467
rect 5089 14433 5123 14467
rect 5365 14433 5399 14467
rect 7481 14433 7515 14467
rect 9045 14433 9079 14467
rect 9137 14433 9171 14467
rect 10057 14433 10091 14467
rect 10885 14433 10919 14467
rect 12725 14433 12759 14467
rect 13369 14433 13403 14467
rect 13553 14433 13587 14467
rect 17509 14433 17543 14467
rect 17601 14433 17635 14467
rect 21005 14433 21039 14467
rect 21189 14433 21223 14467
rect 22569 14433 22603 14467
rect 22753 14433 22787 14467
rect 10241 14365 10275 14399
rect 26433 14365 26467 14399
rect 4261 14297 4295 14331
rect 12173 14297 12207 14331
rect 17325 14297 17359 14331
rect 20821 14297 20855 14331
rect 26801 14297 26835 14331
rect 28181 14297 28215 14331
rect 4905 14229 4939 14263
rect 7573 14229 7607 14263
rect 9689 14229 9723 14263
rect 2329 14025 2363 14059
rect 2881 14025 2915 14059
rect 4721 14025 4755 14059
rect 10977 14025 11011 14059
rect 17141 14025 17175 14059
rect 20545 14025 20579 14059
rect 23765 14025 23799 14059
rect 27353 14025 27387 14059
rect 2237 13957 2271 13991
rect 4629 13957 4663 13991
rect 7941 13957 7975 13991
rect 17049 13957 17083 13991
rect 10517 13889 10551 13923
rect 11437 13889 11471 13923
rect 11621 13889 11655 13923
rect 18889 13889 18923 13923
rect 20729 13889 20763 13923
rect 21097 13889 21131 13923
rect 1869 13821 1903 13855
rect 2421 13821 2455 13855
rect 3065 13821 3099 13855
rect 4261 13821 4295 13855
rect 4813 13821 4847 13855
rect 7113 13821 7147 13855
rect 8033 13821 8067 13855
rect 9781 13821 9815 13855
rect 9873 13821 9907 13855
rect 12173 13821 12207 13855
rect 12357 13821 12391 13855
rect 16681 13821 16715 13855
rect 17601 13821 17635 13855
rect 17693 13821 17727 13855
rect 18797 13821 18831 13855
rect 20821 13821 20855 13855
rect 21189 13821 21223 13855
rect 22385 13821 22419 13855
rect 22641 13821 22675 13855
rect 25789 13821 25823 13855
rect 25973 13821 26007 13855
rect 26709 13821 26743 13855
rect 27261 13821 27295 13855
rect 27997 13821 28031 13855
rect 28181 13821 28215 13855
rect 1961 13753 1995 13787
rect 4353 13753 4387 13787
rect 10011 13753 10045 13787
rect 26525 13753 26559 13787
rect 11345 13685 11379 13719
rect 12265 13685 12299 13719
rect 18337 13685 18371 13719
rect 18705 13685 18739 13719
rect 20913 13685 20947 13719
rect 2697 13481 2731 13515
rect 3249 13481 3283 13515
rect 4077 13481 4111 13515
rect 5089 13481 5123 13515
rect 9137 13481 9171 13515
rect 10517 13481 10551 13515
rect 13553 13481 13587 13515
rect 15485 13481 15519 13515
rect 16313 13481 16347 13515
rect 18153 13481 18187 13515
rect 19993 13481 20027 13515
rect 20821 13481 20855 13515
rect 21005 13481 21039 13515
rect 18858 13413 18892 13447
rect 27997 13413 28031 13447
rect 1869 13345 1903 13379
rect 2605 13345 2639 13379
rect 3433 13345 3467 13379
rect 3985 13345 4019 13379
rect 7665 13345 7699 13379
rect 8309 13345 8343 13379
rect 8953 13345 8987 13379
rect 9137 13345 9171 13379
rect 10425 13345 10459 13379
rect 12440 13345 12474 13379
rect 14361 13345 14395 13379
rect 16129 13345 16163 13379
rect 16405 13345 16439 13379
rect 17785 13345 17819 13379
rect 18613 13345 18647 13379
rect 20729 13345 20763 13379
rect 21097 13345 21131 13379
rect 23857 13345 23891 13379
rect 23949 13345 23983 13379
rect 24133 13345 24167 13379
rect 25217 13345 25251 13379
rect 5181 13277 5215 13311
rect 5365 13277 5399 13311
rect 7757 13277 7791 13311
rect 8493 13277 8527 13311
rect 12173 13277 12207 13311
rect 14105 13277 14139 13311
rect 17693 13277 17727 13311
rect 20913 13277 20947 13311
rect 24961 13277 24995 13311
rect 2053 13209 2087 13243
rect 8217 13209 8251 13243
rect 23949 13209 23983 13243
rect 28181 13209 28215 13243
rect 4721 13141 4755 13175
rect 15945 13141 15979 13175
rect 26341 13141 26375 13175
rect 4353 12937 4387 12971
rect 5089 12937 5123 12971
rect 16773 12937 16807 12971
rect 17693 12937 17727 12971
rect 23857 12937 23891 12971
rect 26709 12937 26743 12971
rect 8493 12869 8527 12903
rect 18797 12869 18831 12903
rect 2053 12801 2087 12835
rect 6653 12801 6687 12835
rect 8217 12801 8251 12835
rect 11069 12801 11103 12835
rect 27905 12801 27939 12835
rect 28089 12801 28123 12835
rect 2513 12733 2547 12767
rect 4261 12733 4295 12767
rect 4997 12733 5031 12767
rect 5917 12733 5951 12767
rect 6009 12733 6043 12767
rect 6193 12733 6227 12767
rect 7205 12733 7239 12767
rect 7481 12733 7515 12767
rect 7849 12733 7883 12767
rect 13645 12733 13679 12767
rect 13829 12733 13863 12767
rect 15761 12733 15795 12767
rect 17417 12733 17451 12767
rect 17509 12733 17543 12767
rect 17877 12733 17911 12767
rect 18521 12733 18555 12767
rect 18809 12733 18843 12767
rect 21741 12733 21775 12767
rect 22937 12733 22971 12767
rect 23305 12733 23339 12767
rect 26157 12733 26191 12767
rect 1869 12665 1903 12699
rect 15485 12665 15519 12699
rect 15853 12665 15887 12699
rect 16221 12665 16255 12699
rect 18705 12665 18739 12699
rect 22845 12665 22879 12699
rect 25421 12665 25455 12699
rect 25697 12665 25731 12699
rect 25789 12665 25823 12699
rect 2697 12597 2731 12631
rect 12081 12597 12115 12631
rect 13829 12597 13863 12631
rect 16589 12597 16623 12631
rect 21557 12597 21591 12631
rect 22569 12597 22603 12631
rect 23673 12597 23707 12631
rect 26525 12597 26559 12631
rect 27445 12597 27479 12631
rect 27813 12597 27847 12631
rect 1593 12393 1627 12427
rect 2881 12393 2915 12427
rect 5825 12393 5859 12427
rect 7205 12393 7239 12427
rect 13829 12393 13863 12427
rect 19165 12393 19199 12427
rect 20453 12393 20487 12427
rect 24501 12393 24535 12427
rect 25329 12393 25363 12427
rect 25421 12393 25455 12427
rect 26893 12393 26927 12427
rect 1869 12325 1903 12359
rect 2697 12325 2731 12359
rect 9413 12325 9447 12359
rect 16037 12325 16071 12359
rect 19533 12325 19567 12359
rect 19901 12325 19935 12359
rect 20269 12325 20303 12359
rect 27997 12325 28031 12359
rect 1961 12257 1995 12291
rect 2329 12257 2363 12291
rect 3433 12257 3467 12291
rect 4077 12257 4111 12291
rect 5733 12257 5767 12291
rect 7573 12257 7607 12291
rect 7665 12257 7699 12291
rect 9229 12257 9263 12291
rect 10241 12257 10275 12291
rect 10977 12257 11011 12291
rect 12613 12257 12647 12291
rect 12725 12257 12759 12291
rect 12817 12257 12851 12291
rect 13001 12257 13035 12291
rect 14105 12257 14139 12291
rect 14197 12257 14231 12291
rect 14289 12257 14323 12291
rect 14473 12257 14507 12291
rect 15393 12257 15427 12291
rect 15577 12257 15611 12291
rect 19441 12257 19475 12291
rect 21281 12257 21315 12291
rect 22017 12257 22051 12291
rect 22753 12257 22787 12291
rect 24133 12257 24167 12291
rect 26525 12257 26559 12291
rect 7389 12189 7423 12223
rect 7481 12189 7515 12223
rect 9505 12189 9539 12223
rect 12357 12189 12391 12223
rect 15301 12189 15335 12223
rect 21189 12189 21223 12223
rect 21373 12189 21407 12223
rect 21465 12189 21499 12223
rect 24225 12189 24259 12223
rect 25605 12189 25639 12223
rect 26433 12189 26467 12223
rect 3617 12121 3651 12155
rect 22017 12121 22051 12155
rect 24961 12121 24995 12155
rect 28181 12121 28215 12155
rect 29009 12121 29043 12155
rect 4721 12053 4755 12087
rect 8953 12053 8987 12087
rect 10333 12053 10367 12087
rect 11069 12053 11103 12087
rect 21005 12053 21039 12087
rect 22569 12053 22603 12087
rect 2605 11849 2639 11883
rect 6377 11849 6411 11883
rect 7573 11849 7607 11883
rect 8309 11849 8343 11883
rect 9597 11849 9631 11883
rect 10793 11849 10827 11883
rect 13001 11849 13035 11883
rect 20545 11849 20579 11883
rect 23765 11849 23799 11883
rect 28181 11849 28215 11883
rect 1777 11781 1811 11815
rect 5825 11781 5859 11815
rect 6929 11713 6963 11747
rect 1961 11645 1995 11679
rect 2421 11645 2455 11679
rect 6745 11645 6779 11679
rect 6837 11645 6871 11679
rect 7573 11645 7607 11679
rect 7849 11645 7883 11679
rect 4813 11577 4847 11611
rect 4905 11577 4939 11611
rect 5273 11577 5307 11611
rect 7757 11577 7791 11611
rect 12357 11781 12391 11815
rect 14749 11781 14783 11815
rect 23581 11781 23615 11815
rect 25605 11781 25639 11815
rect 10149 11713 10183 11747
rect 11253 11713 11287 11747
rect 11437 11713 11471 11747
rect 21465 11713 21499 11747
rect 23305 11713 23339 11747
rect 26341 11713 26375 11747
rect 8401 11645 8435 11679
rect 9965 11645 9999 11679
rect 12265 11645 12299 11679
rect 12449 11645 12483 11679
rect 12909 11645 12943 11679
rect 13737 11645 13771 11679
rect 14197 11645 14231 11679
rect 14933 11645 14967 11679
rect 20729 11645 20763 11679
rect 21005 11645 21039 11679
rect 21721 11645 21755 11679
rect 25421 11645 25455 11679
rect 26801 11645 26835 11679
rect 27068 11645 27102 11679
rect 10057 11577 10091 11611
rect 11161 11577 11195 11611
rect 26157 11577 26191 11611
rect 4537 11509 4571 11543
rect 5641 11509 5675 11543
rect 8309 11509 8343 11543
rect 8493 11509 8527 11543
rect 13553 11509 13587 11543
rect 14197 11509 14231 11543
rect 20913 11509 20947 11543
rect 22845 11509 22879 11543
rect 1777 11305 1811 11339
rect 2421 11305 2455 11339
rect 9965 11305 9999 11339
rect 10793 11305 10827 11339
rect 12081 11305 12115 11339
rect 19717 11305 19751 11339
rect 20269 11305 20303 11339
rect 12449 11237 12483 11271
rect 12541 11237 12575 11271
rect 13829 11237 13863 11271
rect 26709 11237 26743 11271
rect 27997 11237 28031 11271
rect 1961 11169 1995 11203
rect 2605 11169 2639 11203
rect 3249 11169 3283 11203
rect 3433 11169 3467 11203
rect 3525 11169 3559 11203
rect 3985 11169 4019 11203
rect 4997 11169 5031 11203
rect 5089 11169 5123 11203
rect 7573 11169 7607 11203
rect 8217 11169 8251 11203
rect 9873 11169 9907 11203
rect 10701 11169 10735 11203
rect 13645 11169 13679 11203
rect 18061 11169 18095 11203
rect 18889 11169 18923 11203
rect 19625 11169 19659 11203
rect 20453 11169 20487 11203
rect 24225 11169 24259 11203
rect 25053 11169 25087 11203
rect 25973 11169 26007 11203
rect 26157 11169 26191 11203
rect 4077 11101 4111 11135
rect 10057 11101 10091 11135
rect 12633 11101 12667 11135
rect 18153 11101 18187 11135
rect 18337 11101 18371 11135
rect 18981 11101 19015 11135
rect 19165 11101 19199 11135
rect 23581 11101 23615 11135
rect 23949 11101 23983 11135
rect 24041 11101 24075 11135
rect 24869 11101 24903 11135
rect 24961 11101 24995 11135
rect 25145 11101 25179 11135
rect 3065 11033 3099 11067
rect 8401 11033 8435 11067
rect 17693 11033 17727 11067
rect 19073 11033 19107 11067
rect 26893 11033 26927 11067
rect 28181 11033 28215 11067
rect 29009 11033 29043 11067
rect 9505 10965 9539 10999
rect 24685 10965 24719 10999
rect 2053 10761 2087 10795
rect 3065 10761 3099 10795
rect 10885 10761 10919 10795
rect 16405 10761 16439 10795
rect 24225 10761 24259 10795
rect 25697 10761 25731 10795
rect 2881 10693 2915 10727
rect 18429 10693 18463 10727
rect 22753 10693 22787 10727
rect 25605 10693 25639 10727
rect 2605 10625 2639 10659
rect 5273 10625 5307 10659
rect 5457 10625 5491 10659
rect 23581 10625 23615 10659
rect 23949 10625 23983 10659
rect 25237 10625 25271 10659
rect 26801 10625 26835 10659
rect 1961 10557 1995 10591
rect 9505 10557 9539 10591
rect 9772 10557 9806 10591
rect 11529 10557 11563 10591
rect 12771 10557 12805 10591
rect 12890 10557 12924 10591
rect 13001 10557 13035 10591
rect 13197 10557 13231 10591
rect 15485 10557 15519 10591
rect 17509 10557 17543 10591
rect 21741 10557 21775 10591
rect 26157 10557 26191 10591
rect 5181 10489 5215 10523
rect 15393 10489 15427 10523
rect 15899 10489 15933 10523
rect 17141 10489 17175 10523
rect 17417 10489 17451 10523
rect 17877 10489 17911 10523
rect 21833 10489 21867 10523
rect 22201 10489 22235 10523
rect 24066 10489 24100 10523
rect 27068 10489 27102 10523
rect 4813 10421 4847 10455
rect 11345 10421 11379 10455
rect 12541 10421 12575 10455
rect 15117 10421 15151 10455
rect 16221 10421 16255 10455
rect 18245 10421 18279 10455
rect 21465 10421 21499 10455
rect 22569 10421 22603 10455
rect 23857 10421 23891 10455
rect 26249 10421 26283 10455
rect 28181 10421 28215 10455
rect 1409 10217 1443 10251
rect 2973 10217 3007 10251
rect 8125 10217 8159 10251
rect 9229 10217 9263 10251
rect 17877 10217 17911 10251
rect 19717 10217 19751 10251
rect 26801 10217 26835 10251
rect 28089 10217 28123 10251
rect 6929 10149 6963 10183
rect 7113 10149 7147 10183
rect 7665 10149 7699 10183
rect 12694 10149 12728 10183
rect 18613 10149 18647 10183
rect 22845 10149 22879 10183
rect 25666 10149 25700 10183
rect 1593 10081 1627 10115
rect 2053 10081 2087 10115
rect 2237 10081 2271 10115
rect 2973 10081 3007 10115
rect 3433 10081 3467 10115
rect 3709 10081 3743 10115
rect 5181 10081 5215 10115
rect 5365 10081 5399 10115
rect 7205 10081 7239 10115
rect 9045 10081 9079 10115
rect 9229 10081 9263 10115
rect 12449 10081 12483 10115
rect 17509 10081 17543 10115
rect 18889 10081 18923 10115
rect 18981 10081 19015 10115
rect 19395 10081 19429 10115
rect 20453 10081 20487 10115
rect 20729 10081 20763 10115
rect 21097 10081 21131 10115
rect 22753 10081 22787 10115
rect 23673 10081 23707 10115
rect 24225 10081 24259 10115
rect 24501 10081 24535 10115
rect 25421 10081 25455 10115
rect 27905 10081 27939 10115
rect 2421 10013 2455 10047
rect 5089 10013 5123 10047
rect 5825 10013 5859 10047
rect 17601 10013 17635 10047
rect 20821 10013 20855 10047
rect 24777 10013 24811 10047
rect 7941 9945 7975 9979
rect 6929 9877 6963 9911
rect 13829 9877 13863 9911
rect 19901 9877 19935 9911
rect 2881 9673 2915 9707
rect 4721 9673 4755 9707
rect 12449 9673 12483 9707
rect 21925 9673 21959 9707
rect 7021 9605 7055 9639
rect 11161 9605 11195 9639
rect 22937 9605 22971 9639
rect 26801 9605 26835 9639
rect 7665 9537 7699 9571
rect 11805 9537 11839 9571
rect 15761 9537 15795 9571
rect 23397 9537 23431 9571
rect 23581 9537 23615 9571
rect 25789 9537 25823 9571
rect 25973 9537 26007 9571
rect 1869 9469 1903 9503
rect 4261 9469 4295 9503
rect 4813 9469 4847 9503
rect 5641 9469 5675 9503
rect 7757 9469 7791 9503
rect 12357 9469 12391 9503
rect 12541 9469 12575 9503
rect 15025 9469 15059 9503
rect 15117 9469 15151 9503
rect 15301 9469 15335 9503
rect 17325 9469 17359 9503
rect 17592 9469 17626 9503
rect 19993 9469 20027 9503
rect 21833 9469 21867 9503
rect 23305 9469 23339 9503
rect 25697 9469 25731 9503
rect 26617 9469 26651 9503
rect 27169 9469 27203 9503
rect 27445 9469 27479 9503
rect 1961 9401 1995 9435
rect 2329 9401 2363 9435
rect 5908 9401 5942 9435
rect 11529 9401 11563 9435
rect 20238 9401 20272 9435
rect 1593 9333 1627 9367
rect 2697 9333 2731 9367
rect 4353 9333 4387 9367
rect 4537 9333 4571 9367
rect 8125 9333 8159 9367
rect 11621 9333 11655 9367
rect 18705 9333 18739 9367
rect 21373 9333 21407 9367
rect 25329 9333 25363 9367
rect 3249 9129 3283 9163
rect 3433 9129 3467 9163
rect 6837 9129 6871 9163
rect 7205 9129 7239 9163
rect 7297 9129 7331 9163
rect 8953 9129 8987 9163
rect 10425 9129 10459 9163
rect 10793 9129 10827 9163
rect 12173 9129 12207 9163
rect 25789 9129 25823 9163
rect 25881 9129 25915 9163
rect 1869 9061 1903 9095
rect 4353 9061 4387 9095
rect 14381 9061 14415 9095
rect 15209 9061 15243 9095
rect 20545 9061 20579 9095
rect 22661 9061 22695 9095
rect 24041 9061 24075 9095
rect 26617 9061 26651 9095
rect 26801 9061 26835 9095
rect 27997 9061 28031 9095
rect 2513 8993 2547 9027
rect 3157 8993 3191 9027
rect 3525 8993 3559 9027
rect 4261 8993 4295 9027
rect 8769 8993 8803 9027
rect 9597 8993 9631 9027
rect 12081 8993 12115 9027
rect 12725 8993 12759 9027
rect 12817 8993 12851 9027
rect 13737 8993 13771 9027
rect 13921 8993 13955 9027
rect 16037 8993 16071 9027
rect 20453 8993 20487 9027
rect 22569 8993 22603 9027
rect 23305 8993 23339 9027
rect 24777 8993 24811 9027
rect 26893 8993 26927 9027
rect 3341 8925 3375 8959
rect 4169 8925 4203 8959
rect 7481 8925 7515 8959
rect 9045 8925 9079 8959
rect 10885 8925 10919 8959
rect 10977 8925 11011 8959
rect 13645 8925 13679 8959
rect 15301 8925 15335 8959
rect 15485 8925 15519 8959
rect 24225 8925 24259 8959
rect 25973 8925 26007 8959
rect 2605 8857 2639 8891
rect 14841 8857 14875 8891
rect 23397 8857 23431 8891
rect 24961 8857 24995 8891
rect 25421 8857 25455 8891
rect 1961 8789 1995 8823
rect 4169 8789 4203 8823
rect 8493 8789 8527 8823
rect 9781 8789 9815 8823
rect 16129 8789 16163 8823
rect 26893 8789 26927 8823
rect 28089 8789 28123 8823
rect 2605 8585 2639 8619
rect 3065 8585 3099 8619
rect 5641 8585 5675 8619
rect 13369 8585 13403 8619
rect 14841 8585 14875 8619
rect 26985 8585 27019 8619
rect 28181 8585 28215 8619
rect 1777 8517 1811 8551
rect 11805 8517 11839 8551
rect 24225 8517 24259 8551
rect 4261 8449 4295 8483
rect 10057 8449 10091 8483
rect 12265 8449 12299 8483
rect 16129 8449 16163 8483
rect 16865 8449 16899 8483
rect 26341 8449 26375 8483
rect 26709 8449 26743 8483
rect 27537 8449 27571 8483
rect 27905 8449 27939 8483
rect 1961 8381 1995 8415
rect 2421 8381 2455 8415
rect 3249 8381 3283 8415
rect 4528 8381 4562 8415
rect 9965 8381 9999 8415
rect 13277 8381 13311 8415
rect 14749 8381 14783 8415
rect 16221 8381 16255 8415
rect 16405 8381 16439 8415
rect 24133 8381 24167 8415
rect 25697 8381 25731 8415
rect 25881 8381 25915 8415
rect 26801 8381 26835 8415
rect 27997 8381 28031 8415
rect 12219 8313 12253 8347
rect 12357 8313 12391 8347
rect 9505 8245 9539 8279
rect 9873 8245 9907 8279
rect 1777 8041 1811 8075
rect 3249 8041 3283 8075
rect 5181 8041 5215 8075
rect 6929 8041 6963 8075
rect 9137 8041 9171 8075
rect 12081 8041 12115 8075
rect 14473 8041 14507 8075
rect 15669 8041 15703 8075
rect 16129 8041 16163 8075
rect 4261 7973 4295 8007
rect 5273 7973 5307 8007
rect 8033 7973 8067 8007
rect 8953 7973 8987 8007
rect 10425 7973 10459 8007
rect 14841 7973 14875 8007
rect 14933 7973 14967 8007
rect 17877 7973 17911 8007
rect 17969 7973 18003 8007
rect 25973 7973 26007 8007
rect 26157 7973 26191 8007
rect 27997 7973 28031 8007
rect 1961 7905 1995 7939
rect 2421 7905 2455 7939
rect 3065 7905 3099 7939
rect 4169 7905 4203 7939
rect 6837 7905 6871 7939
rect 7941 7905 7975 7939
rect 8125 7905 8159 7939
rect 12449 7905 12483 7939
rect 12541 7905 12575 7939
rect 16037 7905 16071 7939
rect 18705 7905 18739 7939
rect 19349 7905 19383 7939
rect 20729 7905 20763 7939
rect 22937 7905 22971 7939
rect 23949 7905 23983 7939
rect 25237 7905 25271 7939
rect 26709 7905 26743 7939
rect 5365 7837 5399 7871
rect 9229 7837 9263 7871
rect 10333 7837 10367 7871
rect 10517 7837 10551 7871
rect 12725 7837 12759 7871
rect 15025 7837 15059 7871
rect 16221 7837 16255 7871
rect 17785 7837 17819 7871
rect 23029 7837 23063 7871
rect 23121 7837 23155 7871
rect 23857 7837 23891 7871
rect 2605 7769 2639 7803
rect 4813 7769 4847 7803
rect 17417 7769 17451 7803
rect 20913 7769 20947 7803
rect 25329 7769 25363 7803
rect 28181 7769 28215 7803
rect 8677 7701 8711 7735
rect 9965 7701 9999 7735
rect 18797 7701 18831 7735
rect 19441 7701 19475 7735
rect 22569 7701 22603 7735
rect 24225 7701 24259 7735
rect 26801 7701 26835 7735
rect 4997 7497 5031 7531
rect 9597 7497 9631 7531
rect 10425 7497 10459 7531
rect 13645 7497 13679 7531
rect 14197 7497 14231 7531
rect 1685 7429 1719 7463
rect 2329 7361 2363 7395
rect 5641 7361 5675 7395
rect 7297 7361 7331 7395
rect 10977 7361 11011 7395
rect 14197 7361 14231 7395
rect 15853 7497 15887 7531
rect 15945 7497 15979 7531
rect 18521 7497 18555 7531
rect 20637 7497 20671 7531
rect 22661 7497 22695 7531
rect 1593 7293 1627 7327
rect 2237 7293 2271 7327
rect 3065 7293 3099 7327
rect 5457 7293 5491 7327
rect 9505 7293 9539 7327
rect 11621 7293 11655 7327
rect 13461 7293 13495 7327
rect 15025 7293 15059 7327
rect 15114 7293 15148 7327
rect 15209 7293 15243 7327
rect 15393 7293 15427 7327
rect 16497 7361 16531 7395
rect 17141 7361 17175 7395
rect 28089 7361 28123 7395
rect 20545 7293 20579 7327
rect 21649 7293 21683 7327
rect 21741 7293 21775 7327
rect 24225 7293 24259 7327
rect 25329 7293 25363 7327
rect 5365 7225 5399 7259
rect 7113 7225 7147 7259
rect 10793 7225 10827 7259
rect 11713 7225 11747 7259
rect 15853 7225 15887 7259
rect 17386 7225 17420 7259
rect 21373 7225 21407 7259
rect 22109 7225 22143 7259
rect 25596 7225 25630 7259
rect 2881 7157 2915 7191
rect 6745 7157 6779 7191
rect 7205 7157 7239 7191
rect 10885 7157 10919 7191
rect 14749 7157 14783 7191
rect 16313 7157 16347 7191
rect 16405 7157 16439 7191
rect 22477 7157 22511 7191
rect 23949 7157 23983 7191
rect 26709 7157 26743 7191
rect 27445 7157 27479 7191
rect 27813 7157 27847 7191
rect 27905 7157 27939 7191
rect 2697 6953 2731 6987
rect 8769 6953 8803 6987
rect 9597 6953 9631 6987
rect 10609 6953 10643 6987
rect 15669 6953 15703 6987
rect 17325 6953 17359 6987
rect 19993 6953 20027 6987
rect 23121 6953 23155 6987
rect 23857 6953 23891 6987
rect 24961 6953 24995 6987
rect 25697 6953 25731 6987
rect 26065 6953 26099 6987
rect 5549 6885 5583 6919
rect 9689 6885 9723 6919
rect 14556 6885 14590 6919
rect 18705 6885 18739 6919
rect 19441 6885 19475 6919
rect 19809 6885 19843 6919
rect 1501 6817 1535 6851
rect 2329 6817 2363 6851
rect 3157 6817 3191 6851
rect 3249 6817 3283 6851
rect 3985 6817 4019 6851
rect 4445 6817 4479 6851
rect 5641 6817 5675 6851
rect 7389 6817 7423 6851
rect 7656 6817 7690 6851
rect 10425 6817 10459 6851
rect 10609 6817 10643 6851
rect 12265 6817 12299 6851
rect 13277 6817 13311 6851
rect 14289 6817 14323 6851
rect 17601 6817 17635 6851
rect 17693 6817 17727 6851
rect 17785 6817 17819 6851
rect 17969 6817 18003 6851
rect 18981 6817 19015 6851
rect 19073 6817 19107 6851
rect 20821 6817 20855 6851
rect 23029 6817 23063 6851
rect 24133 6817 24167 6851
rect 24225 6817 24259 6851
rect 24593 6817 24627 6851
rect 27997 6817 28031 6851
rect 2237 6749 2271 6783
rect 5825 6749 5859 6783
rect 9781 6749 9815 6783
rect 13369 6749 13403 6783
rect 13553 6749 13587 6783
rect 20913 6749 20947 6783
rect 26157 6749 26191 6783
rect 26249 6749 26283 6783
rect 1593 6681 1627 6715
rect 9229 6681 9263 6715
rect 12909 6681 12943 6715
rect 21189 6681 21223 6715
rect 28181 6681 28215 6715
rect 3801 6613 3835 6647
rect 4629 6613 4663 6647
rect 5181 6613 5215 6647
rect 12357 6613 12391 6647
rect 25145 6613 25179 6647
rect 2881 6409 2915 6443
rect 11253 6409 11287 6443
rect 11345 6409 11379 6443
rect 12173 6409 12207 6443
rect 14933 6409 14967 6443
rect 16037 6409 16071 6443
rect 16773 6409 16807 6443
rect 18797 6409 18831 6443
rect 24225 6409 24259 6443
rect 26249 6409 26283 6443
rect 6561 6341 6595 6375
rect 11253 6273 11287 6307
rect 13461 6273 13495 6307
rect 26065 6273 26099 6307
rect 26801 6273 26835 6307
rect 1869 6205 1903 6239
rect 1961 6205 1995 6239
rect 2329 6205 2363 6239
rect 4261 6205 4295 6239
rect 4905 6205 4939 6239
rect 5825 6205 5859 6239
rect 7113 6205 7147 6239
rect 11437 6205 11471 6239
rect 12081 6205 12115 6239
rect 12725 6205 12759 6239
rect 13553 6205 13587 6239
rect 14841 6205 14875 6239
rect 15025 6205 15059 6239
rect 15945 6205 15979 6239
rect 16681 6205 16715 6239
rect 17601 6205 17635 6239
rect 18705 6205 18739 6239
rect 19993 6205 20027 6239
rect 22017 6205 22051 6239
rect 22284 6205 22318 6239
rect 24133 6205 24167 6239
rect 25973 6205 26007 6239
rect 27068 6205 27102 6239
rect 5917 6137 5951 6171
rect 6837 6137 6871 6171
rect 11069 6137 11103 6171
rect 20238 6137 20272 6171
rect 1593 6069 1627 6103
rect 2697 6069 2731 6103
rect 4445 6069 4479 6103
rect 5089 6069 5123 6103
rect 7021 6069 7055 6103
rect 13829 6069 13863 6103
rect 17693 6069 17727 6103
rect 21373 6069 21407 6103
rect 23397 6069 23431 6103
rect 28181 6069 28215 6103
rect 8585 5865 8619 5899
rect 10977 5865 11011 5899
rect 17509 5865 17543 5899
rect 25329 5865 25363 5899
rect 26065 5865 26099 5899
rect 2237 5797 2271 5831
rect 12326 5797 12360 5831
rect 14013 5797 14047 5831
rect 14749 5797 14783 5831
rect 14933 5797 14967 5831
rect 25237 5797 25271 5831
rect 1593 5729 1627 5763
rect 3433 5729 3467 5763
rect 4261 5729 4295 5763
rect 5365 5729 5399 5763
rect 6837 5729 6871 5763
rect 8401 5729 8435 5763
rect 9689 5729 9723 5763
rect 9873 5729 9907 5763
rect 10517 5729 10551 5763
rect 10977 5729 11011 5763
rect 17325 5729 17359 5763
rect 17509 5729 17543 5763
rect 18521 5729 18555 5763
rect 24041 5729 24075 5763
rect 24685 5729 24719 5763
rect 25973 5729 26007 5763
rect 26709 5729 26743 5763
rect 27997 5729 28031 5763
rect 3341 5661 3375 5695
rect 10057 5661 10091 5695
rect 12081 5661 12115 5695
rect 14197 5661 14231 5695
rect 1685 5593 1719 5627
rect 2513 5593 2547 5627
rect 4445 5593 4479 5627
rect 13461 5593 13495 5627
rect 23857 5593 23891 5627
rect 26893 5593 26927 5627
rect 2697 5525 2731 5559
rect 3801 5525 3835 5559
rect 5549 5525 5583 5559
rect 7021 5525 7055 5559
rect 10655 5525 10689 5559
rect 10793 5525 10827 5559
rect 18337 5525 18371 5559
rect 24501 5525 24535 5559
rect 28089 5525 28123 5559
rect 1777 5321 1811 5355
rect 2697 5321 2731 5355
rect 2973 5321 3007 5355
rect 6561 5321 6595 5355
rect 11161 5321 11195 5355
rect 16497 5321 16531 5355
rect 25789 5321 25823 5355
rect 27169 5321 27203 5355
rect 5825 5253 5859 5287
rect 11529 5253 11563 5287
rect 12173 5253 12207 5287
rect 13829 5253 13863 5287
rect 25605 5253 25639 5287
rect 10701 5185 10735 5219
rect 11621 5185 11655 5219
rect 1961 5117 1995 5151
rect 2973 5117 3007 5151
rect 3157 5117 3191 5151
rect 4445 5117 4479 5151
rect 6377 5117 6411 5151
rect 7021 5117 7055 5151
rect 8217 5117 8251 5151
rect 8401 5117 8435 5151
rect 9965 5117 9999 5151
rect 10425 5117 10459 5151
rect 11345 5117 11379 5151
rect 12081 5117 12115 5151
rect 13645 5117 13679 5151
rect 16405 5117 16439 5151
rect 17601 5117 17635 5151
rect 17785 5117 17819 5151
rect 20177 5117 20211 5151
rect 21281 5117 21315 5151
rect 23673 5117 23707 5151
rect 24133 5117 24167 5151
rect 24317 5117 24351 5151
rect 4690 5049 4724 5083
rect 18337 5049 18371 5083
rect 18521 5049 18555 5083
rect 27537 5185 27571 5219
rect 25697 5117 25731 5151
rect 26433 5049 26467 5083
rect 26617 5049 26651 5083
rect 27721 5049 27755 5083
rect 7205 4981 7239 5015
rect 8309 4981 8343 5015
rect 17785 4981 17819 5015
rect 19993 4981 20027 5015
rect 21097 4981 21131 5015
rect 23489 4981 23523 5015
rect 24317 4981 24351 5015
rect 25605 4981 25639 5015
rect 27629 4981 27663 5015
rect 2421 4777 2455 4811
rect 4537 4777 4571 4811
rect 12449 4777 12483 4811
rect 15209 4777 15243 4811
rect 19625 4777 19659 4811
rect 13829 4709 13863 4743
rect 19993 4709 20027 4743
rect 23397 4709 23431 4743
rect 23581 4709 23615 4743
rect 23673 4709 23707 4743
rect 27997 4709 28031 4743
rect 1961 4641 1995 4675
rect 2605 4641 2639 4675
rect 3249 4641 3283 4675
rect 5549 4641 5583 4675
rect 7021 4641 7055 4675
rect 8125 4641 8159 4675
rect 8769 4641 8803 4675
rect 9045 4641 9079 4675
rect 10149 4641 10183 4675
rect 10609 4641 10643 4675
rect 12357 4641 12391 4675
rect 14473 4641 14507 4675
rect 14657 4641 14691 4675
rect 15117 4641 15151 4675
rect 16037 4641 16071 4675
rect 16129 4641 16163 4675
rect 16221 4641 16255 4675
rect 16405 4641 16439 4675
rect 18153 4641 18187 4675
rect 18245 4641 18279 4675
rect 18337 4641 18371 4675
rect 18521 4641 18555 4675
rect 18981 4641 19015 4675
rect 19165 4641 19199 4675
rect 21281 4641 21315 4675
rect 21370 4641 21404 4675
rect 21465 4641 21499 4675
rect 21649 4641 21683 4675
rect 24501 4641 24535 4675
rect 25677 4641 25711 4675
rect 4629 4573 4663 4607
rect 4721 4573 4755 4607
rect 7113 4573 7147 4607
rect 10885 4573 10919 4607
rect 20085 4573 20119 4607
rect 20177 4573 20211 4607
rect 25421 4573 25455 4607
rect 1777 4505 1811 4539
rect 8309 4505 8343 4539
rect 10057 4505 10091 4539
rect 14013 4505 14047 4539
rect 23121 4505 23155 4539
rect 26801 4505 26835 4539
rect 3065 4437 3099 4471
rect 4169 4437 4203 4471
rect 5365 4437 5399 4471
rect 7389 4437 7423 4471
rect 14565 4437 14599 4471
rect 15761 4437 15795 4471
rect 17877 4437 17911 4471
rect 19073 4437 19107 4471
rect 21005 4437 21039 4471
rect 24593 4437 24627 4471
rect 28089 4437 28123 4471
rect 5641 4233 5675 4267
rect 10885 4233 10919 4267
rect 17325 4233 17359 4267
rect 24225 4233 24259 4267
rect 27445 4233 27479 4267
rect 22017 4165 22051 4199
rect 1685 4097 1719 4131
rect 3249 4097 3283 4131
rect 6653 4097 6687 4131
rect 6837 4097 6871 4131
rect 8585 4097 8619 4131
rect 10057 4097 10091 4131
rect 10241 4097 10275 4131
rect 23029 4097 23063 4131
rect 23121 4097 23155 4131
rect 28089 4097 28123 4131
rect 1593 4029 1627 4063
rect 4261 4029 4295 4063
rect 4517 4029 4551 4063
rect 7941 4029 7975 4063
rect 8217 4029 8251 4063
rect 9965 4029 9999 4063
rect 10793 4029 10827 4063
rect 11713 4029 11747 4063
rect 12265 4029 12299 4063
rect 12449 4029 12483 4063
rect 13139 4029 13173 4063
rect 13277 4029 13311 4063
rect 13369 4029 13403 4063
rect 13553 4029 13587 4063
rect 15025 4029 15059 4063
rect 15114 4029 15148 4063
rect 15209 4029 15243 4063
rect 15393 4029 15427 4063
rect 15945 4029 15979 4063
rect 16201 4029 16235 4063
rect 18659 4029 18693 4063
rect 18797 4029 18831 4063
rect 18889 4029 18923 4063
rect 19073 4029 19107 4063
rect 19993 4029 20027 4063
rect 21925 4029 21959 4063
rect 22109 4029 22143 4063
rect 22293 4029 22327 4063
rect 22937 4029 22971 4063
rect 24133 4029 24167 4063
rect 26065 4029 26099 4063
rect 27997 4029 28031 4063
rect 12357 3961 12391 3995
rect 18429 3961 18463 3995
rect 20238 3961 20272 3995
rect 22385 3961 22419 3995
rect 25421 3961 25455 3995
rect 26310 3961 26344 3995
rect 2605 3893 2639 3927
rect 2973 3893 3007 3927
rect 3065 3893 3099 3927
rect 6193 3893 6227 3927
rect 6561 3893 6595 3927
rect 9597 3893 9631 3927
rect 11529 3893 11563 3927
rect 12909 3893 12943 3927
rect 14749 3893 14783 3927
rect 21373 3893 21407 3927
rect 22293 3893 22327 3927
rect 22569 3893 22603 3927
rect 25513 3893 25547 3927
rect 1685 3689 1719 3723
rect 4169 3689 4203 3723
rect 7205 3689 7239 3723
rect 10701 3689 10735 3723
rect 13829 3689 13863 3723
rect 15761 3689 15795 3723
rect 16405 3689 16439 3723
rect 19717 3689 19751 3723
rect 19901 3689 19935 3723
rect 20361 3689 20395 3723
rect 21281 3689 21315 3723
rect 24593 3689 24627 3723
rect 25329 3689 25363 3723
rect 26801 3689 26835 3723
rect 3034 3621 3068 3655
rect 12716 3621 12750 3655
rect 14648 3621 14682 3655
rect 18214 3621 18248 3655
rect 19533 3621 19567 3655
rect 20269 3621 20303 3655
rect 22661 3621 22695 3655
rect 27997 3621 28031 3655
rect 1593 3553 1627 3587
rect 4997 3553 5031 3587
rect 5089 3553 5123 3587
rect 5457 3553 5491 3587
rect 7297 3553 7331 3587
rect 8401 3553 8435 3587
rect 9413 3553 9447 3587
rect 10609 3553 10643 3587
rect 16221 3553 16255 3587
rect 16405 3553 16439 3587
rect 17325 3553 17359 3587
rect 2789 3485 2823 3519
rect 7481 3485 7515 3519
rect 8493 3485 8527 3519
rect 12449 3485 12483 3519
rect 14381 3485 14415 3519
rect 17969 3485 18003 3519
rect 8769 3417 8803 3451
rect 9505 3417 9539 3451
rect 17417 3417 17451 3451
rect 21097 3553 21131 3587
rect 21281 3553 21315 3587
rect 22569 3553 22603 3587
rect 22753 3553 22787 3587
rect 23469 3553 23503 3587
rect 25559 3553 25593 3587
rect 25678 3553 25712 3587
rect 25794 3553 25828 3587
rect 25973 3553 26007 3587
rect 26709 3553 26743 3587
rect 20453 3485 20487 3519
rect 23213 3485 23247 3519
rect 28181 3417 28215 3451
rect 6837 3349 6871 3383
rect 19349 3349 19383 3383
rect 19533 3349 19567 3383
rect 2881 3145 2915 3179
rect 10885 3145 10919 3179
rect 12817 3145 12851 3179
rect 13553 3145 13587 3179
rect 16405 3145 16439 3179
rect 17049 3145 17083 3179
rect 27445 3145 27479 3179
rect 1869 3077 1903 3111
rect 6469 3077 6503 3111
rect 11529 3077 11563 3111
rect 2605 3009 2639 3043
rect 5089 3009 5123 3043
rect 7021 3009 7055 3043
rect 12173 3009 12207 3043
rect 18981 3077 19015 3111
rect 20085 3077 20119 3111
rect 22385 3077 22419 3111
rect 22937 3077 22971 3111
rect 25329 3077 25363 3111
rect 13737 3009 13771 3043
rect 15393 3009 15427 3043
rect 17693 3009 17727 3043
rect 27905 3009 27939 3043
rect 27997 3009 28031 3043
rect 1685 2941 1719 2975
rect 2513 2941 2547 2975
rect 4261 2941 4295 2975
rect 5356 2941 5390 2975
rect 7277 2941 7311 2975
rect 9505 2941 9539 2975
rect 9761 2941 9795 2975
rect 12725 2941 12759 2975
rect 13553 2941 13587 2975
rect 13645 2941 13679 2975
rect 16313 2941 16347 2975
rect 18245 2941 18279 2975
rect 18337 2941 18371 2975
rect 18889 2941 18923 2975
rect 19993 2941 20027 2975
rect 21005 2941 21039 2975
rect 21261 2941 21295 2975
rect 23167 2941 23201 2975
rect 23305 2941 23339 2975
rect 23397 2941 23431 2975
rect 23581 2941 23615 2975
rect 25585 2941 25619 2975
rect 25678 2941 25712 2975
rect 25794 2941 25828 2975
rect 25973 2941 26007 2975
rect 27813 2941 27847 2975
rect 4353 2873 4387 2907
rect 11897 2873 11931 2907
rect 15209 2873 15243 2907
rect 17417 2873 17451 2907
rect 17509 2873 17543 2907
rect 24133 2873 24167 2907
rect 26801 2873 26835 2907
rect 26985 2873 27019 2907
rect 8401 2805 8435 2839
rect 11989 2805 12023 2839
rect 14841 2805 14875 2839
rect 15301 2805 15335 2839
rect 24225 2805 24259 2839
rect 4353 2601 4387 2635
rect 5089 2601 5123 2635
rect 8401 2601 8435 2635
rect 9597 2601 9631 2635
rect 10241 2601 10275 2635
rect 11253 2601 11287 2635
rect 12357 2601 12391 2635
rect 15025 2601 15059 2635
rect 15577 2601 15611 2635
rect 16221 2601 16255 2635
rect 18245 2601 18279 2635
rect 20269 2601 20303 2635
rect 20913 2601 20947 2635
rect 7941 2533 7975 2567
rect 21649 2533 21683 2567
rect 23121 2533 23155 2567
rect 25697 2533 25731 2567
rect 26433 2533 26467 2567
rect 1869 2465 1903 2499
rect 2605 2465 2639 2499
rect 4261 2465 4295 2499
rect 4905 2465 4939 2499
rect 5733 2465 5767 2499
rect 7573 2465 7607 2499
rect 8585 2465 8619 2499
rect 9781 2465 9815 2499
rect 10425 2465 10459 2499
rect 11161 2465 11195 2499
rect 12265 2465 12299 2499
rect 12909 2465 12943 2499
rect 13829 2465 13863 2499
rect 14933 2465 14967 2499
rect 15761 2465 15795 2499
rect 16405 2465 16439 2499
rect 17785 2465 17819 2499
rect 18429 2465 18463 2499
rect 19349 2465 19383 2499
rect 20453 2465 20487 2499
rect 21105 2465 21139 2499
rect 21557 2465 21591 2499
rect 23029 2465 23063 2499
rect 23765 2465 23799 2499
rect 24501 2465 24535 2499
rect 27169 2465 27203 2499
rect 2789 2397 2823 2431
rect 2053 2329 2087 2363
rect 5917 2329 5951 2363
rect 17601 2329 17635 2363
rect 23949 2329 23983 2363
rect 25881 2329 25915 2363
rect 27353 2329 27387 2363
rect 13001 2261 13035 2295
rect 13921 2261 13955 2295
rect 19165 2261 19199 2295
rect 24593 2261 24627 2295
rect 26525 2261 26559 2295
<< metal1 >>
rect 3878 54000 3884 54052
rect 3936 54040 3942 54052
rect 5902 54040 5908 54052
rect 3936 54012 5908 54040
rect 3936 54000 3942 54012
rect 5902 54000 5908 54012
rect 5960 54000 5966 54052
rect 24026 53864 24032 53916
rect 24084 53904 24090 53916
rect 25038 53904 25044 53916
rect 24084 53876 25044 53904
rect 24084 53864 24090 53876
rect 25038 53864 25044 53876
rect 25096 53864 25102 53916
rect 20714 53728 20720 53780
rect 20772 53768 20778 53780
rect 27062 53768 27068 53780
rect 20772 53740 27068 53768
rect 20772 53728 20778 53740
rect 27062 53728 27068 53740
rect 27120 53728 27126 53780
rect 19150 53660 19156 53712
rect 19208 53700 19214 53712
rect 26694 53700 26700 53712
rect 19208 53672 26700 53700
rect 19208 53660 19214 53672
rect 26694 53660 26700 53672
rect 26752 53660 26758 53712
rect 20898 53592 20904 53644
rect 20956 53632 20962 53644
rect 25682 53632 25688 53644
rect 20956 53604 25688 53632
rect 20956 53592 20962 53604
rect 25682 53592 25688 53604
rect 25740 53592 25746 53644
rect 23198 53524 23204 53576
rect 23256 53564 23262 53576
rect 25498 53564 25504 53576
rect 23256 53536 25504 53564
rect 23256 53524 23262 53536
rect 25498 53524 25504 53536
rect 25556 53524 25562 53576
rect 22830 53456 22836 53508
rect 22888 53496 22894 53508
rect 24854 53496 24860 53508
rect 22888 53468 24860 53496
rect 22888 53456 22894 53468
rect 24854 53456 24860 53468
rect 24912 53456 24918 53508
rect 21174 53388 21180 53440
rect 21232 53428 21238 53440
rect 27246 53428 27252 53440
rect 21232 53400 27252 53428
rect 21232 53388 21238 53400
rect 27246 53388 27252 53400
rect 27304 53388 27310 53440
rect 1104 53338 28888 53360
rect 1104 53286 5614 53338
rect 5666 53286 5678 53338
rect 5730 53286 5742 53338
rect 5794 53286 5806 53338
rect 5858 53286 14878 53338
rect 14930 53286 14942 53338
rect 14994 53286 15006 53338
rect 15058 53286 15070 53338
rect 15122 53286 24142 53338
rect 24194 53286 24206 53338
rect 24258 53286 24270 53338
rect 24322 53286 24334 53338
rect 24386 53286 28888 53338
rect 1104 53264 28888 53286
rect 4338 53184 4344 53236
rect 4396 53224 4402 53236
rect 5169 53227 5227 53233
rect 5169 53224 5181 53227
rect 4396 53196 5181 53224
rect 4396 53184 4402 53196
rect 5169 53193 5181 53196
rect 5215 53193 5227 53227
rect 5169 53187 5227 53193
rect 6086 53184 6092 53236
rect 6144 53224 6150 53236
rect 7101 53227 7159 53233
rect 7101 53224 7113 53227
rect 6144 53196 7113 53224
rect 6144 53184 6150 53196
rect 7101 53193 7113 53196
rect 7147 53193 7159 53227
rect 7101 53187 7159 53193
rect 7834 53184 7840 53236
rect 7892 53224 7898 53236
rect 8021 53227 8079 53233
rect 8021 53224 8033 53227
rect 7892 53196 8033 53224
rect 7892 53184 7898 53196
rect 8021 53193 8033 53196
rect 8067 53193 8079 53227
rect 8021 53187 8079 53193
rect 9582 53184 9588 53236
rect 9640 53224 9646 53236
rect 9769 53227 9827 53233
rect 9769 53224 9781 53227
rect 9640 53196 9781 53224
rect 9640 53184 9646 53196
rect 9769 53193 9781 53196
rect 9815 53193 9827 53227
rect 9769 53187 9827 53193
rect 11422 53184 11428 53236
rect 11480 53224 11486 53236
rect 12437 53227 12495 53233
rect 12437 53224 12449 53227
rect 11480 53196 12449 53224
rect 11480 53184 11486 53196
rect 12437 53193 12449 53196
rect 12483 53193 12495 53227
rect 12437 53187 12495 53193
rect 13170 53184 13176 53236
rect 13228 53224 13234 53236
rect 13357 53227 13415 53233
rect 13357 53224 13369 53227
rect 13228 53196 13369 53224
rect 13228 53184 13234 53196
rect 13357 53193 13369 53196
rect 13403 53193 13415 53227
rect 13357 53187 13415 53193
rect 18414 53184 18420 53236
rect 18472 53224 18478 53236
rect 18601 53227 18659 53233
rect 18601 53224 18613 53227
rect 18472 53196 18613 53224
rect 18472 53184 18478 53196
rect 18601 53193 18613 53196
rect 18647 53193 18659 53227
rect 19150 53224 19156 53236
rect 19111 53196 19156 53224
rect 18601 53187 18659 53193
rect 19150 53184 19156 53196
rect 19208 53184 19214 53236
rect 20162 53184 20168 53236
rect 20220 53224 20226 53236
rect 20441 53227 20499 53233
rect 20441 53224 20453 53227
rect 20220 53196 20453 53224
rect 20220 53184 20226 53196
rect 20441 53193 20453 53196
rect 20487 53193 20499 53227
rect 21174 53224 21180 53236
rect 21135 53196 21180 53224
rect 20441 53187 20499 53193
rect 21174 53184 21180 53196
rect 21232 53184 21238 53236
rect 23198 53224 23204 53236
rect 23159 53196 23204 53224
rect 23198 53184 23204 53196
rect 23256 53184 23262 53236
rect 23750 53184 23756 53236
rect 23808 53224 23814 53236
rect 23937 53227 23995 53233
rect 23937 53224 23949 53227
rect 23808 53196 23949 53224
rect 23808 53184 23814 53196
rect 23937 53193 23949 53196
rect 23983 53193 23995 53227
rect 27890 53224 27896 53236
rect 23937 53187 23995 53193
rect 24504 53196 27896 53224
rect 2590 53116 2596 53168
rect 2648 53156 2654 53168
rect 4525 53159 4583 53165
rect 4525 53156 4537 53159
rect 2648 53128 4537 53156
rect 2648 53116 2654 53128
rect 4525 53125 4537 53128
rect 4571 53125 4583 53159
rect 15194 53156 15200 53168
rect 15155 53128 15200 53156
rect 4525 53119 4583 53125
rect 15194 53116 15200 53128
rect 15252 53116 15258 53168
rect 16666 53156 16672 53168
rect 16627 53128 16672 53156
rect 16666 53116 16672 53128
rect 16724 53116 16730 53168
rect 22002 53156 22008 53168
rect 21963 53128 22008 53156
rect 22002 53116 22008 53128
rect 22060 53116 22066 53168
rect 2774 53088 2780 53100
rect 1872 53060 2780 53088
rect 1872 53029 1900 53060
rect 2774 53048 2780 53060
rect 2832 53048 2838 53100
rect 4062 53048 4068 53100
rect 4120 53088 4126 53100
rect 5997 53091 6055 53097
rect 5997 53088 6009 53091
rect 4120 53060 6009 53088
rect 4120 53048 4126 53060
rect 5997 53057 6009 53060
rect 6043 53057 6055 53091
rect 24026 53088 24032 53100
rect 5997 53051 6055 53057
rect 22066 53060 24032 53088
rect 1857 53023 1915 53029
rect 1857 52989 1869 53023
rect 1903 52989 1915 53023
rect 1857 52983 1915 52989
rect 4341 53023 4399 53029
rect 4341 52989 4353 53023
rect 4387 53020 4399 53023
rect 5350 53020 5356 53032
rect 4387 52992 5356 53020
rect 4387 52989 4399 52992
rect 4341 52983 4399 52989
rect 5350 52980 5356 52992
rect 5408 52980 5414 53032
rect 19337 53023 19395 53029
rect 19337 52989 19349 53023
rect 19383 53020 19395 53023
rect 22066 53020 22094 53060
rect 24026 53048 24032 53060
rect 24084 53048 24090 53100
rect 19383 52992 22094 53020
rect 19383 52989 19395 52992
rect 19337 52983 19395 52989
rect 23290 52980 23296 53032
rect 23348 53020 23354 53032
rect 24504 53020 24532 53196
rect 27890 53184 27896 53196
rect 27948 53184 27954 53236
rect 25593 53159 25651 53165
rect 25593 53125 25605 53159
rect 25639 53156 25651 53159
rect 27982 53156 27988 53168
rect 25639 53128 27988 53156
rect 25639 53125 25651 53128
rect 25593 53119 25651 53125
rect 27982 53116 27988 53128
rect 28040 53116 28046 53168
rect 24854 53048 24860 53100
rect 24912 53088 24918 53100
rect 27246 53088 27252 53100
rect 24912 53060 27252 53088
rect 24912 53048 24918 53060
rect 27246 53048 27252 53060
rect 27304 53048 27310 53100
rect 23348 52992 24532 53020
rect 23348 52980 23354 52992
rect 24578 52980 24584 53032
rect 24636 53020 24642 53032
rect 24673 53023 24731 53029
rect 24673 53020 24685 53023
rect 24636 52992 24685 53020
rect 24636 52980 24642 52992
rect 24673 52989 24685 52992
rect 24719 52989 24731 53023
rect 25774 53020 25780 53032
rect 25735 52992 25780 53020
rect 24673 52983 24731 52989
rect 25774 52980 25780 52992
rect 25832 52980 25838 53032
rect 27062 53020 27068 53032
rect 27023 52992 27068 53020
rect 27062 52980 27068 52992
rect 27120 52980 27126 53032
rect 2777 52955 2835 52961
rect 2777 52921 2789 52955
rect 2823 52952 2835 52955
rect 3970 52952 3976 52964
rect 2823 52924 3976 52952
rect 2823 52921 2835 52924
rect 2777 52915 2835 52921
rect 3970 52912 3976 52924
rect 4028 52912 4034 52964
rect 5077 52955 5135 52961
rect 5077 52921 5089 52955
rect 5123 52921 5135 52955
rect 5810 52952 5816 52964
rect 5771 52924 5816 52952
rect 5077 52915 5135 52921
rect 1949 52887 2007 52893
rect 1949 52853 1961 52887
rect 1995 52884 2007 52887
rect 2038 52884 2044 52896
rect 1995 52856 2044 52884
rect 1995 52853 2007 52856
rect 1949 52847 2007 52853
rect 2038 52844 2044 52856
rect 2096 52844 2102 52896
rect 2866 52884 2872 52896
rect 2827 52856 2872 52884
rect 2866 52844 2872 52856
rect 2924 52844 2930 52896
rect 5092 52884 5120 52915
rect 5810 52912 5816 52924
rect 5868 52912 5874 52964
rect 7006 52952 7012 52964
rect 6967 52924 7012 52952
rect 7006 52912 7012 52924
rect 7064 52912 7070 52964
rect 7834 52912 7840 52964
rect 7892 52952 7898 52964
rect 7929 52955 7987 52961
rect 7929 52952 7941 52955
rect 7892 52924 7941 52952
rect 7892 52912 7898 52924
rect 7929 52921 7941 52924
rect 7975 52921 7987 52955
rect 7929 52915 7987 52921
rect 9677 52955 9735 52961
rect 9677 52921 9689 52955
rect 9723 52952 9735 52955
rect 9950 52952 9956 52964
rect 9723 52924 9956 52952
rect 9723 52921 9735 52924
rect 9677 52915 9735 52921
rect 9950 52912 9956 52924
rect 10008 52912 10014 52964
rect 12066 52912 12072 52964
rect 12124 52952 12130 52964
rect 12345 52955 12403 52961
rect 12345 52952 12357 52955
rect 12124 52924 12357 52952
rect 12124 52912 12130 52924
rect 12345 52921 12357 52924
rect 12391 52921 12403 52955
rect 13262 52952 13268 52964
rect 13223 52924 13268 52952
rect 12345 52915 12403 52921
rect 13262 52912 13268 52924
rect 13320 52912 13326 52964
rect 14366 52912 14372 52964
rect 14424 52952 14430 52964
rect 15013 52955 15071 52961
rect 15013 52952 15025 52955
rect 14424 52924 15025 52952
rect 14424 52912 14430 52924
rect 15013 52921 15025 52924
rect 15059 52921 15071 52955
rect 16482 52952 16488 52964
rect 16443 52924 16488 52952
rect 15013 52915 15071 52921
rect 16482 52912 16488 52924
rect 16540 52912 16546 52964
rect 18506 52952 18512 52964
rect 18467 52924 18512 52952
rect 18506 52912 18512 52924
rect 18564 52912 18570 52964
rect 20346 52952 20352 52964
rect 20307 52924 20352 52952
rect 20346 52912 20352 52924
rect 20404 52912 20410 52964
rect 21085 52955 21143 52961
rect 21085 52921 21097 52955
rect 21131 52921 21143 52955
rect 21085 52915 21143 52921
rect 11514 52884 11520 52896
rect 5092 52856 11520 52884
rect 11514 52844 11520 52856
rect 11572 52844 11578 52896
rect 21100 52884 21128 52915
rect 21634 52912 21640 52964
rect 21692 52952 21698 52964
rect 21821 52955 21879 52961
rect 21821 52952 21833 52955
rect 21692 52924 21833 52952
rect 21692 52912 21698 52924
rect 21821 52921 21833 52924
rect 21867 52921 21879 52955
rect 21821 52915 21879 52921
rect 22094 52912 22100 52964
rect 22152 52952 22158 52964
rect 23109 52955 23167 52961
rect 23109 52952 23121 52955
rect 22152 52924 23121 52952
rect 22152 52912 22158 52924
rect 23109 52921 23121 52924
rect 23155 52921 23167 52955
rect 23109 52915 23167 52921
rect 23750 52912 23756 52964
rect 23808 52952 23814 52964
rect 23845 52955 23903 52961
rect 23845 52952 23857 52955
rect 23808 52924 23857 52952
rect 23808 52912 23814 52924
rect 23845 52921 23857 52924
rect 23891 52921 23903 52955
rect 26234 52952 26240 52964
rect 23845 52915 23903 52921
rect 24412 52924 26240 52952
rect 22002 52884 22008 52896
rect 21100 52856 22008 52884
rect 22002 52844 22008 52856
rect 22060 52844 22066 52896
rect 22646 52844 22652 52896
rect 22704 52884 22710 52896
rect 24412 52884 24440 52924
rect 26234 52912 26240 52924
rect 26292 52912 26298 52964
rect 26329 52955 26387 52961
rect 26329 52921 26341 52955
rect 26375 52952 26387 52955
rect 26602 52952 26608 52964
rect 26375 52924 26608 52952
rect 26375 52921 26387 52924
rect 26329 52915 26387 52921
rect 26602 52912 26608 52924
rect 26660 52912 26666 52964
rect 22704 52856 24440 52884
rect 24489 52887 24547 52893
rect 22704 52844 22710 52856
rect 24489 52853 24501 52887
rect 24535 52884 24547 52887
rect 24670 52884 24676 52896
rect 24535 52856 24676 52884
rect 24535 52853 24547 52856
rect 24489 52847 24547 52853
rect 24670 52844 24676 52856
rect 24728 52844 24734 52896
rect 24762 52844 24768 52896
rect 24820 52884 24826 52896
rect 25498 52884 25504 52896
rect 24820 52856 25504 52884
rect 24820 52844 24826 52856
rect 25498 52844 25504 52856
rect 25556 52844 25562 52896
rect 26418 52884 26424 52896
rect 26379 52856 26424 52884
rect 26418 52844 26424 52856
rect 26476 52844 26482 52896
rect 27154 52884 27160 52896
rect 27115 52856 27160 52884
rect 27154 52844 27160 52856
rect 27212 52844 27218 52896
rect 1104 52794 28888 52816
rect 1104 52742 10246 52794
rect 10298 52742 10310 52794
rect 10362 52742 10374 52794
rect 10426 52742 10438 52794
rect 10490 52742 19510 52794
rect 19562 52742 19574 52794
rect 19626 52742 19638 52794
rect 19690 52742 19702 52794
rect 19754 52742 28888 52794
rect 1104 52720 28888 52742
rect 20073 52683 20131 52689
rect 20073 52649 20085 52683
rect 20119 52649 20131 52683
rect 22646 52680 22652 52692
rect 22607 52652 22652 52680
rect 20073 52643 20131 52649
rect 20088 52612 20116 52643
rect 22646 52640 22652 52652
rect 22704 52640 22710 52692
rect 23290 52680 23296 52692
rect 23251 52652 23296 52680
rect 23290 52640 23296 52652
rect 23348 52640 23354 52692
rect 23937 52683 23995 52689
rect 23937 52649 23949 52683
rect 23983 52680 23995 52683
rect 26510 52680 26516 52692
rect 23983 52652 26516 52680
rect 23983 52649 23995 52652
rect 23937 52643 23995 52649
rect 26510 52640 26516 52652
rect 26568 52640 26574 52692
rect 24854 52612 24860 52624
rect 20088 52584 23428 52612
rect 1854 52544 1860 52556
rect 1815 52516 1860 52544
rect 1854 52504 1860 52516
rect 1912 52504 1918 52556
rect 2590 52544 2596 52556
rect 2551 52516 2596 52544
rect 2590 52504 2596 52516
rect 2648 52504 2654 52556
rect 4062 52553 4068 52556
rect 4056 52507 4068 52553
rect 4120 52544 4126 52556
rect 4120 52516 4156 52544
rect 4062 52504 4068 52507
rect 4120 52504 4126 52516
rect 5166 52504 5172 52556
rect 5224 52544 5230 52556
rect 5629 52547 5687 52553
rect 5629 52544 5641 52547
rect 5224 52516 5641 52544
rect 5224 52504 5230 52516
rect 5629 52513 5641 52516
rect 5675 52513 5687 52547
rect 5629 52507 5687 52513
rect 7377 52547 7435 52553
rect 7377 52513 7389 52547
rect 7423 52544 7435 52547
rect 7558 52544 7564 52556
rect 7423 52516 7564 52544
rect 7423 52513 7435 52516
rect 7377 52507 7435 52513
rect 7558 52504 7564 52516
rect 7616 52504 7622 52556
rect 8205 52547 8263 52553
rect 8205 52513 8217 52547
rect 8251 52513 8263 52547
rect 8205 52507 8263 52513
rect 12529 52547 12587 52553
rect 12529 52513 12541 52547
rect 12575 52544 12587 52547
rect 14090 52544 14096 52556
rect 12575 52516 14096 52544
rect 12575 52513 12587 52516
rect 12529 52507 12587 52513
rect 2774 52436 2780 52488
rect 2832 52476 2838 52488
rect 3786 52476 3792 52488
rect 2832 52448 2877 52476
rect 3747 52448 3792 52476
rect 2832 52436 2838 52448
rect 3786 52436 3792 52448
rect 3844 52436 3850 52488
rect 7469 52479 7527 52485
rect 7469 52445 7481 52479
rect 7515 52476 7527 52479
rect 8018 52476 8024 52488
rect 7515 52448 8024 52476
rect 7515 52445 7527 52448
rect 7469 52439 7527 52445
rect 8018 52436 8024 52448
rect 8076 52436 8082 52488
rect 842 52368 848 52420
rect 900 52408 906 52420
rect 2866 52408 2872 52420
rect 900 52380 2872 52408
rect 900 52368 906 52380
rect 2866 52368 2872 52380
rect 2924 52368 2930 52420
rect 8220 52408 8248 52507
rect 9674 52408 9680 52420
rect 8220 52380 9680 52408
rect 9674 52368 9680 52380
rect 9732 52368 9738 52420
rect 11606 52368 11612 52420
rect 11664 52408 11670 52420
rect 12544 52408 12572 52507
rect 14090 52504 14096 52516
rect 14148 52504 14154 52556
rect 18230 52553 18236 52556
rect 18224 52507 18236 52553
rect 18288 52544 18294 52556
rect 20254 52544 20260 52556
rect 18288 52516 18324 52544
rect 20215 52516 20260 52544
rect 18230 52504 18236 52507
rect 18288 52504 18294 52516
rect 20254 52504 20260 52516
rect 20312 52504 20318 52556
rect 20898 52544 20904 52556
rect 20859 52516 20904 52544
rect 20898 52504 20904 52516
rect 20956 52504 20962 52556
rect 21358 52544 21364 52556
rect 21319 52516 21364 52544
rect 21358 52504 21364 52516
rect 21416 52504 21422 52556
rect 22830 52544 22836 52556
rect 22791 52516 22836 52544
rect 22830 52504 22836 52516
rect 22888 52504 22894 52556
rect 12710 52436 12716 52488
rect 12768 52476 12774 52488
rect 12805 52479 12863 52485
rect 12805 52476 12817 52479
rect 12768 52448 12817 52476
rect 12768 52436 12774 52448
rect 12805 52445 12817 52448
rect 12851 52445 12863 52479
rect 12805 52439 12863 52445
rect 12986 52436 12992 52488
rect 13044 52476 13050 52488
rect 13909 52479 13967 52485
rect 13909 52476 13921 52479
rect 13044 52448 13921 52476
rect 13044 52436 13050 52448
rect 13909 52445 13921 52448
rect 13955 52445 13967 52479
rect 13909 52439 13967 52445
rect 16114 52436 16120 52488
rect 16172 52476 16178 52488
rect 17957 52479 18015 52485
rect 17957 52476 17969 52479
rect 16172 52448 17969 52476
rect 16172 52436 16178 52448
rect 17957 52445 17969 52448
rect 18003 52445 18015 52479
rect 21450 52476 21456 52488
rect 21411 52448 21456 52476
rect 17957 52439 18015 52445
rect 21450 52436 21456 52448
rect 21508 52436 21514 52488
rect 23400 52476 23428 52584
rect 23492 52584 24860 52612
rect 23492 52553 23520 52584
rect 24854 52572 24860 52584
rect 24912 52572 24918 52624
rect 27522 52612 27528 52624
rect 25148 52584 27528 52612
rect 23477 52547 23535 52553
rect 23477 52513 23489 52547
rect 23523 52513 23535 52547
rect 23477 52507 23535 52513
rect 24121 52547 24179 52553
rect 24121 52513 24133 52547
rect 24167 52544 24179 52547
rect 24670 52544 24676 52556
rect 24167 52516 24676 52544
rect 24167 52513 24179 52516
rect 24121 52507 24179 52513
rect 24670 52504 24676 52516
rect 24728 52504 24734 52556
rect 24765 52547 24823 52553
rect 24765 52513 24777 52547
rect 24811 52544 24823 52547
rect 25038 52544 25044 52556
rect 24811 52516 25044 52544
rect 24811 52513 24823 52516
rect 24765 52507 24823 52513
rect 25038 52504 25044 52516
rect 25096 52504 25102 52556
rect 24486 52476 24492 52488
rect 23400 52448 24492 52476
rect 24486 52436 24492 52448
rect 24544 52436 24550 52488
rect 25148 52476 25176 52584
rect 27522 52572 27528 52584
rect 27580 52572 27586 52624
rect 27890 52612 27896 52624
rect 27851 52584 27896 52612
rect 27890 52572 27896 52584
rect 27948 52572 27954 52624
rect 25406 52544 25412 52556
rect 25367 52516 25412 52544
rect 25406 52504 25412 52516
rect 25464 52504 25470 52556
rect 25498 52504 25504 52556
rect 25556 52544 25562 52556
rect 25961 52547 26019 52553
rect 25961 52544 25973 52547
rect 25556 52516 25973 52544
rect 25556 52504 25562 52516
rect 25961 52513 25973 52516
rect 26007 52513 26019 52547
rect 25961 52507 26019 52513
rect 26234 52504 26240 52556
rect 26292 52544 26298 52556
rect 26697 52547 26755 52553
rect 26697 52544 26709 52547
rect 26292 52516 26709 52544
rect 26292 52504 26298 52516
rect 26697 52513 26709 52516
rect 26743 52513 26755 52547
rect 26697 52507 26755 52513
rect 26326 52476 26332 52488
rect 24596 52448 25176 52476
rect 25240 52448 26332 52476
rect 24596 52417 24624 52448
rect 25240 52417 25268 52448
rect 26326 52436 26332 52448
rect 26384 52436 26390 52488
rect 27614 52436 27620 52488
rect 27672 52476 27678 52488
rect 28077 52479 28135 52485
rect 28077 52476 28089 52479
rect 27672 52448 28089 52476
rect 27672 52436 27678 52448
rect 28077 52445 28089 52448
rect 28123 52445 28135 52479
rect 28077 52439 28135 52445
rect 24581 52411 24639 52417
rect 11664 52380 12572 52408
rect 13832 52380 14136 52408
rect 11664 52368 11670 52380
rect 1946 52340 1952 52352
rect 1907 52312 1952 52340
rect 1946 52300 1952 52312
rect 2004 52300 2010 52352
rect 5166 52340 5172 52352
rect 5127 52312 5172 52340
rect 5166 52300 5172 52312
rect 5224 52300 5230 52352
rect 5721 52343 5779 52349
rect 5721 52309 5733 52343
rect 5767 52340 5779 52343
rect 6546 52340 6552 52352
rect 5767 52312 6552 52340
rect 5767 52309 5779 52312
rect 5721 52303 5779 52309
rect 6546 52300 6552 52312
rect 6604 52300 6610 52352
rect 7742 52340 7748 52352
rect 7703 52312 7748 52340
rect 7742 52300 7748 52312
rect 7800 52300 7806 52352
rect 8294 52340 8300 52352
rect 8255 52312 8300 52340
rect 8294 52300 8300 52312
rect 8352 52300 8358 52352
rect 8386 52300 8392 52352
rect 8444 52340 8450 52352
rect 13832 52340 13860 52380
rect 8444 52312 13860 52340
rect 14108 52340 14136 52380
rect 18892 52380 22094 52408
rect 18892 52340 18920 52380
rect 19334 52340 19340 52352
rect 14108 52312 18920 52340
rect 19295 52312 19340 52340
rect 8444 52300 8450 52312
rect 19334 52300 19340 52312
rect 19392 52300 19398 52352
rect 20714 52340 20720 52352
rect 20675 52312 20720 52340
rect 20714 52300 20720 52312
rect 20772 52300 20778 52352
rect 22066 52340 22094 52380
rect 24581 52377 24593 52411
rect 24627 52377 24639 52411
rect 24581 52371 24639 52377
rect 25225 52411 25283 52417
rect 25225 52377 25237 52411
rect 25271 52377 25283 52411
rect 26881 52411 26939 52417
rect 26881 52408 26893 52411
rect 25225 52371 25283 52377
rect 25424 52380 26893 52408
rect 25424 52340 25452 52380
rect 26881 52377 26893 52380
rect 26927 52377 26939 52411
rect 26881 52371 26939 52377
rect 26050 52340 26056 52352
rect 22066 52312 25452 52340
rect 26011 52312 26056 52340
rect 26050 52300 26056 52312
rect 26108 52300 26114 52352
rect 1104 52250 28888 52272
rect 1104 52198 5614 52250
rect 5666 52198 5678 52250
rect 5730 52198 5742 52250
rect 5794 52198 5806 52250
rect 5858 52198 14878 52250
rect 14930 52198 14942 52250
rect 14994 52198 15006 52250
rect 15058 52198 15070 52250
rect 15122 52198 24142 52250
rect 24194 52198 24206 52250
rect 24258 52198 24270 52250
rect 24322 52198 24334 52250
rect 24386 52198 28888 52250
rect 1104 52176 28888 52198
rect 2590 52096 2596 52148
rect 2648 52136 2654 52148
rect 26605 52139 26663 52145
rect 26605 52136 26617 52139
rect 2648 52108 26617 52136
rect 2648 52096 2654 52108
rect 26605 52105 26617 52108
rect 26651 52105 26663 52139
rect 26605 52099 26663 52105
rect 3602 52028 3608 52080
rect 3660 52068 3666 52080
rect 4525 52071 4583 52077
rect 4525 52068 4537 52071
rect 3660 52040 4537 52068
rect 3660 52028 3666 52040
rect 4525 52037 4537 52040
rect 4571 52037 4583 52071
rect 4525 52031 4583 52037
rect 5368 52040 8708 52068
rect 2774 51960 2780 52012
rect 2832 52000 2838 52012
rect 2832 51972 2877 52000
rect 2832 51960 2838 51972
rect 2593 51935 2651 51941
rect 2593 51901 2605 51935
rect 2639 51932 2651 51935
rect 5368 51932 5396 52040
rect 8110 52000 8116 52012
rect 7668 51972 8116 52000
rect 5994 51932 6000 51944
rect 2639 51904 5396 51932
rect 5955 51904 6000 51932
rect 2639 51901 2651 51904
rect 2593 51895 2651 51901
rect 5994 51892 6000 51904
rect 6052 51892 6058 51944
rect 6362 51932 6368 51944
rect 6323 51904 6368 51932
rect 6362 51892 6368 51904
rect 6420 51892 6426 51944
rect 1857 51867 1915 51873
rect 1857 51833 1869 51867
rect 1903 51864 1915 51867
rect 2682 51864 2688 51876
rect 1903 51836 2688 51864
rect 1903 51833 1915 51836
rect 1857 51827 1915 51833
rect 2682 51824 2688 51836
rect 2740 51824 2746 51876
rect 4341 51867 4399 51873
rect 4341 51833 4353 51867
rect 4387 51833 4399 51867
rect 7558 51864 7564 51876
rect 6670 51836 7564 51864
rect 4341 51827 4399 51833
rect 1486 51756 1492 51808
rect 1544 51796 1550 51808
rect 1949 51799 2007 51805
rect 1949 51796 1961 51799
rect 1544 51768 1961 51796
rect 1544 51756 1550 51768
rect 1949 51765 1961 51768
rect 1995 51765 2007 51799
rect 4356 51796 4384 51827
rect 7558 51824 7564 51836
rect 7616 51824 7622 51876
rect 7668 51796 7696 51972
rect 8110 51960 8116 51972
rect 8168 51960 8174 52012
rect 8478 52009 8484 52012
rect 8435 52003 8484 52009
rect 8435 51969 8447 52003
rect 8481 51969 8484 52003
rect 8435 51963 8484 51969
rect 8478 51960 8484 51963
rect 8536 51960 8542 52012
rect 8680 52000 8708 52040
rect 10594 52028 10600 52080
rect 10652 52068 10658 52080
rect 10652 52040 11468 52068
rect 10652 52028 10658 52040
rect 8680 51972 11376 52000
rect 7742 51892 7748 51944
rect 7800 51932 7806 51944
rect 8205 51935 8263 51941
rect 8205 51932 8217 51935
rect 7800 51904 8217 51932
rect 7800 51892 7806 51904
rect 8205 51901 8217 51904
rect 8251 51901 8263 51935
rect 8205 51895 8263 51901
rect 9493 51935 9551 51941
rect 9493 51901 9505 51935
rect 9539 51901 9551 51935
rect 9766 51932 9772 51944
rect 9727 51904 9772 51932
rect 9493 51895 9551 51901
rect 7926 51824 7932 51876
rect 7984 51864 7990 51876
rect 9508 51864 9536 51895
rect 9766 51892 9772 51904
rect 9824 51892 9830 51944
rect 7984 51836 9536 51864
rect 11149 51867 11207 51873
rect 7984 51824 7990 51836
rect 11149 51833 11161 51867
rect 11195 51864 11207 51867
rect 11238 51864 11244 51876
rect 11195 51836 11244 51864
rect 11195 51833 11207 51836
rect 11149 51827 11207 51833
rect 11238 51824 11244 51836
rect 11296 51824 11302 51876
rect 11348 51864 11376 51972
rect 11440 51932 11468 52040
rect 22922 52028 22928 52080
rect 22980 52068 22986 52080
rect 23201 52071 23259 52077
rect 23201 52068 23213 52071
rect 22980 52040 23213 52068
rect 22980 52028 22986 52040
rect 23201 52037 23213 52040
rect 23247 52068 23259 52071
rect 23247 52040 23704 52068
rect 23247 52037 23259 52040
rect 23201 52031 23259 52037
rect 11606 52000 11612 52012
rect 11567 51972 11612 52000
rect 11606 51960 11612 51972
rect 11664 51960 11670 52012
rect 14642 52000 14648 52012
rect 13648 51972 14648 52000
rect 11865 51935 11923 51941
rect 11865 51932 11877 51935
rect 11440 51904 11877 51932
rect 11865 51901 11877 51904
rect 11911 51901 11923 51935
rect 11865 51895 11923 51901
rect 12158 51892 12164 51944
rect 12216 51932 12222 51944
rect 13648 51932 13676 51972
rect 14642 51960 14648 51972
rect 14700 52000 14706 52012
rect 15289 52003 15347 52009
rect 15289 52000 15301 52003
rect 14700 51972 15301 52000
rect 14700 51960 14706 51972
rect 15289 51969 15301 51972
rect 15335 51969 15347 52003
rect 15289 51963 15347 51969
rect 15470 51960 15476 52012
rect 15528 52000 15534 52012
rect 16114 52000 16120 52012
rect 15528 51972 16120 52000
rect 15528 51960 15534 51972
rect 16114 51960 16120 51972
rect 16172 51960 16178 52012
rect 19981 51935 20039 51941
rect 12216 51904 13676 51932
rect 13740 51904 15332 51932
rect 12216 51892 12222 51904
rect 13740 51864 13768 51904
rect 11348 51836 13768 51864
rect 13814 51824 13820 51876
rect 13872 51864 13878 51876
rect 15197 51867 15255 51873
rect 15197 51864 15209 51867
rect 13872 51836 15209 51864
rect 13872 51824 13878 51836
rect 15197 51833 15209 51836
rect 15243 51833 15255 51867
rect 15197 51827 15255 51833
rect 4356 51768 7696 51796
rect 7837 51799 7895 51805
rect 1949 51759 2007 51765
rect 7837 51765 7849 51799
rect 7883 51796 7895 51799
rect 8202 51796 8208 51808
rect 7883 51768 8208 51796
rect 7883 51765 7895 51768
rect 7837 51759 7895 51765
rect 8202 51756 8208 51768
rect 8260 51756 8266 51808
rect 8297 51799 8355 51805
rect 8297 51765 8309 51799
rect 8343 51796 8355 51799
rect 9582 51796 9588 51808
rect 8343 51768 9588 51796
rect 8343 51765 8355 51768
rect 8297 51759 8355 51765
rect 9582 51756 9588 51768
rect 9640 51756 9646 51808
rect 10778 51756 10784 51808
rect 10836 51796 10842 51808
rect 12989 51799 13047 51805
rect 12989 51796 13001 51799
rect 10836 51768 13001 51796
rect 10836 51756 10842 51768
rect 12989 51765 13001 51768
rect 13035 51796 13047 51799
rect 13630 51796 13636 51808
rect 13035 51768 13636 51796
rect 13035 51765 13047 51768
rect 12989 51759 13047 51765
rect 13630 51756 13636 51768
rect 13688 51756 13694 51808
rect 14734 51796 14740 51808
rect 14695 51768 14740 51796
rect 14734 51756 14740 51768
rect 14792 51756 14798 51808
rect 15102 51796 15108 51808
rect 15063 51768 15108 51796
rect 15102 51756 15108 51768
rect 15160 51756 15166 51808
rect 15304 51796 15332 51904
rect 19981 51901 19993 51935
rect 20027 51932 20039 51935
rect 21818 51932 21824 51944
rect 20027 51904 21824 51932
rect 20027 51901 20039 51904
rect 19981 51895 20039 51901
rect 21818 51892 21824 51904
rect 21876 51892 21882 51944
rect 23676 51941 23704 52040
rect 23842 52028 23848 52080
rect 23900 52068 23906 52080
rect 28994 52068 29000 52080
rect 23900 52040 29000 52068
rect 23900 52028 23906 52040
rect 28994 52028 29000 52040
rect 29052 52028 29058 52080
rect 27433 52003 27491 52009
rect 27433 52000 27445 52003
rect 23768 51972 27445 52000
rect 23661 51935 23719 51941
rect 21928 51904 23612 51932
rect 16390 51873 16396 51876
rect 16384 51827 16396 51873
rect 16448 51864 16454 51876
rect 20248 51867 20306 51873
rect 16448 51836 16484 51864
rect 16592 51836 17632 51864
rect 16390 51824 16396 51827
rect 16448 51824 16454 51836
rect 16592 51796 16620 51836
rect 17494 51796 17500 51808
rect 15304 51768 16620 51796
rect 17455 51768 17500 51796
rect 17494 51756 17500 51768
rect 17552 51756 17558 51808
rect 17604 51796 17632 51836
rect 20248 51833 20260 51867
rect 20294 51864 20306 51867
rect 20438 51864 20444 51876
rect 20294 51836 20444 51864
rect 20294 51833 20306 51836
rect 20248 51827 20306 51833
rect 20438 51824 20444 51836
rect 20496 51824 20502 51876
rect 21928 51864 21956 51904
rect 20548 51836 21956 51864
rect 22088 51867 22146 51873
rect 20548 51796 20576 51836
rect 22088 51833 22100 51867
rect 22134 51864 22146 51867
rect 22554 51864 22560 51876
rect 22134 51836 22560 51864
rect 22134 51833 22146 51836
rect 22088 51827 22146 51833
rect 22554 51824 22560 51836
rect 22612 51824 22618 51876
rect 23584 51864 23612 51904
rect 23661 51901 23673 51935
rect 23707 51901 23719 51935
rect 23661 51895 23719 51901
rect 23768 51864 23796 51972
rect 27433 51969 27445 51972
rect 27479 51969 27491 52003
rect 27433 51963 27491 51969
rect 24486 51892 24492 51944
rect 24544 51932 24550 51944
rect 25777 51935 25835 51941
rect 25777 51932 25789 51935
rect 24544 51904 25789 51932
rect 24544 51892 24550 51904
rect 25777 51901 25789 51904
rect 25823 51901 25835 51935
rect 26510 51932 26516 51944
rect 26471 51904 26516 51932
rect 25777 51895 25835 51901
rect 26510 51892 26516 51904
rect 26568 51892 26574 51944
rect 27246 51932 27252 51944
rect 27207 51904 27252 51932
rect 27246 51892 27252 51904
rect 27304 51892 27310 51944
rect 27522 51892 27528 51944
rect 27580 51932 27586 51944
rect 27985 51935 28043 51941
rect 27985 51932 27997 51935
rect 27580 51904 27997 51932
rect 27580 51892 27586 51904
rect 27985 51901 27997 51904
rect 28031 51901 28043 51935
rect 27985 51895 28043 51901
rect 23584 51836 23796 51864
rect 23934 51824 23940 51876
rect 23992 51864 23998 51876
rect 26418 51864 26424 51876
rect 23992 51836 26424 51864
rect 23992 51824 23998 51836
rect 26418 51824 26424 51836
rect 26476 51824 26482 51876
rect 17604 51768 20576 51796
rect 20806 51756 20812 51808
rect 20864 51796 20870 51808
rect 21358 51796 21364 51808
rect 20864 51768 21364 51796
rect 20864 51756 20870 51768
rect 21358 51756 21364 51768
rect 21416 51756 21422 51808
rect 23382 51756 23388 51808
rect 23440 51796 23446 51808
rect 23753 51799 23811 51805
rect 23753 51796 23765 51799
rect 23440 51768 23765 51796
rect 23440 51756 23446 51768
rect 23753 51765 23765 51768
rect 23799 51765 23811 51799
rect 25866 51796 25872 51808
rect 25827 51768 25872 51796
rect 23753 51759 23811 51765
rect 25866 51756 25872 51768
rect 25924 51756 25930 51808
rect 28074 51796 28080 51808
rect 28035 51768 28080 51796
rect 28074 51756 28080 51768
rect 28132 51756 28138 51808
rect 1104 51706 28888 51728
rect 1104 51654 10246 51706
rect 10298 51654 10310 51706
rect 10362 51654 10374 51706
rect 10426 51654 10438 51706
rect 10490 51654 19510 51706
rect 19562 51654 19574 51706
rect 19626 51654 19638 51706
rect 19690 51654 19702 51706
rect 19754 51654 28888 51706
rect 1104 51632 28888 51654
rect 3418 51592 3424 51604
rect 3379 51564 3424 51592
rect 3418 51552 3424 51564
rect 3476 51552 3482 51604
rect 4062 51552 4068 51604
rect 4120 51592 4126 51604
rect 4341 51595 4399 51601
rect 4341 51592 4353 51595
rect 4120 51564 4353 51592
rect 4120 51552 4126 51564
rect 4341 51561 4353 51564
rect 4387 51561 4399 51595
rect 4341 51555 4399 51561
rect 4709 51595 4767 51601
rect 4709 51561 4721 51595
rect 4755 51592 4767 51595
rect 5166 51592 5172 51604
rect 4755 51564 5172 51592
rect 4755 51561 4767 51564
rect 4709 51555 4767 51561
rect 5166 51552 5172 51564
rect 5224 51552 5230 51604
rect 5721 51595 5779 51601
rect 5721 51561 5733 51595
rect 5767 51592 5779 51595
rect 5902 51592 5908 51604
rect 5767 51564 5908 51592
rect 5767 51561 5779 51564
rect 5721 51555 5779 51561
rect 5902 51552 5908 51564
rect 5960 51552 5966 51604
rect 6546 51552 6552 51604
rect 6604 51592 6610 51604
rect 7193 51595 7251 51601
rect 7193 51592 7205 51595
rect 6604 51564 7205 51592
rect 6604 51552 6610 51564
rect 7193 51561 7205 51564
rect 7239 51561 7251 51595
rect 7193 51555 7251 51561
rect 7285 51595 7343 51601
rect 7285 51561 7297 51595
rect 7331 51592 7343 51595
rect 8110 51592 8116 51604
rect 7331 51564 8116 51592
rect 7331 51561 7343 51564
rect 7285 51555 7343 51561
rect 8110 51552 8116 51564
rect 8168 51552 8174 51604
rect 10413 51595 10471 51601
rect 8220 51564 9076 51592
rect 5629 51527 5687 51533
rect 5629 51493 5641 51527
rect 5675 51524 5687 51527
rect 8220 51524 8248 51564
rect 5675 51496 8248 51524
rect 9048 51524 9076 51564
rect 10413 51561 10425 51595
rect 10459 51592 10471 51595
rect 10594 51592 10600 51604
rect 10459 51564 10600 51592
rect 10459 51561 10471 51564
rect 10413 51555 10471 51561
rect 10594 51552 10600 51564
rect 10652 51552 10658 51604
rect 10778 51592 10784 51604
rect 10739 51564 10784 51592
rect 10778 51552 10784 51564
rect 10836 51552 10842 51604
rect 12437 51595 12495 51601
rect 12437 51561 12449 51595
rect 12483 51592 12495 51595
rect 12526 51592 12532 51604
rect 12483 51564 12532 51592
rect 12483 51561 12495 51564
rect 12437 51555 12495 51561
rect 12526 51552 12532 51564
rect 12584 51552 12590 51604
rect 12805 51595 12863 51601
rect 12805 51592 12817 51595
rect 12636 51564 12817 51592
rect 12342 51524 12348 51536
rect 9048 51496 12348 51524
rect 5675 51493 5687 51496
rect 5629 51487 5687 51493
rect 12342 51484 12348 51496
rect 12400 51484 12406 51536
rect 1854 51456 1860 51468
rect 1815 51428 1860 51456
rect 1854 51416 1860 51428
rect 1912 51416 1918 51468
rect 2593 51459 2651 51465
rect 2593 51425 2605 51459
rect 2639 51425 2651 51459
rect 3326 51456 3332 51468
rect 3287 51428 3332 51456
rect 2593 51419 2651 51425
rect 2608 51388 2636 51419
rect 3326 51416 3332 51428
rect 3384 51416 3390 51468
rect 4801 51459 4859 51465
rect 4801 51425 4813 51459
rect 4847 51456 4859 51459
rect 6362 51456 6368 51468
rect 4847 51428 6368 51456
rect 4847 51425 4859 51428
rect 4801 51419 4859 51425
rect 6362 51416 6368 51428
rect 6420 51416 6426 51468
rect 7650 51416 7656 51468
rect 7708 51456 7714 51468
rect 7926 51456 7932 51468
rect 7708 51428 7932 51456
rect 7708 51416 7714 51428
rect 7926 51416 7932 51428
rect 7984 51456 7990 51468
rect 8113 51459 8171 51465
rect 8113 51456 8125 51459
rect 7984 51428 8125 51456
rect 7984 51416 7990 51428
rect 8113 51425 8125 51428
rect 8159 51425 8171 51459
rect 8113 51419 8171 51425
rect 8202 51416 8208 51468
rect 8260 51456 8266 51468
rect 8389 51459 8447 51465
rect 8389 51456 8401 51459
rect 8260 51428 8401 51456
rect 8260 51416 8266 51428
rect 8389 51425 8401 51428
rect 8435 51425 8447 51459
rect 8389 51419 8447 51425
rect 8478 51416 8484 51468
rect 8536 51456 8542 51468
rect 9858 51456 9864 51468
rect 8536 51428 9864 51456
rect 8536 51416 8542 51428
rect 9858 51416 9864 51428
rect 9916 51456 9922 51468
rect 10778 51456 10784 51468
rect 9916 51428 10784 51456
rect 9916 51416 9922 51428
rect 10778 51416 10784 51428
rect 10836 51416 10842 51468
rect 10873 51459 10931 51465
rect 10873 51425 10885 51459
rect 10919 51456 10931 51459
rect 11882 51456 11888 51468
rect 10919 51428 11888 51456
rect 10919 51425 10931 51428
rect 10873 51419 10931 51425
rect 11882 51416 11888 51428
rect 11940 51416 11946 51468
rect 12636 51456 12664 51564
rect 12805 51561 12817 51564
rect 12851 51561 12863 51595
rect 12805 51555 12863 51561
rect 15102 51552 15108 51604
rect 15160 51592 15166 51604
rect 15749 51595 15807 51601
rect 15749 51592 15761 51595
rect 15160 51564 15761 51592
rect 15160 51552 15166 51564
rect 15749 51561 15761 51564
rect 15795 51561 15807 51595
rect 15749 51555 15807 51561
rect 14636 51527 14694 51533
rect 14636 51493 14648 51527
rect 14682 51524 14694 51527
rect 14734 51524 14740 51536
rect 14682 51496 14740 51524
rect 14682 51493 14694 51496
rect 14636 51487 14694 51493
rect 14734 51484 14740 51496
rect 14792 51484 14798 51536
rect 13630 51456 13636 51468
rect 12636 51428 12848 51456
rect 13591 51428 13636 51456
rect 12820 51400 12848 51428
rect 13630 51416 13636 51428
rect 13688 51416 13694 51468
rect 15764 51456 15792 51555
rect 18230 51552 18236 51604
rect 18288 51592 18294 51604
rect 18325 51595 18383 51601
rect 18325 51592 18337 51595
rect 18288 51564 18337 51592
rect 18288 51552 18294 51564
rect 18325 51561 18337 51564
rect 18371 51561 18383 51595
rect 20438 51592 20444 51604
rect 20399 51564 20444 51592
rect 18325 51555 18383 51561
rect 20438 51552 20444 51564
rect 20496 51552 20502 51604
rect 20806 51592 20812 51604
rect 20767 51564 20812 51592
rect 20806 51552 20812 51564
rect 20864 51552 20870 51604
rect 22554 51592 22560 51604
rect 22515 51564 22560 51592
rect 22554 51552 22560 51564
rect 22612 51552 22618 51604
rect 22922 51592 22928 51604
rect 22883 51564 22928 51592
rect 22922 51552 22928 51564
rect 22980 51552 22986 51604
rect 23106 51552 23112 51604
rect 23164 51592 23170 51604
rect 26050 51592 26056 51604
rect 23164 51564 26056 51592
rect 23164 51552 23170 51564
rect 26050 51552 26056 51564
rect 26108 51552 26114 51604
rect 15838 51484 15844 51536
rect 15896 51524 15902 51536
rect 28169 51527 28227 51533
rect 28169 51524 28181 51527
rect 15896 51496 28181 51524
rect 15896 51484 15902 51496
rect 28169 51493 28181 51496
rect 28215 51493 28227 51527
rect 28169 51487 28227 51493
rect 16209 51459 16267 51465
rect 16209 51456 16221 51459
rect 15764 51428 16221 51456
rect 16209 51425 16221 51428
rect 16255 51425 16267 51459
rect 16209 51419 16267 51425
rect 18693 51459 18751 51465
rect 18693 51425 18705 51459
rect 18739 51456 18751 51459
rect 19334 51456 19340 51468
rect 18739 51428 19340 51456
rect 18739 51425 18751 51428
rect 18693 51419 18751 51425
rect 19334 51416 19340 51428
rect 19392 51456 19398 51468
rect 19521 51459 19579 51465
rect 19521 51456 19533 51459
rect 19392 51428 19533 51456
rect 19392 51416 19398 51428
rect 19521 51425 19533 51428
rect 19567 51425 19579 51459
rect 19521 51419 19579 51425
rect 22370 51416 22376 51468
rect 22428 51456 22434 51468
rect 23934 51456 23940 51468
rect 22428 51428 23940 51456
rect 22428 51416 22434 51428
rect 23934 51416 23940 51428
rect 23992 51416 23998 51468
rect 24026 51416 24032 51468
rect 24084 51456 24090 51468
rect 24377 51459 24435 51465
rect 24377 51456 24389 51459
rect 24084 51428 24389 51456
rect 24084 51416 24090 51428
rect 24377 51425 24389 51428
rect 24423 51425 24435 51459
rect 26694 51456 26700 51468
rect 26655 51428 26700 51456
rect 24377 51419 24435 51425
rect 26694 51416 26700 51428
rect 26752 51416 26758 51468
rect 27982 51456 27988 51468
rect 27943 51428 27988 51456
rect 27982 51416 27988 51428
rect 28040 51416 28046 51468
rect 4985 51391 5043 51397
rect 2608 51360 4936 51388
rect 2774 51280 2780 51332
rect 2832 51320 2838 51332
rect 4908 51320 4936 51360
rect 4985 51357 4997 51391
rect 5031 51388 5043 51391
rect 5166 51388 5172 51400
rect 5031 51360 5172 51388
rect 5031 51357 5043 51360
rect 4985 51351 5043 51357
rect 5166 51348 5172 51360
rect 5224 51348 5230 51400
rect 7469 51391 7527 51397
rect 7469 51357 7481 51391
rect 7515 51388 7527 51391
rect 8021 51391 8079 51397
rect 8021 51388 8033 51391
rect 7515 51360 8033 51388
rect 7515 51357 7527 51360
rect 7469 51351 7527 51357
rect 8021 51357 8033 51360
rect 8067 51357 8079 51391
rect 10962 51388 10968 51400
rect 8021 51351 8079 51357
rect 8128 51360 9076 51388
rect 10875 51360 10968 51388
rect 8128 51320 8156 51360
rect 2832 51292 2877 51320
rect 4908 51292 8156 51320
rect 9048 51320 9076 51360
rect 10962 51348 10968 51360
rect 11020 51388 11026 51400
rect 12158 51388 12164 51400
rect 11020 51360 12164 51388
rect 11020 51348 11026 51360
rect 12158 51348 12164 51360
rect 12216 51348 12222 51400
rect 12802 51348 12808 51400
rect 12860 51348 12866 51400
rect 12897 51391 12955 51397
rect 12897 51357 12909 51391
rect 12943 51388 12955 51391
rect 12986 51388 12992 51400
rect 12943 51360 12992 51388
rect 12943 51357 12955 51360
rect 12897 51351 12955 51357
rect 12986 51348 12992 51360
rect 13044 51348 13050 51400
rect 13081 51391 13139 51397
rect 13081 51357 13093 51391
rect 13127 51388 13139 51391
rect 13170 51388 13176 51400
rect 13127 51360 13176 51388
rect 13127 51357 13139 51360
rect 13081 51351 13139 51357
rect 13170 51348 13176 51360
rect 13228 51348 13234 51400
rect 14090 51348 14096 51400
rect 14148 51388 14154 51400
rect 14369 51391 14427 51397
rect 14369 51388 14381 51391
rect 14148 51360 14381 51388
rect 14148 51348 14154 51360
rect 14369 51357 14381 51360
rect 14415 51357 14427 51391
rect 18782 51388 18788 51400
rect 18743 51360 18788 51388
rect 14369 51351 14427 51357
rect 18782 51348 18788 51360
rect 18840 51348 18846 51400
rect 18874 51348 18880 51400
rect 18932 51388 18938 51400
rect 20898 51388 20904 51400
rect 18932 51360 18977 51388
rect 20859 51360 20904 51388
rect 18932 51348 18938 51360
rect 20898 51348 20904 51360
rect 20956 51348 20962 51400
rect 21085 51391 21143 51397
rect 21085 51357 21097 51391
rect 21131 51388 21143 51391
rect 21358 51388 21364 51400
rect 21131 51360 21364 51388
rect 21131 51357 21143 51360
rect 21085 51351 21143 51357
rect 21358 51348 21364 51360
rect 21416 51388 21422 51400
rect 23014 51388 23020 51400
rect 21416 51360 22600 51388
rect 22975 51360 23020 51388
rect 21416 51348 21422 51360
rect 12710 51320 12716 51332
rect 9048 51292 12716 51320
rect 2832 51280 2838 51292
rect 12710 51280 12716 51292
rect 12768 51280 12774 51332
rect 15304 51292 19748 51320
rect 1394 51212 1400 51264
rect 1452 51252 1458 51264
rect 1949 51255 2007 51261
rect 1949 51252 1961 51255
rect 1452 51224 1961 51252
rect 1452 51212 1458 51224
rect 1949 51221 1961 51224
rect 1995 51221 2007 51255
rect 1949 51215 2007 51221
rect 5902 51212 5908 51264
rect 5960 51252 5966 51264
rect 6825 51255 6883 51261
rect 6825 51252 6837 51255
rect 5960 51224 6837 51252
rect 5960 51212 5966 51224
rect 6825 51221 6837 51224
rect 6871 51221 6883 51255
rect 6825 51215 6883 51221
rect 8021 51255 8079 51261
rect 8021 51221 8033 51255
rect 8067 51252 8079 51255
rect 8570 51252 8576 51264
rect 8067 51224 8576 51252
rect 8067 51221 8079 51224
rect 8021 51215 8079 51221
rect 8570 51212 8576 51224
rect 8628 51212 8634 51264
rect 9674 51252 9680 51264
rect 9635 51224 9680 51252
rect 9674 51212 9680 51224
rect 9732 51212 9738 51264
rect 12434 51212 12440 51264
rect 12492 51252 12498 51264
rect 13725 51255 13783 51261
rect 13725 51252 13737 51255
rect 12492 51224 13737 51252
rect 12492 51212 12498 51224
rect 13725 51221 13737 51224
rect 13771 51221 13783 51255
rect 13725 51215 13783 51221
rect 13906 51212 13912 51264
rect 13964 51252 13970 51264
rect 15304 51252 15332 51292
rect 16298 51252 16304 51264
rect 13964 51224 15332 51252
rect 16259 51224 16304 51252
rect 13964 51212 13970 51224
rect 16298 51212 16304 51224
rect 16356 51212 16362 51264
rect 19610 51252 19616 51264
rect 19571 51224 19616 51252
rect 19610 51212 19616 51224
rect 19668 51212 19674 51264
rect 19720 51252 19748 51292
rect 21818 51280 21824 51332
rect 21876 51320 21882 51332
rect 22572 51320 22600 51360
rect 23014 51348 23020 51360
rect 23072 51348 23078 51400
rect 23109 51391 23167 51397
rect 23109 51357 23121 51391
rect 23155 51357 23167 51391
rect 23109 51351 23167 51357
rect 24121 51391 24179 51397
rect 24121 51357 24133 51391
rect 24167 51357 24179 51391
rect 24121 51351 24179 51357
rect 23124 51320 23152 51351
rect 21876 51292 22508 51320
rect 22572 51292 23152 51320
rect 21876 51280 21882 51292
rect 22370 51252 22376 51264
rect 19720 51224 22376 51252
rect 22370 51212 22376 51224
rect 22428 51212 22434 51264
rect 22480 51252 22508 51292
rect 23934 51252 23940 51264
rect 22480 51224 23940 51252
rect 23934 51212 23940 51224
rect 23992 51252 23998 51264
rect 24136 51252 24164 51351
rect 23992 51224 24164 51252
rect 25501 51255 25559 51261
rect 23992 51212 23998 51224
rect 25501 51221 25513 51255
rect 25547 51252 25559 51255
rect 25682 51252 25688 51264
rect 25547 51224 25688 51252
rect 25547 51221 25559 51224
rect 25501 51215 25559 51221
rect 25682 51212 25688 51224
rect 25740 51212 25746 51264
rect 26786 51252 26792 51264
rect 26747 51224 26792 51252
rect 26786 51212 26792 51224
rect 26844 51212 26850 51264
rect 1104 51162 28888 51184
rect 1104 51110 5614 51162
rect 5666 51110 5678 51162
rect 5730 51110 5742 51162
rect 5794 51110 5806 51162
rect 5858 51110 14878 51162
rect 14930 51110 14942 51162
rect 14994 51110 15006 51162
rect 15058 51110 15070 51162
rect 15122 51110 24142 51162
rect 24194 51110 24206 51162
rect 24258 51110 24270 51162
rect 24322 51110 24334 51162
rect 24386 51110 28888 51162
rect 1104 51088 28888 51110
rect 3234 51008 3240 51060
rect 3292 51048 3298 51060
rect 4433 51051 4491 51057
rect 4433 51048 4445 51051
rect 3292 51020 4445 51048
rect 3292 51008 3298 51020
rect 4433 51017 4445 51020
rect 4479 51017 4491 51051
rect 23106 51048 23112 51060
rect 4433 51011 4491 51017
rect 5828 51020 23112 51048
rect 2777 50983 2835 50989
rect 2777 50949 2789 50983
rect 2823 50980 2835 50983
rect 2958 50980 2964 50992
rect 2823 50952 2964 50980
rect 2823 50949 2835 50952
rect 2777 50943 2835 50949
rect 2958 50940 2964 50952
rect 3016 50940 3022 50992
rect 5828 50980 5856 51020
rect 23106 51008 23112 51020
rect 23164 51008 23170 51060
rect 23198 51008 23204 51060
rect 23256 51048 23262 51060
rect 23256 51020 23888 51048
rect 23256 51008 23262 51020
rect 4356 50952 5856 50980
rect 1872 50884 2774 50912
rect 1872 50853 1900 50884
rect 1857 50847 1915 50853
rect 1857 50813 1869 50847
rect 1903 50813 1915 50847
rect 1857 50807 1915 50813
rect 2590 50776 2596 50788
rect 2551 50748 2596 50776
rect 2590 50736 2596 50748
rect 2648 50736 2654 50788
rect 1946 50708 1952 50720
rect 1907 50680 1952 50708
rect 1946 50668 1952 50680
rect 2004 50668 2010 50720
rect 2746 50708 2774 50884
rect 4356 50853 4384 50952
rect 5902 50940 5908 50992
rect 5960 50940 5966 50992
rect 8113 50983 8171 50989
rect 8113 50980 8125 50983
rect 7392 50952 8125 50980
rect 4341 50847 4399 50853
rect 4341 50813 4353 50847
rect 4387 50813 4399 50847
rect 5810 50844 5816 50856
rect 5771 50816 5816 50844
rect 4341 50807 4399 50813
rect 5810 50804 5816 50816
rect 5868 50804 5874 50856
rect 5920 50853 5948 50940
rect 7392 50921 7420 50952
rect 8113 50949 8125 50952
rect 8159 50949 8171 50983
rect 8113 50943 8171 50949
rect 10137 50983 10195 50989
rect 10137 50949 10149 50983
rect 10183 50980 10195 50983
rect 11330 50980 11336 50992
rect 10183 50952 11336 50980
rect 10183 50949 10195 50952
rect 10137 50943 10195 50949
rect 11330 50940 11336 50952
rect 11388 50940 11394 50992
rect 12526 50980 12532 50992
rect 12360 50952 12532 50980
rect 7377 50915 7435 50921
rect 7377 50881 7389 50915
rect 7423 50881 7435 50915
rect 7377 50875 7435 50881
rect 7653 50915 7711 50921
rect 7653 50881 7665 50915
rect 7699 50912 7711 50915
rect 9490 50912 9496 50924
rect 7699 50884 9496 50912
rect 7699 50881 7711 50884
rect 7653 50875 7711 50881
rect 9490 50872 9496 50884
rect 9548 50872 9554 50924
rect 9769 50915 9827 50921
rect 9769 50881 9781 50915
rect 9815 50912 9827 50915
rect 10962 50912 10968 50924
rect 9815 50884 10968 50912
rect 9815 50881 9827 50884
rect 9769 50875 9827 50881
rect 10962 50872 10968 50884
rect 11020 50872 11026 50924
rect 12360 50921 12388 50952
rect 12526 50940 12532 50952
rect 12584 50980 12590 50992
rect 12584 50952 13952 50980
rect 12584 50940 12590 50952
rect 12345 50915 12403 50921
rect 12345 50881 12357 50915
rect 12391 50881 12403 50915
rect 12345 50875 12403 50881
rect 12710 50872 12716 50924
rect 12768 50912 12774 50924
rect 13924 50912 13952 50952
rect 16390 50940 16396 50992
rect 16448 50980 16454 50992
rect 16577 50983 16635 50989
rect 16577 50980 16589 50983
rect 16448 50952 16589 50980
rect 16448 50940 16454 50952
rect 16577 50949 16589 50952
rect 16623 50949 16635 50983
rect 16577 50943 16635 50949
rect 17218 50940 17224 50992
rect 17276 50980 17282 50992
rect 22462 50980 22468 50992
rect 17276 50952 22468 50980
rect 17276 50940 17282 50952
rect 22462 50940 22468 50952
rect 22520 50940 22526 50992
rect 23566 50980 23572 50992
rect 22572 50952 23572 50980
rect 15381 50915 15439 50921
rect 15381 50912 15393 50915
rect 12768 50884 13860 50912
rect 13924 50884 15393 50912
rect 12768 50872 12774 50884
rect 5905 50847 5963 50853
rect 5905 50813 5917 50847
rect 5951 50813 5963 50847
rect 5905 50807 5963 50813
rect 6089 50847 6147 50853
rect 6089 50813 6101 50847
rect 6135 50844 6147 50847
rect 6822 50844 6828 50856
rect 6135 50816 6828 50844
rect 6135 50813 6147 50816
rect 6089 50807 6147 50813
rect 6822 50804 6828 50816
rect 6880 50804 6886 50856
rect 7098 50804 7104 50856
rect 7156 50844 7162 50856
rect 7285 50847 7343 50853
rect 7285 50844 7297 50847
rect 7156 50816 7297 50844
rect 7156 50804 7162 50816
rect 7285 50813 7297 50816
rect 7331 50813 7343 50847
rect 7285 50807 7343 50813
rect 7558 50804 7564 50856
rect 7616 50844 7622 50856
rect 8389 50847 8447 50853
rect 8389 50844 8401 50847
rect 7616 50816 8401 50844
rect 7616 50804 7622 50816
rect 8389 50813 8401 50816
rect 8435 50813 8447 50847
rect 8389 50807 8447 50813
rect 12161 50847 12219 50853
rect 12161 50813 12173 50847
rect 12207 50844 12219 50847
rect 12434 50844 12440 50856
rect 12207 50816 12440 50844
rect 12207 50813 12219 50816
rect 12161 50807 12219 50813
rect 12434 50804 12440 50816
rect 12492 50804 12498 50856
rect 12986 50844 12992 50856
rect 12947 50816 12992 50844
rect 12986 50804 12992 50816
rect 13044 50804 13050 50856
rect 13078 50804 13084 50856
rect 13136 50844 13142 50856
rect 13633 50847 13691 50853
rect 13633 50844 13645 50847
rect 13136 50816 13645 50844
rect 13136 50804 13142 50816
rect 13633 50813 13645 50816
rect 13679 50844 13691 50847
rect 13722 50844 13728 50856
rect 13679 50816 13728 50844
rect 13679 50813 13691 50816
rect 13633 50807 13691 50813
rect 13722 50804 13728 50816
rect 13780 50804 13786 50856
rect 13832 50853 13860 50884
rect 15381 50881 15393 50884
rect 15427 50881 15439 50915
rect 15381 50875 15439 50881
rect 17129 50915 17187 50921
rect 17129 50881 17141 50915
rect 17175 50912 17187 50915
rect 17175 50884 18184 50912
rect 17175 50881 17187 50884
rect 17129 50875 17187 50881
rect 13817 50847 13875 50853
rect 13817 50813 13829 50847
rect 13863 50813 13875 50847
rect 13817 50807 13875 50813
rect 15197 50847 15255 50853
rect 15197 50813 15209 50847
rect 15243 50844 15255 50847
rect 16298 50844 16304 50856
rect 15243 50816 16304 50844
rect 15243 50813 15255 50816
rect 15197 50807 15255 50813
rect 16298 50804 16304 50816
rect 16356 50804 16362 50856
rect 16945 50847 17003 50853
rect 16945 50813 16957 50847
rect 16991 50844 17003 50847
rect 17494 50844 17500 50856
rect 16991 50816 17500 50844
rect 16991 50813 17003 50816
rect 16945 50807 17003 50813
rect 17494 50804 17500 50816
rect 17552 50844 17558 50856
rect 17773 50847 17831 50853
rect 17773 50844 17785 50847
rect 17552 50816 17785 50844
rect 17552 50804 17558 50816
rect 17773 50813 17785 50816
rect 17819 50813 17831 50847
rect 18156 50844 18184 50884
rect 18414 50872 18420 50924
rect 18472 50912 18478 50924
rect 20533 50915 20591 50921
rect 20533 50912 20545 50915
rect 18472 50884 20545 50912
rect 18472 50872 18478 50884
rect 20533 50881 20545 50884
rect 20579 50912 20591 50915
rect 21729 50915 21787 50921
rect 21729 50912 21741 50915
rect 20579 50884 21741 50912
rect 20579 50881 20591 50884
rect 20533 50875 20591 50881
rect 21729 50881 21741 50884
rect 21775 50881 21787 50915
rect 21729 50875 21787 50881
rect 18322 50844 18328 50856
rect 18156 50816 18328 50844
rect 17773 50807 17831 50813
rect 18322 50804 18328 50816
rect 18380 50844 18386 50856
rect 18874 50844 18880 50856
rect 18380 50816 18880 50844
rect 18380 50804 18386 50816
rect 18874 50804 18880 50816
rect 18932 50804 18938 50856
rect 19610 50804 19616 50856
rect 19668 50844 19674 50856
rect 20349 50847 20407 50853
rect 20349 50844 20361 50847
rect 19668 50816 20361 50844
rect 19668 50804 19674 50816
rect 20349 50813 20361 50816
rect 20395 50813 20407 50847
rect 20349 50807 20407 50813
rect 21450 50804 21456 50856
rect 21508 50844 21514 50856
rect 21545 50847 21603 50853
rect 21545 50844 21557 50847
rect 21508 50816 21557 50844
rect 21508 50804 21514 50816
rect 21545 50813 21557 50816
rect 21591 50813 21603 50847
rect 21744 50844 21772 50875
rect 22186 50844 22192 50856
rect 21744 50816 22192 50844
rect 21545 50807 21603 50813
rect 22186 50804 22192 50816
rect 22244 50804 22250 50856
rect 22572 50853 22600 50952
rect 23566 50940 23572 50952
rect 23624 50940 23630 50992
rect 23474 50872 23480 50924
rect 23532 50912 23538 50924
rect 23661 50915 23719 50921
rect 23661 50912 23673 50915
rect 23532 50884 23673 50912
rect 23532 50872 23538 50884
rect 23661 50881 23673 50884
rect 23707 50881 23719 50915
rect 23860 50912 23888 51020
rect 23934 51008 23940 51060
rect 23992 51048 23998 51060
rect 25314 51048 25320 51060
rect 23992 51020 25320 51048
rect 23992 51008 23998 51020
rect 25314 51008 25320 51020
rect 25372 51008 25378 51060
rect 27338 51048 27344 51060
rect 27299 51020 27344 51048
rect 27338 51008 27344 51020
rect 27396 51008 27402 51060
rect 26602 50912 26608 50924
rect 23860 50884 26608 50912
rect 23661 50875 23719 50881
rect 26602 50872 26608 50884
rect 26660 50872 26666 50924
rect 22557 50847 22615 50853
rect 22557 50813 22569 50847
rect 22603 50813 22615 50847
rect 23382 50844 23388 50856
rect 23343 50816 23388 50844
rect 22557 50807 22615 50813
rect 23382 50804 23388 50816
rect 23440 50804 23446 50856
rect 25225 50847 25283 50853
rect 25225 50813 25237 50847
rect 25271 50844 25283 50847
rect 25682 50844 25688 50856
rect 25271 50816 25688 50844
rect 25271 50813 25283 50816
rect 25225 50807 25283 50813
rect 25682 50804 25688 50816
rect 25740 50804 25746 50856
rect 26050 50844 26056 50856
rect 26011 50816 26056 50844
rect 26050 50804 26056 50816
rect 26108 50804 26114 50856
rect 26694 50844 26700 50856
rect 26655 50816 26700 50844
rect 26694 50804 26700 50816
rect 26752 50804 26758 50856
rect 5534 50736 5540 50788
rect 5592 50776 5598 50788
rect 5994 50776 6000 50788
rect 5592 50748 6000 50776
rect 5592 50736 5598 50748
rect 5994 50736 6000 50748
rect 6052 50776 6058 50788
rect 6454 50776 6460 50788
rect 6052 50748 6460 50776
rect 6052 50736 6058 50748
rect 6454 50736 6460 50748
rect 6512 50776 6518 50788
rect 6549 50779 6607 50785
rect 6549 50776 6561 50779
rect 6512 50748 6561 50776
rect 6512 50736 6518 50748
rect 6549 50745 6561 50748
rect 6595 50745 6607 50779
rect 8110 50776 8116 50788
rect 8071 50748 8116 50776
rect 6549 50739 6607 50745
rect 8110 50736 8116 50748
rect 8168 50736 8174 50788
rect 22278 50776 22284 50788
rect 8220 50748 22284 50776
rect 8220 50708 8248 50748
rect 22278 50736 22284 50748
rect 22336 50736 22342 50788
rect 26326 50736 26332 50788
rect 26384 50776 26390 50788
rect 27249 50779 27307 50785
rect 27249 50776 27261 50779
rect 26384 50748 27261 50776
rect 26384 50736 26390 50748
rect 27249 50745 27261 50748
rect 27295 50745 27307 50779
rect 27249 50739 27307 50745
rect 27430 50736 27436 50788
rect 27488 50776 27494 50788
rect 27985 50779 28043 50785
rect 27985 50776 27997 50779
rect 27488 50748 27997 50776
rect 27488 50736 27494 50748
rect 27985 50745 27997 50748
rect 28031 50745 28043 50779
rect 27985 50739 28043 50745
rect 2746 50680 8248 50708
rect 8294 50668 8300 50720
rect 8352 50708 8358 50720
rect 8352 50680 8397 50708
rect 8352 50668 8358 50680
rect 9214 50668 9220 50720
rect 9272 50708 9278 50720
rect 10229 50711 10287 50717
rect 10229 50708 10241 50711
rect 9272 50680 10241 50708
rect 9272 50668 9278 50680
rect 10229 50677 10241 50680
rect 10275 50677 10287 50711
rect 11790 50708 11796 50720
rect 11751 50680 11796 50708
rect 10229 50671 10287 50677
rect 11790 50668 11796 50680
rect 11848 50668 11854 50720
rect 12253 50711 12311 50717
rect 12253 50677 12265 50711
rect 12299 50708 12311 50711
rect 13081 50711 13139 50717
rect 13081 50708 13093 50711
rect 12299 50680 13093 50708
rect 12299 50677 12311 50680
rect 12253 50671 12311 50677
rect 13081 50677 13093 50680
rect 13127 50677 13139 50711
rect 13081 50671 13139 50677
rect 13817 50711 13875 50717
rect 13817 50677 13829 50711
rect 13863 50708 13875 50711
rect 14182 50708 14188 50720
rect 13863 50680 14188 50708
rect 13863 50677 13875 50680
rect 13817 50671 13875 50677
rect 14182 50668 14188 50680
rect 14240 50668 14246 50720
rect 14274 50668 14280 50720
rect 14332 50708 14338 50720
rect 14829 50711 14887 50717
rect 14829 50708 14841 50711
rect 14332 50680 14841 50708
rect 14332 50668 14338 50680
rect 14829 50677 14841 50680
rect 14875 50677 14887 50711
rect 15286 50708 15292 50720
rect 15247 50680 15292 50708
rect 14829 50671 14887 50677
rect 15286 50668 15292 50680
rect 15344 50668 15350 50720
rect 16850 50668 16856 50720
rect 16908 50708 16914 50720
rect 17037 50711 17095 50717
rect 17037 50708 17049 50711
rect 16908 50680 17049 50708
rect 16908 50668 16914 50680
rect 17037 50677 17049 50680
rect 17083 50677 17095 50711
rect 17037 50671 17095 50677
rect 17865 50711 17923 50717
rect 17865 50677 17877 50711
rect 17911 50708 17923 50711
rect 18230 50708 18236 50720
rect 17911 50680 18236 50708
rect 17911 50677 17923 50680
rect 17865 50671 17923 50677
rect 18230 50668 18236 50680
rect 18288 50668 18294 50720
rect 19978 50708 19984 50720
rect 19939 50680 19984 50708
rect 19978 50668 19984 50680
rect 20036 50668 20042 50720
rect 20070 50668 20076 50720
rect 20128 50708 20134 50720
rect 20441 50711 20499 50717
rect 20441 50708 20453 50711
rect 20128 50680 20453 50708
rect 20128 50668 20134 50680
rect 20441 50677 20453 50680
rect 20487 50677 20499 50711
rect 20441 50671 20499 50677
rect 21177 50711 21235 50717
rect 21177 50677 21189 50711
rect 21223 50708 21235 50711
rect 21266 50708 21272 50720
rect 21223 50680 21272 50708
rect 21223 50677 21235 50680
rect 21177 50671 21235 50677
rect 21266 50668 21272 50680
rect 21324 50668 21330 50720
rect 21637 50711 21695 50717
rect 21637 50677 21649 50711
rect 21683 50708 21695 50711
rect 21818 50708 21824 50720
rect 21683 50680 21824 50708
rect 21683 50677 21695 50680
rect 21637 50671 21695 50677
rect 21818 50668 21824 50680
rect 21876 50668 21882 50720
rect 22373 50711 22431 50717
rect 22373 50677 22385 50711
rect 22419 50708 22431 50711
rect 22922 50708 22928 50720
rect 22419 50680 22928 50708
rect 22419 50677 22431 50680
rect 22373 50671 22431 50677
rect 22922 50668 22928 50680
rect 22980 50668 22986 50720
rect 23017 50711 23075 50717
rect 23017 50677 23029 50711
rect 23063 50708 23075 50711
rect 23106 50708 23112 50720
rect 23063 50680 23112 50708
rect 23063 50677 23075 50680
rect 23017 50671 23075 50677
rect 23106 50668 23112 50680
rect 23164 50668 23170 50720
rect 23477 50711 23535 50717
rect 23477 50677 23489 50711
rect 23523 50708 23535 50711
rect 24118 50708 24124 50720
rect 23523 50680 24124 50708
rect 23523 50677 23535 50680
rect 23477 50671 23535 50677
rect 24118 50668 24124 50680
rect 24176 50708 24182 50720
rect 25317 50711 25375 50717
rect 25317 50708 25329 50711
rect 24176 50680 25329 50708
rect 24176 50668 24182 50680
rect 25317 50677 25329 50680
rect 25363 50677 25375 50711
rect 25866 50708 25872 50720
rect 25827 50680 25872 50708
rect 25317 50671 25375 50677
rect 25866 50668 25872 50680
rect 25924 50668 25930 50720
rect 26513 50711 26571 50717
rect 26513 50677 26525 50711
rect 26559 50708 26571 50711
rect 27154 50708 27160 50720
rect 26559 50680 27160 50708
rect 26559 50677 26571 50680
rect 26513 50671 26571 50677
rect 27154 50668 27160 50680
rect 27212 50668 27218 50720
rect 28074 50708 28080 50720
rect 28035 50680 28080 50708
rect 28074 50668 28080 50680
rect 28132 50668 28138 50720
rect 1104 50618 28888 50640
rect 1104 50566 10246 50618
rect 10298 50566 10310 50618
rect 10362 50566 10374 50618
rect 10426 50566 10438 50618
rect 10490 50566 19510 50618
rect 19562 50566 19574 50618
rect 19626 50566 19638 50618
rect 19690 50566 19702 50618
rect 19754 50566 28888 50618
rect 1104 50544 28888 50566
rect 3142 50464 3148 50516
rect 3200 50504 3206 50516
rect 3421 50507 3479 50513
rect 3421 50504 3433 50507
rect 3200 50476 3433 50504
rect 3200 50464 3206 50476
rect 3421 50473 3433 50476
rect 3467 50473 3479 50507
rect 3421 50467 3479 50473
rect 5629 50507 5687 50513
rect 5629 50473 5641 50507
rect 5675 50504 5687 50507
rect 8110 50504 8116 50516
rect 5675 50476 8116 50504
rect 5675 50473 5687 50476
rect 5629 50467 5687 50473
rect 8110 50464 8116 50476
rect 8168 50464 8174 50516
rect 9401 50507 9459 50513
rect 9401 50473 9413 50507
rect 9447 50504 9459 50507
rect 9766 50504 9772 50516
rect 9447 50476 9772 50504
rect 9447 50473 9459 50476
rect 9401 50467 9459 50473
rect 9766 50464 9772 50476
rect 9824 50464 9830 50516
rect 11790 50464 11796 50516
rect 11848 50504 11854 50516
rect 12621 50507 12679 50513
rect 12621 50504 12633 50507
rect 11848 50476 12633 50504
rect 11848 50464 11854 50476
rect 12621 50473 12633 50476
rect 12667 50473 12679 50507
rect 14182 50504 14188 50516
rect 14143 50476 14188 50504
rect 12621 50467 12679 50473
rect 14182 50464 14188 50476
rect 14240 50464 14246 50516
rect 14274 50464 14280 50516
rect 14332 50504 14338 50516
rect 18230 50504 18236 50516
rect 14332 50476 14377 50504
rect 18191 50476 18236 50504
rect 14332 50464 14338 50476
rect 18230 50464 18236 50476
rect 18288 50464 18294 50516
rect 21266 50504 21272 50516
rect 18340 50476 20116 50504
rect 21227 50476 21272 50504
rect 3329 50439 3387 50445
rect 3329 50405 3341 50439
rect 3375 50436 3387 50439
rect 17218 50436 17224 50448
rect 3375 50408 17224 50436
rect 3375 50405 3387 50408
rect 3329 50399 3387 50405
rect 17218 50396 17224 50408
rect 17276 50396 17282 50448
rect 18340 50436 18368 50476
rect 19978 50436 19984 50448
rect 17328 50408 18368 50436
rect 19444 50408 19984 50436
rect 1857 50371 1915 50377
rect 1857 50337 1869 50371
rect 1903 50368 1915 50371
rect 2498 50368 2504 50380
rect 1903 50340 2504 50368
rect 1903 50337 1915 50340
rect 1857 50331 1915 50337
rect 2498 50328 2504 50340
rect 2556 50328 2562 50380
rect 2593 50371 2651 50377
rect 2593 50337 2605 50371
rect 2639 50337 2651 50371
rect 5534 50368 5540 50380
rect 5495 50340 5540 50368
rect 2593 50331 2651 50337
rect 2608 50300 2636 50331
rect 5534 50328 5540 50340
rect 5592 50328 5598 50380
rect 5721 50371 5779 50377
rect 5721 50337 5733 50371
rect 5767 50368 5779 50371
rect 6086 50368 6092 50380
rect 5767 50340 6092 50368
rect 5767 50337 5779 50340
rect 5721 50331 5779 50337
rect 6086 50328 6092 50340
rect 6144 50368 6150 50380
rect 6362 50368 6368 50380
rect 6144 50340 6368 50368
rect 6144 50328 6150 50340
rect 6362 50328 6368 50340
rect 6420 50328 6426 50380
rect 7098 50368 7104 50380
rect 7059 50340 7104 50368
rect 7098 50328 7104 50340
rect 7156 50328 7162 50380
rect 7558 50368 7564 50380
rect 7519 50340 7564 50368
rect 7558 50328 7564 50340
rect 7616 50328 7622 50380
rect 8018 50368 8024 50380
rect 7979 50340 8024 50368
rect 8018 50328 8024 50340
rect 8076 50368 8082 50380
rect 8294 50368 8300 50380
rect 8076 50340 8300 50368
rect 8076 50328 8082 50340
rect 8294 50328 8300 50340
rect 8352 50328 8358 50380
rect 9214 50368 9220 50380
rect 9175 50340 9220 50368
rect 9214 50328 9220 50340
rect 9272 50328 9278 50380
rect 9490 50368 9496 50380
rect 9451 50340 9496 50368
rect 9490 50328 9496 50340
rect 9548 50328 9554 50380
rect 9677 50371 9735 50377
rect 9677 50337 9689 50371
rect 9723 50368 9735 50371
rect 9858 50368 9864 50380
rect 9723 50340 9864 50368
rect 9723 50337 9735 50340
rect 9677 50331 9735 50337
rect 9858 50328 9864 50340
rect 9916 50328 9922 50380
rect 16209 50371 16267 50377
rect 16209 50337 16221 50371
rect 16255 50337 16267 50371
rect 16390 50368 16396 50380
rect 16351 50340 16396 50368
rect 16209 50331 16267 50337
rect 2608 50272 7604 50300
rect 2774 50192 2780 50244
rect 2832 50232 2838 50244
rect 7576 50232 7604 50272
rect 7650 50260 7656 50312
rect 7708 50300 7714 50312
rect 7708 50272 7753 50300
rect 7708 50260 7714 50272
rect 11974 50260 11980 50312
rect 12032 50300 12038 50312
rect 12529 50303 12587 50309
rect 12529 50300 12541 50303
rect 12032 50272 12541 50300
rect 12032 50260 12038 50272
rect 12529 50269 12541 50272
rect 12575 50269 12587 50303
rect 12529 50263 12587 50269
rect 12618 50260 12624 50312
rect 12676 50300 12682 50312
rect 12713 50303 12771 50309
rect 12713 50300 12725 50303
rect 12676 50272 12725 50300
rect 12676 50260 12682 50272
rect 12713 50269 12725 50272
rect 12759 50300 12771 50303
rect 14369 50303 14427 50309
rect 14369 50300 14381 50303
rect 12759 50272 14381 50300
rect 12759 50269 12771 50272
rect 12713 50263 12771 50269
rect 14369 50269 14381 50272
rect 14415 50269 14427 50303
rect 16224 50300 16252 50331
rect 16390 50328 16396 50340
rect 16448 50328 16454 50380
rect 16850 50300 16856 50312
rect 16224 50272 16856 50300
rect 14369 50263 14427 50269
rect 16850 50260 16856 50272
rect 16908 50260 16914 50312
rect 17328 50232 17356 50408
rect 18325 50371 18383 50377
rect 18325 50337 18337 50371
rect 18371 50368 18383 50371
rect 19242 50368 19248 50380
rect 18371 50340 19248 50368
rect 18371 50337 18383 50340
rect 18325 50331 18383 50337
rect 19242 50328 19248 50340
rect 19300 50328 19306 50380
rect 19444 50377 19472 50408
rect 19978 50396 19984 50408
rect 20036 50396 20042 50448
rect 20088 50436 20116 50476
rect 21266 50464 21272 50476
rect 21324 50464 21330 50516
rect 22186 50464 22192 50516
rect 22244 50504 22250 50516
rect 23198 50504 23204 50516
rect 22244 50476 23204 50504
rect 22244 50464 22250 50476
rect 23198 50464 23204 50476
rect 23256 50464 23262 50516
rect 23293 50507 23351 50513
rect 23293 50473 23305 50507
rect 23339 50504 23351 50507
rect 23339 50476 23980 50504
rect 23339 50473 23351 50476
rect 23293 50467 23351 50473
rect 21910 50436 21916 50448
rect 20088 50408 21916 50436
rect 21910 50396 21916 50408
rect 21968 50396 21974 50448
rect 23842 50436 23848 50448
rect 22664 50408 23848 50436
rect 19429 50371 19487 50377
rect 19429 50337 19441 50371
rect 19475 50337 19487 50371
rect 19613 50371 19671 50377
rect 19613 50368 19625 50371
rect 19429 50331 19487 50337
rect 19536 50340 19625 50368
rect 18414 50300 18420 50312
rect 18375 50272 18420 50300
rect 18414 50260 18420 50272
rect 18472 50260 18478 50312
rect 18506 50260 18512 50312
rect 18564 50300 18570 50312
rect 19337 50303 19395 50309
rect 19337 50300 19349 50303
rect 18564 50272 19349 50300
rect 18564 50260 18570 50272
rect 19337 50269 19349 50272
rect 19383 50269 19395 50303
rect 19337 50263 19395 50269
rect 2832 50204 2877 50232
rect 7576 50204 17356 50232
rect 2832 50192 2838 50204
rect 1394 50124 1400 50176
rect 1452 50164 1458 50176
rect 1949 50167 2007 50173
rect 1949 50164 1961 50167
rect 1452 50136 1961 50164
rect 1452 50124 1458 50136
rect 1949 50133 1961 50136
rect 1995 50133 2007 50167
rect 1949 50127 2007 50133
rect 11054 50124 11060 50176
rect 11112 50164 11118 50176
rect 12161 50167 12219 50173
rect 12161 50164 12173 50167
rect 11112 50136 12173 50164
rect 11112 50124 11118 50136
rect 12161 50133 12173 50136
rect 12207 50133 12219 50167
rect 12161 50127 12219 50133
rect 13630 50124 13636 50176
rect 13688 50164 13694 50176
rect 13817 50167 13875 50173
rect 13817 50164 13829 50167
rect 13688 50136 13829 50164
rect 13688 50124 13694 50136
rect 13817 50133 13829 50136
rect 13863 50133 13875 50167
rect 16298 50164 16304 50176
rect 16259 50136 16304 50164
rect 13817 50127 13875 50133
rect 16298 50124 16304 50136
rect 16356 50124 16362 50176
rect 17678 50124 17684 50176
rect 17736 50164 17742 50176
rect 17865 50167 17923 50173
rect 17865 50164 17877 50167
rect 17736 50136 17877 50164
rect 17736 50124 17742 50136
rect 17865 50133 17877 50136
rect 17911 50133 17923 50167
rect 17865 50127 17923 50133
rect 18230 50124 18236 50176
rect 18288 50164 18294 50176
rect 19536 50164 19564 50340
rect 19613 50337 19625 50340
rect 19659 50368 19671 50371
rect 21361 50371 21419 50377
rect 21361 50368 21373 50371
rect 19659 50340 21373 50368
rect 19659 50337 19671 50340
rect 19613 50331 19671 50337
rect 21361 50337 21373 50340
rect 21407 50368 21419 50371
rect 22554 50368 22560 50380
rect 21407 50340 22560 50368
rect 21407 50337 21419 50340
rect 21361 50331 21419 50337
rect 22554 50328 22560 50340
rect 22612 50328 22618 50380
rect 22664 50377 22692 50408
rect 23842 50396 23848 50408
rect 23900 50396 23906 50448
rect 23952 50436 23980 50476
rect 24026 50464 24032 50516
rect 24084 50504 24090 50516
rect 24213 50507 24271 50513
rect 24213 50504 24225 50507
rect 24084 50476 24225 50504
rect 24084 50464 24090 50476
rect 24213 50473 24225 50476
rect 24259 50473 24271 50507
rect 24213 50467 24271 50473
rect 24765 50507 24823 50513
rect 24765 50473 24777 50507
rect 24811 50504 24823 50507
rect 27430 50504 27436 50516
rect 24811 50476 27436 50504
rect 24811 50473 24823 50476
rect 24765 50467 24823 50473
rect 27430 50464 27436 50476
rect 27488 50464 27494 50516
rect 24670 50436 24676 50448
rect 23952 50408 24676 50436
rect 24670 50396 24676 50408
rect 24728 50396 24734 50448
rect 25866 50396 25872 50448
rect 25924 50436 25930 50448
rect 27985 50439 28043 50445
rect 27985 50436 27997 50439
rect 25924 50408 27997 50436
rect 25924 50396 25930 50408
rect 27985 50405 27997 50408
rect 28031 50405 28043 50439
rect 27985 50399 28043 50405
rect 22649 50371 22707 50377
rect 22649 50337 22661 50371
rect 22695 50337 22707 50371
rect 22649 50331 22707 50337
rect 23477 50371 23535 50377
rect 23477 50337 23489 50371
rect 23523 50337 23535 50371
rect 23477 50331 23535 50337
rect 20073 50303 20131 50309
rect 20073 50269 20085 50303
rect 20119 50300 20131 50303
rect 20254 50300 20260 50312
rect 20119 50272 20260 50300
rect 20119 50269 20131 50272
rect 20073 50263 20131 50269
rect 20254 50260 20260 50272
rect 20312 50260 20318 50312
rect 21174 50300 21180 50312
rect 21135 50272 21180 50300
rect 21174 50260 21180 50272
rect 21232 50260 21238 50312
rect 22278 50192 22284 50244
rect 22336 50232 22342 50244
rect 23492 50232 23520 50331
rect 23566 50328 23572 50380
rect 23624 50368 23630 50380
rect 23937 50371 23995 50377
rect 23937 50368 23949 50371
rect 23624 50340 23949 50368
rect 23624 50328 23630 50340
rect 23937 50337 23949 50340
rect 23983 50337 23995 50371
rect 23937 50331 23995 50337
rect 24029 50371 24087 50377
rect 24029 50337 24041 50371
rect 24075 50368 24087 50371
rect 24118 50368 24124 50380
rect 24075 50340 24124 50368
rect 24075 50337 24087 50340
rect 24029 50331 24087 50337
rect 24118 50328 24124 50340
rect 24176 50328 24182 50380
rect 24946 50368 24952 50380
rect 24907 50340 24952 50368
rect 24946 50328 24952 50340
rect 25004 50328 25010 50380
rect 25590 50368 25596 50380
rect 25551 50340 25596 50368
rect 25590 50328 25596 50340
rect 25648 50328 25654 50380
rect 26234 50368 26240 50380
rect 26195 50340 26240 50368
rect 26234 50328 26240 50340
rect 26292 50328 26298 50380
rect 26881 50371 26939 50377
rect 26881 50337 26893 50371
rect 26927 50368 26939 50371
rect 26970 50368 26976 50380
rect 26927 50340 26976 50368
rect 26927 50337 26939 50340
rect 26881 50331 26939 50337
rect 26970 50328 26976 50340
rect 27028 50328 27034 50380
rect 24213 50303 24271 50309
rect 24213 50269 24225 50303
rect 24259 50300 24271 50303
rect 24762 50300 24768 50312
rect 24259 50272 24768 50300
rect 24259 50269 24271 50272
rect 24213 50263 24271 50269
rect 24762 50260 24768 50272
rect 24820 50260 24826 50312
rect 28169 50303 28227 50309
rect 28169 50300 28181 50303
rect 25240 50272 28181 50300
rect 25130 50232 25136 50244
rect 22336 50204 23152 50232
rect 23492 50204 25136 50232
rect 22336 50192 22342 50204
rect 18288 50136 19564 50164
rect 18288 50124 18294 50136
rect 20162 50124 20168 50176
rect 20220 50164 20226 50176
rect 20809 50167 20867 50173
rect 20809 50164 20821 50167
rect 20220 50136 20821 50164
rect 20220 50124 20226 50136
rect 20809 50133 20821 50136
rect 20855 50133 20867 50167
rect 20809 50127 20867 50133
rect 20990 50124 20996 50176
rect 21048 50164 21054 50176
rect 22738 50164 22744 50176
rect 21048 50136 22744 50164
rect 21048 50124 21054 50136
rect 22738 50124 22744 50136
rect 22796 50124 22802 50176
rect 22833 50167 22891 50173
rect 22833 50133 22845 50167
rect 22879 50164 22891 50167
rect 23014 50164 23020 50176
rect 22879 50136 23020 50164
rect 22879 50133 22891 50136
rect 22833 50127 22891 50133
rect 23014 50124 23020 50136
rect 23072 50124 23078 50176
rect 23124 50164 23152 50204
rect 25130 50192 25136 50204
rect 25188 50192 25194 50244
rect 25240 50164 25268 50272
rect 28169 50269 28181 50272
rect 28215 50269 28227 50303
rect 28169 50263 28227 50269
rect 26053 50235 26111 50241
rect 26053 50201 26065 50235
rect 26099 50232 26111 50235
rect 27890 50232 27896 50244
rect 26099 50204 27896 50232
rect 26099 50201 26111 50204
rect 26053 50195 26111 50201
rect 27890 50192 27896 50204
rect 27948 50192 27954 50244
rect 23124 50136 25268 50164
rect 25409 50167 25467 50173
rect 25409 50133 25421 50167
rect 25455 50164 25467 50167
rect 25866 50164 25872 50176
rect 25455 50136 25872 50164
rect 25455 50133 25467 50136
rect 25409 50127 25467 50133
rect 25866 50124 25872 50136
rect 25924 50124 25930 50176
rect 26697 50167 26755 50173
rect 26697 50133 26709 50167
rect 26743 50164 26755 50167
rect 27982 50164 27988 50176
rect 26743 50136 27988 50164
rect 26743 50133 26755 50136
rect 26697 50127 26755 50133
rect 27982 50124 27988 50136
rect 28040 50124 28046 50176
rect 1104 50074 28888 50096
rect 1104 50022 5614 50074
rect 5666 50022 5678 50074
rect 5730 50022 5742 50074
rect 5794 50022 5806 50074
rect 5858 50022 14878 50074
rect 14930 50022 14942 50074
rect 14994 50022 15006 50074
rect 15058 50022 15070 50074
rect 15122 50022 24142 50074
rect 24194 50022 24206 50074
rect 24258 50022 24270 50074
rect 24322 50022 24334 50074
rect 24386 50022 28888 50074
rect 1104 50000 28888 50022
rect 11974 49960 11980 49972
rect 11935 49932 11980 49960
rect 11974 49920 11980 49932
rect 12032 49920 12038 49972
rect 18506 49960 18512 49972
rect 18467 49932 18512 49960
rect 18506 49920 18512 49932
rect 18564 49920 18570 49972
rect 20070 49960 20076 49972
rect 20031 49932 20076 49960
rect 20070 49920 20076 49932
rect 20128 49920 20134 49972
rect 21174 49960 21180 49972
rect 21135 49932 21180 49960
rect 21174 49920 21180 49932
rect 21232 49920 21238 49972
rect 21818 49960 21824 49972
rect 21779 49932 21824 49960
rect 21818 49920 21824 49932
rect 21876 49920 21882 49972
rect 21910 49920 21916 49972
rect 21968 49960 21974 49972
rect 27985 49963 28043 49969
rect 27985 49960 27997 49963
rect 21968 49932 27997 49960
rect 21968 49920 21974 49932
rect 27985 49929 27997 49932
rect 28031 49929 28043 49963
rect 27985 49923 28043 49929
rect 16390 49852 16396 49904
rect 16448 49892 16454 49904
rect 25130 49892 25136 49904
rect 16448 49864 18644 49892
rect 16448 49852 16454 49864
rect 2041 49827 2099 49833
rect 2041 49793 2053 49827
rect 2087 49824 2099 49827
rect 2958 49824 2964 49836
rect 2087 49796 2964 49824
rect 2087 49793 2099 49796
rect 2041 49787 2099 49793
rect 2958 49784 2964 49796
rect 3016 49784 3022 49836
rect 11330 49824 11336 49836
rect 7852 49796 11336 49824
rect 2593 49759 2651 49765
rect 2593 49725 2605 49759
rect 2639 49756 2651 49759
rect 2682 49756 2688 49768
rect 2639 49728 2688 49756
rect 2639 49725 2651 49728
rect 2593 49719 2651 49725
rect 2682 49716 2688 49728
rect 2740 49716 2746 49768
rect 2777 49759 2835 49765
rect 2777 49725 2789 49759
rect 2823 49756 2835 49759
rect 2866 49756 2872 49768
rect 2823 49728 2872 49756
rect 2823 49725 2835 49728
rect 2777 49719 2835 49725
rect 2866 49716 2872 49728
rect 2924 49716 2930 49768
rect 5994 49756 6000 49768
rect 5644 49728 6000 49756
rect 1857 49691 1915 49697
rect 1857 49657 1869 49691
rect 1903 49688 1915 49691
rect 5644 49688 5672 49728
rect 5994 49716 6000 49728
rect 6052 49716 6058 49768
rect 7852 49765 7880 49796
rect 11330 49784 11336 49796
rect 11388 49784 11394 49836
rect 15105 49827 15163 49833
rect 12820 49796 13676 49824
rect 7837 49759 7895 49765
rect 7837 49725 7849 49759
rect 7883 49725 7895 49759
rect 7837 49719 7895 49725
rect 7929 49759 7987 49765
rect 7929 49725 7941 49759
rect 7975 49756 7987 49759
rect 8202 49756 8208 49768
rect 7975 49728 8208 49756
rect 7975 49725 7987 49728
rect 7929 49719 7987 49725
rect 8202 49716 8208 49728
rect 8260 49716 8266 49768
rect 11882 49756 11888 49768
rect 11843 49728 11888 49756
rect 11882 49716 11888 49728
rect 11940 49716 11946 49768
rect 12069 49759 12127 49765
rect 12069 49725 12081 49759
rect 12115 49756 12127 49759
rect 12710 49756 12716 49768
rect 12115 49728 12716 49756
rect 12115 49725 12127 49728
rect 12069 49719 12127 49725
rect 12710 49716 12716 49728
rect 12768 49716 12774 49768
rect 12820 49765 12848 49796
rect 13648 49768 13676 49796
rect 15105 49793 15117 49827
rect 15151 49824 15163 49827
rect 15470 49824 15476 49836
rect 15151 49796 15476 49824
rect 15151 49793 15163 49796
rect 15105 49787 15163 49793
rect 15470 49784 15476 49796
rect 15528 49784 15534 49836
rect 17678 49824 17684 49836
rect 17639 49796 17684 49824
rect 17678 49784 17684 49796
rect 17736 49784 17742 49836
rect 17865 49827 17923 49833
rect 17865 49793 17877 49827
rect 17911 49824 17923 49827
rect 18230 49824 18236 49836
rect 17911 49796 18236 49824
rect 17911 49793 17923 49796
rect 17865 49787 17923 49793
rect 18230 49784 18236 49796
rect 18288 49784 18294 49836
rect 12805 49759 12863 49765
rect 12805 49725 12817 49759
rect 12851 49725 12863 49759
rect 12805 49719 12863 49725
rect 12989 49759 13047 49765
rect 12989 49725 13001 49759
rect 13035 49756 13047 49759
rect 13078 49756 13084 49768
rect 13035 49728 13084 49756
rect 13035 49725 13047 49728
rect 12989 49719 13047 49725
rect 13078 49716 13084 49728
rect 13136 49756 13142 49768
rect 13449 49759 13507 49765
rect 13449 49756 13461 49759
rect 13136 49728 13461 49756
rect 13136 49716 13142 49728
rect 13449 49725 13461 49728
rect 13495 49725 13507 49759
rect 13630 49756 13636 49768
rect 13591 49728 13636 49756
rect 13449 49719 13507 49725
rect 13630 49716 13636 49728
rect 13688 49716 13694 49768
rect 15378 49756 15384 49768
rect 15339 49728 15384 49756
rect 15378 49716 15384 49728
rect 15436 49716 15442 49768
rect 16761 49759 16819 49765
rect 16761 49725 16773 49759
rect 16807 49756 16819 49759
rect 16942 49756 16948 49768
rect 16807 49728 16948 49756
rect 16807 49725 16819 49728
rect 16761 49719 16819 49725
rect 16942 49716 16948 49728
rect 17000 49716 17006 49768
rect 18616 49765 18644 49864
rect 21744 49864 25136 49892
rect 20898 49784 20904 49836
rect 20956 49824 20962 49836
rect 20956 49796 21128 49824
rect 20956 49784 20962 49796
rect 18417 49759 18475 49765
rect 18417 49725 18429 49759
rect 18463 49756 18475 49759
rect 18601 49759 18659 49765
rect 18463 49728 18552 49756
rect 18463 49725 18475 49728
rect 18417 49719 18475 49725
rect 15194 49688 15200 49700
rect 1903 49660 5672 49688
rect 5736 49660 15200 49688
rect 1903 49657 1915 49660
rect 1857 49651 1915 49657
rect 2498 49580 2504 49632
rect 2556 49620 2562 49632
rect 5736 49620 5764 49660
rect 15194 49648 15200 49660
rect 15252 49648 15258 49700
rect 16298 49648 16304 49700
rect 16356 49688 16362 49700
rect 17589 49691 17647 49697
rect 17589 49688 17601 49691
rect 16356 49660 17601 49688
rect 16356 49648 16362 49660
rect 17589 49657 17601 49660
rect 17635 49657 17647 49691
rect 18524 49688 18552 49728
rect 18601 49725 18613 49759
rect 18647 49725 18659 49759
rect 18782 49756 18788 49768
rect 18695 49728 18788 49756
rect 18601 49719 18659 49725
rect 18708 49688 18736 49728
rect 18782 49716 18788 49728
rect 18840 49756 18846 49768
rect 19334 49756 19340 49768
rect 18840 49728 19340 49756
rect 18840 49716 18846 49728
rect 19334 49716 19340 49728
rect 19392 49716 19398 49768
rect 19981 49759 20039 49765
rect 19981 49725 19993 49759
rect 20027 49756 20039 49759
rect 20990 49756 20996 49768
rect 20027 49728 20996 49756
rect 20027 49725 20039 49728
rect 19981 49719 20039 49725
rect 20990 49716 20996 49728
rect 21048 49716 21054 49768
rect 21100 49765 21128 49796
rect 21744 49765 21772 49864
rect 25130 49852 25136 49864
rect 25188 49852 25194 49904
rect 21836 49796 22692 49824
rect 21085 49759 21143 49765
rect 21085 49725 21097 49759
rect 21131 49725 21143 49759
rect 21085 49719 21143 49725
rect 21269 49759 21327 49765
rect 21269 49725 21281 49759
rect 21315 49756 21327 49759
rect 21729 49759 21787 49765
rect 21315 49728 21680 49756
rect 21315 49725 21327 49728
rect 21269 49719 21327 49725
rect 18524 49660 18736 49688
rect 21652 49688 21680 49728
rect 21729 49725 21741 49759
rect 21775 49725 21787 49759
rect 21729 49719 21787 49725
rect 21836 49688 21864 49796
rect 22664 49768 22692 49796
rect 23014 49784 23020 49836
rect 23072 49824 23078 49836
rect 26418 49824 26424 49836
rect 23072 49796 26424 49824
rect 23072 49784 23078 49796
rect 26418 49784 26424 49796
rect 26476 49784 26482 49836
rect 22557 49759 22615 49765
rect 22557 49725 22569 49759
rect 22603 49725 22615 49759
rect 22557 49719 22615 49725
rect 21652 49660 21864 49688
rect 22572 49688 22600 49719
rect 22646 49716 22652 49768
rect 22704 49756 22710 49768
rect 22741 49759 22799 49765
rect 22741 49756 22753 49759
rect 22704 49728 22753 49756
rect 22704 49716 22710 49728
rect 22741 49725 22753 49728
rect 22787 49725 22799 49759
rect 22741 49719 22799 49725
rect 22922 49716 22928 49768
rect 22980 49756 22986 49768
rect 22980 49728 23796 49756
rect 22980 49716 22986 49728
rect 22830 49688 22836 49700
rect 22572 49660 22836 49688
rect 17589 49651 17647 49657
rect 22830 49648 22836 49660
rect 22888 49648 22894 49700
rect 23768 49688 23796 49728
rect 23842 49716 23848 49768
rect 23900 49756 23906 49768
rect 23937 49759 23995 49765
rect 23937 49756 23949 49759
rect 23900 49728 23949 49756
rect 23900 49716 23906 49728
rect 23937 49725 23949 49728
rect 23983 49725 23995 49759
rect 23937 49719 23995 49725
rect 24026 49716 24032 49768
rect 24084 49756 24090 49768
rect 24121 49759 24179 49765
rect 24121 49756 24133 49759
rect 24084 49728 24133 49756
rect 24084 49716 24090 49728
rect 24121 49725 24133 49728
rect 24167 49725 24179 49759
rect 24121 49719 24179 49725
rect 24228 49728 24900 49756
rect 24228 49688 24256 49728
rect 23768 49660 24256 49688
rect 12894 49620 12900 49632
rect 2556 49592 5764 49620
rect 12855 49592 12900 49620
rect 2556 49580 2562 49592
rect 12894 49580 12900 49592
rect 12952 49580 12958 49632
rect 13817 49623 13875 49629
rect 13817 49589 13829 49623
rect 13863 49620 13875 49623
rect 13906 49620 13912 49632
rect 13863 49592 13912 49620
rect 13863 49589 13875 49592
rect 13817 49583 13875 49589
rect 13906 49580 13912 49592
rect 13964 49580 13970 49632
rect 17221 49623 17279 49629
rect 17221 49589 17233 49623
rect 17267 49620 17279 49623
rect 17494 49620 17500 49632
rect 17267 49592 17500 49620
rect 17267 49589 17279 49592
rect 17221 49583 17279 49589
rect 17494 49580 17500 49592
rect 17552 49580 17558 49632
rect 22738 49620 22744 49632
rect 22699 49592 22744 49620
rect 22738 49580 22744 49592
rect 22796 49580 22802 49632
rect 24026 49620 24032 49632
rect 23987 49592 24032 49620
rect 24026 49580 24032 49592
rect 24084 49580 24090 49632
rect 24872 49620 24900 49728
rect 25406 49716 25412 49768
rect 25464 49756 25470 49768
rect 25501 49759 25559 49765
rect 25501 49756 25513 49759
rect 25464 49728 25513 49756
rect 25464 49716 25470 49728
rect 25501 49725 25513 49728
rect 25547 49725 25559 49759
rect 25774 49756 25780 49768
rect 25735 49728 25780 49756
rect 25501 49719 25559 49725
rect 25774 49716 25780 49728
rect 25832 49716 25838 49768
rect 25866 49716 25872 49768
rect 25924 49756 25930 49768
rect 27893 49759 27951 49765
rect 27893 49756 27905 49759
rect 25924 49728 27905 49756
rect 25924 49716 25930 49728
rect 27893 49725 27905 49728
rect 27939 49725 27951 49759
rect 27893 49719 27951 49725
rect 25866 49620 25872 49632
rect 24872 49592 25872 49620
rect 25866 49580 25872 49592
rect 25924 49620 25930 49632
rect 26881 49623 26939 49629
rect 26881 49620 26893 49623
rect 25924 49592 26893 49620
rect 25924 49580 25930 49592
rect 26881 49589 26893 49592
rect 26927 49589 26939 49623
rect 26881 49583 26939 49589
rect 1104 49530 28888 49552
rect 1104 49478 10246 49530
rect 10298 49478 10310 49530
rect 10362 49478 10374 49530
rect 10426 49478 10438 49530
rect 10490 49478 19510 49530
rect 19562 49478 19574 49530
rect 19626 49478 19638 49530
rect 19690 49478 19702 49530
rect 19754 49478 28888 49530
rect 1104 49456 28888 49478
rect 5902 49416 5908 49428
rect 5863 49388 5908 49416
rect 5902 49376 5908 49388
rect 5960 49376 5966 49428
rect 5994 49376 6000 49428
rect 6052 49416 6058 49428
rect 15933 49419 15991 49425
rect 15933 49416 15945 49419
rect 6052 49388 15945 49416
rect 6052 49376 6058 49388
rect 15933 49385 15945 49388
rect 15979 49385 15991 49419
rect 15933 49379 15991 49385
rect 17236 49388 22094 49416
rect 2682 49308 2688 49360
rect 2740 49348 2746 49360
rect 17236 49348 17264 49388
rect 2740 49320 17264 49348
rect 17405 49351 17463 49357
rect 2740 49308 2746 49320
rect 17405 49317 17417 49351
rect 17451 49348 17463 49351
rect 18414 49348 18420 49360
rect 17451 49320 18420 49348
rect 17451 49317 17463 49320
rect 17405 49311 17463 49317
rect 18414 49308 18420 49320
rect 18472 49308 18478 49360
rect 19334 49308 19340 49360
rect 19392 49348 19398 49360
rect 20438 49348 20444 49360
rect 19392 49320 20444 49348
rect 19392 49308 19398 49320
rect 1854 49280 1860 49292
rect 1815 49252 1860 49280
rect 1854 49240 1860 49252
rect 1912 49240 1918 49292
rect 2593 49283 2651 49289
rect 2593 49249 2605 49283
rect 2639 49249 2651 49283
rect 2593 49243 2651 49249
rect 4148 49283 4206 49289
rect 4148 49249 4160 49283
rect 4194 49280 4206 49283
rect 4706 49280 4712 49292
rect 4194 49252 4712 49280
rect 4194 49249 4206 49252
rect 4148 49243 4206 49249
rect 2608 49212 2636 49243
rect 4706 49240 4712 49252
rect 4764 49240 4770 49292
rect 5721 49283 5779 49289
rect 5721 49249 5733 49283
rect 5767 49249 5779 49283
rect 5721 49243 5779 49249
rect 5905 49283 5963 49289
rect 5905 49249 5917 49283
rect 5951 49280 5963 49283
rect 6178 49280 6184 49292
rect 5951 49252 6184 49280
rect 5951 49249 5963 49252
rect 5905 49243 5963 49249
rect 2682 49212 2688 49224
rect 2608 49184 2688 49212
rect 2682 49172 2688 49184
rect 2740 49172 2746 49224
rect 3786 49172 3792 49224
rect 3844 49212 3850 49224
rect 3881 49215 3939 49221
rect 3881 49212 3893 49215
rect 3844 49184 3893 49212
rect 3844 49172 3850 49184
rect 3881 49181 3893 49184
rect 3927 49181 3939 49215
rect 5736 49212 5764 49243
rect 6178 49240 6184 49252
rect 6236 49240 6242 49292
rect 7653 49283 7711 49289
rect 7653 49249 7665 49283
rect 7699 49280 7711 49283
rect 7742 49280 7748 49292
rect 7699 49252 7748 49280
rect 7699 49249 7711 49252
rect 7653 49243 7711 49249
rect 6086 49212 6092 49224
rect 5736 49184 6092 49212
rect 3881 49175 3939 49181
rect 2774 49104 2780 49156
rect 2832 49144 2838 49156
rect 2832 49116 2877 49144
rect 2832 49104 2838 49116
rect 1946 49076 1952 49088
rect 1907 49048 1952 49076
rect 1946 49036 1952 49048
rect 2004 49036 2010 49088
rect 3896 49076 3924 49175
rect 6086 49172 6092 49184
rect 6144 49212 6150 49224
rect 6638 49212 6644 49224
rect 6144 49184 6644 49212
rect 6144 49172 6150 49184
rect 6638 49172 6644 49184
rect 6696 49172 6702 49224
rect 7668 49144 7696 49243
rect 7742 49240 7748 49252
rect 7800 49240 7806 49292
rect 7926 49289 7932 49292
rect 7920 49243 7932 49289
rect 7984 49280 7990 49292
rect 7984 49252 8020 49280
rect 7926 49240 7932 49243
rect 7984 49240 7990 49252
rect 9858 49240 9864 49292
rect 9916 49280 9922 49292
rect 10137 49283 10195 49289
rect 10137 49280 10149 49283
rect 9916 49252 10149 49280
rect 9916 49240 9922 49252
rect 10137 49249 10149 49252
rect 10183 49249 10195 49283
rect 10137 49243 10195 49249
rect 10229 49283 10287 49289
rect 10229 49249 10241 49283
rect 10275 49249 10287 49283
rect 10229 49243 10287 49249
rect 10413 49283 10471 49289
rect 10413 49249 10425 49283
rect 10459 49249 10471 49283
rect 10413 49243 10471 49249
rect 10505 49283 10563 49289
rect 10505 49249 10517 49283
rect 10551 49280 10563 49283
rect 10965 49283 11023 49289
rect 10965 49280 10977 49283
rect 10551 49252 10977 49280
rect 10551 49249 10563 49252
rect 10505 49243 10563 49249
rect 10965 49249 10977 49252
rect 11011 49280 11023 49283
rect 11054 49280 11060 49292
rect 11011 49252 11060 49280
rect 11011 49249 11023 49252
rect 10965 49243 11023 49249
rect 9582 49172 9588 49224
rect 9640 49212 9646 49224
rect 10244 49212 10272 49243
rect 9640 49184 10272 49212
rect 10428 49212 10456 49243
rect 11054 49240 11060 49252
rect 11112 49240 11118 49292
rect 11149 49283 11207 49289
rect 11149 49249 11161 49283
rect 11195 49280 11207 49283
rect 11882 49280 11888 49292
rect 11195 49252 11888 49280
rect 11195 49249 11207 49252
rect 11149 49243 11207 49249
rect 10686 49212 10692 49224
rect 10428 49184 10692 49212
rect 9640 49172 9646 49184
rect 10686 49172 10692 49184
rect 10744 49212 10750 49224
rect 11164 49212 11192 49243
rect 11882 49240 11888 49252
rect 11940 49240 11946 49292
rect 12250 49280 12256 49292
rect 12211 49252 12256 49280
rect 12250 49240 12256 49252
rect 12308 49240 12314 49292
rect 13170 49240 13176 49292
rect 13228 49280 13234 49292
rect 13538 49280 13544 49292
rect 13228 49252 13544 49280
rect 13228 49240 13234 49252
rect 13538 49240 13544 49252
rect 13596 49240 13602 49292
rect 13725 49283 13783 49289
rect 13725 49249 13737 49283
rect 13771 49280 13783 49283
rect 13906 49280 13912 49292
rect 13771 49252 13912 49280
rect 13771 49249 13783 49252
rect 13725 49243 13783 49249
rect 13906 49240 13912 49252
rect 13964 49240 13970 49292
rect 14277 49283 14335 49289
rect 14277 49249 14289 49283
rect 14323 49249 14335 49283
rect 14734 49280 14740 49292
rect 14695 49252 14740 49280
rect 14277 49243 14335 49249
rect 12342 49212 12348 49224
rect 10744 49184 11192 49212
rect 12303 49184 12348 49212
rect 10744 49172 10750 49184
rect 12342 49172 12348 49184
rect 12400 49172 12406 49224
rect 12621 49215 12679 49221
rect 12621 49181 12633 49215
rect 12667 49212 12679 49215
rect 12802 49212 12808 49224
rect 12667 49184 12808 49212
rect 12667 49181 12679 49184
rect 12621 49175 12679 49181
rect 12802 49172 12808 49184
rect 12860 49172 12866 49224
rect 12894 49172 12900 49224
rect 12952 49212 12958 49224
rect 13817 49215 13875 49221
rect 13817 49212 13829 49215
rect 12952 49184 13829 49212
rect 12952 49172 12958 49184
rect 13817 49181 13829 49184
rect 13863 49212 13875 49215
rect 14292 49212 14320 49243
rect 14734 49240 14740 49252
rect 14792 49240 14798 49292
rect 16025 49283 16083 49289
rect 16025 49249 16037 49283
rect 16071 49280 16083 49283
rect 16942 49280 16948 49292
rect 16071 49252 16948 49280
rect 16071 49249 16083 49252
rect 16025 49243 16083 49249
rect 16942 49240 16948 49252
rect 17000 49240 17006 49292
rect 20088 49289 20116 49320
rect 20438 49308 20444 49320
rect 20496 49308 20502 49360
rect 22066 49348 22094 49388
rect 22738 49376 22744 49428
rect 22796 49416 22802 49428
rect 23017 49419 23075 49425
rect 23017 49416 23029 49419
rect 22796 49388 23029 49416
rect 22796 49376 22802 49388
rect 23017 49385 23029 49388
rect 23063 49385 23075 49419
rect 23017 49379 23075 49385
rect 23106 49376 23112 49428
rect 23164 49416 23170 49428
rect 25409 49419 25467 49425
rect 23164 49388 23209 49416
rect 23164 49376 23170 49388
rect 25409 49385 25421 49419
rect 25455 49416 25467 49419
rect 25774 49416 25780 49428
rect 25455 49388 25780 49416
rect 25455 49385 25467 49388
rect 25409 49379 25467 49385
rect 25774 49376 25780 49388
rect 25832 49376 25838 49428
rect 27985 49419 28043 49425
rect 27985 49416 27997 49419
rect 25884 49388 27997 49416
rect 25884 49348 25912 49388
rect 27985 49385 27997 49388
rect 28031 49385 28043 49419
rect 27985 49379 28043 49385
rect 27890 49348 27896 49360
rect 22066 49320 25912 49348
rect 27851 49320 27896 49348
rect 27890 49308 27896 49320
rect 27948 49308 27954 49360
rect 20073 49283 20131 49289
rect 20073 49249 20085 49283
rect 20119 49249 20131 49283
rect 20254 49280 20260 49292
rect 20215 49252 20260 49280
rect 20073 49243 20131 49249
rect 20254 49240 20260 49252
rect 20312 49240 20318 49292
rect 23842 49240 23848 49292
rect 23900 49280 23906 49292
rect 24489 49283 24547 49289
rect 24489 49280 24501 49283
rect 23900 49252 24501 49280
rect 23900 49240 23906 49252
rect 24489 49249 24501 49252
rect 24535 49249 24547 49283
rect 24489 49243 24547 49249
rect 24581 49283 24639 49289
rect 24581 49249 24593 49283
rect 24627 49249 24639 49283
rect 24581 49243 24639 49249
rect 21358 49212 21364 49224
rect 13863 49184 14320 49212
rect 21319 49184 21364 49212
rect 13863 49181 13875 49184
rect 13817 49175 13875 49181
rect 21358 49172 21364 49184
rect 21416 49172 21422 49224
rect 22554 49172 22560 49224
rect 22612 49212 22618 49224
rect 22922 49212 22928 49224
rect 22612 49184 22928 49212
rect 22612 49172 22618 49184
rect 22922 49172 22928 49184
rect 22980 49212 22986 49224
rect 23201 49215 23259 49221
rect 23201 49212 23213 49215
rect 22980 49184 23213 49212
rect 22980 49172 22986 49184
rect 23201 49181 23213 49184
rect 23247 49181 23259 49215
rect 23201 49175 23259 49181
rect 23934 49172 23940 49224
rect 23992 49212 23998 49224
rect 24596 49212 24624 49243
rect 24670 49240 24676 49292
rect 24728 49280 24734 49292
rect 24854 49280 24860 49292
rect 24728 49252 24773 49280
rect 24815 49252 24860 49280
rect 24728 49240 24734 49252
rect 24854 49240 24860 49252
rect 24912 49240 24918 49292
rect 25774 49280 25780 49292
rect 25735 49252 25780 49280
rect 25774 49240 25780 49252
rect 25832 49240 25838 49292
rect 26878 49280 26884 49292
rect 26839 49252 26884 49280
rect 26878 49240 26884 49252
rect 26936 49240 26942 49292
rect 23992 49184 24624 49212
rect 23992 49172 23998 49184
rect 25590 49172 25596 49224
rect 25648 49212 25654 49224
rect 25866 49212 25872 49224
rect 25648 49184 25872 49212
rect 25648 49172 25654 49184
rect 25866 49172 25872 49184
rect 25924 49172 25930 49224
rect 26053 49215 26111 49221
rect 26053 49181 26065 49215
rect 26099 49212 26111 49215
rect 26142 49212 26148 49224
rect 26099 49184 26148 49212
rect 26099 49181 26111 49184
rect 26053 49175 26111 49181
rect 26142 49172 26148 49184
rect 26200 49172 26206 49224
rect 4816 49116 7696 49144
rect 4816 49076 4844 49116
rect 13906 49104 13912 49156
rect 13964 49144 13970 49156
rect 14415 49147 14473 49153
rect 14415 49144 14427 49147
rect 13964 49116 14427 49144
rect 13964 49104 13970 49116
rect 14415 49113 14427 49116
rect 14461 49113 14473 49147
rect 14415 49107 14473 49113
rect 15933 49147 15991 49153
rect 15933 49113 15945 49147
rect 15979 49144 15991 49147
rect 28074 49144 28080 49156
rect 15979 49116 28080 49144
rect 15979 49113 15991 49116
rect 15933 49107 15991 49113
rect 28074 49104 28080 49116
rect 28132 49104 28138 49156
rect 5258 49076 5264 49088
rect 3896 49048 4844 49076
rect 5219 49048 5264 49076
rect 5258 49036 5264 49048
rect 5316 49036 5322 49088
rect 9030 49076 9036 49088
rect 8991 49048 9036 49076
rect 9030 49036 9036 49048
rect 9088 49036 9094 49088
rect 9953 49079 10011 49085
rect 9953 49045 9965 49079
rect 9999 49076 10011 49079
rect 10042 49076 10048 49088
rect 9999 49048 10048 49076
rect 9999 49045 10011 49048
rect 9953 49039 10011 49045
rect 10042 49036 10048 49048
rect 10100 49036 10106 49088
rect 10962 49076 10968 49088
rect 10923 49048 10968 49076
rect 10962 49036 10968 49048
rect 11020 49036 11026 49088
rect 13354 49076 13360 49088
rect 13315 49048 13360 49076
rect 13354 49036 13360 49048
rect 13412 49036 13418 49088
rect 13538 49036 13544 49088
rect 13596 49076 13602 49088
rect 14553 49079 14611 49085
rect 14553 49076 14565 49079
rect 13596 49048 14565 49076
rect 13596 49036 13602 49048
rect 14553 49045 14565 49048
rect 14599 49045 14611 49079
rect 14553 49039 14611 49045
rect 14642 49036 14648 49088
rect 14700 49076 14706 49088
rect 16114 49076 16120 49088
rect 14700 49048 14745 49076
rect 16075 49048 16120 49076
rect 14700 49036 14706 49048
rect 16114 49036 16120 49048
rect 16172 49036 16178 49088
rect 16390 49036 16396 49088
rect 16448 49076 16454 49088
rect 17497 49079 17555 49085
rect 17497 49076 17509 49079
rect 16448 49048 17509 49076
rect 16448 49036 16454 49048
rect 17497 49045 17509 49048
rect 17543 49045 17555 49079
rect 17497 49039 17555 49045
rect 22649 49079 22707 49085
rect 22649 49045 22661 49079
rect 22695 49076 22707 49079
rect 23198 49076 23204 49088
rect 22695 49048 23204 49076
rect 22695 49045 22707 49048
rect 22649 49039 22707 49045
rect 23198 49036 23204 49048
rect 23256 49036 23262 49088
rect 24213 49079 24271 49085
rect 24213 49045 24225 49079
rect 24259 49076 24271 49079
rect 25498 49076 25504 49088
rect 24259 49048 25504 49076
rect 24259 49045 24271 49048
rect 24213 49039 24271 49045
rect 25498 49036 25504 49048
rect 25556 49036 25562 49088
rect 26697 49079 26755 49085
rect 26697 49045 26709 49079
rect 26743 49076 26755 49079
rect 27890 49076 27896 49088
rect 26743 49048 27896 49076
rect 26743 49045 26755 49048
rect 26697 49039 26755 49045
rect 27890 49036 27896 49048
rect 27948 49036 27954 49088
rect 1104 48986 28888 49008
rect 1104 48934 5614 48986
rect 5666 48934 5678 48986
rect 5730 48934 5742 48986
rect 5794 48934 5806 48986
rect 5858 48934 14878 48986
rect 14930 48934 14942 48986
rect 14994 48934 15006 48986
rect 15058 48934 15070 48986
rect 15122 48934 24142 48986
rect 24194 48934 24206 48986
rect 24258 48934 24270 48986
rect 24322 48934 24334 48986
rect 24386 48934 28888 48986
rect 1104 48912 28888 48934
rect 5166 48832 5172 48884
rect 5224 48872 5230 48884
rect 5442 48872 5448 48884
rect 5224 48844 5448 48872
rect 5224 48832 5230 48844
rect 5442 48832 5448 48844
rect 5500 48832 5506 48884
rect 7837 48875 7895 48881
rect 7837 48841 7849 48875
rect 7883 48872 7895 48875
rect 7926 48872 7932 48884
rect 7883 48844 7932 48872
rect 7883 48841 7895 48844
rect 7837 48835 7895 48841
rect 7926 48832 7932 48844
rect 7984 48832 7990 48884
rect 14921 48875 14979 48881
rect 14921 48841 14933 48875
rect 14967 48872 14979 48875
rect 15378 48872 15384 48884
rect 14967 48844 15384 48872
rect 14967 48841 14979 48844
rect 14921 48835 14979 48841
rect 15378 48832 15384 48844
rect 15436 48832 15442 48884
rect 21729 48875 21787 48881
rect 21729 48841 21741 48875
rect 21775 48872 21787 48875
rect 25774 48872 25780 48884
rect 21775 48844 25780 48872
rect 21775 48841 21787 48844
rect 21729 48835 21787 48841
rect 25774 48832 25780 48844
rect 25832 48832 25838 48884
rect 28074 48872 28080 48884
rect 28035 48844 28080 48872
rect 28074 48832 28080 48844
rect 28132 48832 28138 48884
rect 3237 48807 3295 48813
rect 3237 48773 3249 48807
rect 3283 48804 3295 48807
rect 4154 48804 4160 48816
rect 3283 48776 4160 48804
rect 3283 48773 3295 48776
rect 3237 48767 3295 48773
rect 4154 48764 4160 48776
rect 4212 48764 4218 48816
rect 6270 48804 6276 48816
rect 6231 48776 6276 48804
rect 6270 48764 6276 48776
rect 6328 48764 6334 48816
rect 8018 48764 8024 48816
rect 8076 48804 8082 48816
rect 9769 48807 9827 48813
rect 9769 48804 9781 48807
rect 8076 48776 9781 48804
rect 8076 48764 8082 48776
rect 9769 48773 9781 48776
rect 9815 48773 9827 48807
rect 10594 48804 10600 48816
rect 9769 48767 9827 48773
rect 9968 48776 10600 48804
rect 4893 48739 4951 48745
rect 4893 48705 4905 48739
rect 4939 48736 4951 48739
rect 5166 48736 5172 48748
rect 4939 48708 5172 48736
rect 4939 48705 4951 48708
rect 4893 48699 4951 48705
rect 5166 48696 5172 48708
rect 5224 48696 5230 48748
rect 5442 48696 5448 48748
rect 5500 48736 5506 48748
rect 8389 48739 8447 48745
rect 8389 48736 8401 48739
rect 5500 48708 8401 48736
rect 5500 48696 5506 48708
rect 8389 48705 8401 48708
rect 8435 48705 8447 48739
rect 8389 48699 8447 48705
rect 1857 48671 1915 48677
rect 1857 48637 1869 48671
rect 1903 48668 1915 48671
rect 2866 48668 2872 48680
rect 1903 48640 2872 48668
rect 1903 48637 1915 48640
rect 1857 48631 1915 48637
rect 2866 48628 2872 48640
rect 2924 48668 2930 48680
rect 3786 48668 3792 48680
rect 2924 48640 3792 48668
rect 2924 48628 2930 48640
rect 3786 48628 3792 48640
rect 3844 48628 3850 48680
rect 5258 48628 5264 48680
rect 5316 48668 5322 48680
rect 5537 48671 5595 48677
rect 5537 48668 5549 48671
rect 5316 48640 5549 48668
rect 5316 48628 5322 48640
rect 5537 48637 5549 48640
rect 5583 48637 5595 48671
rect 5537 48631 5595 48637
rect 5629 48671 5687 48677
rect 5629 48637 5641 48671
rect 5675 48668 5687 48671
rect 8294 48668 8300 48680
rect 5675 48640 8300 48668
rect 5675 48637 5687 48640
rect 5629 48631 5687 48637
rect 8294 48628 8300 48640
rect 8352 48628 8358 48680
rect 9968 48677 9996 48776
rect 10594 48764 10600 48776
rect 10652 48764 10658 48816
rect 13354 48764 13360 48816
rect 13412 48804 13418 48816
rect 14737 48807 14795 48813
rect 14737 48804 14749 48807
rect 13412 48776 14749 48804
rect 13412 48764 13418 48776
rect 14737 48773 14749 48776
rect 14783 48773 14795 48807
rect 14737 48767 14795 48773
rect 15194 48764 15200 48816
rect 15252 48804 15258 48816
rect 15252 48776 24716 48804
rect 15252 48764 15258 48776
rect 11146 48736 11152 48748
rect 10060 48708 11152 48736
rect 9953 48671 10011 48677
rect 9953 48637 9965 48671
rect 9999 48637 10011 48671
rect 9953 48631 10011 48637
rect 2124 48603 2182 48609
rect 2124 48569 2136 48603
rect 2170 48600 2182 48603
rect 2590 48600 2596 48612
rect 2170 48572 2596 48600
rect 2170 48569 2182 48572
rect 2124 48563 2182 48569
rect 2590 48560 2596 48572
rect 2648 48560 2654 48612
rect 4430 48560 4436 48612
rect 4488 48600 4494 48612
rect 4709 48603 4767 48609
rect 4709 48600 4721 48603
rect 4488 48572 4721 48600
rect 4488 48560 4494 48572
rect 4709 48569 4721 48572
rect 4755 48569 4767 48603
rect 6546 48600 6552 48612
rect 6507 48572 6552 48600
rect 4709 48563 4767 48569
rect 6546 48560 6552 48572
rect 6604 48560 6610 48612
rect 6825 48603 6883 48609
rect 6825 48569 6837 48603
rect 6871 48600 6883 48603
rect 6914 48600 6920 48612
rect 6871 48572 6920 48600
rect 6871 48569 6883 48572
rect 6825 48563 6883 48569
rect 6914 48560 6920 48572
rect 6972 48560 6978 48612
rect 8205 48603 8263 48609
rect 8205 48569 8217 48603
rect 8251 48600 8263 48603
rect 9030 48600 9036 48612
rect 8251 48572 9036 48600
rect 8251 48569 8263 48572
rect 8205 48563 8263 48569
rect 9030 48560 9036 48572
rect 9088 48560 9094 48612
rect 4246 48532 4252 48544
rect 4207 48504 4252 48532
rect 4246 48492 4252 48504
rect 4304 48492 4310 48544
rect 4614 48532 4620 48544
rect 4575 48504 4620 48532
rect 4614 48492 4620 48504
rect 4672 48492 4678 48544
rect 6730 48532 6736 48544
rect 6691 48504 6736 48532
rect 6730 48492 6736 48504
rect 6788 48492 6794 48544
rect 8297 48535 8355 48541
rect 8297 48501 8309 48535
rect 8343 48532 8355 48535
rect 9582 48532 9588 48544
rect 8343 48504 9588 48532
rect 8343 48501 8355 48504
rect 8297 48495 8355 48501
rect 9582 48492 9588 48504
rect 9640 48492 9646 48544
rect 10060 48541 10088 48708
rect 11146 48696 11152 48708
rect 11204 48736 11210 48748
rect 11885 48739 11943 48745
rect 11885 48736 11897 48739
rect 11204 48708 11897 48736
rect 11204 48696 11210 48708
rect 11885 48705 11897 48708
rect 11931 48736 11943 48739
rect 12250 48736 12256 48748
rect 11931 48708 12256 48736
rect 11931 48705 11943 48708
rect 11885 48699 11943 48705
rect 12250 48696 12256 48708
rect 12308 48696 12314 48748
rect 12342 48696 12348 48748
rect 12400 48736 12406 48748
rect 13081 48739 13139 48745
rect 13081 48736 13093 48739
rect 12400 48708 13093 48736
rect 12400 48696 12434 48708
rect 13081 48705 13093 48708
rect 13127 48705 13139 48739
rect 13081 48699 13139 48705
rect 14642 48696 14648 48748
rect 14700 48736 14706 48748
rect 14921 48739 14979 48745
rect 14921 48736 14933 48739
rect 14700 48708 14933 48736
rect 14700 48696 14706 48708
rect 14921 48705 14933 48708
rect 14967 48705 14979 48739
rect 14921 48699 14979 48705
rect 15013 48739 15071 48745
rect 15013 48705 15025 48739
rect 15059 48736 15071 48739
rect 15286 48736 15292 48748
rect 15059 48708 15292 48736
rect 15059 48705 15071 48708
rect 15013 48699 15071 48705
rect 15286 48696 15292 48708
rect 15344 48736 15350 48748
rect 16114 48736 16120 48748
rect 15344 48708 16120 48736
rect 15344 48696 15350 48708
rect 16114 48696 16120 48708
rect 16172 48696 16178 48748
rect 21174 48696 21180 48748
rect 21232 48736 21238 48748
rect 21269 48739 21327 48745
rect 21269 48736 21281 48739
rect 21232 48708 21281 48736
rect 21232 48696 21238 48708
rect 21269 48705 21281 48708
rect 21315 48705 21327 48739
rect 21269 48699 21327 48705
rect 23845 48739 23903 48745
rect 23845 48705 23857 48739
rect 23891 48736 23903 48739
rect 24026 48736 24032 48748
rect 23891 48708 24032 48736
rect 23891 48705 23903 48708
rect 23845 48699 23903 48705
rect 24026 48696 24032 48708
rect 24084 48696 24090 48748
rect 24688 48736 24716 48776
rect 24762 48764 24768 48816
rect 24820 48804 24826 48816
rect 25501 48807 25559 48813
rect 25501 48804 25513 48807
rect 24820 48776 25513 48804
rect 24820 48764 24826 48776
rect 25501 48773 25513 48776
rect 25547 48773 25559 48807
rect 25501 48767 25559 48773
rect 27433 48739 27491 48745
rect 27433 48736 27445 48739
rect 24688 48708 27445 48736
rect 27433 48705 27445 48708
rect 27479 48705 27491 48739
rect 27433 48699 27491 48705
rect 10134 48628 10140 48680
rect 10192 48668 10198 48680
rect 10321 48671 10379 48677
rect 10321 48668 10333 48671
rect 10192 48640 10333 48668
rect 10192 48628 10198 48640
rect 10321 48637 10333 48640
rect 10367 48637 10379 48671
rect 10321 48631 10379 48637
rect 10686 48628 10692 48680
rect 10744 48668 10750 48680
rect 10873 48671 10931 48677
rect 10873 48668 10885 48671
rect 10744 48640 10885 48668
rect 10744 48628 10750 48640
rect 10873 48637 10885 48640
rect 10919 48637 10931 48671
rect 10873 48631 10931 48637
rect 11054 48628 11060 48680
rect 11112 48628 11118 48680
rect 10045 48535 10103 48541
rect 10045 48501 10057 48535
rect 10091 48501 10103 48535
rect 10045 48495 10103 48501
rect 10137 48535 10195 48541
rect 10137 48501 10149 48535
rect 10183 48532 10195 48535
rect 11054 48532 11060 48544
rect 10183 48504 11060 48532
rect 10183 48501 10195 48504
rect 10137 48495 10195 48501
rect 11054 48492 11060 48504
rect 11112 48532 11118 48544
rect 12406 48532 12434 48696
rect 12894 48668 12900 48680
rect 12855 48640 12900 48668
rect 12894 48628 12900 48640
rect 12952 48628 12958 48680
rect 13170 48628 13176 48680
rect 13228 48668 13234 48680
rect 13265 48671 13323 48677
rect 13265 48668 13277 48671
rect 13228 48640 13277 48668
rect 13228 48628 13234 48640
rect 13265 48637 13277 48640
rect 13311 48637 13323 48671
rect 13265 48631 13323 48637
rect 13633 48671 13691 48677
rect 13633 48637 13645 48671
rect 13679 48668 13691 48671
rect 13906 48668 13912 48680
rect 13679 48640 13912 48668
rect 13679 48637 13691 48640
rect 13633 48631 13691 48637
rect 13906 48628 13912 48640
rect 13964 48628 13970 48680
rect 14550 48628 14556 48680
rect 14608 48668 14614 48680
rect 15105 48671 15163 48677
rect 15105 48668 15117 48671
rect 14608 48640 15117 48668
rect 14608 48628 14614 48640
rect 15105 48637 15117 48640
rect 15151 48637 15163 48671
rect 15105 48631 15163 48637
rect 16850 48628 16856 48680
rect 16908 48668 16914 48680
rect 17313 48671 17371 48677
rect 17313 48668 17325 48671
rect 16908 48640 17325 48668
rect 16908 48628 16914 48640
rect 17313 48637 17325 48640
rect 17359 48637 17371 48671
rect 17494 48668 17500 48680
rect 17455 48640 17500 48668
rect 17313 48631 17371 48637
rect 17494 48628 17500 48640
rect 17552 48628 17558 48680
rect 21358 48668 21364 48680
rect 21319 48640 21364 48668
rect 21358 48628 21364 48640
rect 21416 48628 21422 48680
rect 22830 48628 22836 48680
rect 22888 48668 22894 48680
rect 23017 48671 23075 48677
rect 23017 48668 23029 48671
rect 22888 48640 23029 48668
rect 22888 48628 22894 48640
rect 23017 48637 23029 48640
rect 23063 48637 23075 48671
rect 23198 48668 23204 48680
rect 23159 48640 23204 48668
rect 23017 48631 23075 48637
rect 23198 48628 23204 48640
rect 23256 48628 23262 48680
rect 24305 48671 24363 48677
rect 24305 48668 24317 48671
rect 24044 48640 24317 48668
rect 24044 48612 24072 48640
rect 24305 48637 24317 48640
rect 24351 48668 24363 48671
rect 24670 48668 24676 48680
rect 24351 48640 24676 48668
rect 24351 48637 24363 48640
rect 24305 48631 24363 48637
rect 24670 48628 24676 48640
rect 24728 48628 24734 48680
rect 25225 48671 25283 48677
rect 25225 48637 25237 48671
rect 25271 48668 25283 48671
rect 25314 48668 25320 48680
rect 25271 48640 25320 48668
rect 25271 48637 25283 48640
rect 25225 48631 25283 48637
rect 25314 48628 25320 48640
rect 25372 48628 25378 48680
rect 25498 48668 25504 48680
rect 25459 48640 25504 48668
rect 25498 48628 25504 48640
rect 25556 48628 25562 48680
rect 25685 48671 25743 48677
rect 25685 48637 25697 48671
rect 25731 48637 25743 48671
rect 26694 48668 26700 48680
rect 26655 48640 26700 48668
rect 25685 48631 25743 48637
rect 22186 48560 22192 48612
rect 22244 48600 22250 48612
rect 22373 48603 22431 48609
rect 22373 48600 22385 48603
rect 22244 48572 22385 48600
rect 22244 48560 22250 48572
rect 22373 48569 22385 48572
rect 22419 48569 22431 48603
rect 22373 48563 22431 48569
rect 22557 48603 22615 48609
rect 22557 48569 22569 48603
rect 22603 48600 22615 48603
rect 22738 48600 22744 48612
rect 22603 48572 22744 48600
rect 22603 48569 22615 48572
rect 22557 48563 22615 48569
rect 22738 48560 22744 48572
rect 22796 48560 22802 48612
rect 23385 48603 23443 48609
rect 23385 48569 23397 48603
rect 23431 48600 23443 48603
rect 23934 48600 23940 48612
rect 23431 48572 23940 48600
rect 23431 48569 23443 48572
rect 23385 48563 23443 48569
rect 23934 48560 23940 48572
rect 23992 48560 23998 48612
rect 24026 48560 24032 48612
rect 24084 48560 24090 48612
rect 25700 48600 25728 48631
rect 26694 48628 26700 48640
rect 26752 48628 26758 48680
rect 27154 48628 27160 48680
rect 27212 48668 27218 48680
rect 27249 48671 27307 48677
rect 27249 48668 27261 48671
rect 27212 48640 27261 48668
rect 27212 48628 27218 48640
rect 27249 48637 27261 48640
rect 27295 48637 27307 48671
rect 27982 48668 27988 48680
rect 27943 48640 27988 48668
rect 27249 48631 27307 48637
rect 27982 48628 27988 48640
rect 28040 48628 28046 48680
rect 24136 48572 25728 48600
rect 17678 48532 17684 48544
rect 11112 48504 12434 48532
rect 17639 48504 17684 48532
rect 11112 48492 11118 48504
rect 17678 48492 17684 48504
rect 17736 48492 17742 48544
rect 24136 48541 24164 48572
rect 24121 48535 24179 48541
rect 24121 48501 24133 48535
rect 24167 48501 24179 48535
rect 24121 48495 24179 48501
rect 24213 48535 24271 48541
rect 24213 48501 24225 48535
rect 24259 48532 24271 48535
rect 24578 48532 24584 48544
rect 24259 48504 24584 48532
rect 24259 48501 24271 48504
rect 24213 48495 24271 48501
rect 24578 48492 24584 48504
rect 24636 48532 24642 48544
rect 24762 48532 24768 48544
rect 24636 48504 24768 48532
rect 24636 48492 24642 48504
rect 24762 48492 24768 48504
rect 24820 48492 24826 48544
rect 25314 48492 25320 48544
rect 25372 48532 25378 48544
rect 26142 48532 26148 48544
rect 25372 48504 26148 48532
rect 25372 48492 25378 48504
rect 26142 48492 26148 48504
rect 26200 48492 26206 48544
rect 26510 48532 26516 48544
rect 26471 48504 26516 48532
rect 26510 48492 26516 48504
rect 26568 48492 26574 48544
rect 1104 48442 28888 48464
rect 1104 48390 10246 48442
rect 10298 48390 10310 48442
rect 10362 48390 10374 48442
rect 10426 48390 10438 48442
rect 10490 48390 19510 48442
rect 19562 48390 19574 48442
rect 19626 48390 19638 48442
rect 19690 48390 19702 48442
rect 19754 48390 28888 48442
rect 1104 48368 28888 48390
rect 4341 48331 4399 48337
rect 4341 48297 4353 48331
rect 4387 48328 4399 48331
rect 4614 48328 4620 48340
rect 4387 48300 4620 48328
rect 4387 48297 4399 48300
rect 4341 48291 4399 48297
rect 4614 48288 4620 48300
rect 4672 48288 4678 48340
rect 4706 48288 4712 48340
rect 4764 48328 4770 48340
rect 4801 48331 4859 48337
rect 4801 48328 4813 48331
rect 4764 48300 4813 48328
rect 4764 48288 4770 48300
rect 4801 48297 4813 48300
rect 4847 48297 4859 48331
rect 4801 48291 4859 48297
rect 5169 48331 5227 48337
rect 5169 48297 5181 48331
rect 5215 48328 5227 48331
rect 5258 48328 5264 48340
rect 5215 48300 5264 48328
rect 5215 48297 5227 48300
rect 5169 48291 5227 48297
rect 5258 48288 5264 48300
rect 5316 48288 5322 48340
rect 7098 48328 7104 48340
rect 7059 48300 7104 48328
rect 7098 48288 7104 48300
rect 7156 48288 7162 48340
rect 10045 48331 10103 48337
rect 10045 48297 10057 48331
rect 10091 48328 10103 48331
rect 10134 48328 10140 48340
rect 10091 48300 10140 48328
rect 10091 48297 10103 48300
rect 10045 48291 10103 48297
rect 10134 48288 10140 48300
rect 10192 48288 10198 48340
rect 11054 48328 11060 48340
rect 11015 48300 11060 48328
rect 11054 48288 11060 48300
rect 11112 48288 11118 48340
rect 20254 48328 20260 48340
rect 16776 48300 18460 48328
rect 3228 48263 3286 48269
rect 3228 48229 3240 48263
rect 3274 48260 3286 48263
rect 4246 48260 4252 48272
rect 3274 48232 4252 48260
rect 3274 48229 3286 48232
rect 3228 48223 3286 48229
rect 4246 48220 4252 48232
rect 4304 48220 4310 48272
rect 8202 48220 8208 48272
rect 8260 48260 8266 48272
rect 8481 48263 8539 48269
rect 8481 48260 8493 48263
rect 8260 48232 8493 48260
rect 8260 48220 8266 48232
rect 8481 48229 8493 48232
rect 8527 48229 8539 48263
rect 10873 48263 10931 48269
rect 8481 48223 8539 48229
rect 8588 48232 10180 48260
rect 1857 48195 1915 48201
rect 1857 48161 1869 48195
rect 1903 48192 1915 48195
rect 7098 48192 7104 48204
rect 1903 48164 6960 48192
rect 7059 48164 7104 48192
rect 1903 48161 1915 48164
rect 1857 48155 1915 48161
rect 1210 48084 1216 48136
rect 1268 48124 1274 48136
rect 2958 48124 2964 48136
rect 1268 48096 2964 48124
rect 1268 48084 1274 48096
rect 2958 48084 2964 48096
rect 3016 48084 3022 48136
rect 5261 48127 5319 48133
rect 5261 48093 5273 48127
rect 5307 48093 5319 48127
rect 5442 48124 5448 48136
rect 5403 48096 5448 48124
rect 5261 48087 5319 48093
rect 2041 48059 2099 48065
rect 2041 48025 2053 48059
rect 2087 48056 2099 48059
rect 2866 48056 2872 48068
rect 2087 48028 2872 48056
rect 2087 48025 2099 48028
rect 2041 48019 2099 48025
rect 2866 48016 2872 48028
rect 2924 48016 2930 48068
rect 5276 48056 5304 48087
rect 5442 48084 5448 48096
rect 5500 48084 5506 48136
rect 6932 48124 6960 48164
rect 7098 48152 7104 48164
rect 7156 48152 7162 48204
rect 7190 48152 7196 48204
rect 7248 48192 7254 48204
rect 7285 48195 7343 48201
rect 7285 48192 7297 48195
rect 7248 48164 7297 48192
rect 7248 48152 7254 48164
rect 7285 48161 7297 48164
rect 7331 48161 7343 48195
rect 7285 48155 7343 48161
rect 8294 48152 8300 48204
rect 8352 48192 8358 48204
rect 8389 48195 8447 48201
rect 8389 48192 8401 48195
rect 8352 48164 8401 48192
rect 8352 48152 8358 48164
rect 8389 48161 8401 48164
rect 8435 48161 8447 48195
rect 8588 48192 8616 48232
rect 8389 48155 8447 48161
rect 8496 48164 8616 48192
rect 8496 48124 8524 48164
rect 9582 48152 9588 48204
rect 9640 48192 9646 48204
rect 9769 48195 9827 48201
rect 9769 48192 9781 48195
rect 9640 48164 9781 48192
rect 9640 48152 9646 48164
rect 9769 48161 9781 48164
rect 9815 48161 9827 48195
rect 9769 48155 9827 48161
rect 9858 48152 9864 48204
rect 9916 48192 9922 48204
rect 9916 48164 9961 48192
rect 9916 48152 9922 48164
rect 6932 48096 8524 48124
rect 8570 48084 8576 48136
rect 8628 48124 8634 48136
rect 10042 48124 10048 48136
rect 8628 48096 8673 48124
rect 10003 48096 10048 48124
rect 8628 48084 8634 48096
rect 10042 48084 10048 48096
rect 10100 48084 10106 48136
rect 10152 48124 10180 48232
rect 10873 48229 10885 48263
rect 10919 48260 10931 48263
rect 10962 48260 10968 48272
rect 10919 48232 10968 48260
rect 10919 48229 10931 48232
rect 10873 48223 10931 48229
rect 10962 48220 10968 48232
rect 11020 48220 11026 48272
rect 11146 48192 11152 48204
rect 11107 48164 11152 48192
rect 11146 48152 11152 48164
rect 11204 48152 11210 48204
rect 16776 48124 16804 48300
rect 16850 48220 16856 48272
rect 16908 48260 16914 48272
rect 16908 48232 17540 48260
rect 16908 48220 16914 48232
rect 17313 48195 17371 48201
rect 17313 48161 17325 48195
rect 17359 48192 17371 48195
rect 17402 48192 17408 48204
rect 17359 48164 17408 48192
rect 17359 48161 17371 48164
rect 17313 48155 17371 48161
rect 17402 48152 17408 48164
rect 17460 48152 17466 48204
rect 17512 48201 17540 48232
rect 17678 48220 17684 48272
rect 17736 48260 17742 48272
rect 18432 48260 18460 48300
rect 20088 48300 20260 48328
rect 17736 48232 18368 48260
rect 18432 48232 19380 48260
rect 17736 48220 17742 48232
rect 17497 48195 17555 48201
rect 17497 48161 17509 48195
rect 17543 48161 17555 48195
rect 18138 48192 18144 48204
rect 18099 48164 18144 48192
rect 17497 48155 17555 48161
rect 18138 48152 18144 48164
rect 18196 48152 18202 48204
rect 18340 48201 18368 48232
rect 18325 48195 18383 48201
rect 18325 48161 18337 48195
rect 18371 48161 18383 48195
rect 18325 48155 18383 48161
rect 18874 48152 18880 48204
rect 18932 48192 18938 48204
rect 19245 48195 19303 48201
rect 19245 48192 19257 48195
rect 18932 48164 19257 48192
rect 18932 48152 18938 48164
rect 19245 48161 19257 48164
rect 19291 48161 19303 48195
rect 19245 48155 19303 48161
rect 18046 48124 18052 48136
rect 10152 48096 16804 48124
rect 17328 48096 18052 48124
rect 5902 48056 5908 48068
rect 5276 48028 5908 48056
rect 5902 48016 5908 48028
rect 5960 48016 5966 48068
rect 6730 48016 6736 48068
rect 6788 48056 6794 48068
rect 17328 48065 17356 48096
rect 18046 48084 18052 48096
rect 18104 48124 18110 48136
rect 18417 48127 18475 48133
rect 18417 48124 18429 48127
rect 18104 48096 18429 48124
rect 18104 48084 18110 48096
rect 18417 48093 18429 48096
rect 18463 48093 18475 48127
rect 18417 48087 18475 48093
rect 18506 48084 18512 48136
rect 18564 48124 18570 48136
rect 19061 48127 19119 48133
rect 19061 48124 19073 48127
rect 18564 48096 19073 48124
rect 18564 48084 18570 48096
rect 19061 48093 19073 48096
rect 19107 48093 19119 48127
rect 19061 48087 19119 48093
rect 8021 48059 8079 48065
rect 8021 48056 8033 48059
rect 6788 48028 8033 48056
rect 6788 48016 6794 48028
rect 8021 48025 8033 48028
rect 8067 48025 8079 48059
rect 17313 48059 17371 48065
rect 8021 48019 8079 48025
rect 8128 48028 12434 48056
rect 2682 47948 2688 48000
rect 2740 47988 2746 48000
rect 8128 47988 8156 48028
rect 10870 47988 10876 48000
rect 2740 47960 8156 47988
rect 10831 47960 10876 47988
rect 2740 47948 2746 47960
rect 10870 47948 10876 47960
rect 10928 47948 10934 48000
rect 12406 47988 12434 48028
rect 17313 48025 17325 48059
rect 17359 48025 17371 48059
rect 17313 48019 17371 48025
rect 17957 48059 18015 48065
rect 17957 48025 17969 48059
rect 18003 48056 18015 48059
rect 18877 48059 18935 48065
rect 18877 48056 18889 48059
rect 18003 48028 18889 48056
rect 18003 48025 18015 48028
rect 17957 48019 18015 48025
rect 18877 48025 18889 48028
rect 18923 48025 18935 48059
rect 19352 48056 19380 48232
rect 20088 48201 20116 48300
rect 20254 48288 20260 48300
rect 20312 48288 20318 48340
rect 24397 48331 24455 48337
rect 24397 48297 24409 48331
rect 24443 48328 24455 48331
rect 24578 48328 24584 48340
rect 24443 48300 24584 48328
rect 24443 48297 24455 48300
rect 24397 48291 24455 48297
rect 24578 48288 24584 48300
rect 24636 48288 24642 48340
rect 20165 48263 20223 48269
rect 20165 48229 20177 48263
rect 20211 48260 20223 48263
rect 20717 48263 20775 48269
rect 20717 48260 20729 48263
rect 20211 48232 20729 48260
rect 20211 48229 20223 48232
rect 20165 48223 20223 48229
rect 20717 48229 20729 48232
rect 20763 48229 20775 48263
rect 20717 48223 20775 48229
rect 23934 48220 23940 48272
rect 23992 48260 23998 48272
rect 23992 48232 24624 48260
rect 23992 48220 23998 48232
rect 20073 48195 20131 48201
rect 20073 48161 20085 48195
rect 20119 48161 20131 48195
rect 20073 48155 20131 48161
rect 20257 48195 20315 48201
rect 20257 48161 20269 48195
rect 20303 48192 20315 48195
rect 20438 48192 20444 48204
rect 20303 48164 20444 48192
rect 20303 48161 20315 48164
rect 20257 48155 20315 48161
rect 20438 48152 20444 48164
rect 20496 48192 20502 48204
rect 20622 48192 20628 48204
rect 20496 48164 20628 48192
rect 20496 48152 20502 48164
rect 20622 48152 20628 48164
rect 20680 48152 20686 48204
rect 20901 48195 20959 48201
rect 20901 48161 20913 48195
rect 20947 48161 20959 48195
rect 20901 48155 20959 48161
rect 20993 48195 21051 48201
rect 20993 48161 21005 48195
rect 21039 48192 21051 48195
rect 21082 48192 21088 48204
rect 21039 48164 21088 48192
rect 21039 48161 21051 48164
rect 20993 48155 21051 48161
rect 19978 48084 19984 48136
rect 20036 48124 20042 48136
rect 20916 48124 20944 48155
rect 21082 48152 21088 48164
rect 21140 48192 21146 48204
rect 21358 48192 21364 48204
rect 21140 48164 21364 48192
rect 21140 48152 21146 48164
rect 21358 48152 21364 48164
rect 21416 48152 21422 48204
rect 23198 48192 23204 48204
rect 23159 48164 23204 48192
rect 23198 48152 23204 48164
rect 23256 48152 23262 48204
rect 24026 48152 24032 48204
rect 24084 48192 24090 48204
rect 24213 48195 24271 48201
rect 24213 48192 24225 48195
rect 24084 48164 24225 48192
rect 24084 48152 24090 48164
rect 24213 48161 24225 48164
rect 24259 48161 24271 48195
rect 24213 48155 24271 48161
rect 24351 48195 24409 48201
rect 24351 48161 24363 48195
rect 24397 48192 24409 48195
rect 24486 48192 24492 48204
rect 24397 48164 24492 48192
rect 24397 48161 24409 48164
rect 24351 48155 24409 48161
rect 24486 48152 24492 48164
rect 24544 48152 24550 48204
rect 24596 48201 24624 48232
rect 27890 48220 27896 48272
rect 27948 48260 27954 48272
rect 27985 48263 28043 48269
rect 27985 48260 27997 48263
rect 27948 48232 27997 48260
rect 27948 48220 27954 48232
rect 27985 48229 27997 48232
rect 28031 48229 28043 48263
rect 27985 48223 28043 48229
rect 24581 48195 24639 48201
rect 24581 48161 24593 48195
rect 24627 48161 24639 48195
rect 25590 48192 25596 48204
rect 25551 48164 25596 48192
rect 24581 48155 24639 48161
rect 25590 48152 25596 48164
rect 25648 48152 25654 48204
rect 26234 48192 26240 48204
rect 26195 48164 26240 48192
rect 26234 48152 26240 48164
rect 26292 48152 26298 48204
rect 26881 48195 26939 48201
rect 26881 48161 26893 48195
rect 26927 48192 26939 48195
rect 26970 48192 26976 48204
rect 26927 48164 26976 48192
rect 26927 48161 26939 48164
rect 26881 48155 26939 48161
rect 26970 48152 26976 48164
rect 27028 48152 27034 48204
rect 21174 48124 21180 48136
rect 20036 48096 21180 48124
rect 20036 48084 20042 48096
rect 21174 48084 21180 48096
rect 21232 48084 21238 48136
rect 22830 48084 22836 48136
rect 22888 48124 22894 48136
rect 23017 48127 23075 48133
rect 23017 48124 23029 48127
rect 22888 48096 23029 48124
rect 22888 48084 22894 48096
rect 23017 48093 23029 48096
rect 23063 48093 23075 48127
rect 24670 48124 24676 48136
rect 23017 48087 23075 48093
rect 24044 48096 24676 48124
rect 21358 48056 21364 48068
rect 19352 48028 21364 48056
rect 18877 48019 18935 48025
rect 21358 48016 21364 48028
rect 21416 48016 21422 48068
rect 24044 48065 24072 48096
rect 24670 48084 24676 48096
rect 24728 48084 24734 48136
rect 24029 48059 24087 48065
rect 24029 48025 24041 48059
rect 24075 48025 24087 48059
rect 28169 48059 28227 48065
rect 28169 48056 28181 48059
rect 24029 48019 24087 48025
rect 24136 48028 28181 48056
rect 18782 47988 18788 48000
rect 12406 47960 18788 47988
rect 18782 47948 18788 47960
rect 18840 47948 18846 48000
rect 19058 47988 19064 48000
rect 19019 47960 19064 47988
rect 19058 47948 19064 47960
rect 19116 47948 19122 48000
rect 19153 47991 19211 47997
rect 19153 47957 19165 47991
rect 19199 47988 19211 47991
rect 19242 47988 19248 48000
rect 19199 47960 19248 47988
rect 19199 47957 19211 47960
rect 19153 47951 19211 47957
rect 19242 47948 19248 47960
rect 19300 47948 19306 48000
rect 20254 47948 20260 48000
rect 20312 47988 20318 48000
rect 20438 47988 20444 48000
rect 20312 47960 20444 47988
rect 20312 47948 20318 47960
rect 20438 47948 20444 47960
rect 20496 47948 20502 48000
rect 20717 47991 20775 47997
rect 20717 47957 20729 47991
rect 20763 47988 20775 47991
rect 21266 47988 21272 48000
rect 20763 47960 21272 47988
rect 20763 47957 20775 47960
rect 20717 47951 20775 47957
rect 21266 47948 21272 47960
rect 21324 47948 21330 48000
rect 23385 47991 23443 47997
rect 23385 47957 23397 47991
rect 23431 47988 23443 47991
rect 23842 47988 23848 48000
rect 23431 47960 23848 47988
rect 23431 47957 23443 47960
rect 23385 47951 23443 47957
rect 23842 47948 23848 47960
rect 23900 47948 23906 48000
rect 23934 47948 23940 48000
rect 23992 47988 23998 48000
rect 24136 47988 24164 48028
rect 28169 48025 28181 48028
rect 28215 48025 28227 48059
rect 28169 48019 28227 48025
rect 23992 47960 24164 47988
rect 25409 47991 25467 47997
rect 23992 47948 23998 47960
rect 25409 47957 25421 47991
rect 25455 47988 25467 47991
rect 25958 47988 25964 48000
rect 25455 47960 25964 47988
rect 25455 47957 25467 47960
rect 25409 47951 25467 47957
rect 25958 47948 25964 47960
rect 26016 47948 26022 48000
rect 26050 47948 26056 48000
rect 26108 47988 26114 48000
rect 26697 47991 26755 47997
rect 26108 47960 26153 47988
rect 26108 47948 26114 47960
rect 26697 47957 26709 47991
rect 26743 47988 26755 47991
rect 27890 47988 27896 48000
rect 26743 47960 27896 47988
rect 26743 47957 26755 47960
rect 26697 47951 26755 47957
rect 27890 47948 27896 47960
rect 27948 47948 27954 48000
rect 1104 47898 28888 47920
rect 1104 47846 5614 47898
rect 5666 47846 5678 47898
rect 5730 47846 5742 47898
rect 5794 47846 5806 47898
rect 5858 47846 14878 47898
rect 14930 47846 14942 47898
rect 14994 47846 15006 47898
rect 15058 47846 15070 47898
rect 15122 47846 24142 47898
rect 24194 47846 24206 47898
rect 24258 47846 24270 47898
rect 24322 47846 24334 47898
rect 24386 47846 28888 47898
rect 1104 47824 28888 47846
rect 2590 47784 2596 47796
rect 2551 47756 2596 47784
rect 2590 47744 2596 47756
rect 2648 47744 2654 47796
rect 23934 47784 23940 47796
rect 2746 47756 23940 47784
rect 1854 47676 1860 47728
rect 1912 47716 1918 47728
rect 2746 47716 2774 47756
rect 23934 47744 23940 47756
rect 23992 47744 23998 47796
rect 24213 47787 24271 47793
rect 24213 47753 24225 47787
rect 24259 47784 24271 47787
rect 24486 47784 24492 47796
rect 24259 47756 24492 47784
rect 24259 47753 24271 47756
rect 24213 47747 24271 47753
rect 24486 47744 24492 47756
rect 24544 47744 24550 47796
rect 1912 47688 2774 47716
rect 6641 47719 6699 47725
rect 1912 47676 1918 47688
rect 6641 47685 6653 47719
rect 6687 47716 6699 47719
rect 7282 47716 7288 47728
rect 6687 47688 7288 47716
rect 6687 47685 6699 47688
rect 6641 47679 6699 47685
rect 7282 47676 7288 47688
rect 7340 47676 7346 47728
rect 18509 47719 18567 47725
rect 18509 47685 18521 47719
rect 18555 47716 18567 47719
rect 19978 47716 19984 47728
rect 18555 47688 19984 47716
rect 18555 47685 18567 47688
rect 18509 47679 18567 47685
rect 19978 47676 19984 47688
rect 20036 47676 20042 47728
rect 20073 47719 20131 47725
rect 20073 47685 20085 47719
rect 20119 47716 20131 47719
rect 20162 47716 20168 47728
rect 20119 47688 20168 47716
rect 20119 47685 20131 47688
rect 20073 47679 20131 47685
rect 20162 47676 20168 47688
rect 20220 47676 20226 47728
rect 3237 47651 3295 47657
rect 3237 47617 3249 47651
rect 3283 47648 3295 47651
rect 5166 47648 5172 47660
rect 3283 47620 5172 47648
rect 3283 47617 3295 47620
rect 3237 47611 3295 47617
rect 5166 47608 5172 47620
rect 5224 47608 5230 47660
rect 6578 47620 6684 47648
rect 6656 47592 6684 47620
rect 9030 47608 9036 47660
rect 9088 47648 9094 47660
rect 9088 47620 11008 47648
rect 9088 47608 9094 47620
rect 4525 47583 4583 47589
rect 4525 47549 4537 47583
rect 4571 47580 4583 47583
rect 4614 47580 4620 47592
rect 4571 47552 4620 47580
rect 4571 47549 4583 47552
rect 4525 47543 4583 47549
rect 4614 47540 4620 47552
rect 4672 47540 4678 47592
rect 5810 47580 5816 47592
rect 5771 47552 5816 47580
rect 5810 47540 5816 47552
rect 5868 47540 5874 47592
rect 5905 47583 5963 47589
rect 5905 47549 5917 47583
rect 5951 47549 5963 47583
rect 6454 47580 6460 47592
rect 6415 47552 6460 47580
rect 5905 47543 5963 47549
rect 1857 47515 1915 47521
rect 1857 47481 1869 47515
rect 1903 47512 1915 47515
rect 2590 47512 2596 47524
rect 1903 47484 2596 47512
rect 1903 47481 1915 47484
rect 1857 47475 1915 47481
rect 2590 47472 2596 47484
rect 2648 47472 2654 47524
rect 2961 47515 3019 47521
rect 2961 47481 2973 47515
rect 3007 47512 3019 47515
rect 4154 47512 4160 47524
rect 3007 47484 4160 47512
rect 3007 47481 3019 47484
rect 2961 47475 3019 47481
rect 4154 47472 4160 47484
rect 4212 47512 4218 47524
rect 4890 47512 4896 47524
rect 4212 47484 4896 47512
rect 4212 47472 4218 47484
rect 4890 47472 4896 47484
rect 4948 47472 4954 47524
rect 5718 47472 5724 47524
rect 5776 47512 5782 47524
rect 5920 47512 5948 47543
rect 6454 47540 6460 47552
rect 6512 47540 6518 47592
rect 6638 47540 6644 47592
rect 6696 47540 6702 47592
rect 6822 47540 6828 47592
rect 6880 47580 6886 47592
rect 7101 47583 7159 47589
rect 7101 47580 7113 47583
rect 6880 47552 7113 47580
rect 6880 47540 6886 47552
rect 7101 47549 7113 47552
rect 7147 47549 7159 47583
rect 7101 47543 7159 47549
rect 7561 47583 7619 47589
rect 7561 47549 7573 47583
rect 7607 47549 7619 47583
rect 7561 47543 7619 47549
rect 6270 47512 6276 47524
rect 5776 47484 6276 47512
rect 5776 47472 5782 47484
rect 6270 47472 6276 47484
rect 6328 47512 6334 47524
rect 7576 47512 7604 47543
rect 8938 47540 8944 47592
rect 8996 47580 9002 47592
rect 9493 47583 9551 47589
rect 9493 47580 9505 47583
rect 8996 47552 9505 47580
rect 8996 47540 9002 47552
rect 9493 47549 9505 47552
rect 9539 47549 9551 47583
rect 9493 47543 9551 47549
rect 9677 47583 9735 47589
rect 9677 47549 9689 47583
rect 9723 47580 9735 47583
rect 9858 47580 9864 47592
rect 9723 47552 9864 47580
rect 9723 47549 9735 47552
rect 9677 47543 9735 47549
rect 9858 47540 9864 47552
rect 9916 47580 9922 47592
rect 10980 47589 11008 47620
rect 15194 47608 15200 47660
rect 15252 47648 15258 47660
rect 15470 47648 15476 47660
rect 15252 47620 15476 47648
rect 15252 47608 15258 47620
rect 15470 47608 15476 47620
rect 15528 47648 15534 47660
rect 15657 47651 15715 47657
rect 15657 47648 15669 47651
rect 15528 47620 15669 47648
rect 15528 47608 15534 47620
rect 15657 47617 15669 47620
rect 15703 47617 15715 47651
rect 15657 47611 15715 47617
rect 17678 47608 17684 47660
rect 17736 47648 17742 47660
rect 17736 47620 18736 47648
rect 17736 47608 17742 47620
rect 10321 47583 10379 47589
rect 10321 47580 10333 47583
rect 9916 47552 10333 47580
rect 9916 47540 9922 47552
rect 10321 47549 10333 47552
rect 10367 47549 10379 47583
rect 10321 47543 10379 47549
rect 10505 47583 10563 47589
rect 10505 47549 10517 47583
rect 10551 47549 10563 47583
rect 10505 47543 10563 47549
rect 10965 47583 11023 47589
rect 10965 47549 10977 47583
rect 11011 47549 11023 47583
rect 18046 47580 18052 47592
rect 18007 47552 18052 47580
rect 10965 47543 11023 47549
rect 8386 47512 8392 47524
rect 6328 47484 7604 47512
rect 8347 47484 8392 47512
rect 6328 47472 6334 47484
rect 8386 47472 8392 47484
rect 8444 47472 8450 47524
rect 8570 47472 8576 47524
rect 8628 47512 8634 47524
rect 9582 47512 9588 47524
rect 8628 47484 9588 47512
rect 8628 47472 8634 47484
rect 9582 47472 9588 47484
rect 9640 47512 9646 47524
rect 10520 47512 10548 47543
rect 18046 47540 18052 47552
rect 18104 47540 18110 47592
rect 18138 47540 18144 47592
rect 18196 47580 18202 47592
rect 18708 47589 18736 47620
rect 19794 47608 19800 47660
rect 19852 47648 19858 47660
rect 20257 47651 20315 47657
rect 20257 47648 20269 47651
rect 19852 47620 20269 47648
rect 19852 47608 19858 47620
rect 20257 47617 20269 47620
rect 20303 47617 20315 47651
rect 21266 47648 21272 47660
rect 21227 47620 21272 47648
rect 20257 47611 20315 47617
rect 21266 47608 21272 47620
rect 21324 47608 21330 47660
rect 27985 47651 28043 47657
rect 27985 47648 27997 47651
rect 22066 47620 27997 47648
rect 18417 47583 18475 47589
rect 18417 47580 18429 47583
rect 18196 47552 18429 47580
rect 18196 47540 18202 47552
rect 18417 47549 18429 47552
rect 18463 47549 18475 47583
rect 18417 47543 18475 47549
rect 18693 47583 18751 47589
rect 18693 47549 18705 47583
rect 18739 47549 18751 47583
rect 18693 47543 18751 47549
rect 19981 47583 20039 47589
rect 19981 47549 19993 47583
rect 20027 47580 20039 47583
rect 20070 47580 20076 47592
rect 20027 47552 20076 47580
rect 20027 47549 20039 47552
rect 19981 47543 20039 47549
rect 20070 47540 20076 47552
rect 20128 47580 20134 47592
rect 20898 47580 20904 47592
rect 20128 47552 20904 47580
rect 20128 47540 20134 47552
rect 20898 47540 20904 47552
rect 20956 47540 20962 47592
rect 20990 47540 20996 47592
rect 21048 47580 21054 47592
rect 21361 47583 21419 47589
rect 21361 47580 21373 47583
rect 21048 47552 21373 47580
rect 21048 47540 21054 47552
rect 21361 47549 21373 47552
rect 21407 47549 21419 47583
rect 21361 47543 21419 47549
rect 9640 47484 10548 47512
rect 15924 47515 15982 47521
rect 9640 47472 9646 47484
rect 15924 47481 15936 47515
rect 15970 47512 15982 47515
rect 16206 47512 16212 47524
rect 15970 47484 16212 47512
rect 15970 47481 15982 47484
rect 15924 47475 15982 47481
rect 16206 47472 16212 47484
rect 16264 47472 16270 47524
rect 18782 47472 18788 47524
rect 18840 47512 18846 47524
rect 22066 47512 22094 47620
rect 27985 47617 27997 47620
rect 28031 47617 28043 47651
rect 27985 47611 28043 47617
rect 23842 47540 23848 47592
rect 23900 47580 23906 47592
rect 24121 47583 24179 47589
rect 24121 47580 24133 47583
rect 23900 47552 24133 47580
rect 23900 47540 23906 47552
rect 24121 47549 24133 47552
rect 24167 47549 24179 47583
rect 24121 47543 24179 47549
rect 25406 47540 25412 47592
rect 25464 47580 25470 47592
rect 25593 47583 25651 47589
rect 25593 47580 25605 47583
rect 25464 47552 25605 47580
rect 25464 47540 25470 47552
rect 25593 47549 25605 47552
rect 25639 47549 25651 47583
rect 25866 47580 25872 47592
rect 25827 47552 25872 47580
rect 25593 47543 25651 47549
rect 25866 47540 25872 47552
rect 25924 47540 25930 47592
rect 25958 47540 25964 47592
rect 26016 47580 26022 47592
rect 27801 47583 27859 47589
rect 27801 47580 27813 47583
rect 26016 47552 27813 47580
rect 26016 47540 26022 47552
rect 27801 47549 27813 47552
rect 27847 47549 27859 47583
rect 27801 47543 27859 47549
rect 18840 47484 22094 47512
rect 18840 47472 18846 47484
rect 1946 47444 1952 47456
rect 1907 47416 1952 47444
rect 1946 47404 1952 47416
rect 2004 47404 2010 47456
rect 3050 47444 3056 47456
rect 3011 47416 3056 47444
rect 3050 47404 3056 47416
rect 3108 47404 3114 47456
rect 4614 47444 4620 47456
rect 4575 47416 4620 47444
rect 4614 47404 4620 47416
rect 4672 47404 4678 47456
rect 7098 47404 7104 47456
rect 7156 47444 7162 47456
rect 7193 47447 7251 47453
rect 7193 47444 7205 47447
rect 7156 47416 7205 47444
rect 7156 47404 7162 47416
rect 7193 47413 7205 47416
rect 7239 47413 7251 47447
rect 7193 47407 7251 47413
rect 8481 47447 8539 47453
rect 8481 47413 8493 47447
rect 8527 47444 8539 47447
rect 8662 47444 8668 47456
rect 8527 47416 8668 47444
rect 8527 47413 8539 47416
rect 8481 47407 8539 47413
rect 8662 47404 8668 47416
rect 8720 47404 8726 47456
rect 9858 47444 9864 47456
rect 9819 47416 9864 47444
rect 9858 47404 9864 47416
rect 9916 47404 9922 47456
rect 10134 47404 10140 47456
rect 10192 47444 10198 47456
rect 10413 47447 10471 47453
rect 10413 47444 10425 47447
rect 10192 47416 10425 47444
rect 10192 47404 10198 47416
rect 10413 47413 10425 47416
rect 10459 47413 10471 47447
rect 11054 47444 11060 47456
rect 11015 47416 11060 47444
rect 10413 47407 10471 47413
rect 11054 47404 11060 47416
rect 11112 47404 11118 47456
rect 17034 47444 17040 47456
rect 16995 47416 17040 47444
rect 17034 47404 17040 47416
rect 17092 47404 17098 47456
rect 20257 47447 20315 47453
rect 20257 47413 20269 47447
rect 20303 47444 20315 47447
rect 21266 47444 21272 47456
rect 20303 47416 21272 47444
rect 20303 47413 20315 47416
rect 20257 47407 20315 47413
rect 21266 47404 21272 47416
rect 21324 47404 21330 47456
rect 21726 47444 21732 47456
rect 21687 47416 21732 47444
rect 21726 47404 21732 47416
rect 21784 47404 21790 47456
rect 25958 47404 25964 47456
rect 26016 47444 26022 47456
rect 26973 47447 27031 47453
rect 26973 47444 26985 47447
rect 26016 47416 26985 47444
rect 26016 47404 26022 47416
rect 26973 47413 26985 47416
rect 27019 47413 27031 47447
rect 26973 47407 27031 47413
rect 1104 47354 28888 47376
rect 1104 47302 10246 47354
rect 10298 47302 10310 47354
rect 10362 47302 10374 47354
rect 10426 47302 10438 47354
rect 10490 47302 19510 47354
rect 19562 47302 19574 47354
rect 19626 47302 19638 47354
rect 19690 47302 19702 47354
rect 19754 47302 28888 47354
rect 1104 47280 28888 47302
rect 3786 47200 3792 47252
rect 3844 47240 3850 47252
rect 4893 47243 4951 47249
rect 4893 47240 4905 47243
rect 3844 47212 4905 47240
rect 3844 47200 3850 47212
rect 4893 47209 4905 47212
rect 4939 47209 4951 47243
rect 4893 47203 4951 47209
rect 5905 47243 5963 47249
rect 5905 47209 5917 47243
rect 5951 47240 5963 47243
rect 7190 47240 7196 47252
rect 5951 47212 7196 47240
rect 5951 47209 5963 47212
rect 5905 47203 5963 47209
rect 7190 47200 7196 47212
rect 7248 47200 7254 47252
rect 18325 47243 18383 47249
rect 9324 47212 18276 47240
rect 2041 47175 2099 47181
rect 2041 47141 2053 47175
rect 2087 47172 2099 47175
rect 2958 47172 2964 47184
rect 2087 47144 2964 47172
rect 2087 47141 2099 47144
rect 2041 47135 2099 47141
rect 2958 47132 2964 47144
rect 3016 47132 3022 47184
rect 4801 47175 4859 47181
rect 4801 47141 4813 47175
rect 4847 47172 4859 47175
rect 9324 47172 9352 47212
rect 9582 47172 9588 47184
rect 4847 47144 9352 47172
rect 9543 47144 9588 47172
rect 4847 47141 4859 47144
rect 4801 47135 4859 47141
rect 9582 47132 9588 47144
rect 9640 47132 9646 47184
rect 9858 47132 9864 47184
rect 9916 47172 9922 47184
rect 10594 47172 10600 47184
rect 9916 47144 10456 47172
rect 10555 47144 10600 47172
rect 9916 47132 9922 47144
rect 1857 47107 1915 47113
rect 1857 47073 1869 47107
rect 1903 47104 1915 47107
rect 2498 47104 2504 47116
rect 1903 47076 2504 47104
rect 1903 47073 1915 47076
rect 1857 47067 1915 47073
rect 2498 47064 2504 47076
rect 2556 47064 2562 47116
rect 2593 47107 2651 47113
rect 2593 47073 2605 47107
rect 2639 47104 2651 47107
rect 2682 47104 2688 47116
rect 2639 47076 2688 47104
rect 2639 47073 2651 47076
rect 2593 47067 2651 47073
rect 2682 47064 2688 47076
rect 2740 47064 2746 47116
rect 3326 47104 3332 47116
rect 3287 47076 3332 47104
rect 3326 47064 3332 47076
rect 3384 47064 3390 47116
rect 4065 47107 4123 47113
rect 4065 47073 4077 47107
rect 4111 47073 4123 47107
rect 5718 47104 5724 47116
rect 5679 47076 5724 47104
rect 4065 47067 4123 47073
rect 2774 46928 2780 46980
rect 2832 46968 2838 46980
rect 4080 46968 4108 47067
rect 5718 47064 5724 47076
rect 5776 47064 5782 47116
rect 7098 47104 7104 47116
rect 7059 47076 7104 47104
rect 7098 47064 7104 47076
rect 7156 47064 7162 47116
rect 7282 47104 7288 47116
rect 7243 47076 7288 47104
rect 7282 47064 7288 47076
rect 7340 47064 7346 47116
rect 8389 47107 8447 47113
rect 8389 47073 8401 47107
rect 8435 47104 8447 47107
rect 8938 47104 8944 47116
rect 8435 47076 8944 47104
rect 8435 47073 8447 47076
rect 8389 47067 8447 47073
rect 8938 47064 8944 47076
rect 8996 47064 9002 47116
rect 9398 47104 9404 47116
rect 9359 47076 9404 47104
rect 9398 47064 9404 47076
rect 9456 47064 9462 47116
rect 10134 47064 10140 47116
rect 10192 47104 10198 47116
rect 10428 47113 10456 47144
rect 10594 47132 10600 47144
rect 10652 47132 10658 47184
rect 12820 47144 13860 47172
rect 10229 47107 10287 47113
rect 10229 47104 10241 47107
rect 10192 47076 10241 47104
rect 10192 47064 10198 47076
rect 10229 47073 10241 47076
rect 10275 47073 10287 47107
rect 10229 47067 10287 47073
rect 10413 47107 10471 47113
rect 10413 47073 10425 47107
rect 10459 47073 10471 47107
rect 10413 47067 10471 47073
rect 10502 47064 10508 47116
rect 10560 47104 10566 47116
rect 12434 47104 12440 47116
rect 10560 47076 12440 47104
rect 10560 47064 10566 47076
rect 12434 47064 12440 47076
rect 12492 47104 12498 47116
rect 12618 47104 12624 47116
rect 12492 47076 12624 47104
rect 12492 47064 12498 47076
rect 12618 47064 12624 47076
rect 12676 47064 12682 47116
rect 12820 47048 12848 47144
rect 13832 47113 13860 47144
rect 13633 47107 13691 47113
rect 13633 47073 13645 47107
rect 13679 47073 13691 47107
rect 13633 47067 13691 47073
rect 13817 47107 13875 47113
rect 13817 47073 13829 47107
rect 13863 47073 13875 47107
rect 13817 47067 13875 47073
rect 5537 47039 5595 47045
rect 5537 47005 5549 47039
rect 5583 47036 5595 47039
rect 5902 47036 5908 47048
rect 5583 47008 5908 47036
rect 5583 47005 5595 47008
rect 5537 46999 5595 47005
rect 5902 46996 5908 47008
rect 5960 47036 5966 47048
rect 6822 47036 6828 47048
rect 5960 47008 6828 47036
rect 5960 46996 5966 47008
rect 6822 46996 6828 47008
rect 6880 46996 6886 47048
rect 7558 47036 7564 47048
rect 7519 47008 7564 47036
rect 7558 46996 7564 47008
rect 7616 46996 7622 47048
rect 9677 47039 9735 47045
rect 9677 47005 9689 47039
rect 9723 47036 9735 47039
rect 10962 47036 10968 47048
rect 9723 47008 10968 47036
rect 9723 47005 9735 47008
rect 9677 46999 9735 47005
rect 10962 46996 10968 47008
rect 11020 47036 11026 47048
rect 12526 47036 12532 47048
rect 11020 47008 12532 47036
rect 11020 46996 11026 47008
rect 12526 46996 12532 47008
rect 12584 46996 12590 47048
rect 12802 47036 12808 47048
rect 12763 47008 12808 47036
rect 12802 46996 12808 47008
rect 12860 46996 12866 47048
rect 13648 47036 13676 47067
rect 14090 47064 14096 47116
rect 14148 47104 14154 47116
rect 14642 47113 14648 47116
rect 14369 47107 14427 47113
rect 14369 47104 14381 47107
rect 14148 47076 14381 47104
rect 14148 47064 14154 47076
rect 14369 47073 14381 47076
rect 14415 47073 14427 47107
rect 14369 47067 14427 47073
rect 14636 47067 14648 47113
rect 14700 47104 14706 47116
rect 17865 47107 17923 47113
rect 14700 47076 14736 47104
rect 14642 47064 14648 47067
rect 14700 47064 14706 47076
rect 17865 47073 17877 47107
rect 17911 47104 17923 47107
rect 18046 47104 18052 47116
rect 17911 47076 18052 47104
rect 17911 47073 17923 47076
rect 17865 47067 17923 47073
rect 18046 47064 18052 47076
rect 18104 47064 18110 47116
rect 14182 47036 14188 47048
rect 13648 47008 14188 47036
rect 14182 46996 14188 47008
rect 14240 46996 14246 47048
rect 9125 46971 9183 46977
rect 2832 46940 2877 46968
rect 4080 46940 4292 46968
rect 2832 46928 2838 46940
rect 3418 46900 3424 46912
rect 3379 46872 3424 46900
rect 3418 46860 3424 46872
rect 3476 46860 3482 46912
rect 3510 46860 3516 46912
rect 3568 46900 3574 46912
rect 4157 46903 4215 46909
rect 4157 46900 4169 46903
rect 3568 46872 4169 46900
rect 3568 46860 3574 46872
rect 4157 46869 4169 46872
rect 4203 46869 4215 46903
rect 4264 46900 4292 46940
rect 9125 46937 9137 46971
rect 9171 46968 9183 46971
rect 9766 46968 9772 46980
rect 9171 46940 9772 46968
rect 9171 46937 9183 46940
rect 9125 46931 9183 46937
rect 9766 46928 9772 46940
rect 9824 46928 9830 46980
rect 11146 46928 11152 46980
rect 11204 46968 11210 46980
rect 14090 46968 14096 46980
rect 11204 46940 14096 46968
rect 11204 46928 11210 46940
rect 14090 46928 14096 46940
rect 14148 46928 14154 46980
rect 17678 46928 17684 46980
rect 17736 46968 17742 46980
rect 18003 46971 18061 46977
rect 18003 46968 18015 46971
rect 17736 46940 18015 46968
rect 17736 46928 17742 46940
rect 18003 46937 18015 46940
rect 18049 46937 18061 46971
rect 18138 46968 18144 46980
rect 18099 46940 18144 46968
rect 18003 46931 18061 46937
rect 18138 46928 18144 46940
rect 18196 46928 18202 46980
rect 18248 46968 18276 47212
rect 18325 47209 18337 47243
rect 18371 47240 18383 47243
rect 18506 47240 18512 47252
rect 18371 47212 18512 47240
rect 18371 47209 18383 47212
rect 18325 47203 18383 47209
rect 18506 47200 18512 47212
rect 18564 47200 18570 47252
rect 19794 47240 19800 47252
rect 19755 47212 19800 47240
rect 19794 47200 19800 47212
rect 19852 47200 19858 47252
rect 20162 47200 20168 47252
rect 20220 47200 20226 47252
rect 20809 47243 20867 47249
rect 20809 47209 20821 47243
rect 20855 47240 20867 47243
rect 23658 47240 23664 47252
rect 20855 47212 23664 47240
rect 20855 47209 20867 47212
rect 20809 47203 20867 47209
rect 23658 47200 23664 47212
rect 23716 47200 23722 47252
rect 24026 47200 24032 47252
rect 24084 47240 24090 47252
rect 24305 47243 24363 47249
rect 24305 47240 24317 47243
rect 24084 47212 24317 47240
rect 24084 47200 24090 47212
rect 24305 47209 24317 47212
rect 24351 47209 24363 47243
rect 24305 47203 24363 47209
rect 25409 47243 25467 47249
rect 25409 47209 25421 47243
rect 25455 47240 25467 47243
rect 25866 47240 25872 47252
rect 25455 47212 25872 47240
rect 25455 47209 25467 47212
rect 25409 47203 25467 47209
rect 25866 47200 25872 47212
rect 25924 47200 25930 47252
rect 20180 47172 20208 47200
rect 19168 47144 20208 47172
rect 18322 47064 18328 47116
rect 18380 47104 18386 47116
rect 19168 47113 19196 47144
rect 19153 47107 19211 47113
rect 18380 47076 18425 47104
rect 18380 47064 18386 47076
rect 19153 47073 19165 47107
rect 19199 47073 19211 47107
rect 19153 47067 19211 47073
rect 19337 47107 19395 47113
rect 19337 47073 19349 47107
rect 19383 47104 19395 47107
rect 19886 47104 19892 47116
rect 19383 47076 19892 47104
rect 19383 47073 19395 47076
rect 19337 47067 19395 47073
rect 19886 47064 19892 47076
rect 19944 47064 19950 47116
rect 19996 47113 20024 47144
rect 21726 47132 21732 47184
rect 21784 47172 21790 47184
rect 25777 47175 25835 47181
rect 25777 47172 25789 47175
rect 21784 47144 25789 47172
rect 21784 47132 21790 47144
rect 25777 47141 25789 47144
rect 25823 47141 25835 47175
rect 25777 47135 25835 47141
rect 26510 47132 26516 47184
rect 26568 47172 26574 47184
rect 26697 47175 26755 47181
rect 26697 47172 26709 47175
rect 26568 47144 26709 47172
rect 26568 47132 26574 47144
rect 26697 47141 26709 47144
rect 26743 47141 26755 47175
rect 27890 47172 27896 47184
rect 27851 47144 27896 47172
rect 26697 47135 26755 47141
rect 27890 47132 27896 47144
rect 27948 47132 27954 47184
rect 19981 47107 20039 47113
rect 19981 47073 19993 47107
rect 20027 47073 20039 47107
rect 19981 47067 20039 47073
rect 20070 47064 20076 47116
rect 20128 47104 20134 47116
rect 20254 47104 20260 47116
rect 20128 47076 20173 47104
rect 20215 47076 20260 47104
rect 20128 47064 20134 47076
rect 20254 47064 20260 47076
rect 20312 47064 20318 47116
rect 20349 47107 20407 47113
rect 20349 47073 20361 47107
rect 20395 47104 20407 47107
rect 20438 47104 20444 47116
rect 20395 47076 20444 47104
rect 20395 47073 20407 47076
rect 20349 47067 20407 47073
rect 20438 47064 20444 47076
rect 20496 47064 20502 47116
rect 20990 47104 20996 47116
rect 20951 47076 20996 47104
rect 20990 47064 20996 47076
rect 21048 47064 21054 47116
rect 21082 47064 21088 47116
rect 21140 47104 21146 47116
rect 21266 47104 21272 47116
rect 21140 47076 21185 47104
rect 21227 47076 21272 47104
rect 21140 47064 21146 47076
rect 21266 47064 21272 47076
rect 21324 47064 21330 47116
rect 22554 47064 22560 47116
rect 22612 47104 22618 47116
rect 22925 47107 22983 47113
rect 22925 47104 22937 47107
rect 22612 47076 22937 47104
rect 22612 47064 22618 47076
rect 22925 47073 22937 47076
rect 22971 47073 22983 47107
rect 22925 47067 22983 47073
rect 24213 47107 24271 47113
rect 24213 47073 24225 47107
rect 24259 47104 24271 47107
rect 24302 47104 24308 47116
rect 24259 47076 24308 47104
rect 24259 47073 24271 47076
rect 24213 47067 24271 47073
rect 24302 47064 24308 47076
rect 24360 47064 24366 47116
rect 26881 47107 26939 47113
rect 26881 47104 26893 47107
rect 24412 47076 26893 47104
rect 19245 47039 19303 47045
rect 19245 47005 19257 47039
rect 19291 47036 19303 47039
rect 20898 47036 20904 47048
rect 19291 47008 20904 47036
rect 19291 47005 19303 47008
rect 19245 46999 19303 47005
rect 20898 46996 20904 47008
rect 20956 46996 20962 47048
rect 21174 47036 21180 47048
rect 21135 47008 21180 47036
rect 21174 46996 21180 47008
rect 21232 46996 21238 47048
rect 24412 47036 24440 47076
rect 26881 47073 26893 47076
rect 26927 47073 26939 47107
rect 26881 47067 26939 47073
rect 21284 47008 24440 47036
rect 21284 46968 21312 47008
rect 25038 46996 25044 47048
rect 25096 47036 25102 47048
rect 25869 47039 25927 47045
rect 25869 47036 25881 47039
rect 25096 47008 25881 47036
rect 25096 46996 25102 47008
rect 25869 47005 25881 47008
rect 25915 47036 25927 47039
rect 25958 47036 25964 47048
rect 25915 47008 25964 47036
rect 25915 47005 25927 47008
rect 25869 46999 25927 47005
rect 25958 46996 25964 47008
rect 26016 46996 26022 47048
rect 26053 47039 26111 47045
rect 26053 47005 26065 47039
rect 26099 47036 26111 47039
rect 26142 47036 26148 47048
rect 26099 47008 26148 47036
rect 26099 47005 26111 47008
rect 26053 46999 26111 47005
rect 26142 46996 26148 47008
rect 26200 46996 26206 47048
rect 18248 46940 21312 46968
rect 21358 46928 21364 46980
rect 21416 46968 21422 46980
rect 28077 46971 28135 46977
rect 28077 46968 28089 46971
rect 21416 46940 28089 46968
rect 21416 46928 21422 46940
rect 28077 46937 28089 46940
rect 28123 46937 28135 46971
rect 28077 46931 28135 46937
rect 8202 46900 8208 46912
rect 4264 46872 8208 46900
rect 4157 46863 4215 46869
rect 8202 46860 8208 46872
rect 8260 46860 8266 46912
rect 8478 46860 8484 46912
rect 8536 46900 8542 46912
rect 8573 46903 8631 46909
rect 8573 46900 8585 46903
rect 8536 46872 8585 46900
rect 8536 46860 8542 46872
rect 8573 46869 8585 46872
rect 8619 46869 8631 46903
rect 13722 46900 13728 46912
rect 13683 46872 13728 46900
rect 8573 46863 8631 46869
rect 13722 46860 13728 46872
rect 13780 46860 13786 46912
rect 15746 46900 15752 46912
rect 15707 46872 15752 46900
rect 15746 46860 15752 46872
rect 15804 46860 15810 46912
rect 20254 46860 20260 46912
rect 20312 46900 20318 46912
rect 20622 46900 20628 46912
rect 20312 46872 20628 46900
rect 20312 46860 20318 46872
rect 20622 46860 20628 46872
rect 20680 46860 20686 46912
rect 23017 46903 23075 46909
rect 23017 46869 23029 46903
rect 23063 46900 23075 46903
rect 23382 46900 23388 46912
rect 23063 46872 23388 46900
rect 23063 46869 23075 46872
rect 23017 46863 23075 46869
rect 23382 46860 23388 46872
rect 23440 46860 23446 46912
rect 1104 46810 28888 46832
rect 1104 46758 5614 46810
rect 5666 46758 5678 46810
rect 5730 46758 5742 46810
rect 5794 46758 5806 46810
rect 5858 46758 14878 46810
rect 14930 46758 14942 46810
rect 14994 46758 15006 46810
rect 15058 46758 15070 46810
rect 15122 46758 24142 46810
rect 24194 46758 24206 46810
rect 24258 46758 24270 46810
rect 24322 46758 24334 46810
rect 24386 46758 28888 46810
rect 1104 46736 28888 46758
rect 6089 46699 6147 46705
rect 6089 46665 6101 46699
rect 6135 46696 6147 46699
rect 6546 46696 6552 46708
rect 6135 46668 6552 46696
rect 6135 46665 6147 46668
rect 6089 46659 6147 46665
rect 6546 46656 6552 46668
rect 6604 46656 6610 46708
rect 8481 46699 8539 46705
rect 8481 46665 8493 46699
rect 8527 46696 8539 46699
rect 9398 46696 9404 46708
rect 8527 46668 9404 46696
rect 8527 46665 8539 46668
rect 8481 46659 8539 46665
rect 9398 46656 9404 46668
rect 9456 46656 9462 46708
rect 9582 46696 9588 46708
rect 9543 46668 9588 46696
rect 9582 46656 9588 46668
rect 9640 46656 9646 46708
rect 27985 46699 28043 46705
rect 27985 46696 27997 46699
rect 12406 46668 27997 46696
rect 3326 46588 3332 46640
rect 3384 46628 3390 46640
rect 12406 46628 12434 46668
rect 27985 46665 27997 46668
rect 28031 46665 28043 46699
rect 27985 46659 28043 46665
rect 3384 46600 12434 46628
rect 13173 46631 13231 46637
rect 3384 46588 3390 46600
rect 13173 46597 13185 46631
rect 13219 46628 13231 46631
rect 13262 46628 13268 46640
rect 13219 46600 13268 46628
rect 13219 46597 13231 46600
rect 13173 46591 13231 46597
rect 13262 46588 13268 46600
rect 13320 46588 13326 46640
rect 14642 46588 14648 46640
rect 14700 46628 14706 46640
rect 14737 46631 14795 46637
rect 14737 46628 14749 46631
rect 14700 46600 14749 46628
rect 14700 46588 14706 46600
rect 14737 46597 14749 46600
rect 14783 46597 14795 46631
rect 16206 46628 16212 46640
rect 16167 46600 16212 46628
rect 14737 46591 14795 46597
rect 16206 46588 16212 46600
rect 16264 46588 16270 46640
rect 20809 46631 20867 46637
rect 20809 46597 20821 46631
rect 20855 46628 20867 46631
rect 20990 46628 20996 46640
rect 20855 46600 20996 46628
rect 20855 46597 20867 46600
rect 20809 46591 20867 46597
rect 20990 46588 20996 46600
rect 21048 46588 21054 46640
rect 22741 46631 22799 46637
rect 22741 46597 22753 46631
rect 22787 46628 22799 46631
rect 23198 46628 23204 46640
rect 22787 46600 23204 46628
rect 22787 46597 22799 46600
rect 22741 46591 22799 46597
rect 23198 46588 23204 46600
rect 23256 46628 23262 46640
rect 25777 46631 25835 46637
rect 23256 46600 24164 46628
rect 23256 46588 23262 46600
rect 2590 46520 2596 46572
rect 2648 46560 2654 46572
rect 2648 46532 7604 46560
rect 2648 46520 2654 46532
rect 1210 46452 1216 46504
rect 1268 46492 1274 46504
rect 1397 46495 1455 46501
rect 1397 46492 1409 46495
rect 1268 46464 1409 46492
rect 1268 46452 1274 46464
rect 1397 46461 1409 46464
rect 1443 46461 1455 46495
rect 1397 46455 1455 46461
rect 3970 46452 3976 46504
rect 4028 46492 4034 46504
rect 4249 46495 4307 46501
rect 4249 46492 4261 46495
rect 4028 46464 4261 46492
rect 4028 46452 4034 46464
rect 4249 46461 4261 46464
rect 4295 46461 4307 46495
rect 4430 46492 4436 46504
rect 4391 46464 4436 46492
rect 4249 46455 4307 46461
rect 4430 46452 4436 46464
rect 4488 46452 4494 46504
rect 4890 46492 4896 46504
rect 4851 46464 4896 46492
rect 4890 46452 4896 46464
rect 4948 46452 4954 46504
rect 5902 46452 5908 46504
rect 5960 46492 5966 46504
rect 5997 46495 6055 46501
rect 5997 46492 6009 46495
rect 5960 46464 6009 46492
rect 5960 46452 5966 46464
rect 5997 46461 6009 46464
rect 6043 46461 6055 46495
rect 5997 46455 6055 46461
rect 6181 46495 6239 46501
rect 6181 46461 6193 46495
rect 6227 46492 6239 46495
rect 6270 46492 6276 46504
rect 6227 46464 6276 46492
rect 6227 46461 6239 46464
rect 6181 46455 6239 46461
rect 6270 46452 6276 46464
rect 6328 46452 6334 46504
rect 1578 46384 1584 46436
rect 1636 46433 1642 46436
rect 1636 46427 1700 46433
rect 1636 46393 1654 46427
rect 1688 46393 1700 46427
rect 7576 46424 7604 46532
rect 8294 46520 8300 46572
rect 8352 46560 8358 46572
rect 10137 46563 10195 46569
rect 10137 46560 10149 46563
rect 8352 46532 10149 46560
rect 8352 46520 8358 46532
rect 10137 46529 10149 46532
rect 10183 46560 10195 46563
rect 10502 46560 10508 46572
rect 10183 46532 10508 46560
rect 10183 46529 10195 46532
rect 10137 46523 10195 46529
rect 10502 46520 10508 46532
rect 10560 46520 10566 46572
rect 10778 46520 10784 46572
rect 10836 46560 10842 46572
rect 11793 46563 11851 46569
rect 11793 46560 11805 46563
rect 10836 46532 11805 46560
rect 10836 46520 10842 46532
rect 11793 46529 11805 46532
rect 11839 46529 11851 46563
rect 11793 46523 11851 46529
rect 13633 46563 13691 46569
rect 13633 46529 13645 46563
rect 13679 46560 13691 46563
rect 13722 46560 13728 46572
rect 13679 46532 13728 46560
rect 13679 46529 13691 46532
rect 13633 46523 13691 46529
rect 13722 46520 13728 46532
rect 13780 46520 13786 46572
rect 14826 46520 14832 46572
rect 14884 46560 14890 46572
rect 15289 46563 15347 46569
rect 15289 46560 15301 46563
rect 14884 46532 15301 46560
rect 14884 46520 14890 46532
rect 15289 46529 15301 46532
rect 15335 46529 15347 46563
rect 15289 46523 15347 46529
rect 16853 46563 16911 46569
rect 16853 46529 16865 46563
rect 16899 46560 16911 46563
rect 18322 46560 18328 46572
rect 16899 46532 18328 46560
rect 16899 46529 16911 46532
rect 16853 46523 16911 46529
rect 18322 46520 18328 46532
rect 18380 46520 18386 46572
rect 23014 46520 23020 46572
rect 23072 46560 23078 46572
rect 23293 46563 23351 46569
rect 23293 46560 23305 46563
rect 23072 46532 23305 46560
rect 23072 46520 23078 46532
rect 23293 46529 23305 46532
rect 23339 46529 23351 46563
rect 23293 46523 23351 46529
rect 8389 46495 8447 46501
rect 8389 46461 8401 46495
rect 8435 46492 8447 46495
rect 8478 46492 8484 46504
rect 8435 46464 8484 46492
rect 8435 46461 8447 46464
rect 8389 46455 8447 46461
rect 8478 46452 8484 46464
rect 8536 46452 8542 46504
rect 8573 46495 8631 46501
rect 8573 46461 8585 46495
rect 8619 46492 8631 46495
rect 8662 46492 8668 46504
rect 8619 46464 8668 46492
rect 8619 46461 8631 46464
rect 8573 46455 8631 46461
rect 8662 46452 8668 46464
rect 8720 46452 8726 46504
rect 9953 46495 10011 46501
rect 9953 46461 9965 46495
rect 9999 46492 10011 46495
rect 11054 46492 11060 46504
rect 9999 46464 11060 46492
rect 9999 46461 10011 46464
rect 9953 46455 10011 46461
rect 11054 46452 11060 46464
rect 11112 46452 11118 46504
rect 13538 46452 13544 46504
rect 13596 46492 13602 46504
rect 16577 46495 16635 46501
rect 13596 46464 15884 46492
rect 13596 46452 13602 46464
rect 11790 46424 11796 46436
rect 7576 46396 11796 46424
rect 1636 46387 1700 46393
rect 1636 46384 1642 46387
rect 11790 46384 11796 46396
rect 11848 46384 11854 46436
rect 12526 46384 12532 46436
rect 12584 46424 12590 46436
rect 13725 46427 13783 46433
rect 13725 46424 13737 46427
rect 12584 46396 13737 46424
rect 12584 46384 12590 46396
rect 13725 46393 13737 46396
rect 13771 46393 13783 46427
rect 13725 46387 13783 46393
rect 15105 46427 15163 46433
rect 15105 46393 15117 46427
rect 15151 46424 15163 46427
rect 15746 46424 15752 46436
rect 15151 46396 15752 46424
rect 15151 46393 15163 46396
rect 15105 46387 15163 46393
rect 15746 46384 15752 46396
rect 15804 46384 15810 46436
rect 15856 46424 15884 46464
rect 16577 46461 16589 46495
rect 16623 46492 16635 46495
rect 17034 46492 17040 46504
rect 16623 46464 17040 46492
rect 16623 46461 16635 46464
rect 16577 46455 16635 46461
rect 17034 46452 17040 46464
rect 17092 46492 17098 46504
rect 17405 46495 17463 46501
rect 17405 46492 17417 46495
rect 17092 46464 17417 46492
rect 17092 46452 17098 46464
rect 17405 46461 17417 46464
rect 17451 46461 17463 46495
rect 17405 46455 17463 46461
rect 19886 46452 19892 46504
rect 19944 46492 19950 46504
rect 19981 46495 20039 46501
rect 19981 46492 19993 46495
rect 19944 46464 19993 46492
rect 19944 46452 19950 46464
rect 19981 46461 19993 46464
rect 20027 46461 20039 46495
rect 20162 46492 20168 46504
rect 20123 46464 20168 46492
rect 19981 46455 20039 46461
rect 20162 46452 20168 46464
rect 20220 46452 20226 46504
rect 20349 46495 20407 46501
rect 20349 46461 20361 46495
rect 20395 46492 20407 46495
rect 20809 46495 20867 46501
rect 20809 46492 20821 46495
rect 20395 46464 20821 46492
rect 20395 46461 20407 46464
rect 20349 46455 20407 46461
rect 20809 46461 20821 46464
rect 20855 46461 20867 46495
rect 20809 46455 20867 46461
rect 20898 46452 20904 46504
rect 20956 46492 20962 46504
rect 20993 46495 21051 46501
rect 20993 46492 21005 46495
rect 20956 46464 21005 46492
rect 20956 46452 20962 46464
rect 20993 46461 21005 46464
rect 21039 46461 21051 46495
rect 20993 46455 21051 46461
rect 23842 46452 23848 46504
rect 23900 46492 23906 46504
rect 24136 46501 24164 46600
rect 25777 46597 25789 46631
rect 25823 46628 25835 46631
rect 25823 46600 27936 46628
rect 25823 46597 25835 46600
rect 25777 46591 25835 46597
rect 27341 46563 27399 46569
rect 27341 46560 27353 46563
rect 24688 46532 27353 46560
rect 23937 46495 23995 46501
rect 23937 46492 23949 46495
rect 23900 46464 23949 46492
rect 23900 46452 23906 46464
rect 23937 46461 23949 46464
rect 23983 46461 23995 46495
rect 23937 46455 23995 46461
rect 24121 46495 24179 46501
rect 24121 46461 24133 46495
rect 24167 46461 24179 46495
rect 24121 46455 24179 46461
rect 24688 46424 24716 46532
rect 27341 46529 27353 46532
rect 27387 46529 27399 46563
rect 27341 46523 27399 46529
rect 25958 46492 25964 46504
rect 25919 46464 25964 46492
rect 25958 46452 25964 46464
rect 26016 46452 26022 46504
rect 26418 46492 26424 46504
rect 26379 46464 26424 46492
rect 26418 46452 26424 46464
rect 26476 46452 26482 46504
rect 27908 46501 27936 46600
rect 27893 46495 27951 46501
rect 27893 46461 27905 46495
rect 27939 46461 27951 46495
rect 27893 46455 27951 46461
rect 15856 46396 24716 46424
rect 26050 46384 26056 46436
rect 26108 46424 26114 46436
rect 27157 46427 27215 46433
rect 27157 46424 27169 46427
rect 26108 46396 27169 46424
rect 26108 46384 26114 46396
rect 27157 46393 27169 46396
rect 27203 46393 27215 46427
rect 27157 46387 27215 46393
rect 2777 46359 2835 46365
rect 2777 46325 2789 46359
rect 2823 46356 2835 46359
rect 3142 46356 3148 46368
rect 2823 46328 3148 46356
rect 2823 46325 2835 46328
rect 2777 46319 2835 46325
rect 3142 46316 3148 46328
rect 3200 46316 3206 46368
rect 4338 46356 4344 46368
rect 4299 46328 4344 46356
rect 4338 46316 4344 46328
rect 4396 46316 4402 46368
rect 4982 46356 4988 46368
rect 4943 46328 4988 46356
rect 4982 46316 4988 46328
rect 5040 46316 5046 46368
rect 6270 46316 6276 46368
rect 6328 46356 6334 46368
rect 8662 46356 8668 46368
rect 6328 46328 8668 46356
rect 6328 46316 6334 46328
rect 8662 46316 8668 46328
rect 8720 46316 8726 46368
rect 10042 46316 10048 46368
rect 10100 46356 10106 46368
rect 11241 46359 11299 46365
rect 10100 46328 10145 46356
rect 10100 46316 10106 46328
rect 11241 46325 11253 46359
rect 11287 46356 11299 46359
rect 11422 46356 11428 46368
rect 11287 46328 11428 46356
rect 11287 46325 11299 46328
rect 11241 46319 11299 46325
rect 11422 46316 11428 46328
rect 11480 46316 11486 46368
rect 11606 46356 11612 46368
rect 11567 46328 11612 46356
rect 11606 46316 11612 46328
rect 11664 46316 11670 46368
rect 11698 46316 11704 46368
rect 11756 46356 11762 46368
rect 13630 46356 13636 46368
rect 11756 46328 11801 46356
rect 13591 46328 13636 46356
rect 11756 46316 11762 46328
rect 13630 46316 13636 46328
rect 13688 46316 13694 46368
rect 14182 46316 14188 46368
rect 14240 46356 14246 46368
rect 15197 46359 15255 46365
rect 15197 46356 15209 46359
rect 14240 46328 15209 46356
rect 14240 46316 14246 46328
rect 15197 46325 15209 46328
rect 15243 46325 15255 46359
rect 15197 46319 15255 46325
rect 16669 46359 16727 46365
rect 16669 46325 16681 46359
rect 16715 46356 16727 46359
rect 17310 46356 17316 46368
rect 16715 46328 17316 46356
rect 16715 46325 16727 46328
rect 16669 46319 16727 46325
rect 17310 46316 17316 46328
rect 17368 46316 17374 46368
rect 17494 46356 17500 46368
rect 17455 46328 17500 46356
rect 17494 46316 17500 46328
rect 17552 46316 17558 46368
rect 23106 46356 23112 46368
rect 23067 46328 23112 46356
rect 23106 46316 23112 46328
rect 23164 46316 23170 46368
rect 23198 46316 23204 46368
rect 23256 46356 23262 46368
rect 24305 46359 24363 46365
rect 23256 46328 23301 46356
rect 23256 46316 23262 46328
rect 24305 46325 24317 46359
rect 24351 46356 24363 46359
rect 24486 46356 24492 46368
rect 24351 46328 24492 46356
rect 24351 46325 24363 46328
rect 24305 46319 24363 46325
rect 24486 46316 24492 46328
rect 24544 46316 24550 46368
rect 25866 46316 25872 46368
rect 25924 46356 25930 46368
rect 26513 46359 26571 46365
rect 26513 46356 26525 46359
rect 25924 46328 26525 46356
rect 25924 46316 25930 46328
rect 26513 46325 26525 46328
rect 26559 46325 26571 46359
rect 26513 46319 26571 46325
rect 1104 46266 28888 46288
rect 1104 46214 10246 46266
rect 10298 46214 10310 46266
rect 10362 46214 10374 46266
rect 10426 46214 10438 46266
rect 10490 46214 19510 46266
rect 19562 46214 19574 46266
rect 19626 46214 19638 46266
rect 19690 46214 19702 46266
rect 19754 46214 28888 46266
rect 1104 46192 28888 46214
rect 4614 46112 4620 46164
rect 4672 46152 4678 46164
rect 4893 46155 4951 46161
rect 4893 46152 4905 46155
rect 4672 46124 4905 46152
rect 4672 46112 4678 46124
rect 4893 46121 4905 46124
rect 4939 46121 4951 46155
rect 4893 46115 4951 46121
rect 4985 46155 5043 46161
rect 4985 46121 4997 46155
rect 5031 46152 5043 46155
rect 6086 46152 6092 46164
rect 5031 46124 6092 46152
rect 5031 46121 5043 46124
rect 4985 46115 5043 46121
rect 6086 46112 6092 46124
rect 6144 46112 6150 46164
rect 10042 46152 10048 46164
rect 10003 46124 10048 46152
rect 10042 46112 10048 46124
rect 10100 46112 10106 46164
rect 11149 46155 11207 46161
rect 11149 46121 11161 46155
rect 11195 46152 11207 46155
rect 11606 46152 11612 46164
rect 11195 46124 11612 46152
rect 11195 46121 11207 46124
rect 11149 46115 11207 46121
rect 11606 46112 11612 46124
rect 11664 46112 11670 46164
rect 11790 46112 11796 46164
rect 11848 46152 11854 46164
rect 23017 46155 23075 46161
rect 11848 46124 22094 46152
rect 11848 46112 11854 46124
rect 3421 46087 3479 46093
rect 3421 46053 3433 46087
rect 3467 46084 3479 46087
rect 4246 46084 4252 46096
rect 3467 46056 4252 46084
rect 3467 46053 3479 46056
rect 3421 46047 3479 46053
rect 4246 46044 4252 46056
rect 4304 46044 4310 46096
rect 8202 46044 8208 46096
rect 8260 46084 8266 46096
rect 13538 46084 13544 46096
rect 8260 46056 13544 46084
rect 8260 46044 8266 46056
rect 13538 46044 13544 46056
rect 13596 46044 13602 46096
rect 13722 46084 13728 46096
rect 13648 46056 13728 46084
rect 1762 45976 1768 46028
rect 1820 46016 1826 46028
rect 1857 46019 1915 46025
rect 1857 46016 1869 46019
rect 1820 45988 1869 46016
rect 1820 45976 1826 45988
rect 1857 45985 1869 45988
rect 1903 45985 1915 46019
rect 1857 45979 1915 45985
rect 3142 45976 3148 46028
rect 3200 46016 3206 46028
rect 3326 46016 3332 46028
rect 3200 45988 3332 46016
rect 3200 45976 3206 45988
rect 3326 45976 3332 45988
rect 3384 46016 3390 46028
rect 5721 46019 5779 46025
rect 5721 46016 5733 46019
rect 3384 45988 5733 46016
rect 3384 45976 3390 45988
rect 5721 45985 5733 45988
rect 5767 45985 5779 46019
rect 5721 45979 5779 45985
rect 9953 46019 10011 46025
rect 9953 45985 9965 46019
rect 9999 45985 10011 46019
rect 9953 45979 10011 45985
rect 3510 45948 3516 45960
rect 3471 45920 3516 45948
rect 3510 45908 3516 45920
rect 3568 45908 3574 45960
rect 3602 45908 3608 45960
rect 3660 45948 3666 45960
rect 3660 45920 3705 45948
rect 3660 45908 3666 45920
rect 4798 45908 4804 45960
rect 4856 45948 4862 45960
rect 5077 45951 5135 45957
rect 5077 45948 5089 45951
rect 4856 45920 5089 45948
rect 4856 45908 4862 45920
rect 5077 45917 5089 45920
rect 5123 45917 5135 45951
rect 5077 45911 5135 45917
rect 2041 45883 2099 45889
rect 2041 45849 2053 45883
rect 2087 45880 2099 45883
rect 2774 45880 2780 45892
rect 2087 45852 2780 45880
rect 2087 45849 2099 45852
rect 2041 45843 2099 45849
rect 2774 45840 2780 45852
rect 2832 45840 2838 45892
rect 4154 45840 4160 45892
rect 4212 45880 4218 45892
rect 5813 45883 5871 45889
rect 5813 45880 5825 45883
rect 4212 45852 5825 45880
rect 4212 45840 4218 45852
rect 5813 45849 5825 45852
rect 5859 45849 5871 45883
rect 9968 45880 9996 45979
rect 10594 45976 10600 46028
rect 10652 46016 10658 46028
rect 13648 46025 13676 46056
rect 13722 46044 13728 46056
rect 13780 46044 13786 46096
rect 19978 46084 19984 46096
rect 19939 46056 19984 46084
rect 19978 46044 19984 46056
rect 20036 46044 20042 46096
rect 22066 46084 22094 46124
rect 23017 46121 23029 46155
rect 23063 46152 23075 46155
rect 23198 46152 23204 46164
rect 23063 46124 23204 46152
rect 23063 46121 23075 46124
rect 23017 46115 23075 46121
rect 23198 46112 23204 46124
rect 23256 46112 23262 46164
rect 23382 46152 23388 46164
rect 23343 46124 23388 46152
rect 23382 46112 23388 46124
rect 23440 46112 23446 46164
rect 24578 46152 24584 46164
rect 24320 46124 24584 46152
rect 24320 46093 24348 46124
rect 24578 46112 24584 46124
rect 24636 46112 24642 46164
rect 25409 46155 25467 46161
rect 25409 46121 25421 46155
rect 25455 46121 25467 46155
rect 25409 46115 25467 46121
rect 24305 46087 24363 46093
rect 22066 46056 23888 46084
rect 10781 46019 10839 46025
rect 10781 46016 10793 46019
rect 10652 45988 10793 46016
rect 10652 45976 10658 45988
rect 10781 45985 10793 45988
rect 10827 45985 10839 46019
rect 10781 45979 10839 45985
rect 12253 46019 12311 46025
rect 12253 45985 12265 46019
rect 12299 46016 12311 46019
rect 13081 46019 13139 46025
rect 13081 46016 13093 46019
rect 12299 45988 13093 46016
rect 12299 45985 12311 45988
rect 12253 45979 12311 45985
rect 13081 45985 13093 45988
rect 13127 45985 13139 46019
rect 13081 45979 13139 45985
rect 13633 46019 13691 46025
rect 13633 45985 13645 46019
rect 13679 45985 13691 46019
rect 13633 45979 13691 45985
rect 10870 45948 10876 45960
rect 10831 45920 10876 45948
rect 10870 45908 10876 45920
rect 10928 45908 10934 45960
rect 11698 45880 11704 45892
rect 9968 45852 11704 45880
rect 5813 45843 5871 45849
rect 11698 45840 11704 45852
rect 11756 45840 11762 45892
rect 12989 45883 13047 45889
rect 12989 45849 13001 45883
rect 13035 45849 13047 45883
rect 13096 45880 13124 45979
rect 14182 45976 14188 46028
rect 14240 46016 14246 46028
rect 14461 46019 14519 46025
rect 14461 46016 14473 46019
rect 14240 45988 14473 46016
rect 14240 45976 14246 45988
rect 14461 45985 14473 45988
rect 14507 45985 14519 46019
rect 14461 45979 14519 45985
rect 14921 46019 14979 46025
rect 14921 45985 14933 46019
rect 14967 46016 14979 46019
rect 15657 46019 15715 46025
rect 14967 45988 15148 46016
rect 14967 45985 14979 45988
rect 14921 45979 14979 45985
rect 13538 45908 13544 45960
rect 13596 45948 13602 45960
rect 13725 45951 13783 45957
rect 13725 45948 13737 45951
rect 13596 45920 13737 45948
rect 13596 45908 13602 45920
rect 13725 45917 13737 45920
rect 13771 45917 13783 45951
rect 13725 45911 13783 45917
rect 15013 45951 15071 45957
rect 15013 45917 15025 45951
rect 15059 45917 15071 45951
rect 15013 45911 15071 45917
rect 15028 45880 15056 45911
rect 13096 45852 15056 45880
rect 12989 45843 13047 45849
rect 3053 45815 3111 45821
rect 3053 45781 3065 45815
rect 3099 45812 3111 45815
rect 3142 45812 3148 45824
rect 3099 45784 3148 45812
rect 3099 45781 3111 45784
rect 3053 45775 3111 45781
rect 3142 45772 3148 45784
rect 3200 45772 3206 45824
rect 4522 45812 4528 45824
rect 4483 45784 4528 45812
rect 4522 45772 4528 45784
rect 4580 45772 4586 45824
rect 12342 45812 12348 45824
rect 12303 45784 12348 45812
rect 12342 45772 12348 45784
rect 12400 45772 12406 45824
rect 13004 45812 13032 45843
rect 13170 45812 13176 45824
rect 13004 45784 13176 45812
rect 13170 45772 13176 45784
rect 13228 45772 13234 45824
rect 13262 45772 13268 45824
rect 13320 45812 13326 45824
rect 15120 45812 15148 45988
rect 15657 45985 15669 46019
rect 15703 46016 15715 46019
rect 15746 46016 15752 46028
rect 15703 45988 15752 46016
rect 15703 45985 15715 45988
rect 15657 45979 15715 45985
rect 15746 45976 15752 45988
rect 15804 45976 15810 46028
rect 17126 45976 17132 46028
rect 17184 46016 17190 46028
rect 17313 46019 17371 46025
rect 17313 46016 17325 46019
rect 17184 45988 17325 46016
rect 17184 45976 17190 45988
rect 17313 45985 17325 45988
rect 17359 45985 17371 46019
rect 17313 45979 17371 45985
rect 17402 45976 17408 46028
rect 17460 46016 17466 46028
rect 17497 46019 17555 46025
rect 17497 46016 17509 46019
rect 17460 45988 17509 46016
rect 17460 45976 17466 45988
rect 17497 45985 17509 45988
rect 17543 45985 17555 46019
rect 17497 45979 17555 45985
rect 17681 46019 17739 46025
rect 17681 45985 17693 46019
rect 17727 46016 17739 46019
rect 18138 46016 18144 46028
rect 17727 45988 18144 46016
rect 17727 45985 17739 45988
rect 17681 45979 17739 45985
rect 18138 45976 18144 45988
rect 18196 45976 18202 46028
rect 19797 46019 19855 46025
rect 19797 45985 19809 46019
rect 19843 46016 19855 46019
rect 19886 46016 19892 46028
rect 19843 45988 19892 46016
rect 19843 45985 19855 45988
rect 19797 45979 19855 45985
rect 19886 45976 19892 45988
rect 19944 45976 19950 46028
rect 23474 45948 23480 45960
rect 23435 45920 23480 45948
rect 23474 45908 23480 45920
rect 23532 45908 23538 45960
rect 23569 45951 23627 45957
rect 23569 45917 23581 45951
rect 23615 45917 23627 45951
rect 23860 45948 23888 46056
rect 24305 46053 24317 46087
rect 24351 46053 24363 46087
rect 25424 46084 25452 46115
rect 27893 46087 27951 46093
rect 27893 46084 27905 46087
rect 25424 46056 27905 46084
rect 24305 46047 24363 46053
rect 27893 46053 27905 46056
rect 27939 46053 27951 46087
rect 27893 46047 27951 46053
rect 24026 45976 24032 46028
rect 24084 46016 24090 46028
rect 24213 46019 24271 46025
rect 24213 46016 24225 46019
rect 24084 45988 24225 46016
rect 24084 45976 24090 45988
rect 24213 45985 24225 45988
rect 24259 45985 24271 46019
rect 24578 46016 24584 46028
rect 24539 45988 24584 46016
rect 24213 45979 24271 45985
rect 24578 45976 24584 45988
rect 24636 45976 24642 46028
rect 24765 46019 24823 46025
rect 24765 45985 24777 46019
rect 24811 46016 24823 46019
rect 24854 46016 24860 46028
rect 24811 45988 24860 46016
rect 24811 45985 24823 45988
rect 24765 45979 24823 45985
rect 24854 45976 24860 45988
rect 24912 45976 24918 46028
rect 25590 46016 25596 46028
rect 25551 45988 25596 46016
rect 25590 45976 25596 45988
rect 25648 45976 25654 46028
rect 26234 46016 26240 46028
rect 26195 45988 26240 46016
rect 26234 45976 26240 45988
rect 26292 45976 26298 46028
rect 26881 46019 26939 46025
rect 26881 45985 26893 46019
rect 26927 46016 26939 46019
rect 26970 46016 26976 46028
rect 26927 45988 26976 46016
rect 26927 45985 26939 45988
rect 26881 45979 26939 45985
rect 26970 45976 26976 45988
rect 27028 45976 27034 46028
rect 28077 45951 28135 45957
rect 28077 45948 28089 45951
rect 23860 45920 28089 45948
rect 23569 45911 23627 45917
rect 28077 45917 28089 45920
rect 28123 45917 28135 45951
rect 28077 45911 28135 45917
rect 22186 45840 22192 45892
rect 22244 45880 22250 45892
rect 23584 45880 23612 45911
rect 22244 45852 23612 45880
rect 26053 45883 26111 45889
rect 22244 45840 22250 45852
rect 26053 45849 26065 45883
rect 26099 45880 26111 45883
rect 27614 45880 27620 45892
rect 26099 45852 27620 45880
rect 26099 45849 26111 45852
rect 26053 45843 26111 45849
rect 27614 45840 27620 45852
rect 27672 45840 27678 45892
rect 15746 45812 15752 45824
rect 13320 45784 15148 45812
rect 15707 45784 15752 45812
rect 13320 45772 13326 45784
rect 15746 45772 15752 45784
rect 15804 45772 15810 45824
rect 18230 45812 18236 45824
rect 18191 45784 18236 45812
rect 18230 45772 18236 45784
rect 18288 45772 18294 45824
rect 26697 45815 26755 45821
rect 26697 45781 26709 45815
rect 26743 45812 26755 45815
rect 27890 45812 27896 45824
rect 26743 45784 27896 45812
rect 26743 45781 26755 45784
rect 26697 45775 26755 45781
rect 27890 45772 27896 45784
rect 27948 45772 27954 45824
rect 1104 45722 28888 45744
rect 1104 45670 5614 45722
rect 5666 45670 5678 45722
rect 5730 45670 5742 45722
rect 5794 45670 5806 45722
rect 5858 45670 14878 45722
rect 14930 45670 14942 45722
rect 14994 45670 15006 45722
rect 15058 45670 15070 45722
rect 15122 45670 24142 45722
rect 24194 45670 24206 45722
rect 24258 45670 24270 45722
rect 24322 45670 24334 45722
rect 24386 45670 28888 45722
rect 1104 45648 28888 45670
rect 1578 45608 1584 45620
rect 1539 45580 1584 45608
rect 1578 45568 1584 45580
rect 1636 45568 1642 45620
rect 3326 45608 3332 45620
rect 2792 45580 3332 45608
rect 2498 45540 2504 45552
rect 2148 45512 2504 45540
rect 2148 45484 2176 45512
rect 2498 45500 2504 45512
rect 2556 45500 2562 45552
rect 2130 45432 2136 45484
rect 2188 45432 2194 45484
rect 2225 45475 2283 45481
rect 2225 45441 2237 45475
rect 2271 45472 2283 45475
rect 2314 45472 2320 45484
rect 2271 45444 2320 45472
rect 2271 45441 2283 45444
rect 2225 45435 2283 45441
rect 2314 45432 2320 45444
rect 2372 45432 2378 45484
rect 1949 45407 2007 45413
rect 1949 45373 1961 45407
rect 1995 45404 2007 45407
rect 2792 45404 2820 45580
rect 3326 45568 3332 45580
rect 3384 45568 3390 45620
rect 7558 45568 7564 45620
rect 7616 45608 7622 45620
rect 8113 45611 8171 45617
rect 8113 45608 8125 45611
rect 7616 45580 8125 45608
rect 7616 45568 7622 45580
rect 8113 45577 8125 45580
rect 8159 45577 8171 45611
rect 8113 45571 8171 45577
rect 13630 45568 13636 45620
rect 13688 45608 13694 45620
rect 13688 45580 13768 45608
rect 13688 45568 13694 45580
rect 1995 45376 2820 45404
rect 3068 45512 3464 45540
rect 1995 45373 2007 45376
rect 1949 45367 2007 45373
rect 2041 45339 2099 45345
rect 2041 45305 2053 45339
rect 2087 45336 2099 45339
rect 3068 45336 3096 45512
rect 3436 45472 3464 45512
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 4249 45543 4307 45549
rect 4249 45540 4261 45543
rect 3568 45512 4261 45540
rect 3568 45500 3574 45512
rect 4249 45509 4261 45512
rect 4295 45509 4307 45543
rect 4249 45503 4307 45509
rect 4614 45500 4620 45552
rect 4672 45500 4678 45552
rect 9677 45543 9735 45549
rect 9677 45509 9689 45543
rect 9723 45540 9735 45543
rect 10778 45540 10784 45552
rect 9723 45512 10784 45540
rect 9723 45509 9735 45512
rect 9677 45503 9735 45509
rect 10778 45500 10784 45512
rect 10836 45500 10842 45552
rect 12342 45500 12348 45552
rect 12400 45540 12406 45552
rect 13740 45540 13768 45580
rect 21450 45568 21456 45620
rect 21508 45608 21514 45620
rect 23017 45611 23075 45617
rect 23017 45608 23029 45611
rect 21508 45580 23029 45608
rect 21508 45568 21514 45580
rect 23017 45577 23029 45580
rect 23063 45577 23075 45611
rect 23017 45571 23075 45577
rect 14829 45543 14887 45549
rect 14829 45540 14841 45543
rect 12400 45512 13676 45540
rect 13740 45512 14841 45540
rect 12400 45500 12406 45512
rect 4632 45472 4660 45500
rect 4798 45472 4804 45484
rect 3436 45444 4660 45472
rect 4759 45444 4804 45472
rect 4798 45432 4804 45444
rect 4856 45432 4862 45484
rect 6457 45475 6515 45481
rect 6457 45441 6469 45475
rect 6503 45472 6515 45475
rect 6914 45472 6920 45484
rect 6503 45444 6920 45472
rect 6503 45441 6515 45444
rect 6457 45435 6515 45441
rect 6914 45432 6920 45444
rect 6972 45472 6978 45484
rect 7466 45472 7472 45484
rect 6972 45444 7472 45472
rect 6972 45432 6978 45444
rect 7466 45432 7472 45444
rect 7524 45432 7530 45484
rect 11146 45472 11152 45484
rect 11107 45444 11152 45472
rect 11146 45432 11152 45444
rect 11204 45432 11210 45484
rect 11422 45472 11428 45484
rect 11383 45444 11428 45472
rect 11422 45432 11428 45444
rect 11480 45432 11486 45484
rect 3145 45407 3203 45413
rect 3145 45373 3157 45407
rect 3191 45404 3203 45407
rect 3234 45404 3240 45416
rect 3191 45376 3240 45404
rect 3191 45373 3203 45376
rect 3145 45367 3203 45373
rect 3234 45364 3240 45376
rect 3292 45364 3298 45416
rect 4617 45407 4675 45413
rect 4617 45373 4629 45407
rect 4663 45404 4675 45407
rect 4982 45404 4988 45416
rect 4663 45376 4988 45404
rect 4663 45373 4675 45376
rect 4617 45367 4675 45373
rect 4982 45364 4988 45376
rect 5040 45364 5046 45416
rect 9306 45364 9312 45416
rect 9364 45404 9370 45416
rect 9493 45407 9551 45413
rect 9493 45404 9505 45407
rect 9364 45376 9505 45404
rect 9364 45364 9370 45376
rect 9493 45373 9505 45376
rect 9539 45373 9551 45407
rect 9493 45367 9551 45373
rect 13449 45407 13507 45413
rect 13449 45373 13461 45407
rect 13495 45404 13507 45407
rect 13538 45404 13544 45416
rect 13495 45376 13544 45404
rect 13495 45373 13507 45376
rect 13449 45367 13507 45373
rect 13538 45364 13544 45376
rect 13596 45364 13602 45416
rect 13648 45413 13676 45512
rect 14829 45509 14841 45512
rect 14875 45509 14887 45543
rect 14829 45503 14887 45509
rect 16301 45543 16359 45549
rect 16301 45509 16313 45543
rect 16347 45540 16359 45543
rect 17126 45540 17132 45552
rect 16347 45512 17132 45540
rect 16347 45509 16359 45512
rect 16301 45503 16359 45509
rect 17126 45500 17132 45512
rect 17184 45500 17190 45552
rect 17865 45543 17923 45549
rect 17865 45509 17877 45543
rect 17911 45540 17923 45543
rect 18046 45540 18052 45552
rect 17911 45512 18052 45540
rect 17911 45509 17923 45512
rect 17865 45503 17923 45509
rect 18046 45500 18052 45512
rect 18104 45500 18110 45552
rect 22554 45540 22560 45552
rect 22515 45512 22560 45540
rect 22554 45500 22560 45512
rect 22612 45500 22618 45552
rect 24578 45500 24584 45552
rect 24636 45540 24642 45552
rect 25317 45543 25375 45549
rect 25317 45540 25329 45543
rect 24636 45512 25329 45540
rect 24636 45500 24642 45512
rect 25317 45509 25329 45512
rect 25363 45509 25375 45543
rect 25317 45503 25375 45509
rect 25682 45500 25688 45552
rect 25740 45540 25746 45552
rect 25740 45512 26096 45540
rect 25740 45500 25746 45512
rect 14274 45432 14280 45484
rect 14332 45472 14338 45484
rect 15381 45475 15439 45481
rect 15381 45472 15393 45475
rect 14332 45444 15393 45472
rect 14332 45432 14338 45444
rect 15381 45441 15393 45444
rect 15427 45441 15439 45475
rect 23569 45475 23627 45481
rect 15381 45435 15439 45441
rect 16868 45444 21312 45472
rect 13633 45407 13691 45413
rect 13633 45373 13645 45407
rect 13679 45373 13691 45407
rect 13633 45367 13691 45373
rect 13722 45364 13728 45416
rect 13780 45404 13786 45416
rect 15197 45407 15255 45413
rect 13780 45376 13825 45404
rect 13780 45364 13786 45376
rect 15197 45373 15209 45407
rect 15243 45404 15255 45407
rect 15746 45404 15752 45416
rect 15243 45376 15752 45404
rect 15243 45373 15255 45376
rect 15197 45367 15255 45373
rect 15746 45364 15752 45376
rect 15804 45364 15810 45416
rect 16022 45364 16028 45416
rect 16080 45404 16086 45416
rect 16868 45413 16896 45444
rect 16853 45407 16911 45413
rect 16853 45404 16865 45407
rect 16080 45376 16865 45404
rect 16080 45364 16086 45376
rect 16853 45373 16865 45376
rect 16899 45373 16911 45407
rect 16853 45367 16911 45373
rect 17773 45407 17831 45413
rect 17773 45373 17785 45407
rect 17819 45373 17831 45407
rect 18138 45404 18144 45416
rect 18099 45376 18144 45404
rect 17773 45367 17831 45373
rect 3602 45336 3608 45348
rect 2087 45308 3096 45336
rect 3160 45308 3608 45336
rect 2087 45305 2099 45308
rect 2041 45299 2099 45305
rect 2222 45228 2228 45280
rect 2280 45268 2286 45280
rect 3160 45268 3188 45308
rect 3602 45296 3608 45308
rect 3660 45296 3666 45348
rect 7650 45296 7656 45348
rect 7708 45336 7714 45348
rect 7929 45339 7987 45345
rect 7929 45336 7941 45339
rect 7708 45308 7941 45336
rect 7708 45296 7714 45308
rect 7929 45305 7941 45308
rect 7975 45336 7987 45339
rect 8018 45336 8024 45348
rect 7975 45308 8024 45336
rect 7975 45305 7987 45308
rect 7929 45299 7987 45305
rect 8018 45296 8024 45308
rect 8076 45296 8082 45348
rect 13265 45339 13323 45345
rect 13265 45305 13277 45339
rect 13311 45336 13323 45339
rect 14090 45336 14096 45348
rect 13311 45308 14096 45336
rect 13311 45305 13323 45308
rect 13265 45299 13323 45305
rect 14090 45296 14096 45308
rect 14148 45296 14154 45348
rect 16114 45296 16120 45348
rect 16172 45336 16178 45348
rect 16577 45339 16635 45345
rect 16577 45336 16589 45339
rect 16172 45308 16589 45336
rect 16172 45296 16178 45308
rect 16577 45305 16589 45308
rect 16623 45305 16635 45339
rect 17788 45336 17816 45367
rect 18138 45364 18144 45376
rect 18196 45364 18202 45416
rect 18414 45404 18420 45416
rect 18375 45376 18420 45404
rect 18414 45364 18420 45376
rect 18472 45364 18478 45416
rect 21174 45404 21180 45416
rect 21135 45376 21180 45404
rect 21174 45364 21180 45376
rect 21232 45364 21238 45416
rect 21284 45404 21312 45444
rect 23569 45441 23581 45475
rect 23615 45441 23627 45475
rect 23569 45435 23627 45441
rect 21284 45376 21588 45404
rect 21450 45345 21456 45348
rect 21444 45336 21456 45345
rect 17788 45308 18184 45336
rect 21411 45308 21456 45336
rect 16577 45299 16635 45305
rect 18156 45280 18184 45308
rect 21444 45299 21456 45308
rect 21450 45296 21456 45299
rect 21508 45296 21514 45348
rect 21560 45336 21588 45376
rect 22554 45364 22560 45416
rect 22612 45404 22618 45416
rect 23385 45407 23443 45413
rect 23385 45404 23397 45407
rect 22612 45376 23397 45404
rect 22612 45364 22618 45376
rect 23385 45373 23397 45376
rect 23431 45373 23443 45407
rect 23385 45367 23443 45373
rect 23014 45336 23020 45348
rect 21560 45308 23020 45336
rect 23014 45296 23020 45308
rect 23072 45296 23078 45348
rect 23584 45336 23612 45435
rect 24486 45432 24492 45484
rect 24544 45472 24550 45484
rect 24544 45444 25912 45472
rect 24544 45432 24550 45444
rect 24118 45364 24124 45416
rect 24176 45404 24182 45416
rect 25225 45407 25283 45413
rect 25225 45404 25237 45407
rect 24176 45376 25237 45404
rect 24176 45364 24182 45376
rect 25225 45373 25237 45376
rect 25271 45404 25283 45407
rect 25590 45404 25596 45416
rect 25271 45376 25596 45404
rect 25271 45373 25283 45376
rect 25225 45367 25283 45373
rect 25590 45364 25596 45376
rect 25648 45364 25654 45416
rect 25884 45413 25912 45444
rect 26068 45413 26096 45512
rect 25869 45407 25927 45413
rect 25869 45373 25881 45407
rect 25915 45373 25927 45407
rect 25869 45367 25927 45373
rect 26053 45407 26111 45413
rect 26053 45373 26065 45407
rect 26099 45373 26111 45407
rect 27062 45404 27068 45416
rect 27023 45376 27068 45404
rect 26053 45367 26111 45373
rect 27062 45364 27068 45376
rect 27120 45364 27126 45416
rect 27614 45404 27620 45416
rect 27575 45376 27620 45404
rect 27614 45364 27620 45376
rect 27672 45364 27678 45416
rect 23308 45308 23612 45336
rect 2280 45240 3188 45268
rect 3237 45271 3295 45277
rect 2280 45228 2286 45240
rect 3237 45237 3249 45271
rect 3283 45268 3295 45271
rect 3326 45268 3332 45280
rect 3283 45240 3332 45268
rect 3283 45237 3295 45240
rect 3237 45231 3295 45237
rect 3326 45228 3332 45240
rect 3384 45268 3390 45280
rect 3970 45268 3976 45280
rect 3384 45240 3976 45268
rect 3384 45228 3390 45240
rect 3970 45228 3976 45240
rect 4028 45228 4034 45280
rect 4706 45228 4712 45280
rect 4764 45268 4770 45280
rect 5813 45271 5871 45277
rect 4764 45240 4809 45268
rect 4764 45228 4770 45240
rect 5813 45237 5825 45271
rect 5859 45268 5871 45271
rect 5994 45268 6000 45280
rect 5859 45240 6000 45268
rect 5859 45237 5871 45240
rect 5813 45231 5871 45237
rect 5994 45228 6000 45240
rect 6052 45228 6058 45280
rect 6178 45268 6184 45280
rect 6139 45240 6184 45268
rect 6178 45228 6184 45240
rect 6236 45228 6242 45280
rect 6273 45271 6331 45277
rect 6273 45237 6285 45271
rect 6319 45268 6331 45271
rect 6454 45268 6460 45280
rect 6319 45240 6460 45268
rect 6319 45237 6331 45240
rect 6273 45231 6331 45237
rect 6454 45228 6460 45240
rect 6512 45228 6518 45280
rect 7742 45228 7748 45280
rect 7800 45268 7806 45280
rect 8134 45271 8192 45277
rect 8134 45268 8146 45271
rect 7800 45240 8146 45268
rect 7800 45228 7806 45240
rect 8134 45237 8146 45240
rect 8180 45237 8192 45271
rect 8134 45231 8192 45237
rect 8297 45271 8355 45277
rect 8297 45237 8309 45271
rect 8343 45268 8355 45271
rect 9490 45268 9496 45280
rect 8343 45240 9496 45268
rect 8343 45237 8355 45240
rect 8297 45231 8355 45237
rect 9490 45228 9496 45240
rect 9548 45228 9554 45280
rect 11790 45228 11796 45280
rect 11848 45268 11854 45280
rect 12529 45271 12587 45277
rect 12529 45268 12541 45271
rect 11848 45240 12541 45268
rect 11848 45228 11854 45240
rect 12529 45237 12541 45240
rect 12575 45237 12587 45271
rect 12529 45231 12587 45237
rect 12618 45228 12624 45280
rect 12676 45268 12682 45280
rect 14274 45268 14280 45280
rect 12676 45240 14280 45268
rect 12676 45228 12682 45240
rect 14274 45228 14280 45240
rect 14332 45228 14338 45280
rect 15289 45271 15347 45277
rect 15289 45237 15301 45271
rect 15335 45268 15347 45271
rect 15562 45268 15568 45280
rect 15335 45240 15568 45268
rect 15335 45237 15347 45240
rect 15289 45231 15347 45237
rect 15562 45228 15568 45240
rect 15620 45228 15626 45280
rect 15654 45228 15660 45280
rect 15712 45268 15718 45280
rect 16761 45271 16819 45277
rect 16761 45268 16773 45271
rect 15712 45240 16773 45268
rect 15712 45228 15718 45240
rect 16761 45237 16773 45240
rect 16807 45237 16819 45271
rect 16761 45231 16819 45237
rect 18138 45228 18144 45280
rect 18196 45228 18202 45280
rect 21542 45228 21548 45280
rect 21600 45268 21606 45280
rect 23308 45268 23336 45308
rect 23934 45296 23940 45348
rect 23992 45336 23998 45348
rect 27801 45339 27859 45345
rect 27801 45336 27813 45339
rect 23992 45308 27813 45336
rect 23992 45296 23998 45308
rect 27801 45305 27813 45308
rect 27847 45305 27859 45339
rect 27801 45299 27859 45305
rect 21600 45240 23336 45268
rect 21600 45228 21606 45240
rect 23382 45228 23388 45280
rect 23440 45268 23446 45280
rect 23477 45271 23535 45277
rect 23477 45268 23489 45271
rect 23440 45240 23489 45268
rect 23440 45228 23446 45240
rect 23477 45237 23489 45240
rect 23523 45268 23535 45271
rect 23842 45268 23848 45280
rect 23523 45240 23848 45268
rect 23523 45237 23535 45240
rect 23477 45231 23535 45237
rect 23842 45228 23848 45240
rect 23900 45228 23906 45280
rect 24302 45228 24308 45280
rect 24360 45268 24366 45280
rect 25961 45271 26019 45277
rect 25961 45268 25973 45271
rect 24360 45240 25973 45268
rect 24360 45228 24366 45240
rect 25961 45237 25973 45240
rect 26007 45237 26019 45271
rect 26878 45268 26884 45280
rect 26839 45240 26884 45268
rect 25961 45231 26019 45237
rect 26878 45228 26884 45240
rect 26936 45228 26942 45280
rect 1104 45178 28888 45200
rect 1104 45126 10246 45178
rect 10298 45126 10310 45178
rect 10362 45126 10374 45178
rect 10426 45126 10438 45178
rect 10490 45126 19510 45178
rect 19562 45126 19574 45178
rect 19626 45126 19638 45178
rect 19690 45126 19702 45178
rect 19754 45126 28888 45178
rect 1104 45104 28888 45126
rect 2869 45067 2927 45073
rect 2869 45033 2881 45067
rect 2915 45064 2927 45067
rect 4154 45064 4160 45076
rect 2915 45036 4160 45064
rect 2915 45033 2927 45036
rect 2869 45027 2927 45033
rect 4154 45024 4160 45036
rect 4212 45024 4218 45076
rect 4338 45064 4344 45076
rect 4299 45036 4344 45064
rect 4338 45024 4344 45036
rect 4396 45024 4402 45076
rect 4433 45067 4491 45073
rect 4433 45033 4445 45067
rect 4479 45064 4491 45067
rect 4522 45064 4528 45076
rect 4479 45036 4528 45064
rect 4479 45033 4491 45036
rect 4433 45027 4491 45033
rect 4522 45024 4528 45036
rect 4580 45024 4586 45076
rect 22833 45067 22891 45073
rect 12406 45036 22094 45064
rect 2130 44956 2136 45008
rect 2188 44996 2194 45008
rect 12406 44996 12434 45036
rect 2188 44968 12434 44996
rect 16025 44999 16083 45005
rect 2188 44956 2194 44968
rect 16025 44965 16037 44999
rect 16071 44996 16083 44999
rect 17494 44996 17500 45008
rect 16071 44968 17500 44996
rect 16071 44965 16083 44968
rect 16025 44959 16083 44965
rect 17494 44956 17500 44968
rect 17552 44956 17558 45008
rect 18322 44956 18328 45008
rect 18380 44996 18386 45008
rect 18380 44968 19012 44996
rect 18380 44956 18386 44968
rect 18984 44940 19012 44968
rect 19058 44956 19064 45008
rect 19116 44996 19122 45008
rect 19858 44999 19916 45005
rect 19858 44996 19870 44999
rect 19116 44968 19870 44996
rect 19116 44956 19122 44968
rect 19858 44965 19870 44968
rect 19904 44965 19916 44999
rect 19858 44959 19916 44965
rect 20070 44956 20076 45008
rect 20128 44956 20134 45008
rect 22066 44996 22094 45036
rect 22833 45033 22845 45067
rect 22879 45064 22891 45067
rect 23106 45064 23112 45076
rect 22879 45036 23112 45064
rect 22879 45033 22891 45036
rect 22833 45027 22891 45033
rect 23106 45024 23112 45036
rect 23164 45024 23170 45076
rect 23385 45067 23443 45073
rect 23385 45033 23397 45067
rect 23431 45064 23443 45067
rect 24118 45064 24124 45076
rect 23431 45036 24124 45064
rect 23431 45033 23443 45036
rect 23385 45027 23443 45033
rect 24118 45024 24124 45036
rect 24176 45024 24182 45076
rect 24397 45067 24455 45073
rect 24397 45033 24409 45067
rect 24443 45033 24455 45067
rect 24397 45027 24455 45033
rect 23934 44996 23940 45008
rect 22066 44968 23940 44996
rect 23934 44956 23940 44968
rect 23992 44956 23998 45008
rect 24026 44956 24032 45008
rect 24084 44996 24090 45008
rect 24302 45005 24308 45008
rect 24245 44999 24308 45005
rect 24084 44968 24129 44996
rect 24084 44956 24090 44968
rect 24245 44965 24257 44999
rect 24291 44965 24308 44999
rect 24245 44959 24308 44965
rect 24302 44956 24308 44959
rect 24360 44956 24366 45008
rect 1857 44931 1915 44937
rect 1857 44897 1869 44931
rect 1903 44928 1915 44931
rect 2590 44928 2596 44940
rect 1903 44900 2596 44928
rect 1903 44897 1915 44900
rect 1857 44891 1915 44897
rect 2590 44888 2596 44900
rect 2648 44888 2654 44940
rect 2961 44931 3019 44937
rect 2961 44897 2973 44931
rect 3007 44928 3019 44931
rect 5074 44928 5080 44940
rect 3007 44900 5080 44928
rect 3007 44897 3019 44900
rect 2961 44891 3019 44897
rect 5074 44888 5080 44900
rect 5132 44888 5138 44940
rect 5718 44928 5724 44940
rect 5679 44900 5724 44928
rect 5718 44888 5724 44900
rect 5776 44888 5782 44940
rect 5994 44888 6000 44940
rect 6052 44928 6058 44940
rect 6822 44928 6828 44940
rect 6052 44900 6828 44928
rect 6052 44888 6058 44900
rect 6822 44888 6828 44900
rect 6880 44888 6886 44940
rect 7009 44931 7067 44937
rect 7009 44897 7021 44931
rect 7055 44897 7067 44931
rect 7558 44928 7564 44940
rect 7519 44900 7564 44928
rect 7009 44891 7067 44897
rect 3145 44863 3203 44869
rect 3145 44829 3157 44863
rect 3191 44860 3203 44863
rect 3234 44860 3240 44872
rect 3191 44832 3240 44860
rect 3191 44829 3203 44832
rect 3145 44823 3203 44829
rect 3234 44820 3240 44832
rect 3292 44860 3298 44872
rect 3510 44860 3516 44872
rect 3292 44832 3516 44860
rect 3292 44820 3298 44832
rect 3510 44820 3516 44832
rect 3568 44820 3574 44872
rect 3602 44820 3608 44872
rect 3660 44860 3666 44872
rect 4525 44863 4583 44869
rect 4525 44860 4537 44863
rect 3660 44832 4537 44860
rect 3660 44820 3666 44832
rect 4525 44829 4537 44832
rect 4571 44829 4583 44863
rect 4525 44823 4583 44829
rect 6362 44820 6368 44872
rect 6420 44860 6426 44872
rect 7024 44860 7052 44891
rect 7558 44888 7564 44900
rect 7616 44888 7622 44940
rect 7926 44928 7932 44940
rect 7887 44900 7932 44928
rect 7926 44888 7932 44900
rect 7984 44888 7990 44940
rect 8018 44888 8024 44940
rect 8076 44928 8082 44940
rect 8297 44931 8355 44937
rect 8297 44928 8309 44931
rect 8076 44900 8309 44928
rect 8076 44888 8082 44900
rect 8297 44897 8309 44900
rect 8343 44897 8355 44931
rect 9490 44928 9496 44940
rect 9451 44900 9496 44928
rect 8297 44891 8355 44897
rect 9490 44888 9496 44900
rect 9548 44888 9554 44940
rect 9674 44928 9680 44940
rect 9635 44900 9680 44928
rect 9674 44888 9680 44900
rect 9732 44888 9738 44940
rect 12342 44888 12348 44940
rect 12400 44928 12406 44940
rect 13173 44931 13231 44937
rect 13173 44928 13185 44931
rect 12400 44900 13185 44928
rect 12400 44888 12406 44900
rect 13173 44897 13185 44900
rect 13219 44897 13231 44931
rect 13173 44891 13231 44897
rect 13449 44931 13507 44937
rect 13449 44897 13461 44931
rect 13495 44928 13507 44931
rect 14277 44931 14335 44937
rect 14277 44928 14289 44931
rect 13495 44900 14289 44928
rect 13495 44897 13507 44900
rect 13449 44891 13507 44897
rect 14277 44897 14289 44900
rect 14323 44897 14335 44931
rect 14277 44891 14335 44897
rect 14921 44931 14979 44937
rect 14921 44897 14933 44931
rect 14967 44928 14979 44931
rect 15562 44928 15568 44940
rect 14967 44900 15568 44928
rect 14967 44897 14979 44900
rect 14921 44891 14979 44897
rect 15562 44888 15568 44900
rect 15620 44888 15626 44940
rect 17586 44888 17592 44940
rect 17644 44928 17650 44940
rect 17681 44931 17739 44937
rect 17681 44928 17693 44931
rect 17644 44900 17693 44928
rect 17644 44888 17650 44900
rect 17681 44897 17693 44900
rect 17727 44897 17739 44931
rect 18138 44928 18144 44940
rect 18099 44900 18144 44928
rect 17681 44891 17739 44897
rect 18138 44888 18144 44900
rect 18196 44888 18202 44940
rect 18230 44888 18236 44940
rect 18288 44928 18294 44940
rect 18417 44931 18475 44937
rect 18417 44928 18429 44931
rect 18288 44900 18429 44928
rect 18288 44888 18294 44900
rect 18417 44897 18429 44900
rect 18463 44897 18475 44931
rect 18966 44928 18972 44940
rect 18879 44900 18972 44928
rect 18417 44891 18475 44897
rect 18966 44888 18972 44900
rect 19024 44888 19030 44940
rect 19613 44931 19671 44937
rect 19613 44897 19625 44931
rect 19659 44928 19671 44931
rect 20088 44928 20116 44956
rect 19659 44900 20116 44928
rect 19659 44897 19671 44900
rect 19613 44891 19671 44897
rect 22554 44888 22560 44940
rect 22612 44928 22618 44940
rect 22649 44931 22707 44937
rect 22649 44928 22661 44931
rect 22612 44900 22661 44928
rect 22612 44888 22618 44900
rect 22649 44897 22661 44900
rect 22695 44897 22707 44931
rect 22649 44891 22707 44897
rect 8754 44860 8760 44872
rect 6420 44832 7052 44860
rect 8715 44832 8760 44860
rect 6420 44820 6426 44832
rect 8754 44820 8760 44832
rect 8812 44820 8818 44872
rect 12894 44860 12900 44872
rect 12855 44832 12900 44860
rect 12894 44820 12900 44832
rect 12952 44820 12958 44872
rect 13081 44863 13139 44869
rect 13081 44829 13093 44863
rect 13127 44860 13139 44863
rect 13538 44860 13544 44872
rect 13127 44832 13544 44860
rect 13127 44829 13139 44832
rect 13081 44823 13139 44829
rect 13538 44820 13544 44832
rect 13596 44820 13602 44872
rect 13633 44863 13691 44869
rect 13633 44829 13645 44863
rect 13679 44829 13691 44863
rect 14090 44860 14096 44872
rect 14051 44832 14096 44860
rect 13633 44823 13691 44829
rect 3528 44792 3556 44820
rect 4798 44792 4804 44804
rect 3528 44764 4804 44792
rect 4798 44752 4804 44764
rect 4856 44752 4862 44804
rect 6638 44752 6644 44804
rect 6696 44792 6702 44804
rect 6825 44795 6883 44801
rect 6825 44792 6837 44795
rect 6696 44764 6837 44792
rect 6696 44752 6702 44764
rect 6825 44761 6837 44764
rect 6871 44761 6883 44795
rect 6825 44755 6883 44761
rect 10778 44752 10784 44804
rect 10836 44792 10842 44804
rect 13648 44792 13676 44823
rect 14090 44820 14096 44832
rect 14148 44820 14154 44872
rect 14550 44820 14556 44872
rect 14608 44860 14614 44872
rect 14829 44863 14887 44869
rect 14829 44860 14841 44863
rect 14608 44832 14841 44860
rect 14608 44820 14614 44832
rect 14829 44829 14841 44832
rect 14875 44829 14887 44863
rect 14829 44823 14887 44829
rect 16117 44863 16175 44869
rect 16117 44829 16129 44863
rect 16163 44829 16175 44863
rect 16117 44823 16175 44829
rect 16301 44863 16359 44869
rect 16301 44829 16313 44863
rect 16347 44860 16359 44863
rect 22664 44860 22692 44891
rect 22738 44888 22744 44940
rect 22796 44928 22802 44940
rect 22833 44931 22891 44937
rect 22833 44928 22845 44931
rect 22796 44900 22845 44928
rect 22796 44888 22802 44900
rect 22833 44897 22845 44900
rect 22879 44897 22891 44931
rect 23290 44928 23296 44940
rect 23251 44900 23296 44928
rect 22833 44891 22891 44897
rect 23290 44888 23296 44900
rect 23348 44888 23354 44940
rect 23477 44931 23535 44937
rect 23477 44897 23489 44931
rect 23523 44897 23535 44931
rect 24412 44928 24440 45027
rect 27890 44996 27896 45008
rect 27851 44968 27896 44996
rect 27890 44956 27896 44968
rect 27948 44956 27954 45008
rect 25133 44931 25191 44937
rect 25133 44928 25145 44931
rect 24412 44900 25145 44928
rect 23477 44891 23535 44897
rect 25133 44897 25145 44900
rect 25179 44897 25191 44931
rect 25314 44928 25320 44940
rect 25275 44900 25320 44928
rect 25133 44891 25191 44897
rect 23382 44860 23388 44872
rect 16347 44832 19288 44860
rect 22664 44832 23388 44860
rect 16347 44829 16359 44832
rect 16301 44823 16359 44829
rect 10836 44764 13676 44792
rect 10836 44752 10842 44764
rect 14458 44752 14464 44804
rect 14516 44792 14522 44804
rect 14645 44795 14703 44801
rect 14645 44792 14657 44795
rect 14516 44764 14657 44792
rect 14516 44752 14522 44764
rect 14645 44761 14657 44764
rect 14691 44761 14703 44795
rect 15654 44792 15660 44804
rect 15615 44764 15660 44792
rect 14645 44755 14703 44761
rect 15654 44752 15660 44764
rect 15712 44752 15718 44804
rect 16132 44792 16160 44823
rect 18782 44792 18788 44804
rect 16132 44764 18788 44792
rect 18782 44752 18788 44764
rect 18840 44752 18846 44804
rect 1946 44724 1952 44736
rect 1907 44696 1952 44724
rect 1946 44684 1952 44696
rect 2004 44684 2010 44736
rect 2406 44684 2412 44736
rect 2464 44724 2470 44736
rect 2501 44727 2559 44733
rect 2501 44724 2513 44727
rect 2464 44696 2513 44724
rect 2464 44684 2470 44696
rect 2501 44693 2513 44696
rect 2547 44693 2559 44727
rect 2501 44687 2559 44693
rect 3602 44684 3608 44736
rect 3660 44724 3666 44736
rect 3973 44727 4031 44733
rect 3973 44724 3985 44727
rect 3660 44696 3985 44724
rect 3660 44684 3666 44696
rect 3973 44693 3985 44696
rect 4019 44693 4031 44727
rect 3973 44687 4031 44693
rect 5813 44727 5871 44733
rect 5813 44693 5825 44727
rect 5859 44724 5871 44727
rect 6730 44724 6736 44736
rect 5859 44696 6736 44724
rect 5859 44693 5871 44696
rect 5813 44687 5871 44693
rect 6730 44684 6736 44696
rect 6788 44684 6794 44736
rect 7098 44684 7104 44736
rect 7156 44724 7162 44736
rect 8386 44724 8392 44736
rect 7156 44696 8392 44724
rect 7156 44684 7162 44696
rect 8386 44684 8392 44696
rect 8444 44684 8450 44736
rect 9217 44727 9275 44733
rect 9217 44693 9229 44727
rect 9263 44724 9275 44727
rect 9306 44724 9312 44736
rect 9263 44696 9312 44724
rect 9263 44693 9275 44696
rect 9217 44687 9275 44693
rect 9306 44684 9312 44696
rect 9364 44684 9370 44736
rect 9493 44727 9551 44733
rect 9493 44693 9505 44727
rect 9539 44724 9551 44727
rect 9766 44724 9772 44736
rect 9539 44696 9772 44724
rect 9539 44693 9551 44696
rect 9493 44687 9551 44693
rect 9766 44684 9772 44696
rect 9824 44684 9830 44736
rect 19150 44724 19156 44736
rect 19111 44696 19156 44724
rect 19150 44684 19156 44696
rect 19208 44684 19214 44736
rect 19260 44724 19288 44832
rect 23382 44820 23388 44832
rect 23440 44860 23446 44872
rect 23492 44860 23520 44891
rect 25314 44888 25320 44900
rect 25372 44888 25378 44940
rect 26142 44888 26148 44940
rect 26200 44928 26206 44940
rect 26237 44931 26295 44937
rect 26237 44928 26249 44931
rect 26200 44900 26249 44928
rect 26200 44888 26206 44900
rect 26237 44897 26249 44900
rect 26283 44897 26295 44931
rect 26237 44891 26295 44897
rect 26881 44931 26939 44937
rect 26881 44897 26893 44931
rect 26927 44928 26939 44931
rect 27154 44928 27160 44940
rect 26927 44900 27160 44928
rect 26927 44897 26939 44900
rect 26881 44891 26939 44897
rect 27154 44888 27160 44900
rect 27212 44888 27218 44940
rect 23440 44832 23520 44860
rect 23440 44820 23446 44832
rect 22186 44792 22192 44804
rect 20548 44764 22192 44792
rect 20548 44724 20576 44764
rect 22186 44752 22192 44764
rect 22244 44752 22250 44804
rect 23934 44752 23940 44804
rect 23992 44792 23998 44804
rect 28077 44795 28135 44801
rect 28077 44792 28089 44795
rect 23992 44764 28089 44792
rect 23992 44752 23998 44764
rect 28077 44761 28089 44764
rect 28123 44761 28135 44795
rect 28077 44755 28135 44761
rect 19260 44696 20576 44724
rect 20993 44727 21051 44733
rect 20993 44693 21005 44727
rect 21039 44724 21051 44727
rect 21634 44724 21640 44736
rect 21039 44696 21640 44724
rect 21039 44693 21051 44696
rect 20993 44687 21051 44693
rect 21634 44684 21640 44696
rect 21692 44684 21698 44736
rect 24213 44727 24271 44733
rect 24213 44693 24225 44727
rect 24259 44724 24271 44727
rect 24762 44724 24768 44736
rect 24259 44696 24768 44724
rect 24259 44693 24271 44696
rect 24213 44687 24271 44693
rect 24762 44684 24768 44696
rect 24820 44684 24826 44736
rect 24857 44727 24915 44733
rect 24857 44693 24869 44727
rect 24903 44724 24915 44727
rect 24946 44724 24952 44736
rect 24903 44696 24952 44724
rect 24903 44693 24915 44696
rect 24857 44687 24915 44693
rect 24946 44684 24952 44696
rect 25004 44684 25010 44736
rect 25130 44724 25136 44736
rect 25091 44696 25136 44724
rect 25130 44684 25136 44696
rect 25188 44684 25194 44736
rect 26050 44724 26056 44736
rect 26011 44696 26056 44724
rect 26050 44684 26056 44696
rect 26108 44684 26114 44736
rect 26694 44724 26700 44736
rect 26655 44696 26700 44724
rect 26694 44684 26700 44696
rect 26752 44684 26758 44736
rect 1104 44634 28888 44656
rect 1104 44582 5614 44634
rect 5666 44582 5678 44634
rect 5730 44582 5742 44634
rect 5794 44582 5806 44634
rect 5858 44582 14878 44634
rect 14930 44582 14942 44634
rect 14994 44582 15006 44634
rect 15058 44582 15070 44634
rect 15122 44582 24142 44634
rect 24194 44582 24206 44634
rect 24258 44582 24270 44634
rect 24322 44582 24334 44634
rect 24386 44582 28888 44634
rect 1104 44560 28888 44582
rect 3050 44480 3056 44532
rect 3108 44520 3114 44532
rect 3145 44523 3203 44529
rect 3145 44520 3157 44523
rect 3108 44492 3157 44520
rect 3108 44480 3114 44492
rect 3145 44489 3157 44492
rect 3191 44520 3203 44523
rect 4982 44520 4988 44532
rect 3191 44492 4988 44520
rect 3191 44489 3203 44492
rect 3145 44483 3203 44489
rect 4982 44480 4988 44492
rect 5040 44480 5046 44532
rect 6454 44520 6460 44532
rect 6415 44492 6460 44520
rect 6454 44480 6460 44492
rect 6512 44480 6518 44532
rect 23934 44520 23940 44532
rect 7576 44492 23940 44520
rect 1854 44412 1860 44464
rect 1912 44452 1918 44464
rect 1949 44455 2007 44461
rect 1949 44452 1961 44455
rect 1912 44424 1961 44452
rect 1912 44412 1918 44424
rect 1949 44421 1961 44424
rect 1995 44421 2007 44455
rect 1949 44415 2007 44421
rect 2682 44412 2688 44464
rect 2740 44452 2746 44464
rect 7576 44452 7604 44492
rect 23934 44480 23940 44492
rect 23992 44480 23998 44532
rect 24029 44523 24087 44529
rect 24029 44489 24041 44523
rect 24075 44520 24087 44523
rect 25314 44520 25320 44532
rect 24075 44492 25320 44520
rect 24075 44489 24087 44492
rect 24029 44483 24087 44489
rect 25314 44480 25320 44492
rect 25372 44480 25378 44532
rect 2740 44424 7604 44452
rect 7745 44455 7803 44461
rect 2740 44412 2746 44424
rect 7745 44421 7757 44455
rect 7791 44452 7803 44455
rect 9674 44452 9680 44464
rect 7791 44424 9680 44452
rect 7791 44421 7803 44424
rect 7745 44415 7803 44421
rect 9674 44412 9680 44424
rect 9732 44412 9738 44464
rect 11146 44452 11152 44464
rect 11107 44424 11152 44452
rect 11146 44412 11152 44424
rect 11204 44412 11210 44464
rect 16114 44452 16120 44464
rect 16075 44424 16120 44452
rect 16114 44412 16120 44424
rect 16172 44412 16178 44464
rect 18230 44452 18236 44464
rect 18191 44424 18236 44452
rect 18230 44412 18236 44424
rect 18288 44412 18294 44464
rect 18690 44412 18696 44464
rect 18748 44452 18754 44464
rect 19981 44455 20039 44461
rect 19981 44452 19993 44455
rect 18748 44424 19993 44452
rect 18748 44412 18754 44424
rect 19981 44421 19993 44424
rect 20027 44421 20039 44455
rect 19981 44415 20039 44421
rect 2409 44387 2467 44393
rect 2409 44353 2421 44387
rect 2455 44384 2467 44387
rect 4338 44384 4344 44396
rect 2455 44356 4344 44384
rect 2455 44353 2467 44356
rect 2409 44347 2467 44353
rect 4338 44344 4344 44356
rect 4396 44344 4402 44396
rect 5442 44384 5448 44396
rect 5403 44356 5448 44384
rect 5442 44344 5448 44356
rect 5500 44344 5506 44396
rect 7098 44384 7104 44396
rect 7059 44356 7104 44384
rect 7098 44344 7104 44356
rect 7156 44344 7162 44396
rect 9585 44387 9643 44393
rect 9585 44384 9597 44387
rect 7484 44356 9597 44384
rect 2222 44276 2228 44328
rect 2280 44316 2286 44328
rect 2501 44319 2559 44325
rect 2501 44316 2513 44319
rect 2280 44288 2513 44316
rect 2280 44276 2286 44288
rect 2501 44285 2513 44288
rect 2547 44285 2559 44319
rect 3050 44316 3056 44328
rect 3011 44288 3056 44316
rect 2501 44279 2559 44285
rect 3050 44276 3056 44288
rect 3108 44276 3114 44328
rect 6730 44276 6736 44328
rect 6788 44316 6794 44328
rect 6825 44319 6883 44325
rect 6825 44316 6837 44319
rect 6788 44288 6837 44316
rect 6788 44276 6794 44288
rect 6825 44285 6837 44288
rect 6871 44285 6883 44319
rect 6825 44279 6883 44285
rect 6917 44319 6975 44325
rect 6917 44285 6929 44319
rect 6963 44316 6975 44319
rect 7484 44316 7512 44356
rect 9585 44353 9597 44356
rect 9631 44353 9643 44387
rect 9766 44384 9772 44396
rect 9727 44356 9772 44384
rect 9585 44347 9643 44353
rect 6963 44288 7512 44316
rect 6963 44285 6975 44288
rect 6917 44279 6975 44285
rect 7558 44276 7564 44328
rect 7616 44316 7622 44328
rect 8021 44319 8079 44325
rect 8021 44316 8033 44319
rect 7616 44288 8033 44316
rect 7616 44276 7622 44288
rect 8021 44285 8033 44288
rect 8067 44285 8079 44319
rect 8021 44279 8079 44285
rect 9398 44276 9404 44328
rect 9456 44316 9462 44328
rect 9493 44319 9551 44325
rect 9493 44316 9505 44319
rect 9456 44288 9505 44316
rect 9456 44276 9462 44288
rect 9493 44285 9505 44288
rect 9539 44285 9551 44319
rect 9493 44279 9551 44285
rect 2406 44248 2412 44260
rect 2367 44220 2412 44248
rect 2406 44208 2412 44220
rect 2464 44208 2470 44260
rect 5169 44251 5227 44257
rect 5169 44217 5181 44251
rect 5215 44248 5227 44251
rect 5902 44248 5908 44260
rect 5215 44220 5908 44248
rect 5215 44217 5227 44220
rect 5169 44211 5227 44217
rect 5902 44208 5908 44220
rect 5960 44208 5966 44260
rect 7742 44248 7748 44260
rect 7703 44220 7748 44248
rect 7742 44208 7748 44220
rect 7800 44248 7806 44260
rect 8202 44248 8208 44260
rect 7800 44220 8208 44248
rect 7800 44208 7806 44220
rect 8202 44208 8208 44220
rect 8260 44208 8266 44260
rect 9600 44248 9628 44347
rect 9766 44344 9772 44356
rect 9824 44344 9830 44396
rect 12894 44344 12900 44396
rect 12952 44384 12958 44396
rect 13541 44387 13599 44393
rect 13541 44384 13553 44387
rect 12952 44356 13553 44384
rect 12952 44344 12958 44356
rect 13541 44353 13553 44356
rect 13587 44384 13599 44387
rect 13722 44384 13728 44396
rect 13587 44356 13728 44384
rect 13587 44353 13599 44356
rect 13541 44347 13599 44353
rect 13722 44344 13728 44356
rect 13780 44344 13786 44396
rect 15470 44344 15476 44396
rect 15528 44384 15534 44396
rect 16390 44384 16396 44396
rect 15528 44356 16396 44384
rect 15528 44344 15534 44356
rect 16390 44344 16396 44356
rect 16448 44344 16454 44396
rect 17405 44387 17463 44393
rect 17405 44353 17417 44387
rect 17451 44384 17463 44387
rect 18138 44384 18144 44396
rect 17451 44356 18144 44384
rect 17451 44353 17463 44356
rect 17405 44347 17463 44353
rect 18138 44344 18144 44356
rect 18196 44384 18202 44396
rect 18325 44387 18383 44393
rect 18325 44384 18337 44387
rect 18196 44356 18337 44384
rect 18196 44344 18202 44356
rect 18325 44353 18337 44356
rect 18371 44353 18383 44387
rect 19996 44384 20024 44415
rect 20070 44412 20076 44464
rect 20128 44452 20134 44464
rect 21174 44452 21180 44464
rect 20128 44424 21180 44452
rect 20128 44412 20134 44424
rect 21174 44412 21180 44424
rect 21232 44452 21238 44464
rect 22005 44455 22063 44461
rect 22005 44452 22017 44455
rect 21232 44424 22017 44452
rect 21232 44412 21238 44424
rect 22005 44421 22017 44424
rect 22051 44421 22063 44455
rect 23474 44452 23480 44464
rect 23435 44424 23480 44452
rect 22005 44415 22063 44421
rect 22020 44384 22048 44415
rect 23474 44412 23480 44424
rect 23532 44412 23538 44464
rect 25406 44452 25412 44464
rect 23952 44424 25412 44452
rect 19996 44356 21956 44384
rect 22020 44356 23520 44384
rect 18325 44347 18383 44353
rect 10042 44276 10048 44328
rect 10100 44316 10106 44328
rect 10229 44319 10287 44325
rect 10229 44316 10241 44319
rect 10100 44288 10241 44316
rect 10100 44276 10106 44288
rect 10229 44285 10241 44288
rect 10275 44285 10287 44319
rect 10229 44279 10287 44285
rect 10686 44276 10692 44328
rect 10744 44316 10750 44328
rect 11333 44319 11391 44325
rect 11333 44316 11345 44319
rect 10744 44288 11345 44316
rect 10744 44276 10750 44288
rect 11333 44285 11345 44288
rect 11379 44285 11391 44319
rect 13262 44316 13268 44328
rect 13223 44288 13268 44316
rect 11333 44279 11391 44285
rect 13262 44276 13268 44288
rect 13320 44276 13326 44328
rect 13449 44319 13507 44325
rect 13449 44285 13461 44319
rect 13495 44316 13507 44319
rect 14090 44316 14096 44328
rect 13495 44288 14096 44316
rect 13495 44285 13507 44288
rect 13449 44279 13507 44285
rect 14090 44276 14096 44288
rect 14148 44276 14154 44328
rect 16025 44319 16083 44325
rect 16025 44285 16037 44319
rect 16071 44285 16083 44319
rect 16025 44279 16083 44285
rect 16209 44319 16267 44325
rect 16209 44285 16221 44319
rect 16255 44316 16267 44319
rect 16408 44316 16436 44344
rect 16255 44288 16436 44316
rect 16945 44319 17003 44325
rect 16255 44285 16267 44288
rect 16209 44279 16267 44285
rect 16945 44285 16957 44319
rect 16991 44285 17003 44319
rect 17126 44316 17132 44328
rect 17087 44288 17132 44316
rect 16945 44279 17003 44285
rect 10321 44251 10379 44257
rect 10321 44248 10333 44251
rect 9600 44220 10333 44248
rect 10321 44217 10333 44220
rect 10367 44217 10379 44251
rect 16040 44248 16068 44279
rect 16960 44248 16988 44279
rect 17126 44276 17132 44288
rect 17184 44276 17190 44328
rect 17586 44276 17592 44328
rect 17644 44316 17650 44328
rect 18049 44319 18107 44325
rect 18049 44316 18061 44319
rect 17644 44288 18061 44316
rect 17644 44276 17650 44288
rect 18049 44285 18061 44288
rect 18095 44285 18107 44319
rect 18049 44279 18107 44285
rect 18785 44319 18843 44325
rect 18785 44285 18797 44319
rect 18831 44316 18843 44319
rect 19794 44316 19800 44328
rect 18831 44288 19800 44316
rect 18831 44285 18843 44288
rect 18785 44279 18843 44285
rect 19794 44276 19800 44288
rect 19852 44276 19858 44328
rect 20165 44319 20223 44325
rect 20165 44285 20177 44319
rect 20211 44316 20223 44319
rect 20714 44316 20720 44328
rect 20211 44288 20720 44316
rect 20211 44285 20223 44288
rect 20165 44279 20223 44285
rect 20714 44276 20720 44288
rect 20772 44276 20778 44328
rect 21266 44316 21272 44328
rect 21227 44288 21272 44316
rect 21266 44276 21272 44288
rect 21324 44316 21330 44328
rect 21818 44316 21824 44328
rect 21324 44288 21824 44316
rect 21324 44276 21330 44288
rect 21818 44276 21824 44288
rect 21876 44276 21882 44328
rect 21928 44316 21956 44356
rect 22189 44319 22247 44325
rect 22189 44316 22201 44319
rect 21928 44288 22201 44316
rect 22189 44285 22201 44288
rect 22235 44285 22247 44319
rect 22189 44279 22247 44285
rect 23385 44319 23443 44325
rect 23385 44285 23397 44319
rect 23431 44285 23443 44319
rect 23492 44316 23520 44356
rect 23566 44344 23572 44396
rect 23624 44384 23630 44396
rect 23842 44384 23848 44396
rect 23624 44356 23848 44384
rect 23624 44344 23630 44356
rect 23842 44344 23848 44356
rect 23900 44344 23906 44396
rect 23952 44316 23980 44424
rect 25406 44412 25412 44424
rect 25464 44452 25470 44464
rect 25464 44424 25544 44452
rect 25464 44412 25470 44424
rect 24486 44384 24492 44396
rect 24044 44356 24492 44384
rect 24044 44325 24072 44356
rect 24486 44344 24492 44356
rect 24544 44344 24550 44396
rect 24854 44344 24860 44396
rect 24912 44344 24918 44396
rect 25516 44393 25544 44424
rect 25501 44387 25559 44393
rect 25501 44353 25513 44387
rect 25547 44353 25559 44387
rect 25501 44347 25559 44353
rect 23492 44288 23980 44316
rect 24029 44319 24087 44325
rect 23385 44279 23443 44285
rect 24029 44285 24041 44319
rect 24075 44285 24087 44319
rect 24029 44279 24087 44285
rect 24305 44319 24363 44325
rect 24305 44285 24317 44319
rect 24351 44316 24363 44319
rect 24872 44316 24900 44344
rect 25406 44316 25412 44328
rect 24351 44288 25412 44316
rect 24351 44285 24363 44288
rect 24305 44279 24363 44285
rect 17310 44248 17316 44260
rect 16040 44220 17316 44248
rect 10321 44211 10379 44217
rect 17310 44208 17316 44220
rect 17368 44208 17374 44260
rect 17865 44251 17923 44257
rect 17865 44217 17877 44251
rect 17911 44248 17923 44251
rect 19334 44248 19340 44260
rect 17911 44220 19340 44248
rect 17911 44217 17923 44220
rect 17865 44211 17923 44217
rect 19334 44208 19340 44220
rect 19392 44208 19398 44260
rect 23400 44248 23428 44279
rect 25406 44276 25412 44288
rect 25464 44276 25470 44328
rect 25516 44316 25544 44347
rect 25590 44316 25596 44328
rect 25516 44288 25596 44316
rect 25590 44276 25596 44288
rect 25648 44276 25654 44328
rect 26878 44276 26884 44328
rect 26936 44316 26942 44328
rect 27985 44319 28043 44325
rect 27985 44316 27997 44319
rect 26936 44288 27997 44316
rect 26936 44276 26942 44288
rect 27985 44285 27997 44288
rect 28031 44285 28043 44319
rect 27985 44279 28043 44285
rect 23566 44248 23572 44260
rect 23400 44220 23572 44248
rect 23566 44208 23572 44220
rect 23624 44248 23630 44260
rect 23624 44220 24348 44248
rect 23624 44208 23630 44220
rect 4798 44180 4804 44192
rect 4759 44152 4804 44180
rect 4798 44140 4804 44152
rect 4856 44140 4862 44192
rect 5261 44183 5319 44189
rect 5261 44149 5273 44183
rect 5307 44180 5319 44183
rect 6362 44180 6368 44192
rect 5307 44152 6368 44180
rect 5307 44149 5319 44152
rect 5261 44143 5319 44149
rect 6362 44140 6368 44152
rect 6420 44140 6426 44192
rect 7929 44183 7987 44189
rect 7929 44149 7941 44183
rect 7975 44180 7987 44183
rect 8018 44180 8024 44192
rect 7975 44152 8024 44180
rect 7975 44149 7987 44152
rect 7929 44143 7987 44149
rect 8018 44140 8024 44152
rect 8076 44140 8082 44192
rect 9766 44180 9772 44192
rect 9727 44152 9772 44180
rect 9766 44140 9772 44152
rect 9824 44140 9830 44192
rect 12802 44140 12808 44192
rect 12860 44180 12866 44192
rect 13262 44180 13268 44192
rect 12860 44152 13268 44180
rect 12860 44140 12866 44152
rect 13262 44140 13268 44152
rect 13320 44140 13326 44192
rect 18966 44180 18972 44192
rect 18927 44152 18972 44180
rect 18966 44140 18972 44152
rect 19024 44140 19030 44192
rect 19794 44140 19800 44192
rect 19852 44180 19858 44192
rect 21266 44180 21272 44192
rect 19852 44152 21272 44180
rect 19852 44140 19858 44152
rect 21266 44140 21272 44152
rect 21324 44140 21330 44192
rect 21453 44183 21511 44189
rect 21453 44149 21465 44183
rect 21499 44180 21511 44183
rect 21542 44180 21548 44192
rect 21499 44152 21548 44180
rect 21499 44149 21511 44152
rect 21453 44143 21511 44149
rect 21542 44140 21548 44152
rect 21600 44140 21606 44192
rect 23934 44140 23940 44192
rect 23992 44180 23998 44192
rect 24213 44183 24271 44189
rect 24213 44180 24225 44183
rect 23992 44152 24225 44180
rect 23992 44140 23998 44152
rect 24213 44149 24225 44152
rect 24259 44149 24271 44183
rect 24320 44180 24348 44220
rect 24854 44208 24860 44260
rect 24912 44248 24918 44260
rect 25746 44251 25804 44257
rect 25746 44248 25758 44251
rect 24912 44220 25758 44248
rect 24912 44208 24918 44220
rect 25746 44217 25758 44220
rect 25792 44217 25804 44251
rect 25746 44211 25804 44217
rect 26881 44183 26939 44189
rect 26881 44180 26893 44183
rect 24320 44152 26893 44180
rect 24213 44143 24271 44149
rect 26881 44149 26893 44152
rect 26927 44149 26939 44183
rect 28074 44180 28080 44192
rect 28035 44152 28080 44180
rect 26881 44143 26939 44149
rect 28074 44140 28080 44152
rect 28132 44140 28138 44192
rect 1104 44090 28888 44112
rect 1104 44038 10246 44090
rect 10298 44038 10310 44090
rect 10362 44038 10374 44090
rect 10426 44038 10438 44090
rect 10490 44038 19510 44090
rect 19562 44038 19574 44090
rect 19626 44038 19638 44090
rect 19690 44038 19702 44090
rect 19754 44038 28888 44090
rect 1104 44016 28888 44038
rect 3418 43976 3424 43988
rect 3379 43948 3424 43976
rect 3418 43936 3424 43948
rect 3476 43936 3482 43988
rect 5629 43979 5687 43985
rect 5629 43945 5641 43979
rect 5675 43976 5687 43979
rect 5902 43976 5908 43988
rect 5675 43948 5908 43976
rect 5675 43945 5687 43948
rect 5629 43939 5687 43945
rect 5902 43936 5908 43948
rect 5960 43936 5966 43988
rect 6638 43936 6644 43988
rect 6696 43976 6702 43988
rect 7745 43979 7803 43985
rect 6696 43948 7604 43976
rect 6696 43936 6702 43948
rect 1857 43911 1915 43917
rect 1857 43877 1869 43911
rect 1903 43908 1915 43911
rect 4516 43911 4574 43917
rect 1903 43880 3096 43908
rect 1903 43877 1915 43880
rect 1857 43871 1915 43877
rect 2593 43843 2651 43849
rect 2593 43809 2605 43843
rect 2639 43840 2651 43843
rect 2682 43840 2688 43852
rect 2639 43812 2688 43840
rect 2639 43809 2651 43812
rect 2593 43803 2651 43809
rect 2682 43800 2688 43812
rect 2740 43800 2746 43852
rect 2774 43664 2780 43716
rect 2832 43704 2838 43716
rect 2832 43676 2877 43704
rect 2832 43664 2838 43676
rect 1394 43596 1400 43648
rect 1452 43636 1458 43648
rect 1949 43639 2007 43645
rect 1949 43636 1961 43639
rect 1452 43608 1961 43636
rect 1452 43596 1458 43608
rect 1949 43605 1961 43608
rect 1995 43605 2007 43639
rect 3068 43636 3096 43880
rect 4516 43877 4528 43911
rect 4562 43908 4574 43911
rect 4798 43908 4804 43920
rect 4562 43880 4804 43908
rect 4562 43877 4574 43880
rect 4516 43871 4574 43877
rect 4798 43868 4804 43880
rect 4856 43868 4862 43920
rect 6822 43868 6828 43920
rect 6880 43868 6886 43920
rect 7576 43908 7604 43948
rect 7745 43945 7757 43979
rect 7791 43976 7803 43979
rect 7926 43976 7932 43988
rect 7791 43948 7932 43976
rect 7791 43945 7803 43948
rect 7745 43939 7803 43945
rect 7926 43936 7932 43948
rect 7984 43936 7990 43988
rect 8202 43936 8208 43988
rect 8260 43976 8266 43988
rect 8389 43979 8447 43985
rect 8389 43976 8401 43979
rect 8260 43948 8401 43976
rect 8260 43936 8266 43948
rect 8389 43945 8401 43948
rect 8435 43945 8447 43979
rect 8389 43939 8447 43945
rect 8588 43948 9996 43976
rect 7576 43880 8524 43908
rect 3145 43843 3203 43849
rect 3145 43809 3157 43843
rect 3191 43840 3203 43843
rect 3329 43843 3387 43849
rect 3329 43840 3341 43843
rect 3191 43812 3341 43840
rect 3191 43809 3203 43812
rect 3145 43803 3203 43809
rect 3329 43809 3341 43812
rect 3375 43840 3387 43843
rect 6840 43840 6868 43868
rect 7009 43843 7067 43849
rect 7009 43840 7021 43843
rect 3375 43812 6316 43840
rect 6840 43812 7021 43840
rect 3375 43809 3387 43812
rect 3329 43803 3387 43809
rect 3970 43732 3976 43784
rect 4028 43772 4034 43784
rect 4249 43775 4307 43781
rect 4249 43772 4261 43775
rect 4028 43744 4261 43772
rect 4028 43732 4034 43744
rect 4249 43741 4261 43744
rect 4295 43741 4307 43775
rect 4249 43735 4307 43741
rect 6288 43704 6316 43812
rect 7009 43809 7021 43812
rect 7055 43809 7067 43843
rect 7576 43840 7604 43880
rect 8496 43849 8524 43880
rect 7653 43843 7711 43849
rect 7653 43840 7665 43843
rect 7576 43812 7665 43840
rect 7009 43803 7067 43809
rect 7653 43809 7665 43812
rect 7699 43809 7711 43843
rect 7653 43803 7711 43809
rect 8297 43843 8355 43849
rect 8297 43809 8309 43843
rect 8343 43809 8355 43843
rect 8297 43803 8355 43809
rect 8481 43843 8539 43849
rect 8481 43809 8493 43843
rect 8527 43809 8539 43843
rect 8481 43803 8539 43809
rect 6362 43732 6368 43784
rect 6420 43772 6426 43784
rect 6825 43775 6883 43781
rect 6825 43772 6837 43775
rect 6420 43744 6837 43772
rect 6420 43732 6426 43744
rect 6825 43741 6837 43744
rect 6871 43741 6883 43775
rect 6825 43735 6883 43741
rect 7193 43775 7251 43781
rect 7193 43741 7205 43775
rect 7239 43772 7251 43775
rect 7742 43772 7748 43784
rect 7239 43744 7748 43772
rect 7239 43741 7251 43744
rect 7193 43735 7251 43741
rect 7742 43732 7748 43744
rect 7800 43772 7806 43784
rect 8312 43772 8340 43803
rect 7800 43744 8340 43772
rect 7800 43732 7806 43744
rect 8588 43704 8616 43948
rect 9766 43868 9772 43920
rect 9824 43917 9830 43920
rect 9824 43911 9888 43917
rect 9824 43877 9842 43911
rect 9876 43877 9888 43911
rect 9968 43908 9996 43948
rect 10042 43936 10048 43988
rect 10100 43976 10106 43988
rect 10965 43979 11023 43985
rect 10965 43976 10977 43979
rect 10100 43948 10977 43976
rect 10100 43936 10106 43948
rect 10965 43945 10977 43948
rect 11011 43945 11023 43979
rect 24673 43979 24731 43985
rect 10965 43939 11023 43945
rect 12406 43948 24624 43976
rect 12406 43908 12434 43948
rect 9968 43880 12434 43908
rect 13357 43911 13415 43917
rect 9824 43871 9888 43877
rect 13357 43877 13369 43911
rect 13403 43908 13415 43911
rect 13538 43908 13544 43920
rect 13403 43880 13544 43908
rect 13403 43877 13415 43880
rect 13357 43871 13415 43877
rect 9824 43868 9830 43871
rect 13538 43868 13544 43880
rect 13596 43868 13602 43920
rect 14734 43868 14740 43920
rect 14792 43908 14798 43920
rect 15013 43911 15071 43917
rect 15013 43908 15025 43911
rect 14792 43880 15025 43908
rect 14792 43868 14798 43880
rect 15013 43877 15025 43880
rect 15059 43877 15071 43911
rect 15013 43871 15071 43877
rect 17681 43911 17739 43917
rect 17681 43877 17693 43911
rect 17727 43908 17739 43911
rect 18414 43908 18420 43920
rect 17727 43880 18420 43908
rect 17727 43877 17739 43880
rect 17681 43871 17739 43877
rect 18414 43868 18420 43880
rect 18472 43868 18478 43920
rect 20717 43911 20775 43917
rect 20717 43877 20729 43911
rect 20763 43908 20775 43911
rect 21358 43908 21364 43920
rect 20763 43880 21364 43908
rect 20763 43877 20775 43880
rect 20717 43871 20775 43877
rect 21358 43868 21364 43880
rect 21416 43868 21422 43920
rect 21450 43868 21456 43920
rect 21508 43908 21514 43920
rect 23842 43908 23848 43920
rect 21508 43880 23848 43908
rect 21508 43868 21514 43880
rect 23842 43868 23848 43880
rect 23900 43908 23906 43920
rect 23900 43880 24440 43908
rect 23900 43868 23906 43880
rect 9125 43843 9183 43849
rect 9125 43809 9137 43843
rect 9171 43840 9183 43843
rect 10686 43840 10692 43852
rect 9171 43812 10692 43840
rect 9171 43809 9183 43812
rect 9125 43803 9183 43809
rect 10686 43800 10692 43812
rect 10744 43800 10750 43852
rect 12618 43800 12624 43852
rect 12676 43840 12682 43852
rect 13265 43843 13323 43849
rect 13265 43840 13277 43843
rect 12676 43812 13277 43840
rect 12676 43800 12682 43812
rect 13265 43809 13277 43812
rect 13311 43809 13323 43843
rect 13265 43803 13323 43809
rect 14642 43800 14648 43852
rect 14700 43840 14706 43852
rect 14829 43843 14887 43849
rect 14829 43840 14841 43843
rect 14700 43812 14841 43840
rect 14700 43800 14706 43812
rect 14829 43809 14841 43812
rect 14875 43809 14887 43843
rect 17586 43840 17592 43852
rect 17547 43812 17592 43840
rect 14829 43803 14887 43809
rect 17586 43800 17592 43812
rect 17644 43800 17650 43852
rect 18782 43840 18788 43852
rect 18743 43812 18788 43840
rect 18782 43800 18788 43812
rect 18840 43840 18846 43852
rect 19058 43840 19064 43852
rect 18840 43812 19064 43840
rect 18840 43800 18846 43812
rect 19058 43800 19064 43812
rect 19116 43800 19122 43852
rect 19150 43800 19156 43852
rect 19208 43840 19214 43852
rect 19429 43843 19487 43849
rect 19429 43840 19441 43843
rect 19208 43812 19441 43840
rect 19208 43800 19214 43812
rect 19429 43809 19441 43812
rect 19475 43809 19487 43843
rect 19429 43803 19487 43809
rect 20809 43843 20867 43849
rect 20809 43809 20821 43843
rect 20855 43840 20867 43843
rect 21913 43843 21971 43849
rect 21913 43840 21925 43843
rect 20855 43812 21925 43840
rect 20855 43809 20867 43812
rect 20809 43803 20867 43809
rect 21913 43809 21925 43812
rect 21959 43809 21971 43843
rect 23382 43840 23388 43852
rect 21913 43803 21971 43809
rect 22112 43812 23388 43840
rect 9214 43732 9220 43784
rect 9272 43772 9278 43784
rect 9585 43775 9643 43781
rect 9585 43772 9597 43775
rect 9272 43744 9597 43772
rect 9272 43732 9278 43744
rect 9585 43741 9597 43744
rect 9631 43741 9643 43775
rect 18874 43772 18880 43784
rect 18835 43744 18880 43772
rect 9585 43735 9643 43741
rect 18874 43732 18880 43744
rect 18932 43732 18938 43784
rect 19334 43772 19340 43784
rect 19295 43744 19340 43772
rect 19334 43732 19340 43744
rect 19392 43732 19398 43784
rect 20990 43772 20996 43784
rect 20903 43744 20996 43772
rect 20990 43732 20996 43744
rect 21048 43772 21054 43784
rect 21542 43772 21548 43784
rect 21048 43744 21548 43772
rect 21048 43732 21054 43744
rect 21542 43732 21548 43744
rect 21600 43732 21606 43784
rect 21818 43732 21824 43784
rect 21876 43772 21882 43784
rect 22112 43772 22140 43812
rect 23382 43800 23388 43812
rect 23440 43840 23446 43852
rect 24412 43849 24440 43880
rect 23569 43843 23627 43849
rect 23569 43840 23581 43843
rect 23440 43812 23581 43840
rect 23440 43800 23446 43812
rect 23569 43809 23581 43812
rect 23615 43809 23627 43843
rect 23569 43803 23627 43809
rect 24397 43843 24455 43849
rect 24397 43809 24409 43843
rect 24443 43809 24455 43843
rect 24596 43840 24624 43948
rect 24673 43945 24685 43979
rect 24719 43976 24731 43979
rect 24854 43976 24860 43988
rect 24719 43948 24860 43976
rect 24719 43945 24731 43948
rect 24673 43939 24731 43945
rect 24854 43936 24860 43948
rect 24912 43936 24918 43988
rect 25498 43936 25504 43988
rect 25556 43976 25562 43988
rect 25682 43976 25688 43988
rect 25556 43948 25688 43976
rect 25556 43936 25562 43948
rect 25682 43936 25688 43948
rect 25740 43936 25746 43988
rect 24946 43868 24952 43920
rect 25004 43908 25010 43920
rect 25314 43908 25320 43920
rect 25004 43880 25320 43908
rect 25004 43868 25010 43880
rect 25314 43868 25320 43880
rect 25372 43868 25378 43920
rect 26050 43868 26056 43920
rect 26108 43908 26114 43920
rect 26697 43911 26755 43917
rect 26697 43908 26709 43911
rect 26108 43880 26709 43908
rect 26108 43868 26114 43880
rect 26697 43877 26709 43880
rect 26743 43877 26755 43911
rect 26697 43871 26755 43877
rect 25501 43843 25559 43849
rect 24596 43812 25268 43840
rect 24397 43803 24455 43809
rect 21876 43744 22140 43772
rect 21876 43732 21882 43744
rect 23474 43732 23480 43784
rect 23532 43772 23538 43784
rect 24489 43775 24547 43781
rect 24489 43772 24501 43775
rect 23532 43744 24501 43772
rect 23532 43732 23538 43744
rect 24489 43741 24501 43744
rect 24535 43741 24547 43775
rect 24489 43735 24547 43741
rect 24673 43775 24731 43781
rect 24673 43741 24685 43775
rect 24719 43772 24731 43775
rect 25130 43772 25136 43784
rect 24719 43744 25136 43772
rect 24719 43741 24731 43744
rect 24673 43735 24731 43741
rect 25130 43732 25136 43744
rect 25188 43732 25194 43784
rect 25240 43772 25268 43812
rect 25501 43809 25513 43843
rect 25547 43840 25559 43843
rect 25958 43840 25964 43852
rect 25547 43812 25964 43840
rect 25547 43809 25559 43812
rect 25501 43803 25559 43809
rect 25958 43800 25964 43812
rect 26016 43800 26022 43852
rect 26142 43840 26148 43852
rect 26103 43812 26148 43840
rect 26142 43800 26148 43812
rect 26200 43800 26206 43852
rect 26234 43800 26240 43852
rect 26292 43840 26298 43852
rect 27985 43843 28043 43849
rect 27985 43840 27997 43843
rect 26292 43812 27997 43840
rect 26292 43800 26298 43812
rect 27985 43809 27997 43812
rect 28031 43809 28043 43843
rect 27985 43803 28043 43809
rect 28074 43772 28080 43784
rect 25240 43744 28080 43772
rect 28074 43732 28080 43744
rect 28132 43732 28138 43784
rect 6288 43676 8616 43704
rect 8680 43676 9168 43704
rect 8680 43636 8708 43676
rect 3068 43608 8708 43636
rect 8941 43639 8999 43645
rect 1949 43599 2007 43605
rect 8941 43605 8953 43639
rect 8987 43636 8999 43639
rect 9030 43636 9036 43648
rect 8987 43608 9036 43636
rect 8987 43605 8999 43608
rect 8941 43599 8999 43605
rect 9030 43596 9036 43608
rect 9088 43596 9094 43648
rect 9140 43636 9168 43676
rect 10594 43664 10600 43716
rect 10652 43704 10658 43716
rect 10652 43676 17816 43704
rect 10652 43664 10658 43676
rect 10778 43636 10784 43648
rect 9140 43608 10784 43636
rect 10778 43596 10784 43608
rect 10836 43596 10842 43648
rect 17788 43636 17816 43676
rect 18322 43664 18328 43716
rect 18380 43704 18386 43716
rect 18785 43707 18843 43713
rect 18785 43704 18797 43707
rect 18380 43676 18797 43704
rect 18380 43664 18386 43676
rect 18785 43673 18797 43676
rect 18831 43673 18843 43707
rect 25961 43707 26019 43713
rect 18785 43667 18843 43673
rect 18892 43676 25544 43704
rect 18892 43636 18920 43676
rect 17788 43608 18920 43636
rect 20254 43596 20260 43648
rect 20312 43636 20318 43648
rect 20349 43639 20407 43645
rect 20349 43636 20361 43639
rect 20312 43608 20361 43636
rect 20312 43596 20318 43608
rect 20349 43605 20361 43608
rect 20395 43605 20407 43639
rect 20349 43599 20407 43605
rect 21913 43639 21971 43645
rect 21913 43605 21925 43639
rect 21959 43636 21971 43639
rect 22370 43636 22376 43648
rect 21959 43608 22376 43636
rect 21959 43605 21971 43608
rect 21913 43599 21971 43605
rect 22370 43596 22376 43608
rect 22428 43596 22434 43648
rect 23753 43639 23811 43645
rect 23753 43605 23765 43639
rect 23799 43636 23811 43639
rect 23842 43636 23848 43648
rect 23799 43608 23848 43636
rect 23799 43605 23811 43608
rect 23753 43599 23811 43605
rect 23842 43596 23848 43608
rect 23900 43596 23906 43648
rect 25516 43636 25544 43676
rect 25961 43673 25973 43707
rect 26007 43704 26019 43707
rect 27246 43704 27252 43716
rect 26007 43676 27252 43704
rect 26007 43673 26019 43676
rect 25961 43667 26019 43673
rect 27246 43664 27252 43676
rect 27304 43664 27310 43716
rect 26789 43639 26847 43645
rect 26789 43636 26801 43639
rect 25516 43608 26801 43636
rect 26789 43605 26801 43608
rect 26835 43605 26847 43639
rect 28074 43636 28080 43648
rect 28035 43608 28080 43636
rect 26789 43599 26847 43605
rect 28074 43596 28080 43608
rect 28132 43596 28138 43648
rect 1104 43546 28888 43568
rect 1104 43494 5614 43546
rect 5666 43494 5678 43546
rect 5730 43494 5742 43546
rect 5794 43494 5806 43546
rect 5858 43494 14878 43546
rect 14930 43494 14942 43546
rect 14994 43494 15006 43546
rect 15058 43494 15070 43546
rect 15122 43494 24142 43546
rect 24194 43494 24206 43546
rect 24258 43494 24270 43546
rect 24322 43494 24334 43546
rect 24386 43494 28888 43546
rect 1104 43472 28888 43494
rect 1302 43392 1308 43444
rect 1360 43432 1366 43444
rect 2685 43435 2743 43441
rect 2685 43432 2697 43435
rect 1360 43404 2697 43432
rect 1360 43392 1366 43404
rect 2685 43401 2697 43404
rect 2731 43401 2743 43435
rect 2685 43395 2743 43401
rect 4341 43435 4399 43441
rect 4341 43401 4353 43435
rect 4387 43432 4399 43435
rect 4430 43432 4436 43444
rect 4387 43404 4436 43432
rect 4387 43401 4399 43404
rect 4341 43395 4399 43401
rect 4430 43392 4436 43404
rect 4488 43392 4494 43444
rect 4614 43392 4620 43444
rect 4672 43432 4678 43444
rect 4985 43435 5043 43441
rect 4985 43432 4997 43435
rect 4672 43404 4997 43432
rect 4672 43392 4678 43404
rect 4985 43401 4997 43404
rect 5031 43401 5043 43435
rect 4985 43395 5043 43401
rect 5813 43435 5871 43441
rect 5813 43401 5825 43435
rect 5859 43432 5871 43435
rect 6178 43432 6184 43444
rect 5859 43404 6184 43432
rect 5859 43401 5871 43404
rect 5813 43395 5871 43401
rect 6178 43392 6184 43404
rect 6236 43392 6242 43444
rect 10137 43435 10195 43441
rect 10137 43401 10149 43435
rect 10183 43432 10195 43435
rect 10686 43432 10692 43444
rect 10183 43404 10692 43432
rect 10183 43401 10195 43404
rect 10137 43395 10195 43401
rect 10686 43392 10692 43404
rect 10744 43392 10750 43444
rect 10778 43392 10784 43444
rect 10836 43432 10842 43444
rect 21358 43432 21364 43444
rect 10836 43404 20944 43432
rect 21319 43404 21364 43432
rect 10836 43392 10842 43404
rect 1762 43324 1768 43376
rect 1820 43364 1826 43376
rect 10594 43364 10600 43376
rect 1820 43336 10600 43364
rect 1820 43324 1826 43336
rect 10594 43324 10600 43336
rect 10652 43324 10658 43376
rect 12894 43324 12900 43376
rect 12952 43364 12958 43376
rect 13078 43364 13084 43376
rect 12952 43336 13084 43364
rect 12952 43324 12958 43336
rect 13078 43324 13084 43336
rect 13136 43324 13142 43376
rect 20916 43364 20944 43404
rect 21358 43392 21364 43404
rect 21416 43432 21422 43444
rect 23014 43432 23020 43444
rect 21416 43404 23020 43432
rect 21416 43392 21422 43404
rect 23014 43392 23020 43404
rect 23072 43392 23078 43444
rect 25314 43432 25320 43444
rect 25275 43404 25320 43432
rect 25314 43392 25320 43404
rect 25372 43392 25378 43444
rect 28077 43435 28135 43441
rect 28077 43432 28089 43435
rect 25424 43404 28089 43432
rect 25424 43364 25452 43404
rect 28077 43401 28089 43404
rect 28123 43401 28135 43435
rect 28077 43395 28135 43401
rect 20916 43336 25452 43364
rect 26513 43367 26571 43373
rect 26513 43333 26525 43367
rect 26559 43364 26571 43367
rect 27982 43364 27988 43376
rect 26559 43336 27988 43364
rect 26559 43333 26571 43336
rect 26513 43327 26571 43333
rect 27982 43324 27988 43336
rect 28040 43324 28046 43376
rect 4080 43268 11008 43296
rect 2593 43231 2651 43237
rect 2593 43197 2605 43231
rect 2639 43228 2651 43231
rect 4080 43228 4108 43268
rect 2639 43200 4108 43228
rect 2639 43197 2651 43200
rect 2593 43191 2651 43197
rect 4154 43188 4160 43240
rect 4212 43228 4218 43240
rect 4249 43231 4307 43237
rect 4249 43228 4261 43231
rect 4212 43200 4261 43228
rect 4212 43188 4218 43200
rect 4249 43197 4261 43200
rect 4295 43228 4307 43231
rect 4614 43228 4620 43240
rect 4295 43200 4620 43228
rect 4295 43197 4307 43200
rect 4249 43191 4307 43197
rect 4614 43188 4620 43200
rect 4672 43188 4678 43240
rect 4890 43228 4896 43240
rect 4851 43200 4896 43228
rect 4890 43188 4896 43200
rect 4948 43188 4954 43240
rect 5721 43231 5779 43237
rect 5721 43197 5733 43231
rect 5767 43197 5779 43231
rect 5721 43191 5779 43197
rect 5905 43231 5963 43237
rect 5905 43197 5917 43231
rect 5951 43228 5963 43231
rect 6178 43228 6184 43240
rect 5951 43200 6184 43228
rect 5951 43197 5963 43200
rect 5905 43191 5963 43197
rect 1857 43163 1915 43169
rect 1857 43129 1869 43163
rect 1903 43160 1915 43163
rect 2498 43160 2504 43172
rect 1903 43132 2504 43160
rect 1903 43129 1915 43132
rect 1857 43123 1915 43129
rect 2498 43120 2504 43132
rect 2556 43120 2562 43172
rect 3326 43120 3332 43172
rect 3384 43160 3390 43172
rect 4430 43160 4436 43172
rect 3384 43132 4436 43160
rect 3384 43120 3390 43132
rect 4430 43120 4436 43132
rect 4488 43120 4494 43172
rect 5736 43160 5764 43191
rect 6178 43188 6184 43200
rect 6236 43228 6242 43240
rect 6546 43228 6552 43240
rect 6236 43200 6552 43228
rect 6236 43188 6242 43200
rect 6546 43188 6552 43200
rect 6604 43188 6610 43240
rect 9490 43228 9496 43240
rect 9451 43200 9496 43228
rect 9490 43188 9496 43200
rect 9548 43188 9554 43240
rect 10321 43231 10379 43237
rect 10321 43197 10333 43231
rect 10367 43228 10379 43231
rect 10686 43228 10692 43240
rect 10367 43200 10692 43228
rect 10367 43197 10379 43200
rect 10321 43191 10379 43197
rect 10686 43188 10692 43200
rect 10744 43188 10750 43240
rect 10873 43231 10931 43237
rect 10873 43197 10885 43231
rect 10919 43197 10931 43231
rect 10980 43228 11008 43268
rect 16040 43268 19104 43296
rect 15013 43231 15071 43237
rect 10980 43200 12434 43228
rect 10873 43191 10931 43197
rect 6270 43160 6276 43172
rect 5736 43132 6276 43160
rect 6270 43120 6276 43132
rect 6328 43120 6334 43172
rect 10888 43160 10916 43191
rect 11146 43169 11152 43172
rect 10888 43132 11100 43160
rect 11072 43104 11100 43132
rect 11140 43123 11152 43169
rect 11204 43160 11210 43172
rect 12406 43160 12434 43200
rect 15013 43197 15025 43231
rect 15059 43228 15071 43231
rect 15102 43228 15108 43240
rect 15059 43200 15108 43228
rect 15059 43197 15071 43200
rect 15013 43191 15071 43197
rect 15102 43188 15108 43200
rect 15160 43188 15166 43240
rect 16040 43228 16068 43268
rect 15212 43200 16068 43228
rect 17589 43231 17647 43237
rect 15212 43160 15240 43200
rect 17589 43197 17601 43231
rect 17635 43228 17647 43231
rect 18690 43228 18696 43240
rect 17635 43200 18696 43228
rect 17635 43197 17647 43200
rect 17589 43191 17647 43197
rect 18690 43188 18696 43200
rect 18748 43188 18754 43240
rect 18782 43188 18788 43240
rect 18840 43228 18846 43240
rect 18840 43200 18885 43228
rect 18840 43188 18846 43200
rect 15286 43169 15292 43172
rect 11204 43132 11240 43160
rect 12406 43132 15240 43160
rect 11146 43120 11152 43123
rect 11204 43120 11210 43132
rect 15280 43123 15292 43169
rect 15344 43160 15350 43172
rect 18601 43163 18659 43169
rect 15344 43132 15380 43160
rect 16224 43132 17448 43160
rect 15286 43120 15292 43123
rect 15344 43120 15350 43132
rect 1949 43095 2007 43101
rect 1949 43061 1961 43095
rect 1995 43092 2007 43095
rect 2958 43092 2964 43104
rect 1995 43064 2964 43092
rect 1995 43061 2007 43064
rect 1949 43055 2007 43061
rect 2958 43052 2964 43064
rect 3016 43052 3022 43104
rect 9306 43052 9312 43104
rect 9364 43092 9370 43104
rect 9585 43095 9643 43101
rect 9585 43092 9597 43095
rect 9364 43064 9597 43092
rect 9364 43052 9370 43064
rect 9585 43061 9597 43064
rect 9631 43061 9643 43095
rect 9585 43055 9643 43061
rect 11054 43052 11060 43104
rect 11112 43092 11118 43104
rect 11606 43092 11612 43104
rect 11112 43064 11612 43092
rect 11112 43052 11118 43064
rect 11606 43052 11612 43064
rect 11664 43052 11670 43104
rect 12253 43095 12311 43101
rect 12253 43061 12265 43095
rect 12299 43092 12311 43095
rect 12342 43092 12348 43104
rect 12299 43064 12348 43092
rect 12299 43061 12311 43064
rect 12253 43055 12311 43061
rect 12342 43052 12348 43064
rect 12400 43052 12406 43104
rect 15194 43052 15200 43104
rect 15252 43092 15258 43104
rect 15378 43092 15384 43104
rect 15252 43064 15384 43092
rect 15252 43052 15258 43064
rect 15378 43052 15384 43064
rect 15436 43092 15442 43104
rect 16224 43092 16252 43132
rect 16390 43092 16396 43104
rect 15436 43064 16252 43092
rect 16351 43064 16396 43092
rect 15436 43052 15442 43064
rect 16390 43052 16396 43064
rect 16448 43052 16454 43104
rect 17420 43101 17448 43132
rect 18601 43129 18613 43163
rect 18647 43129 18659 43163
rect 18966 43160 18972 43172
rect 18927 43132 18972 43160
rect 18601 43123 18659 43129
rect 17405 43095 17463 43101
rect 17405 43061 17417 43095
rect 17451 43092 17463 43095
rect 18414 43092 18420 43104
rect 17451 43064 18420 43092
rect 17451 43061 17463 43064
rect 17405 43055 17463 43061
rect 18414 43052 18420 43064
rect 18472 43052 18478 43104
rect 18616 43092 18644 43123
rect 18966 43120 18972 43132
rect 19024 43120 19030 43172
rect 19076 43160 19104 43268
rect 22278 43256 22284 43308
rect 22336 43296 22342 43308
rect 22373 43299 22431 43305
rect 22373 43296 22385 43299
rect 22336 43268 22385 43296
rect 22336 43256 22342 43268
rect 22373 43265 22385 43268
rect 22419 43265 22431 43299
rect 27433 43299 27491 43305
rect 27433 43296 27445 43299
rect 22373 43259 22431 43265
rect 22480 43268 27445 43296
rect 19981 43231 20039 43237
rect 19981 43197 19993 43231
rect 20027 43228 20039 43231
rect 20070 43228 20076 43240
rect 20027 43200 20076 43228
rect 20027 43197 20039 43200
rect 19981 43191 20039 43197
rect 20070 43188 20076 43200
rect 20128 43188 20134 43240
rect 20254 43237 20260 43240
rect 20248 43228 20260 43237
rect 20215 43200 20260 43228
rect 20248 43191 20260 43200
rect 20254 43188 20260 43191
rect 20312 43188 20318 43240
rect 22480 43228 22508 43268
rect 27433 43265 27445 43268
rect 27479 43265 27491 43299
rect 27433 43259 27491 43265
rect 23014 43228 23020 43240
rect 22066 43200 22508 43228
rect 22975 43200 23020 43228
rect 22066 43160 22094 43200
rect 23014 43188 23020 43200
rect 23072 43188 23078 43240
rect 24305 43231 24363 43237
rect 24305 43197 24317 43231
rect 24351 43228 24363 43231
rect 24854 43228 24860 43240
rect 24351 43200 24860 43228
rect 24351 43197 24363 43200
rect 24305 43191 24363 43197
rect 24854 43188 24860 43200
rect 24912 43188 24918 43240
rect 25130 43188 25136 43240
rect 25188 43228 25194 43240
rect 25225 43231 25283 43237
rect 25225 43228 25237 43231
rect 25188 43200 25237 43228
rect 25188 43188 25194 43200
rect 25225 43197 25237 43200
rect 25271 43197 25283 43231
rect 26050 43228 26056 43240
rect 26011 43200 26056 43228
rect 25225 43191 25283 43197
rect 26050 43188 26056 43200
rect 26108 43188 26114 43240
rect 26697 43231 26755 43237
rect 26697 43197 26709 43231
rect 26743 43228 26755 43231
rect 26786 43228 26792 43240
rect 26743 43200 26792 43228
rect 26743 43197 26755 43200
rect 26697 43191 26755 43197
rect 26786 43188 26792 43200
rect 26844 43188 26850 43240
rect 19076 43132 22094 43160
rect 22189 43163 22247 43169
rect 22189 43129 22201 43163
rect 22235 43160 22247 43163
rect 23109 43163 23167 43169
rect 23109 43160 23121 43163
rect 22235 43132 23121 43160
rect 22235 43129 22247 43132
rect 22189 43123 22247 43129
rect 23109 43129 23121 43132
rect 23155 43129 23167 43163
rect 26234 43160 26240 43172
rect 23109 43123 23167 43129
rect 24136 43132 26240 43160
rect 18874 43092 18880 43104
rect 18616 43064 18880 43092
rect 18874 43052 18880 43064
rect 18932 43092 18938 43104
rect 21450 43092 21456 43104
rect 18932 43064 21456 43092
rect 18932 43052 18938 43064
rect 21450 43052 21456 43064
rect 21508 43052 21514 43104
rect 21818 43092 21824 43104
rect 21779 43064 21824 43092
rect 21818 43052 21824 43064
rect 21876 43052 21882 43104
rect 22278 43092 22284 43104
rect 22239 43064 22284 43092
rect 22278 43052 22284 43064
rect 22336 43052 22342 43104
rect 24136 43101 24164 43132
rect 26234 43120 26240 43132
rect 26292 43120 26298 43172
rect 27246 43160 27252 43172
rect 27207 43132 27252 43160
rect 27246 43120 27252 43132
rect 27304 43120 27310 43172
rect 27985 43163 28043 43169
rect 27985 43129 27997 43163
rect 28031 43129 28043 43163
rect 27985 43123 28043 43129
rect 24121 43095 24179 43101
rect 24121 43061 24133 43095
rect 24167 43061 24179 43095
rect 24121 43055 24179 43061
rect 25869 43095 25927 43101
rect 25869 43061 25881 43095
rect 25915 43092 25927 43095
rect 28000 43092 28028 43123
rect 25915 43064 28028 43092
rect 25915 43061 25927 43064
rect 25869 43055 25927 43061
rect 1104 43002 28888 43024
rect 1104 42950 10246 43002
rect 10298 42950 10310 43002
rect 10362 42950 10374 43002
rect 10426 42950 10438 43002
rect 10490 42950 19510 43002
rect 19562 42950 19574 43002
rect 19626 42950 19638 43002
rect 19690 42950 19702 43002
rect 19754 42950 28888 43002
rect 1104 42928 28888 42950
rect 2590 42848 2596 42900
rect 2648 42888 2654 42900
rect 28074 42888 28080 42900
rect 2648 42860 28080 42888
rect 2648 42848 2654 42860
rect 28074 42848 28080 42860
rect 28132 42848 28138 42900
rect 1578 42780 1584 42832
rect 1636 42820 1642 42832
rect 4890 42820 4896 42832
rect 1636 42792 4896 42820
rect 1636 42780 1642 42792
rect 4890 42780 4896 42792
rect 4948 42780 4954 42832
rect 11146 42820 11152 42832
rect 11107 42792 11152 42820
rect 11146 42780 11152 42792
rect 11204 42780 11210 42832
rect 11238 42780 11244 42832
rect 11296 42820 11302 42832
rect 12437 42823 12495 42829
rect 12437 42820 12449 42823
rect 11296 42792 12449 42820
rect 11296 42780 11302 42792
rect 12437 42789 12449 42792
rect 12483 42789 12495 42823
rect 12437 42783 12495 42789
rect 12526 42780 12532 42832
rect 12584 42820 12590 42832
rect 18684 42823 18742 42829
rect 12584 42792 12629 42820
rect 12584 42780 12590 42792
rect 18684 42789 18696 42823
rect 18730 42820 18742 42823
rect 18966 42820 18972 42832
rect 18730 42792 18972 42820
rect 18730 42789 18742 42792
rect 18684 42783 18742 42789
rect 18966 42780 18972 42792
rect 19024 42780 19030 42832
rect 21818 42780 21824 42832
rect 21876 42820 21882 42832
rect 23109 42823 23167 42829
rect 23109 42820 23121 42823
rect 21876 42792 23121 42820
rect 21876 42780 21882 42792
rect 23109 42789 23121 42792
rect 23155 42789 23167 42823
rect 23109 42783 23167 42789
rect 23382 42780 23388 42832
rect 23440 42820 23446 42832
rect 25130 42820 25136 42832
rect 23440 42792 25136 42820
rect 23440 42780 23446 42792
rect 25130 42780 25136 42792
rect 25188 42780 25194 42832
rect 1857 42755 1915 42761
rect 1857 42721 1869 42755
rect 1903 42752 1915 42755
rect 2406 42752 2412 42764
rect 1903 42724 2412 42752
rect 1903 42721 1915 42724
rect 1857 42715 1915 42721
rect 2406 42712 2412 42724
rect 2464 42712 2470 42764
rect 2590 42752 2596 42764
rect 2551 42724 2596 42752
rect 2590 42712 2596 42724
rect 2648 42712 2654 42764
rect 3697 42755 3755 42761
rect 3697 42721 3709 42755
rect 3743 42721 3755 42755
rect 3697 42715 3755 42721
rect 4525 42755 4583 42761
rect 4525 42721 4537 42755
rect 4571 42721 4583 42755
rect 4525 42715 4583 42721
rect 4709 42755 4767 42761
rect 4709 42721 4721 42755
rect 4755 42752 4767 42755
rect 4982 42752 4988 42764
rect 4755 42724 4988 42752
rect 4755 42721 4767 42724
rect 4709 42715 4767 42721
rect 3602 42684 3608 42696
rect 3563 42656 3608 42684
rect 3602 42644 3608 42656
rect 3660 42644 3666 42696
rect 3712 42684 3740 42715
rect 4154 42684 4160 42696
rect 3712 42656 4160 42684
rect 4154 42644 4160 42656
rect 4212 42644 4218 42696
rect 4430 42644 4436 42696
rect 4488 42684 4494 42696
rect 4540 42684 4568 42715
rect 4982 42712 4988 42724
rect 5040 42712 5046 42764
rect 7653 42755 7711 42761
rect 7653 42721 7665 42755
rect 7699 42752 7711 42755
rect 7742 42752 7748 42764
rect 7699 42724 7748 42752
rect 7699 42721 7711 42724
rect 7653 42715 7711 42721
rect 7742 42712 7748 42724
rect 7800 42712 7806 42764
rect 8849 42755 8907 42761
rect 8849 42721 8861 42755
rect 8895 42752 8907 42755
rect 9490 42752 9496 42764
rect 8895 42724 9496 42752
rect 8895 42721 8907 42724
rect 8849 42715 8907 42721
rect 9490 42712 9496 42724
rect 9548 42752 9554 42764
rect 9861 42755 9919 42761
rect 9861 42752 9873 42755
rect 9548 42724 9873 42752
rect 9548 42712 9554 42724
rect 9861 42721 9873 42724
rect 9907 42721 9919 42755
rect 10778 42752 10784 42764
rect 10739 42724 10784 42752
rect 9861 42715 9919 42721
rect 10778 42712 10784 42724
rect 10836 42712 10842 42764
rect 10965 42755 11023 42761
rect 10965 42721 10977 42755
rect 11011 42752 11023 42755
rect 12342 42752 12348 42764
rect 11011 42724 12348 42752
rect 11011 42721 11023 42724
rect 10965 42715 11023 42721
rect 12342 42712 12348 42724
rect 12400 42712 12406 42764
rect 14274 42752 14280 42764
rect 12636 42724 14280 42752
rect 4488 42656 4568 42684
rect 4488 42644 4494 42656
rect 9398 42644 9404 42696
rect 9456 42684 9462 42696
rect 10045 42687 10103 42693
rect 10045 42684 10057 42687
rect 9456 42656 10057 42684
rect 9456 42644 9462 42656
rect 10045 42653 10057 42656
rect 10091 42684 10103 42687
rect 12636 42684 12664 42724
rect 14274 42712 14280 42724
rect 14332 42712 14338 42764
rect 18414 42752 18420 42764
rect 18375 42724 18420 42752
rect 18414 42712 18420 42724
rect 18472 42712 18478 42764
rect 21453 42755 21511 42761
rect 21453 42721 21465 42755
rect 21499 42721 21511 42755
rect 21453 42715 21511 42721
rect 21545 42755 21603 42761
rect 21545 42721 21557 42755
rect 21591 42752 21603 42755
rect 22278 42752 22284 42764
rect 21591 42724 22284 42752
rect 21591 42721 21603 42724
rect 21545 42715 21603 42721
rect 10091 42656 12664 42684
rect 12713 42687 12771 42693
rect 10091 42653 10103 42656
rect 10045 42647 10103 42653
rect 12713 42653 12725 42687
rect 12759 42684 12771 42687
rect 13630 42684 13636 42696
rect 12759 42656 13636 42684
rect 12759 42653 12771 42656
rect 12713 42647 12771 42653
rect 13630 42644 13636 42656
rect 13688 42644 13694 42696
rect 13722 42644 13728 42696
rect 13780 42684 13786 42696
rect 13998 42684 14004 42696
rect 13780 42656 13825 42684
rect 13959 42656 14004 42684
rect 13780 42644 13786 42656
rect 13998 42644 14004 42656
rect 14056 42644 14062 42696
rect 14182 42644 14188 42696
rect 14240 42684 14246 42696
rect 15105 42687 15163 42693
rect 15105 42684 15117 42687
rect 14240 42656 15117 42684
rect 14240 42644 14246 42656
rect 15105 42653 15117 42656
rect 15151 42653 15163 42687
rect 15105 42647 15163 42653
rect 2774 42576 2780 42628
rect 2832 42616 2838 42628
rect 3620 42616 3648 42644
rect 4890 42616 4896 42628
rect 2832 42588 2877 42616
rect 3620 42588 4896 42616
rect 2832 42576 2838 42588
rect 4890 42576 4896 42588
rect 4948 42576 4954 42628
rect 5442 42576 5448 42628
rect 5500 42616 5506 42628
rect 7374 42616 7380 42628
rect 5500 42588 7380 42616
rect 5500 42576 5506 42588
rect 7374 42576 7380 42588
rect 7432 42616 7438 42628
rect 9033 42619 9091 42625
rect 9033 42616 9045 42619
rect 7432 42588 9045 42616
rect 7432 42576 7438 42588
rect 9033 42585 9045 42588
rect 9079 42585 9091 42619
rect 11606 42616 11612 42628
rect 9033 42579 9091 42585
rect 11072 42588 11612 42616
rect 11072 42560 11100 42588
rect 11606 42576 11612 42588
rect 11664 42616 11670 42628
rect 12250 42616 12256 42628
rect 11664 42588 12256 42616
rect 11664 42576 11670 42588
rect 12250 42576 12256 42588
rect 12308 42616 12314 42628
rect 13740 42616 13768 42644
rect 12308 42588 13768 42616
rect 21468 42616 21496 42715
rect 22278 42712 22284 42724
rect 22336 42712 22342 42764
rect 23842 42752 23848 42764
rect 23803 42724 23848 42752
rect 23842 42712 23848 42724
rect 23900 42712 23906 42764
rect 24026 42752 24032 42764
rect 23987 42724 24032 42752
rect 24026 42712 24032 42724
rect 24084 42712 24090 42764
rect 26694 42752 26700 42764
rect 26655 42724 26700 42752
rect 26694 42712 26700 42724
rect 26752 42712 26758 42764
rect 27982 42752 27988 42764
rect 27943 42724 27988 42752
rect 27982 42712 27988 42724
rect 28040 42712 28046 42764
rect 22186 42644 22192 42696
rect 22244 42684 22250 42696
rect 23017 42687 23075 42693
rect 23017 42684 23029 42687
rect 22244 42656 23029 42684
rect 22244 42644 22250 42656
rect 23017 42653 23029 42656
rect 23063 42653 23075 42687
rect 23198 42684 23204 42696
rect 23159 42656 23204 42684
rect 23017 42647 23075 42653
rect 23198 42644 23204 42656
rect 23256 42644 23262 42696
rect 24121 42687 24179 42693
rect 24121 42653 24133 42687
rect 24167 42684 24179 42687
rect 24486 42684 24492 42696
rect 24167 42656 24492 42684
rect 24167 42653 24179 42656
rect 24121 42647 24179 42653
rect 24486 42644 24492 42656
rect 24544 42644 24550 42696
rect 25409 42619 25467 42625
rect 25409 42616 25421 42619
rect 21468 42588 25421 42616
rect 12308 42576 12314 42588
rect 25409 42585 25421 42588
rect 25455 42616 25467 42619
rect 25498 42616 25504 42628
rect 25455 42588 25504 42616
rect 25455 42585 25467 42588
rect 25409 42579 25467 42585
rect 25498 42576 25504 42588
rect 25556 42576 25562 42628
rect 1946 42548 1952 42560
rect 1907 42520 1952 42548
rect 1946 42508 1952 42520
rect 2004 42508 2010 42560
rect 3878 42508 3884 42560
rect 3936 42548 3942 42560
rect 3973 42551 4031 42557
rect 3973 42548 3985 42551
rect 3936 42520 3985 42548
rect 3936 42508 3942 42520
rect 3973 42517 3985 42520
rect 4019 42517 4031 42551
rect 3973 42511 4031 42517
rect 4246 42508 4252 42560
rect 4304 42548 4310 42560
rect 4617 42551 4675 42557
rect 4617 42548 4629 42551
rect 4304 42520 4629 42548
rect 4304 42508 4310 42520
rect 4617 42517 4629 42520
rect 4663 42517 4675 42551
rect 4617 42511 4675 42517
rect 7745 42551 7803 42557
rect 7745 42517 7757 42551
rect 7791 42548 7803 42551
rect 8846 42548 8852 42560
rect 7791 42520 8852 42548
rect 7791 42517 7803 42520
rect 7745 42511 7803 42517
rect 8846 42508 8852 42520
rect 8904 42508 8910 42560
rect 11054 42508 11060 42560
rect 11112 42508 11118 42560
rect 12069 42551 12127 42557
rect 12069 42517 12081 42551
rect 12115 42548 12127 42551
rect 13170 42548 13176 42560
rect 12115 42520 13176 42548
rect 12115 42517 12127 42520
rect 12069 42511 12127 42517
rect 13170 42508 13176 42520
rect 13228 42508 13234 42560
rect 19794 42548 19800 42560
rect 19755 42520 19800 42548
rect 19794 42508 19800 42520
rect 19852 42508 19858 42560
rect 22649 42551 22707 42557
rect 22649 42517 22661 42551
rect 22695 42548 22707 42551
rect 23290 42548 23296 42560
rect 22695 42520 23296 42548
rect 22695 42517 22707 42520
rect 22649 42511 22707 42517
rect 23290 42508 23296 42520
rect 23348 42508 23354 42560
rect 25593 42551 25651 42557
rect 25593 42517 25605 42551
rect 25639 42548 25651 42551
rect 26142 42548 26148 42560
rect 25639 42520 26148 42548
rect 25639 42517 25651 42520
rect 25593 42511 25651 42517
rect 26142 42508 26148 42520
rect 26200 42508 26206 42560
rect 26602 42508 26608 42560
rect 26660 42548 26666 42560
rect 26789 42551 26847 42557
rect 26789 42548 26801 42551
rect 26660 42520 26801 42548
rect 26660 42508 26666 42520
rect 26789 42517 26801 42520
rect 26835 42517 26847 42551
rect 28074 42548 28080 42560
rect 28035 42520 28080 42548
rect 26789 42511 26847 42517
rect 28074 42508 28080 42520
rect 28132 42508 28138 42560
rect 1104 42458 28888 42480
rect 1104 42406 5614 42458
rect 5666 42406 5678 42458
rect 5730 42406 5742 42458
rect 5794 42406 5806 42458
rect 5858 42406 14878 42458
rect 14930 42406 14942 42458
rect 14994 42406 15006 42458
rect 15058 42406 15070 42458
rect 15122 42406 24142 42458
rect 24194 42406 24206 42458
rect 24258 42406 24270 42458
rect 24322 42406 24334 42458
rect 24386 42406 28888 42458
rect 1104 42384 28888 42406
rect 2590 42304 2596 42356
rect 2648 42344 2654 42356
rect 22186 42344 22192 42356
rect 2648 42316 22094 42344
rect 22147 42316 22192 42344
rect 2648 42304 2654 42316
rect 2777 42279 2835 42285
rect 2777 42245 2789 42279
rect 2823 42276 2835 42279
rect 2866 42276 2872 42288
rect 2823 42248 2872 42276
rect 2823 42245 2835 42248
rect 2777 42239 2835 42245
rect 2866 42236 2872 42248
rect 2924 42276 2930 42288
rect 13630 42276 13636 42288
rect 2924 42248 4936 42276
rect 13591 42248 13636 42276
rect 2924 42236 2930 42248
rect 4338 42208 4344 42220
rect 4299 42180 4344 42208
rect 4338 42168 4344 42180
rect 4396 42168 4402 42220
rect 1210 42100 1216 42152
rect 1268 42140 1274 42152
rect 1397 42143 1455 42149
rect 1397 42140 1409 42143
rect 1268 42112 1409 42140
rect 1268 42100 1274 42112
rect 1397 42109 1409 42112
rect 1443 42140 1455 42143
rect 3970 42140 3976 42152
rect 1443 42112 3976 42140
rect 1443 42109 1455 42112
rect 1397 42103 1455 42109
rect 3970 42100 3976 42112
rect 4028 42100 4034 42152
rect 4246 42140 4252 42152
rect 4207 42112 4252 42140
rect 4246 42100 4252 42112
rect 4304 42100 4310 42152
rect 4433 42143 4491 42149
rect 4433 42109 4445 42143
rect 4479 42140 4491 42143
rect 4522 42140 4528 42152
rect 4479 42112 4528 42140
rect 4479 42109 4491 42112
rect 4433 42103 4491 42109
rect 4522 42100 4528 42112
rect 4580 42100 4586 42152
rect 4908 42149 4936 42248
rect 13630 42236 13636 42248
rect 13688 42236 13694 42288
rect 15286 42276 15292 42288
rect 15247 42248 15292 42276
rect 15286 42236 15292 42248
rect 15344 42236 15350 42288
rect 17313 42279 17371 42285
rect 16500 42248 16804 42276
rect 7650 42168 7656 42220
rect 7708 42208 7714 42220
rect 9585 42211 9643 42217
rect 9585 42208 9597 42211
rect 7708 42180 9597 42208
rect 7708 42168 7714 42180
rect 9585 42177 9597 42180
rect 9631 42177 9643 42211
rect 9585 42171 9643 42177
rect 4893 42143 4951 42149
rect 4893 42109 4905 42143
rect 4939 42109 4951 42143
rect 4893 42103 4951 42109
rect 9398 42100 9404 42152
rect 9456 42140 9462 42152
rect 9493 42143 9551 42149
rect 9493 42140 9505 42143
rect 9456 42112 9505 42140
rect 9456 42100 9462 42112
rect 9493 42109 9505 42112
rect 9539 42109 9551 42143
rect 9600 42140 9628 42171
rect 9674 42168 9680 42220
rect 9732 42208 9738 42220
rect 9769 42211 9827 42217
rect 9769 42208 9781 42211
rect 9732 42180 9781 42208
rect 9732 42168 9738 42180
rect 9769 42177 9781 42180
rect 9815 42177 9827 42211
rect 12250 42208 12256 42220
rect 12211 42180 12256 42208
rect 9769 42171 9827 42177
rect 12250 42168 12256 42180
rect 12308 42168 12314 42220
rect 16500 42208 16528 42248
rect 16666 42208 16672 42220
rect 15120 42180 16528 42208
rect 16627 42180 16672 42208
rect 10134 42140 10140 42152
rect 9600 42112 10140 42140
rect 9493 42103 9551 42109
rect 10134 42100 10140 42112
rect 10192 42100 10198 42152
rect 12342 42100 12348 42152
rect 12400 42140 12406 42152
rect 15120 42149 15148 42180
rect 16666 42168 16672 42180
rect 16724 42168 16730 42220
rect 16776 42208 16804 42248
rect 17313 42245 17325 42279
rect 17359 42276 17371 42279
rect 19334 42276 19340 42288
rect 17359 42248 19340 42276
rect 17359 42245 17371 42248
rect 17313 42239 17371 42245
rect 19334 42236 19340 42248
rect 19392 42276 19398 42288
rect 19702 42276 19708 42288
rect 19392 42248 19708 42276
rect 19392 42236 19398 42248
rect 19702 42236 19708 42248
rect 19760 42236 19766 42288
rect 22066 42276 22094 42316
rect 22186 42304 22192 42316
rect 22244 42304 22250 42356
rect 24026 42304 24032 42356
rect 24084 42344 24090 42356
rect 24305 42347 24363 42353
rect 24305 42344 24317 42347
rect 24084 42316 24317 42344
rect 24084 42304 24090 42316
rect 24305 42313 24317 42316
rect 24351 42313 24363 42347
rect 28074 42344 28080 42356
rect 24305 42307 24363 42313
rect 24392 42316 28080 42344
rect 24392 42276 24420 42316
rect 28074 42304 28080 42316
rect 28132 42304 28138 42356
rect 22066 42248 24420 42276
rect 25406 42236 25412 42288
rect 25464 42276 25470 42288
rect 25501 42279 25559 42285
rect 25501 42276 25513 42279
rect 25464 42248 25513 42276
rect 25464 42236 25470 42248
rect 25501 42245 25513 42248
rect 25547 42245 25559 42279
rect 25501 42239 25559 42245
rect 18693 42211 18751 42217
rect 18693 42208 18705 42211
rect 16776 42180 18705 42208
rect 18693 42177 18705 42180
rect 18739 42208 18751 42211
rect 18782 42208 18788 42220
rect 18739 42180 18788 42208
rect 18739 42177 18751 42180
rect 18693 42171 18751 42177
rect 18782 42168 18788 42180
rect 18840 42168 18846 42220
rect 22370 42208 22376 42220
rect 22112 42180 22376 42208
rect 22112 42149 22140 42180
rect 22370 42168 22376 42180
rect 22428 42208 22434 42220
rect 23014 42208 23020 42220
rect 22428 42180 23020 42208
rect 22428 42168 22434 42180
rect 23014 42168 23020 42180
rect 23072 42208 23078 42220
rect 23477 42211 23535 42217
rect 23072 42180 23428 42208
rect 23072 42168 23078 42180
rect 15105 42143 15163 42149
rect 15105 42140 15117 42143
rect 12400 42112 15117 42140
rect 12400 42100 12406 42112
rect 15105 42109 15117 42112
rect 15151 42109 15163 42143
rect 22097 42143 22155 42149
rect 15105 42103 15163 42109
rect 15948 42112 18000 42140
rect 1486 42032 1492 42084
rect 1544 42072 1550 42084
rect 1642 42075 1700 42081
rect 1642 42072 1654 42075
rect 1544 42044 1654 42072
rect 1544 42032 1550 42044
rect 1642 42041 1654 42044
rect 1688 42041 1700 42075
rect 1642 42035 1700 42041
rect 2682 42032 2688 42084
rect 2740 42072 2746 42084
rect 2740 42044 9904 42072
rect 2740 42032 2746 42044
rect 4982 42004 4988 42016
rect 4943 41976 4988 42004
rect 4982 41964 4988 41976
rect 5040 41964 5046 42016
rect 9766 42004 9772 42016
rect 9727 41976 9772 42004
rect 9766 41964 9772 41976
rect 9824 41964 9830 42016
rect 9876 42004 9904 42044
rect 12434 42032 12440 42084
rect 12492 42081 12498 42084
rect 12492 42075 12556 42081
rect 12492 42041 12510 42075
rect 12544 42041 12556 42075
rect 12492 42035 12556 42041
rect 12492 42032 12498 42035
rect 14274 42032 14280 42084
rect 14332 42072 14338 42084
rect 14550 42072 14556 42084
rect 14332 42044 14556 42072
rect 14332 42032 14338 42044
rect 14550 42032 14556 42044
rect 14608 42072 14614 42084
rect 14921 42075 14979 42081
rect 14921 42072 14933 42075
rect 14608 42044 14933 42072
rect 14608 42032 14614 42044
rect 14921 42041 14933 42044
rect 14967 42041 14979 42075
rect 14921 42035 14979 42041
rect 15948 42004 15976 42112
rect 16040 42044 16988 42072
rect 16040 42013 16068 42044
rect 9876 41976 15976 42004
rect 16025 42007 16083 42013
rect 16025 41973 16037 42007
rect 16071 41973 16083 42007
rect 16390 42004 16396 42016
rect 16351 41976 16396 42004
rect 16025 41967 16083 41973
rect 16390 41964 16396 41976
rect 16448 41964 16454 42016
rect 16485 42007 16543 42013
rect 16485 41973 16497 42007
rect 16531 42004 16543 42007
rect 16574 42004 16580 42016
rect 16531 41976 16580 42004
rect 16531 41973 16543 41976
rect 16485 41967 16543 41973
rect 16574 41964 16580 41976
rect 16632 41964 16638 42016
rect 16960 42004 16988 42044
rect 17494 42032 17500 42084
rect 17552 42072 17558 42084
rect 17589 42075 17647 42081
rect 17589 42072 17601 42075
rect 17552 42044 17601 42072
rect 17552 42032 17558 42044
rect 17589 42041 17601 42044
rect 17635 42041 17647 42075
rect 17862 42072 17868 42084
rect 17823 42044 17868 42072
rect 17589 42035 17647 42041
rect 17862 42032 17868 42044
rect 17920 42032 17926 42084
rect 17773 42007 17831 42013
rect 17773 42004 17785 42007
rect 16960 41976 17785 42004
rect 17773 41973 17785 41976
rect 17819 41973 17831 42007
rect 17972 42004 18000 42112
rect 22097 42109 22109 42143
rect 22143 42109 22155 42143
rect 22097 42103 22155 42109
rect 22186 42100 22192 42152
rect 22244 42140 22250 42152
rect 22281 42143 22339 42149
rect 22281 42140 22293 42143
rect 22244 42112 22293 42140
rect 22244 42100 22250 42112
rect 22281 42109 22293 42112
rect 22327 42140 22339 42143
rect 22738 42140 22744 42152
rect 22327 42112 22744 42140
rect 22327 42109 22339 42112
rect 22281 42103 22339 42109
rect 22738 42100 22744 42112
rect 22796 42100 22802 42152
rect 23124 42149 23152 42180
rect 23109 42143 23167 42149
rect 23109 42109 23121 42143
rect 23155 42109 23167 42143
rect 23290 42140 23296 42152
rect 23251 42112 23296 42140
rect 23109 42103 23167 42109
rect 23290 42100 23296 42112
rect 23348 42100 23354 42152
rect 23400 42140 23428 42180
rect 23477 42177 23489 42211
rect 23523 42208 23535 42211
rect 23842 42208 23848 42220
rect 23523 42180 23848 42208
rect 23523 42177 23535 42180
rect 23477 42171 23535 42177
rect 23842 42168 23848 42180
rect 23900 42208 23906 42220
rect 23900 42180 25268 42208
rect 23900 42168 23906 42180
rect 25240 42149 25268 42180
rect 25590 42168 25596 42220
rect 25648 42208 25654 42220
rect 26053 42211 26111 42217
rect 26053 42208 26065 42211
rect 25648 42180 26065 42208
rect 25648 42168 25654 42180
rect 26053 42177 26065 42180
rect 26099 42177 26111 42211
rect 26053 42171 26111 42177
rect 23937 42143 23995 42149
rect 23937 42140 23949 42143
rect 23400 42112 23949 42140
rect 23937 42109 23949 42112
rect 23983 42109 23995 42143
rect 23937 42103 23995 42109
rect 24121 42143 24179 42149
rect 24121 42109 24133 42143
rect 24167 42109 24179 42143
rect 24121 42103 24179 42109
rect 25225 42143 25283 42149
rect 25225 42109 25237 42143
rect 25271 42109 25283 42143
rect 25406 42140 25412 42152
rect 25367 42112 25412 42140
rect 25225 42103 25283 42109
rect 18414 42032 18420 42084
rect 18472 42072 18478 42084
rect 18509 42075 18567 42081
rect 18509 42072 18521 42075
rect 18472 42044 18521 42072
rect 18472 42032 18478 42044
rect 18509 42041 18521 42044
rect 18555 42041 18567 42075
rect 23308 42072 23336 42100
rect 24136 42072 24164 42103
rect 25406 42100 25412 42112
rect 25464 42100 25470 42152
rect 26602 42140 26608 42152
rect 26160 42112 26608 42140
rect 26160 42072 26188 42112
rect 26602 42100 26608 42112
rect 26660 42100 26666 42152
rect 27430 42100 27436 42152
rect 27488 42140 27494 42152
rect 28169 42143 28227 42149
rect 28169 42140 28181 42143
rect 27488 42112 28181 42140
rect 27488 42100 27494 42112
rect 28169 42109 28181 42112
rect 28215 42109 28227 42143
rect 28169 42103 28227 42109
rect 26326 42081 26332 42084
rect 23308 42044 24164 42072
rect 24412 42044 26188 42072
rect 18509 42035 18567 42041
rect 24412 42004 24440 42044
rect 26320 42035 26332 42081
rect 26384 42072 26390 42084
rect 26384 42044 26420 42072
rect 26326 42032 26332 42035
rect 26384 42032 26390 42044
rect 17972 41976 24440 42004
rect 17773 41967 17831 41973
rect 25590 41964 25596 42016
rect 25648 42004 25654 42016
rect 27433 42007 27491 42013
rect 27433 42004 27445 42007
rect 25648 41976 27445 42004
rect 25648 41964 25654 41976
rect 27433 41973 27445 41976
rect 27479 41973 27491 42007
rect 27433 41967 27491 41973
rect 27890 41964 27896 42016
rect 27948 42004 27954 42016
rect 27985 42007 28043 42013
rect 27985 42004 27997 42007
rect 27948 41976 27997 42004
rect 27948 41964 27954 41976
rect 27985 41973 27997 41976
rect 28031 41973 28043 42007
rect 27985 41967 28043 41973
rect 1104 41914 28888 41936
rect 1104 41862 10246 41914
rect 10298 41862 10310 41914
rect 10362 41862 10374 41914
rect 10426 41862 10438 41914
rect 10490 41862 19510 41914
rect 19562 41862 19574 41914
rect 19626 41862 19638 41914
rect 19690 41862 19702 41914
rect 19754 41862 28888 41914
rect 1104 41840 28888 41862
rect 1486 41800 1492 41812
rect 1447 41772 1492 41800
rect 1486 41760 1492 41772
rect 1544 41760 1550 41812
rect 1857 41803 1915 41809
rect 1857 41769 1869 41803
rect 1903 41800 1915 41803
rect 2866 41800 2872 41812
rect 1903 41772 2872 41800
rect 1903 41769 1915 41772
rect 1857 41763 1915 41769
rect 2866 41760 2872 41772
rect 2924 41760 2930 41812
rect 4246 41760 4252 41812
rect 4304 41800 4310 41812
rect 5350 41800 5356 41812
rect 4304 41772 5356 41800
rect 4304 41760 4310 41772
rect 5350 41760 5356 41772
rect 5408 41760 5414 41812
rect 7650 41800 7656 41812
rect 7611 41772 7656 41800
rect 7650 41760 7656 41772
rect 7708 41760 7714 41812
rect 8754 41800 8760 41812
rect 8715 41772 8760 41800
rect 8754 41760 8760 41772
rect 8812 41760 8818 41812
rect 9493 41803 9551 41809
rect 9493 41769 9505 41803
rect 9539 41800 9551 41803
rect 9674 41800 9680 41812
rect 9539 41772 9680 41800
rect 9539 41769 9551 41772
rect 9493 41763 9551 41769
rect 9674 41760 9680 41772
rect 9732 41760 9738 41812
rect 10134 41760 10140 41812
rect 10192 41800 10198 41812
rect 10321 41803 10379 41809
rect 10321 41800 10333 41803
rect 10192 41772 10333 41800
rect 10192 41760 10198 41772
rect 10321 41769 10333 41772
rect 10367 41769 10379 41803
rect 17494 41800 17500 41812
rect 10321 41763 10379 41769
rect 12406 41772 15700 41800
rect 17455 41772 17500 41800
rect 2498 41692 2504 41744
rect 2556 41732 2562 41744
rect 12406 41732 12434 41772
rect 13170 41732 13176 41744
rect 2556 41704 12434 41732
rect 13131 41704 13176 41732
rect 2556 41692 2562 41704
rect 13170 41692 13176 41704
rect 13228 41692 13234 41744
rect 15672 41732 15700 41772
rect 17494 41760 17500 41772
rect 17552 41760 17558 41812
rect 19334 41760 19340 41812
rect 19392 41800 19398 41812
rect 19521 41803 19579 41809
rect 19521 41800 19533 41803
rect 19392 41772 19533 41800
rect 19392 41760 19398 41772
rect 19521 41769 19533 41772
rect 19567 41769 19579 41803
rect 19521 41763 19579 41769
rect 19613 41803 19671 41809
rect 19613 41769 19625 41803
rect 19659 41800 19671 41803
rect 19794 41800 19800 41812
rect 19659 41772 19800 41800
rect 19659 41769 19671 41772
rect 19613 41763 19671 41769
rect 19794 41760 19800 41772
rect 19852 41760 19858 41812
rect 26326 41800 26332 41812
rect 26287 41772 26332 41800
rect 26326 41760 26332 41772
rect 26384 41760 26390 41812
rect 28169 41735 28227 41741
rect 28169 41732 28181 41735
rect 13464 41704 14044 41732
rect 15672 41704 28181 41732
rect 2869 41667 2927 41673
rect 2869 41633 2881 41667
rect 2915 41664 2927 41667
rect 3050 41664 3056 41676
rect 2915 41636 3056 41664
rect 2915 41633 2927 41636
rect 2869 41627 2927 41633
rect 3050 41624 3056 41636
rect 3108 41664 3114 41676
rect 3694 41664 3700 41676
rect 3108 41636 3700 41664
rect 3108 41624 3114 41636
rect 3694 41624 3700 41636
rect 3752 41624 3758 41676
rect 7561 41667 7619 41673
rect 7561 41633 7573 41667
rect 7607 41664 7619 41667
rect 8110 41664 8116 41676
rect 7607 41636 8116 41664
rect 7607 41633 7619 41636
rect 7561 41627 7619 41633
rect 8110 41624 8116 41636
rect 8168 41624 8174 41676
rect 8478 41624 8484 41676
rect 8536 41664 8542 41676
rect 8846 41664 8852 41676
rect 8536 41636 8852 41664
rect 8536 41624 8542 41636
rect 8846 41624 8852 41636
rect 8904 41624 8910 41676
rect 9306 41664 9312 41676
rect 9267 41636 9312 41664
rect 9306 41624 9312 41636
rect 9364 41624 9370 41676
rect 9582 41664 9588 41676
rect 9543 41636 9588 41664
rect 9582 41624 9588 41636
rect 9640 41624 9646 41676
rect 9769 41667 9827 41673
rect 9769 41633 9781 41667
rect 9815 41633 9827 41667
rect 9769 41627 9827 41633
rect 1949 41599 2007 41605
rect 1949 41565 1961 41599
rect 1995 41565 2007 41599
rect 1949 41559 2007 41565
rect 2133 41599 2191 41605
rect 2133 41565 2145 41599
rect 2179 41596 2191 41599
rect 2314 41596 2320 41608
rect 2179 41568 2320 41596
rect 2179 41565 2191 41568
rect 2133 41559 2191 41565
rect 1964 41460 1992 41559
rect 2314 41556 2320 41568
rect 2372 41556 2378 41608
rect 2961 41599 3019 41605
rect 2961 41565 2973 41599
rect 3007 41596 3019 41599
rect 3142 41596 3148 41608
rect 3007 41568 3148 41596
rect 3007 41565 3019 41568
rect 2961 41559 3019 41565
rect 3142 41556 3148 41568
rect 3200 41596 3206 41608
rect 3786 41596 3792 41608
rect 3200 41568 3792 41596
rect 3200 41556 3206 41568
rect 3786 41556 3792 41568
rect 3844 41556 3850 41608
rect 4614 41596 4620 41608
rect 4575 41568 4620 41596
rect 4614 41556 4620 41568
rect 4672 41556 4678 41608
rect 6178 41596 6184 41608
rect 4724 41568 6184 41596
rect 3237 41531 3295 41537
rect 3237 41497 3249 41531
rect 3283 41528 3295 41531
rect 3510 41528 3516 41540
rect 3283 41500 3516 41528
rect 3283 41497 3295 41500
rect 3237 41491 3295 41497
rect 3510 41488 3516 41500
rect 3568 41488 3574 41540
rect 3804 41528 3832 41556
rect 3973 41531 4031 41537
rect 3973 41528 3985 41531
rect 3804 41500 3985 41528
rect 3973 41497 3985 41500
rect 4019 41497 4031 41531
rect 4724 41528 4752 41568
rect 6178 41556 6184 41568
rect 6236 41556 6242 41608
rect 7098 41556 7104 41608
rect 7156 41596 7162 41608
rect 7745 41599 7803 41605
rect 7745 41596 7757 41599
rect 7156 41568 7757 41596
rect 7156 41556 7162 41568
rect 7745 41565 7757 41568
rect 7791 41565 7803 41599
rect 7745 41559 7803 41565
rect 8294 41556 8300 41608
rect 8352 41596 8358 41608
rect 8389 41599 8447 41605
rect 8389 41596 8401 41599
rect 8352 41568 8401 41596
rect 8352 41556 8358 41568
rect 8389 41565 8401 41568
rect 8435 41565 8447 41599
rect 8389 41559 8447 41565
rect 8573 41599 8631 41605
rect 8573 41565 8585 41599
rect 8619 41596 8631 41599
rect 9784 41596 9812 41627
rect 9858 41624 9864 41676
rect 9916 41664 9922 41676
rect 10134 41664 10140 41676
rect 9916 41636 10140 41664
rect 9916 41624 9922 41636
rect 10134 41624 10140 41636
rect 10192 41624 10198 41676
rect 10229 41667 10287 41673
rect 10229 41633 10241 41667
rect 10275 41633 10287 41667
rect 10229 41627 10287 41633
rect 10244 41596 10272 41627
rect 12526 41624 12532 41676
rect 12584 41664 12590 41676
rect 13464 41664 13492 41704
rect 12584 41636 13492 41664
rect 12584 41624 12590 41636
rect 13630 41624 13636 41676
rect 13688 41664 13694 41676
rect 14016 41673 14044 41704
rect 28169 41701 28181 41704
rect 28215 41701 28227 41735
rect 28169 41695 28227 41701
rect 13817 41667 13875 41673
rect 13817 41664 13829 41667
rect 13688 41636 13829 41664
rect 13688 41624 13694 41636
rect 13817 41633 13829 41636
rect 13863 41633 13875 41667
rect 13817 41627 13875 41633
rect 14001 41667 14059 41673
rect 14001 41633 14013 41667
rect 14047 41633 14059 41667
rect 14001 41627 14059 41633
rect 8619 41568 9812 41596
rect 9876 41568 10272 41596
rect 13173 41599 13231 41605
rect 8619 41565 8631 41568
rect 8573 41559 8631 41565
rect 9876 41540 9904 41568
rect 13173 41565 13185 41599
rect 13219 41565 13231 41599
rect 13173 41559 13231 41565
rect 13265 41599 13323 41605
rect 13265 41565 13277 41599
rect 13311 41596 13323 41599
rect 13538 41596 13544 41608
rect 13311 41568 13544 41596
rect 13311 41565 13323 41568
rect 13265 41559 13323 41565
rect 4890 41528 4896 41540
rect 3973 41491 4031 41497
rect 4080 41500 4752 41528
rect 4851 41500 4896 41528
rect 4080 41460 4108 41500
rect 4890 41488 4896 41500
rect 4948 41488 4954 41540
rect 9858 41488 9864 41540
rect 9916 41488 9922 41540
rect 13188 41528 13216 41559
rect 13538 41556 13544 41568
rect 13596 41556 13602 41608
rect 14016 41596 14044 41627
rect 16114 41624 16120 41676
rect 16172 41664 16178 41676
rect 16666 41664 16672 41676
rect 16172 41636 16672 41664
rect 16172 41624 16178 41636
rect 16666 41624 16672 41636
rect 16724 41664 16730 41676
rect 17313 41667 17371 41673
rect 17313 41664 17325 41667
rect 16724 41636 17325 41664
rect 16724 41624 16730 41636
rect 17313 41633 17325 41636
rect 17359 41633 17371 41667
rect 17313 41627 17371 41633
rect 17497 41667 17555 41673
rect 17497 41633 17509 41667
rect 17543 41633 17555 41667
rect 21450 41664 21456 41676
rect 21411 41636 21456 41664
rect 17497 41627 17555 41633
rect 17512 41596 17540 41627
rect 21450 41624 21456 41636
rect 21508 41624 21514 41676
rect 23658 41624 23664 41676
rect 23716 41664 23722 41676
rect 24029 41667 24087 41673
rect 24029 41664 24041 41667
rect 23716 41636 24041 41664
rect 23716 41624 23722 41636
rect 24029 41633 24041 41636
rect 24075 41633 24087 41667
rect 24029 41627 24087 41633
rect 24118 41624 24124 41676
rect 24176 41664 24182 41676
rect 24213 41667 24271 41673
rect 24213 41664 24225 41667
rect 24176 41636 24225 41664
rect 24176 41624 24182 41636
rect 24213 41633 24225 41636
rect 24259 41633 24271 41667
rect 24486 41664 24492 41676
rect 24447 41636 24492 41664
rect 24213 41627 24271 41633
rect 24486 41624 24492 41636
rect 24544 41664 24550 41676
rect 25317 41667 25375 41673
rect 25317 41664 25329 41667
rect 24544 41636 25329 41664
rect 24544 41624 24550 41636
rect 25317 41633 25329 41636
rect 25363 41633 25375 41667
rect 26421 41667 26479 41673
rect 26421 41664 26433 41667
rect 25317 41627 25375 41633
rect 25700 41636 26433 41664
rect 18046 41596 18052 41608
rect 14016 41568 18052 41596
rect 18046 41556 18052 41568
rect 18104 41556 18110 41608
rect 19334 41556 19340 41608
rect 19392 41596 19398 41608
rect 19705 41599 19763 41605
rect 19705 41596 19717 41599
rect 19392 41568 19717 41596
rect 19392 41556 19398 41568
rect 19705 41565 19717 41568
rect 19751 41565 19763 41599
rect 25222 41596 25228 41608
rect 25183 41568 25228 41596
rect 19705 41559 19763 41565
rect 25222 41556 25228 41568
rect 25280 41556 25286 41608
rect 25700 41605 25728 41636
rect 26421 41633 26433 41636
rect 26467 41633 26479 41667
rect 26421 41627 26479 41633
rect 26605 41667 26663 41673
rect 26605 41633 26617 41667
rect 26651 41633 26663 41667
rect 26605 41627 26663 41633
rect 25685 41599 25743 41605
rect 25685 41565 25697 41599
rect 25731 41565 25743 41599
rect 26142 41596 26148 41608
rect 26103 41568 26148 41596
rect 25685 41559 25743 41565
rect 26142 41556 26148 41568
rect 26200 41556 26206 41608
rect 13909 41531 13967 41537
rect 13909 41528 13921 41531
rect 13188 41500 13921 41528
rect 13909 41497 13921 41500
rect 13955 41497 13967 41531
rect 13909 41491 13967 41497
rect 16390 41488 16396 41540
rect 16448 41488 16454 41540
rect 23934 41488 23940 41540
rect 23992 41528 23998 41540
rect 24121 41531 24179 41537
rect 24121 41528 24133 41531
rect 23992 41500 24133 41528
rect 23992 41488 23998 41500
rect 24121 41497 24133 41500
rect 24167 41497 24179 41531
rect 24121 41491 24179 41497
rect 25958 41488 25964 41540
rect 26016 41528 26022 41540
rect 26620 41528 26648 41627
rect 27062 41624 27068 41676
rect 27120 41664 27126 41676
rect 27985 41667 28043 41673
rect 27985 41664 27997 41667
rect 27120 41636 27997 41664
rect 27120 41624 27126 41636
rect 27985 41633 27997 41636
rect 28031 41633 28043 41667
rect 27985 41627 28043 41633
rect 26016 41500 26648 41528
rect 26016 41488 26022 41500
rect 1964 41432 4108 41460
rect 4157 41463 4215 41469
rect 4157 41429 4169 41463
rect 4203 41460 4215 41463
rect 4246 41460 4252 41472
rect 4203 41432 4252 41460
rect 4203 41429 4215 41432
rect 4157 41423 4215 41429
rect 4246 41420 4252 41432
rect 4304 41420 4310 41472
rect 5077 41463 5135 41469
rect 5077 41429 5089 41463
rect 5123 41460 5135 41463
rect 5902 41460 5908 41472
rect 5123 41432 5908 41460
rect 5123 41429 5135 41432
rect 5077 41423 5135 41429
rect 5902 41420 5908 41432
rect 5960 41420 5966 41472
rect 7190 41460 7196 41472
rect 7151 41432 7196 41460
rect 7190 41420 7196 41432
rect 7248 41420 7254 41472
rect 9490 41420 9496 41472
rect 9548 41460 9554 41472
rect 12713 41463 12771 41469
rect 12713 41460 12725 41463
rect 9548 41432 12725 41460
rect 9548 41420 9554 41432
rect 12713 41429 12725 41432
rect 12759 41460 12771 41463
rect 14642 41460 14648 41472
rect 12759 41432 14648 41460
rect 12759 41429 12771 41432
rect 12713 41423 12771 41429
rect 14642 41420 14648 41432
rect 14700 41460 14706 41472
rect 16408 41460 16436 41488
rect 14700 41432 16436 41460
rect 14700 41420 14706 41432
rect 18874 41420 18880 41472
rect 18932 41460 18938 41472
rect 19153 41463 19211 41469
rect 19153 41460 19165 41463
rect 18932 41432 19165 41460
rect 18932 41420 18938 41432
rect 19153 41429 19165 41432
rect 19199 41429 19211 41463
rect 19153 41423 19211 41429
rect 21082 41420 21088 41472
rect 21140 41460 21146 41472
rect 21545 41463 21603 41469
rect 21545 41460 21557 41463
rect 21140 41432 21557 41460
rect 21140 41420 21146 41432
rect 21545 41429 21557 41432
rect 21591 41429 21603 41463
rect 21545 41423 21603 41429
rect 1104 41370 28888 41392
rect 1104 41318 5614 41370
rect 5666 41318 5678 41370
rect 5730 41318 5742 41370
rect 5794 41318 5806 41370
rect 5858 41318 14878 41370
rect 14930 41318 14942 41370
rect 14994 41318 15006 41370
rect 15058 41318 15070 41370
rect 15122 41318 24142 41370
rect 24194 41318 24206 41370
rect 24258 41318 24270 41370
rect 24322 41318 24334 41370
rect 24386 41318 28888 41370
rect 1104 41296 28888 41318
rect 2406 41216 2412 41268
rect 2464 41256 2470 41268
rect 8110 41256 8116 41268
rect 2464 41228 7604 41256
rect 8071 41228 8116 41256
rect 2464 41216 2470 41228
rect 1486 41148 1492 41200
rect 1544 41188 1550 41200
rect 1857 41191 1915 41197
rect 1857 41188 1869 41191
rect 1544 41160 1869 41188
rect 1544 41148 1550 41160
rect 1857 41157 1869 41160
rect 1903 41157 1915 41191
rect 1857 41151 1915 41157
rect 6365 41191 6423 41197
rect 6365 41157 6377 41191
rect 6411 41157 6423 41191
rect 6365 41151 6423 41157
rect 3970 41080 3976 41132
rect 4028 41120 4034 41132
rect 4028 41092 5028 41120
rect 4028 41080 4034 41092
rect 4246 41052 4252 41064
rect 4207 41024 4252 41052
rect 4246 41012 4252 41024
rect 4304 41012 4310 41064
rect 5000 41061 5028 41092
rect 4985 41055 5043 41061
rect 4985 41021 4997 41055
rect 5031 41052 5043 41055
rect 5534 41052 5540 41064
rect 5031 41024 5540 41052
rect 5031 41021 5043 41024
rect 4985 41015 5043 41021
rect 5534 41012 5540 41024
rect 5592 41012 5598 41064
rect 6380 41052 6408 41151
rect 6638 41148 6644 41200
rect 6696 41188 6702 41200
rect 6825 41191 6883 41197
rect 6825 41188 6837 41191
rect 6696 41160 6837 41188
rect 6696 41148 6702 41160
rect 6825 41157 6837 41160
rect 6871 41157 6883 41191
rect 7576 41188 7604 41228
rect 8110 41216 8116 41228
rect 8168 41216 8174 41268
rect 25225 41259 25283 41265
rect 25225 41256 25237 41259
rect 8220 41228 25237 41256
rect 8220 41188 8248 41228
rect 25225 41225 25237 41228
rect 25271 41225 25283 41259
rect 25225 41219 25283 41225
rect 25317 41259 25375 41265
rect 25317 41225 25329 41259
rect 25363 41256 25375 41259
rect 27062 41256 27068 41268
rect 25363 41228 27068 41256
rect 25363 41225 25375 41228
rect 25317 41219 25375 41225
rect 27062 41216 27068 41228
rect 27120 41216 27126 41268
rect 13446 41188 13452 41200
rect 7576 41160 8248 41188
rect 13096 41160 13452 41188
rect 6825 41151 6883 41157
rect 7374 41120 7380 41132
rect 7335 41092 7380 41120
rect 7374 41080 7380 41092
rect 7432 41080 7438 41132
rect 9214 41080 9220 41132
rect 9272 41120 9278 41132
rect 9493 41123 9551 41129
rect 9493 41120 9505 41123
rect 9272 41092 9505 41120
rect 9272 41080 9278 41092
rect 9493 41089 9505 41092
rect 9539 41089 9551 41123
rect 9493 41083 9551 41089
rect 9766 41061 9772 41064
rect 7193 41055 7251 41061
rect 7193 41052 7205 41055
rect 6380 41024 7205 41052
rect 7193 41021 7205 41024
rect 7239 41052 7251 41055
rect 8021 41055 8079 41061
rect 8021 41052 8033 41055
rect 7239 41024 8033 41052
rect 7239 41021 7251 41024
rect 7193 41015 7251 41021
rect 8021 41021 8033 41024
rect 8067 41021 8079 41055
rect 8021 41015 8079 41021
rect 9760 41015 9772 41061
rect 9824 41052 9830 41064
rect 9824 41024 9860 41052
rect 9766 41012 9772 41015
rect 9824 41012 9830 41024
rect 12802 41012 12808 41064
rect 12860 41052 12866 41064
rect 13096 41061 13124 41160
rect 13446 41148 13452 41160
rect 13504 41148 13510 41200
rect 24121 41191 24179 41197
rect 24121 41157 24133 41191
rect 24167 41188 24179 41191
rect 25406 41188 25412 41200
rect 24167 41160 25412 41188
rect 24167 41157 24179 41160
rect 24121 41151 24179 41157
rect 25406 41148 25412 41160
rect 25464 41148 25470 41200
rect 27525 41191 27583 41197
rect 27525 41157 27537 41191
rect 27571 41157 27583 41191
rect 27525 41151 27583 41157
rect 13630 41120 13636 41132
rect 12897 41055 12955 41061
rect 12897 41052 12909 41055
rect 12860 41024 12909 41052
rect 12860 41012 12866 41024
rect 12897 41021 12909 41024
rect 12943 41021 12955 41055
rect 12897 41015 12955 41021
rect 13045 41055 13124 41061
rect 13045 41021 13057 41055
rect 13091 41024 13124 41055
rect 13280 41092 13636 41120
rect 13280 41052 13308 41092
rect 13630 41080 13636 41092
rect 13688 41080 13694 41132
rect 15194 41080 15200 41132
rect 15252 41120 15258 41132
rect 15749 41123 15807 41129
rect 15749 41120 15761 41123
rect 15252 41092 15761 41120
rect 15252 41080 15258 41092
rect 15749 41089 15761 41092
rect 15795 41089 15807 41123
rect 15749 41083 15807 41089
rect 16114 41080 16120 41132
rect 16172 41120 16178 41132
rect 16482 41120 16488 41132
rect 16172 41092 16488 41120
rect 16172 41080 16178 41092
rect 16482 41080 16488 41092
rect 16540 41120 16546 41132
rect 16540 41092 17724 41120
rect 16540 41080 16546 41092
rect 13188 41024 13308 41052
rect 13403 41055 13461 41061
rect 13091 41021 13103 41024
rect 13045 41015 13103 41021
rect 2130 40984 2136 40996
rect 2091 40956 2136 40984
rect 2130 40944 2136 40956
rect 2188 40944 2194 40996
rect 2222 40944 2228 40996
rect 2280 40984 2286 40996
rect 2409 40987 2467 40993
rect 2409 40984 2421 40987
rect 2280 40956 2421 40984
rect 2280 40944 2286 40956
rect 2409 40953 2421 40956
rect 2455 40953 2467 40987
rect 3050 40984 3056 40996
rect 3011 40956 3056 40984
rect 2409 40947 2467 40953
rect 3050 40944 3056 40956
rect 3108 40944 3114 40996
rect 5252 40987 5310 40993
rect 5252 40953 5264 40987
rect 5298 40984 5310 40987
rect 6638 40984 6644 40996
rect 5298 40956 6644 40984
rect 5298 40953 5310 40956
rect 5252 40947 5310 40953
rect 6638 40944 6644 40956
rect 6696 40944 6702 40996
rect 7834 40944 7840 40996
rect 7892 40984 7898 40996
rect 7892 40956 12434 40984
rect 7892 40944 7898 40956
rect 2317 40919 2375 40925
rect 2317 40885 2329 40919
rect 2363 40916 2375 40919
rect 2498 40916 2504 40928
rect 2363 40888 2504 40916
rect 2363 40885 2375 40888
rect 2317 40879 2375 40885
rect 2498 40876 2504 40888
rect 2556 40876 2562 40928
rect 3142 40916 3148 40928
rect 3103 40888 3148 40916
rect 3142 40876 3148 40888
rect 3200 40876 3206 40928
rect 4338 40916 4344 40928
rect 4299 40888 4344 40916
rect 4338 40876 4344 40888
rect 4396 40876 4402 40928
rect 7098 40876 7104 40928
rect 7156 40916 7162 40928
rect 7285 40919 7343 40925
rect 7285 40916 7297 40919
rect 7156 40888 7297 40916
rect 7156 40876 7162 40888
rect 7285 40885 7297 40888
rect 7331 40885 7343 40919
rect 7285 40879 7343 40885
rect 9858 40876 9864 40928
rect 9916 40916 9922 40928
rect 10873 40919 10931 40925
rect 10873 40916 10885 40919
rect 9916 40888 10885 40916
rect 9916 40876 9922 40888
rect 10873 40885 10885 40888
rect 10919 40885 10931 40919
rect 12406 40916 12434 40956
rect 12710 40944 12716 40996
rect 12768 40984 12774 40996
rect 13188 40993 13216 41024
rect 13403 41021 13415 41055
rect 13449 41052 13461 41055
rect 14642 41052 14648 41064
rect 13449 41024 14648 41052
rect 13449 41021 13461 41024
rect 13403 41015 13461 41021
rect 14642 41012 14648 41024
rect 14700 41012 14706 41064
rect 15378 41012 15384 41064
rect 15436 41052 15442 41064
rect 15473 41055 15531 41061
rect 15473 41052 15485 41055
rect 15436 41024 15485 41052
rect 15436 41012 15442 41024
rect 15473 41021 15485 41024
rect 15519 41052 15531 41055
rect 17589 41055 17647 41061
rect 17589 41052 17601 41055
rect 15519 41024 17601 41052
rect 15519 41021 15531 41024
rect 15473 41015 15531 41021
rect 17589 41021 17601 41024
rect 17635 41021 17647 41055
rect 17696 41052 17724 41092
rect 20990 41080 20996 41132
rect 21048 41120 21054 41132
rect 21085 41123 21143 41129
rect 21085 41120 21097 41123
rect 21048 41092 21097 41120
rect 21048 41080 21054 41092
rect 21085 41089 21097 41092
rect 21131 41089 21143 41123
rect 23290 41120 23296 41132
rect 23251 41092 23296 41120
rect 21085 41083 21143 41089
rect 23290 41080 23296 41092
rect 23348 41080 23354 41132
rect 23658 41080 23664 41132
rect 23716 41080 23722 41132
rect 25225 41123 25283 41129
rect 25225 41089 25237 41123
rect 25271 41120 25283 41123
rect 27540 41120 27568 41151
rect 25271 41092 27568 41120
rect 25271 41089 25283 41092
rect 25225 41083 25283 41089
rect 22005 41055 22063 41061
rect 17696 41024 19012 41052
rect 17589 41015 17647 41021
rect 13173 40987 13231 40993
rect 13173 40984 13185 40987
rect 12768 40956 13185 40984
rect 12768 40944 12774 40956
rect 13173 40953 13185 40956
rect 13219 40953 13231 40987
rect 13173 40947 13231 40953
rect 13262 40944 13268 40996
rect 13320 40984 13326 40996
rect 13320 40956 13365 40984
rect 13320 40944 13326 40956
rect 16758 40944 16764 40996
rect 16816 40984 16822 40996
rect 17834 40987 17892 40993
rect 17834 40984 17846 40987
rect 16816 40956 17846 40984
rect 16816 40944 16822 40956
rect 17834 40953 17846 40956
rect 17880 40953 17892 40987
rect 17834 40947 17892 40953
rect 13541 40919 13599 40925
rect 13541 40916 13553 40919
rect 12406 40888 13553 40916
rect 10873 40879 10931 40885
rect 13541 40885 13553 40888
rect 13587 40885 13599 40919
rect 17034 40916 17040 40928
rect 16995 40888 17040 40916
rect 13541 40879 13599 40885
rect 17034 40876 17040 40888
rect 17092 40876 17098 40928
rect 18984 40925 19012 41024
rect 22005 41021 22017 41055
rect 22051 41021 22063 41055
rect 22186 41052 22192 41064
rect 22147 41024 22192 41052
rect 22005 41015 22063 41021
rect 20993 40987 21051 40993
rect 20993 40953 21005 40987
rect 21039 40984 21051 40987
rect 22020 40984 22048 41015
rect 22186 41012 22192 41024
rect 22244 41012 22250 41064
rect 23014 41012 23020 41064
rect 23072 41052 23078 41064
rect 23109 41055 23167 41061
rect 23109 41052 23121 41055
rect 23072 41024 23121 41052
rect 23072 41012 23078 41024
rect 23109 41021 23121 41024
rect 23155 41021 23167 41055
rect 23842 41052 23848 41064
rect 23803 41024 23848 41052
rect 23109 41015 23167 41021
rect 23842 41012 23848 41024
rect 23900 41012 23906 41064
rect 24946 41012 24952 41064
rect 25004 41052 25010 41064
rect 25314 41052 25320 41064
rect 25004 41024 25320 41052
rect 25004 41012 25010 41024
rect 25314 41012 25320 41024
rect 25372 41012 25378 41064
rect 25498 41052 25504 41064
rect 25459 41024 25504 41052
rect 25498 41012 25504 41024
rect 25556 41012 25562 41064
rect 26142 41052 26148 41064
rect 26103 41024 26148 41052
rect 26142 41012 26148 41024
rect 26200 41012 26206 41064
rect 26786 41052 26792 41064
rect 26747 41024 26792 41052
rect 26786 41012 26792 41024
rect 26844 41012 26850 41064
rect 27522 41012 27528 41064
rect 27580 41052 27586 41064
rect 28169 41055 28227 41061
rect 28169 41052 28181 41055
rect 27580 41024 28181 41052
rect 27580 41012 27586 41024
rect 28169 41021 28181 41024
rect 28215 41021 28227 41055
rect 28169 41015 28227 41021
rect 23658 40984 23664 40996
rect 21039 40956 23664 40984
rect 21039 40953 21051 40956
rect 20993 40947 21051 40953
rect 23658 40944 23664 40956
rect 23716 40944 23722 40996
rect 27341 40987 27399 40993
rect 27341 40984 27353 40987
rect 25976 40956 27353 40984
rect 18969 40919 19027 40925
rect 18969 40885 18981 40919
rect 19015 40885 19027 40919
rect 20530 40916 20536 40928
rect 20491 40888 20536 40916
rect 18969 40879 19027 40885
rect 20530 40876 20536 40888
rect 20588 40876 20594 40928
rect 20901 40919 20959 40925
rect 20901 40885 20913 40919
rect 20947 40916 20959 40919
rect 21450 40916 21456 40928
rect 20947 40888 21456 40916
rect 20947 40885 20959 40888
rect 20901 40879 20959 40885
rect 21450 40876 21456 40888
rect 21508 40876 21514 40928
rect 22186 40916 22192 40928
rect 22147 40888 22192 40916
rect 22186 40876 22192 40888
rect 22244 40876 22250 40928
rect 25976 40925 26004 40956
rect 27341 40953 27353 40956
rect 27387 40953 27399 40987
rect 27341 40947 27399 40953
rect 25961 40919 26019 40925
rect 25961 40885 25973 40919
rect 26007 40885 26019 40919
rect 26602 40916 26608 40928
rect 26563 40888 26608 40916
rect 25961 40879 26019 40885
rect 26602 40876 26608 40888
rect 26660 40876 26666 40928
rect 27246 40876 27252 40928
rect 27304 40916 27310 40928
rect 27985 40919 28043 40925
rect 27985 40916 27997 40919
rect 27304 40888 27997 40916
rect 27304 40876 27310 40888
rect 27985 40885 27997 40888
rect 28031 40885 28043 40919
rect 27985 40879 28043 40885
rect 1104 40826 28888 40848
rect 1104 40774 10246 40826
rect 10298 40774 10310 40826
rect 10362 40774 10374 40826
rect 10426 40774 10438 40826
rect 10490 40774 19510 40826
rect 19562 40774 19574 40826
rect 19626 40774 19638 40826
rect 19690 40774 19702 40826
rect 19754 40774 28888 40826
rect 1104 40752 28888 40774
rect 2498 40712 2504 40724
rect 2459 40684 2504 40712
rect 2498 40672 2504 40684
rect 2556 40672 2562 40724
rect 5721 40715 5779 40721
rect 5721 40712 5733 40715
rect 2746 40684 5733 40712
rect 2130 40604 2136 40656
rect 2188 40644 2194 40656
rect 2746 40644 2774 40684
rect 5721 40681 5733 40684
rect 5767 40681 5779 40715
rect 5721 40675 5779 40681
rect 7190 40672 7196 40724
rect 7248 40712 7254 40724
rect 7377 40715 7435 40721
rect 7377 40712 7389 40715
rect 7248 40684 7389 40712
rect 7248 40672 7254 40684
rect 7377 40681 7389 40684
rect 7423 40681 7435 40715
rect 7650 40712 7656 40724
rect 7377 40675 7435 40681
rect 7484 40684 7656 40712
rect 2188 40616 2774 40644
rect 2869 40647 2927 40653
rect 2188 40604 2194 40616
rect 2869 40613 2881 40647
rect 2915 40644 2927 40647
rect 4709 40647 4767 40653
rect 2915 40616 3924 40644
rect 2915 40613 2927 40616
rect 2869 40607 2927 40613
rect 1857 40579 1915 40585
rect 1857 40545 1869 40579
rect 1903 40576 1915 40579
rect 2682 40576 2688 40588
rect 1903 40548 2688 40576
rect 1903 40545 1915 40548
rect 1857 40539 1915 40545
rect 2682 40536 2688 40548
rect 2740 40536 2746 40588
rect 3694 40576 3700 40588
rect 3655 40548 3700 40576
rect 3694 40536 3700 40548
rect 3752 40536 3758 40588
rect 3896 40576 3924 40616
rect 4709 40613 4721 40647
rect 4755 40644 4767 40647
rect 4890 40644 4896 40656
rect 4755 40616 4896 40644
rect 4755 40613 4767 40616
rect 4709 40607 4767 40613
rect 4890 40604 4896 40616
rect 4948 40604 4954 40656
rect 7484 40653 7512 40684
rect 7650 40672 7656 40684
rect 7708 40712 7714 40724
rect 10962 40712 10968 40724
rect 7708 40684 10968 40712
rect 7708 40672 7714 40684
rect 10962 40672 10968 40684
rect 11020 40712 11026 40724
rect 13814 40712 13820 40724
rect 11020 40684 13820 40712
rect 11020 40672 11026 40684
rect 13814 40672 13820 40684
rect 13872 40712 13878 40724
rect 15381 40715 15439 40721
rect 15381 40712 15393 40715
rect 13872 40684 15393 40712
rect 13872 40672 13878 40684
rect 15381 40681 15393 40684
rect 15427 40681 15439 40715
rect 15381 40675 15439 40681
rect 21361 40715 21419 40721
rect 21361 40681 21373 40715
rect 21407 40712 21419 40715
rect 21450 40712 21456 40724
rect 21407 40684 21456 40712
rect 21407 40681 21419 40684
rect 21361 40675 21419 40681
rect 21450 40672 21456 40684
rect 21508 40672 21514 40724
rect 7469 40647 7527 40653
rect 7469 40613 7481 40647
rect 7515 40613 7527 40647
rect 19426 40644 19432 40656
rect 7469 40607 7527 40613
rect 12544 40616 14136 40644
rect 4982 40576 4988 40588
rect 3896 40548 4988 40576
rect 4982 40536 4988 40548
rect 5040 40536 5046 40588
rect 5350 40536 5356 40588
rect 5408 40576 5414 40588
rect 5629 40579 5687 40585
rect 5629 40576 5641 40579
rect 5408 40548 5641 40576
rect 5408 40536 5414 40548
rect 5629 40545 5641 40548
rect 5675 40545 5687 40579
rect 5629 40539 5687 40545
rect 5813 40579 5871 40585
rect 5813 40545 5825 40579
rect 5859 40576 5871 40579
rect 6178 40576 6184 40588
rect 5859 40548 6184 40576
rect 5859 40545 5871 40548
rect 5813 40539 5871 40545
rect 6178 40536 6184 40548
rect 6236 40536 6242 40588
rect 7190 40576 7196 40588
rect 7151 40548 7196 40576
rect 7190 40536 7196 40548
rect 7248 40536 7254 40588
rect 11149 40579 11207 40585
rect 11149 40545 11161 40579
rect 11195 40576 11207 40579
rect 12544 40576 12572 40616
rect 12710 40576 12716 40588
rect 11195 40548 12572 40576
rect 12671 40548 12716 40576
rect 11195 40545 11207 40548
rect 11149 40539 11207 40545
rect 12710 40536 12716 40548
rect 12768 40536 12774 40588
rect 12805 40579 12863 40585
rect 12805 40545 12817 40579
rect 12851 40545 12863 40579
rect 12805 40539 12863 40545
rect 12897 40579 12955 40585
rect 12897 40545 12909 40579
rect 12943 40545 12955 40579
rect 13078 40576 13084 40588
rect 13039 40548 13084 40576
rect 12897 40539 12955 40545
rect 2961 40511 3019 40517
rect 2961 40477 2973 40511
rect 3007 40477 3019 40511
rect 2961 40471 3019 40477
rect 3145 40511 3203 40517
rect 3145 40477 3157 40511
rect 3191 40508 3203 40511
rect 3326 40508 3332 40520
rect 3191 40480 3332 40508
rect 3191 40477 3203 40480
rect 3145 40471 3203 40477
rect 2976 40440 3004 40471
rect 3326 40468 3332 40480
rect 3384 40508 3390 40520
rect 3602 40508 3608 40520
rect 3384 40480 3608 40508
rect 3384 40468 3390 40480
rect 3602 40468 3608 40480
rect 3660 40468 3666 40520
rect 4890 40468 4896 40520
rect 4948 40508 4954 40520
rect 5258 40508 5264 40520
rect 4948 40480 5264 40508
rect 4948 40468 4954 40480
rect 5258 40468 5264 40480
rect 5316 40468 5322 40520
rect 9950 40468 9956 40520
rect 10008 40508 10014 40520
rect 11882 40508 11888 40520
rect 10008 40480 11888 40508
rect 10008 40468 10014 40480
rect 11882 40468 11888 40480
rect 11940 40468 11946 40520
rect 12434 40468 12440 40520
rect 12492 40508 12498 40520
rect 12820 40508 12848 40539
rect 12492 40480 12848 40508
rect 12492 40468 12498 40480
rect 4246 40440 4252 40452
rect 2976 40412 4252 40440
rect 4246 40400 4252 40412
rect 4304 40400 4310 40452
rect 4614 40400 4620 40452
rect 4672 40440 4678 40452
rect 4982 40440 4988 40452
rect 4672 40412 4988 40440
rect 4672 40400 4678 40412
rect 4982 40400 4988 40412
rect 5040 40400 5046 40452
rect 7006 40400 7012 40452
rect 7064 40440 7070 40452
rect 9766 40440 9772 40452
rect 7064 40412 9772 40440
rect 7064 40400 7070 40412
rect 9766 40400 9772 40412
rect 9824 40400 9830 40452
rect 12710 40400 12716 40452
rect 12768 40440 12774 40452
rect 12912 40440 12940 40539
rect 13078 40536 13084 40548
rect 13136 40536 13142 40588
rect 13722 40536 13728 40588
rect 13780 40576 13786 40588
rect 14001 40579 14059 40585
rect 14001 40576 14013 40579
rect 13780 40548 14013 40576
rect 13780 40536 13786 40548
rect 14001 40545 14013 40548
rect 14047 40545 14059 40579
rect 14108 40576 14136 40616
rect 17880 40616 19432 40644
rect 14734 40576 14740 40588
rect 14108 40548 14740 40576
rect 14001 40539 14059 40545
rect 14734 40536 14740 40548
rect 14792 40536 14798 40588
rect 17880 40585 17908 40616
rect 19426 40604 19432 40616
rect 19484 40604 19490 40656
rect 20248 40647 20306 40653
rect 20248 40613 20260 40647
rect 20294 40644 20306 40647
rect 20530 40644 20536 40656
rect 20294 40616 20536 40644
rect 20294 40613 20306 40616
rect 20248 40607 20306 40613
rect 20530 40604 20536 40616
rect 20588 40604 20594 40656
rect 24026 40604 24032 40656
rect 24084 40604 24090 40656
rect 26602 40604 26608 40656
rect 26660 40644 26666 40656
rect 27893 40647 27951 40653
rect 27893 40644 27905 40647
rect 26660 40616 27905 40644
rect 26660 40604 26666 40616
rect 27893 40613 27905 40616
rect 27939 40613 27951 40647
rect 27893 40607 27951 40613
rect 17865 40579 17923 40585
rect 17865 40545 17877 40579
rect 17911 40545 17923 40579
rect 18046 40576 18052 40588
rect 18007 40548 18052 40576
rect 17865 40539 17923 40545
rect 18046 40536 18052 40548
rect 18104 40536 18110 40588
rect 18874 40576 18880 40588
rect 18835 40548 18880 40576
rect 18874 40536 18880 40548
rect 18932 40536 18938 40588
rect 18966 40536 18972 40588
rect 19024 40576 19030 40588
rect 19061 40579 19119 40585
rect 19061 40576 19073 40579
rect 19024 40548 19073 40576
rect 19024 40536 19030 40548
rect 19061 40545 19073 40548
rect 19107 40545 19119 40579
rect 19061 40539 19119 40545
rect 19981 40579 20039 40585
rect 19981 40545 19993 40579
rect 20027 40576 20039 40579
rect 20070 40576 20076 40588
rect 20027 40548 20076 40576
rect 20027 40545 20039 40548
rect 19981 40539 20039 40545
rect 20070 40536 20076 40548
rect 20128 40536 20134 40588
rect 23385 40579 23443 40585
rect 23385 40545 23397 40579
rect 23431 40576 23443 40579
rect 23658 40576 23664 40588
rect 23431 40548 23664 40576
rect 23431 40545 23443 40548
rect 23385 40539 23443 40545
rect 23658 40536 23664 40548
rect 23716 40536 23722 40588
rect 23842 40576 23848 40588
rect 23803 40548 23848 40576
rect 23842 40536 23848 40548
rect 23900 40536 23906 40588
rect 24854 40536 24860 40588
rect 24912 40576 24918 40588
rect 25961 40579 26019 40585
rect 25961 40576 25973 40579
rect 24912 40548 25973 40576
rect 24912 40536 24918 40548
rect 25961 40545 25973 40548
rect 26007 40545 26019 40579
rect 25961 40539 26019 40545
rect 14274 40508 14280 40520
rect 14235 40480 14280 40508
rect 14274 40468 14280 40480
rect 14332 40468 14338 40520
rect 17957 40511 18015 40517
rect 17957 40477 17969 40511
rect 18003 40508 18015 40511
rect 18785 40511 18843 40517
rect 18785 40508 18797 40511
rect 18003 40480 18797 40508
rect 18003 40477 18015 40480
rect 17957 40471 18015 40477
rect 18785 40477 18797 40480
rect 18831 40477 18843 40511
rect 19518 40508 19524 40520
rect 19479 40480 19524 40508
rect 18785 40471 18843 40477
rect 19518 40468 19524 40480
rect 19576 40468 19582 40520
rect 24486 40468 24492 40520
rect 24544 40508 24550 40520
rect 26053 40511 26111 40517
rect 26053 40508 26065 40511
rect 24544 40480 26065 40508
rect 24544 40468 24550 40480
rect 26053 40477 26065 40480
rect 26099 40477 26111 40511
rect 26053 40471 26111 40477
rect 26142 40468 26148 40520
rect 26200 40508 26206 40520
rect 26200 40480 26245 40508
rect 26200 40468 26206 40480
rect 12768 40412 14044 40440
rect 12768 40400 12774 40412
rect 1946 40372 1952 40384
rect 1907 40344 1952 40372
rect 1946 40332 1952 40344
rect 2004 40332 2010 40384
rect 3786 40372 3792 40384
rect 3747 40344 3792 40372
rect 3786 40332 3792 40344
rect 3844 40332 3850 40384
rect 4154 40372 4160 40384
rect 4115 40344 4160 40372
rect 4154 40332 4160 40344
rect 4212 40332 4218 40384
rect 5169 40375 5227 40381
rect 5169 40341 5181 40375
rect 5215 40372 5227 40375
rect 5442 40372 5448 40384
rect 5215 40344 5448 40372
rect 5215 40341 5227 40344
rect 5169 40335 5227 40341
rect 5442 40332 5448 40344
rect 5500 40332 5506 40384
rect 6914 40372 6920 40384
rect 6875 40344 6920 40372
rect 6914 40332 6920 40344
rect 6972 40332 6978 40384
rect 9490 40332 9496 40384
rect 9548 40372 9554 40384
rect 10686 40372 10692 40384
rect 9548 40344 10692 40372
rect 9548 40332 9554 40344
rect 10686 40332 10692 40344
rect 10744 40372 10750 40384
rect 10965 40375 11023 40381
rect 10965 40372 10977 40375
rect 10744 40344 10977 40372
rect 10744 40332 10750 40344
rect 10965 40341 10977 40344
rect 11011 40341 11023 40375
rect 10965 40335 11023 40341
rect 12342 40332 12348 40384
rect 12400 40372 12406 40384
rect 12437 40375 12495 40381
rect 12437 40372 12449 40375
rect 12400 40344 12449 40372
rect 12400 40332 12406 40344
rect 12437 40341 12449 40344
rect 12483 40341 12495 40375
rect 12437 40335 12495 40341
rect 12802 40332 12808 40384
rect 12860 40372 12866 40384
rect 13170 40372 13176 40384
rect 12860 40344 13176 40372
rect 12860 40332 12866 40344
rect 13170 40332 13176 40344
rect 13228 40332 13234 40384
rect 14016 40372 14044 40412
rect 16666 40372 16672 40384
rect 14016 40344 16672 40372
rect 16666 40332 16672 40344
rect 16724 40332 16730 40384
rect 25593 40375 25651 40381
rect 25593 40341 25605 40375
rect 25639 40372 25651 40375
rect 25958 40372 25964 40384
rect 25639 40344 25964 40372
rect 25639 40341 25651 40344
rect 25593 40335 25651 40341
rect 25958 40332 25964 40344
rect 26016 40332 26022 40384
rect 27982 40372 27988 40384
rect 27943 40344 27988 40372
rect 27982 40332 27988 40344
rect 28040 40332 28046 40384
rect 1104 40282 28888 40304
rect 1104 40230 5614 40282
rect 5666 40230 5678 40282
rect 5730 40230 5742 40282
rect 5794 40230 5806 40282
rect 5858 40230 14878 40282
rect 14930 40230 14942 40282
rect 14994 40230 15006 40282
rect 15058 40230 15070 40282
rect 15122 40230 24142 40282
rect 24194 40230 24206 40282
rect 24258 40230 24270 40282
rect 24322 40230 24334 40282
rect 24386 40230 28888 40282
rect 1104 40208 28888 40230
rect 3050 40128 3056 40180
rect 3108 40168 3114 40180
rect 27982 40168 27988 40180
rect 3108 40140 27988 40168
rect 3108 40128 3114 40140
rect 27982 40128 27988 40140
rect 28040 40128 28046 40180
rect 13446 40060 13452 40112
rect 13504 40100 13510 40112
rect 15102 40100 15108 40112
rect 13504 40072 15108 40100
rect 13504 40060 13510 40072
rect 15102 40060 15108 40072
rect 15160 40060 15166 40112
rect 17034 40060 17040 40112
rect 17092 40100 17098 40112
rect 22462 40100 22468 40112
rect 17092 40072 22468 40100
rect 17092 40060 17098 40072
rect 5442 39992 5448 40044
rect 5500 40032 5506 40044
rect 5537 40035 5595 40041
rect 5537 40032 5549 40035
rect 5500 40004 5549 40032
rect 5500 39992 5506 40004
rect 5537 40001 5549 40004
rect 5583 40001 5595 40035
rect 5537 39995 5595 40001
rect 6457 40035 6515 40041
rect 6457 40001 6469 40035
rect 6503 40032 6515 40035
rect 7190 40032 7196 40044
rect 6503 40004 7196 40032
rect 6503 40001 6515 40004
rect 6457 39995 6515 40001
rect 7190 39992 7196 40004
rect 7248 39992 7254 40044
rect 7929 40035 7987 40041
rect 7929 40001 7941 40035
rect 7975 40032 7987 40035
rect 9582 40032 9588 40044
rect 7975 40004 9588 40032
rect 7975 40001 7987 40004
rect 7929 39995 7987 40001
rect 9582 39992 9588 40004
rect 9640 39992 9646 40044
rect 9858 39992 9864 40044
rect 9916 40032 9922 40044
rect 13173 40035 13231 40041
rect 9916 40004 10824 40032
rect 9916 39992 9922 40004
rect 10796 39976 10824 40004
rect 13173 40001 13185 40035
rect 13219 40032 13231 40035
rect 13998 40032 14004 40044
rect 13219 40004 14004 40032
rect 13219 40001 13231 40004
rect 13173 39995 13231 40001
rect 13998 39992 14004 40004
rect 14056 39992 14062 40044
rect 16209 40035 16267 40041
rect 14292 40004 15332 40032
rect 4338 39924 4344 39976
rect 4396 39964 4402 39976
rect 4433 39967 4491 39973
rect 4433 39964 4445 39967
rect 4396 39936 4445 39964
rect 4396 39924 4402 39936
rect 4433 39933 4445 39936
rect 4479 39933 4491 39967
rect 5074 39964 5080 39976
rect 5035 39936 5080 39964
rect 4433 39927 4491 39933
rect 5074 39924 5080 39936
rect 5132 39924 5138 39976
rect 5169 39967 5227 39973
rect 5169 39933 5181 39967
rect 5215 39933 5227 39967
rect 6362 39964 6368 39976
rect 6323 39936 6368 39964
rect 5169 39927 5227 39933
rect 1857 39899 1915 39905
rect 1857 39865 1869 39899
rect 1903 39896 1915 39899
rect 2406 39896 2412 39908
rect 1903 39868 2412 39896
rect 1903 39865 1915 39868
rect 1857 39859 1915 39865
rect 2406 39856 2412 39868
rect 2464 39856 2470 39908
rect 2590 39896 2596 39908
rect 2551 39868 2596 39896
rect 2590 39856 2596 39868
rect 2648 39856 2654 39908
rect 2774 39856 2780 39908
rect 2832 39896 2838 39908
rect 2832 39868 2877 39896
rect 2832 39856 2838 39868
rect 4522 39856 4528 39908
rect 4580 39896 4586 39908
rect 5184 39896 5212 39927
rect 6362 39924 6368 39936
rect 6420 39924 6426 39976
rect 6546 39964 6552 39976
rect 6507 39936 6552 39964
rect 6546 39924 6552 39936
rect 6604 39924 6610 39976
rect 7742 39924 7748 39976
rect 7800 39964 7806 39976
rect 8159 39967 8217 39973
rect 8159 39964 8171 39967
rect 7800 39936 8171 39964
rect 7800 39924 7806 39936
rect 8159 39933 8171 39936
rect 8205 39933 8217 39967
rect 8159 39927 8217 39933
rect 8297 39967 8355 39973
rect 8297 39933 8309 39967
rect 8343 39933 8355 39967
rect 8297 39927 8355 39933
rect 8389 39967 8447 39973
rect 8389 39933 8401 39967
rect 8435 39964 8447 39967
rect 8478 39964 8484 39976
rect 8435 39936 8484 39964
rect 8435 39933 8447 39936
rect 8389 39927 8447 39933
rect 4580 39868 5212 39896
rect 5813 39899 5871 39905
rect 4580 39856 4586 39868
rect 5813 39865 5825 39899
rect 5859 39896 5871 39899
rect 8312 39896 8340 39927
rect 8478 39924 8484 39936
rect 8536 39924 8542 39976
rect 8573 39967 8631 39973
rect 8573 39933 8585 39967
rect 8619 39964 8631 39967
rect 8662 39964 8668 39976
rect 8619 39936 8668 39964
rect 8619 39933 8631 39936
rect 8573 39927 8631 39933
rect 8662 39924 8668 39936
rect 8720 39924 8726 39976
rect 10689 39967 10747 39973
rect 10689 39933 10701 39967
rect 10735 39933 10747 39967
rect 10689 39927 10747 39933
rect 5859 39868 6592 39896
rect 5859 39865 5871 39868
rect 5813 39859 5871 39865
rect 6564 39840 6592 39868
rect 8266 39868 8340 39896
rect 1394 39788 1400 39840
rect 1452 39828 1458 39840
rect 1949 39831 2007 39837
rect 1949 39828 1961 39831
rect 1452 39800 1961 39828
rect 1452 39788 1458 39800
rect 1949 39797 1961 39800
rect 1995 39797 2007 39831
rect 1949 39791 2007 39797
rect 6546 39788 6552 39840
rect 6604 39788 6610 39840
rect 8110 39788 8116 39840
rect 8168 39828 8174 39840
rect 8266 39828 8294 39868
rect 8168 39800 8294 39828
rect 10704 39828 10732 39927
rect 10778 39924 10784 39976
rect 10836 39964 10842 39976
rect 12526 39964 12532 39976
rect 10836 39936 12532 39964
rect 10836 39924 10842 39936
rect 12526 39924 12532 39936
rect 12584 39924 12590 39976
rect 13262 39924 13268 39976
rect 13320 39964 13326 39976
rect 13449 39967 13507 39973
rect 13449 39964 13461 39967
rect 13320 39936 13461 39964
rect 13320 39924 13326 39936
rect 13449 39933 13461 39936
rect 13495 39933 13507 39967
rect 13449 39927 13507 39933
rect 13541 39967 13599 39973
rect 13541 39933 13553 39967
rect 13587 39933 13599 39967
rect 13541 39927 13599 39933
rect 10956 39899 11014 39905
rect 10956 39865 10968 39899
rect 11002 39896 11014 39899
rect 11974 39896 11980 39908
rect 11002 39868 11980 39896
rect 11002 39865 11014 39868
rect 10956 39859 11014 39865
rect 11974 39856 11980 39868
rect 12032 39856 12038 39908
rect 13556 39896 13584 39927
rect 13630 39924 13636 39976
rect 13688 39964 13694 39976
rect 13817 39967 13875 39973
rect 13688 39936 13733 39964
rect 13688 39924 13694 39936
rect 13817 39933 13829 39967
rect 13863 39964 13875 39967
rect 13906 39964 13912 39976
rect 13863 39936 13912 39964
rect 13863 39933 13875 39936
rect 13817 39927 13875 39933
rect 13906 39924 13912 39936
rect 13964 39924 13970 39976
rect 13722 39896 13728 39908
rect 13556 39868 13728 39896
rect 13722 39856 13728 39868
rect 13780 39896 13786 39908
rect 14292 39896 14320 40004
rect 15304 39973 15332 40004
rect 16209 40001 16221 40035
rect 16255 40032 16267 40035
rect 16758 40032 16764 40044
rect 16255 40004 16764 40032
rect 16255 40001 16267 40004
rect 16209 39995 16267 40001
rect 16758 39992 16764 40004
rect 16816 39992 16822 40044
rect 18046 39992 18052 40044
rect 18104 40032 18110 40044
rect 21284 40041 21312 40072
rect 22462 40060 22468 40072
rect 22520 40060 22526 40112
rect 20257 40035 20315 40041
rect 20257 40032 20269 40035
rect 18104 40004 20269 40032
rect 18104 39992 18110 40004
rect 20257 40001 20269 40004
rect 20303 40001 20315 40035
rect 20257 39995 20315 40001
rect 21269 40035 21327 40041
rect 21269 40001 21281 40035
rect 21315 40001 21327 40035
rect 22186 40032 22192 40044
rect 22147 40004 22192 40032
rect 21269 39995 21327 40001
rect 22186 39992 22192 40004
rect 22244 39992 22250 40044
rect 22925 40035 22983 40041
rect 22925 40001 22937 40035
rect 22971 40032 22983 40035
rect 23842 40032 23848 40044
rect 22971 40004 23848 40032
rect 22971 40001 22983 40004
rect 22925 39995 22983 40001
rect 15197 39967 15255 39973
rect 15197 39933 15209 39967
rect 15243 39933 15255 39967
rect 15197 39927 15255 39933
rect 15289 39967 15347 39973
rect 15289 39933 15301 39967
rect 15335 39933 15347 39967
rect 15289 39927 15347 39933
rect 13780 39868 14320 39896
rect 15212 39896 15240 39927
rect 15378 39924 15384 39976
rect 15436 39964 15442 39976
rect 15565 39967 15623 39973
rect 15436 39936 15481 39964
rect 15436 39924 15442 39936
rect 15565 39933 15577 39967
rect 15611 39964 15623 39967
rect 16114 39964 16120 39976
rect 15611 39936 16120 39964
rect 15611 39933 15623 39936
rect 15565 39927 15623 39933
rect 16114 39924 16120 39936
rect 16172 39924 16178 39976
rect 16482 39964 16488 39976
rect 16443 39936 16488 39964
rect 16482 39924 16488 39936
rect 16540 39924 16546 39976
rect 16577 39967 16635 39973
rect 16577 39933 16589 39967
rect 16623 39933 16635 39967
rect 16577 39927 16635 39933
rect 15470 39896 15476 39908
rect 15212 39868 15476 39896
rect 13780 39856 13786 39868
rect 15470 39856 15476 39868
rect 15528 39856 15534 39908
rect 11054 39828 11060 39840
rect 10704 39800 11060 39828
rect 8168 39788 8174 39800
rect 11054 39788 11060 39800
rect 11112 39788 11118 39840
rect 12066 39828 12072 39840
rect 12027 39800 12072 39828
rect 12066 39788 12072 39800
rect 12124 39788 12130 39840
rect 14366 39788 14372 39840
rect 14424 39828 14430 39840
rect 14826 39828 14832 39840
rect 14424 39800 14832 39828
rect 14424 39788 14430 39800
rect 14826 39788 14832 39800
rect 14884 39788 14890 39840
rect 14921 39831 14979 39837
rect 14921 39797 14933 39831
rect 14967 39828 14979 39831
rect 15194 39828 15200 39840
rect 14967 39800 15200 39828
rect 14967 39797 14979 39800
rect 14921 39791 14979 39797
rect 15194 39788 15200 39800
rect 15252 39788 15258 39840
rect 15286 39788 15292 39840
rect 15344 39828 15350 39840
rect 16500 39828 16528 39924
rect 16592 39896 16620 39927
rect 16666 39924 16672 39976
rect 16724 39964 16730 39976
rect 16853 39967 16911 39973
rect 16724 39936 16769 39964
rect 16724 39924 16730 39936
rect 16853 39933 16865 39967
rect 16899 39964 16911 39967
rect 16942 39964 16948 39976
rect 16899 39936 16948 39964
rect 16899 39933 16911 39936
rect 16853 39927 16911 39933
rect 16942 39924 16948 39936
rect 17000 39924 17006 39976
rect 18414 39964 18420 39976
rect 18064 39936 18420 39964
rect 18064 39908 18092 39936
rect 18414 39924 18420 39936
rect 18472 39924 18478 39976
rect 21082 39964 21088 39976
rect 21043 39936 21088 39964
rect 21082 39924 21088 39936
rect 21140 39924 21146 39976
rect 22281 39967 22339 39973
rect 22281 39964 22293 39967
rect 22066 39936 22293 39964
rect 16758 39896 16764 39908
rect 16592 39868 16764 39896
rect 16758 39856 16764 39868
rect 16816 39856 16822 39908
rect 18046 39856 18052 39908
rect 18104 39856 18110 39908
rect 18233 39899 18291 39905
rect 18233 39865 18245 39899
rect 18279 39865 18291 39899
rect 18598 39896 18604 39908
rect 18559 39868 18604 39896
rect 18233 39859 18291 39865
rect 15344 39800 16528 39828
rect 18248 39828 18276 39859
rect 18598 39856 18604 39868
rect 18656 39856 18662 39908
rect 19518 39896 19524 39908
rect 19306 39868 19524 39896
rect 18414 39828 18420 39840
rect 18248 39800 18420 39828
rect 15344 39788 15350 39800
rect 18414 39788 18420 39800
rect 18472 39828 18478 39840
rect 19306 39828 19334 39868
rect 19518 39856 19524 39868
rect 19576 39856 19582 39908
rect 20073 39899 20131 39905
rect 20073 39865 20085 39899
rect 20119 39896 20131 39899
rect 20162 39896 20168 39908
rect 20119 39868 20168 39896
rect 20119 39865 20131 39868
rect 20073 39859 20131 39865
rect 20162 39856 20168 39868
rect 20220 39856 20226 39908
rect 22066 39896 22094 39936
rect 22281 39933 22293 39936
rect 22327 39933 22339 39967
rect 22281 39927 22339 39933
rect 22465 39967 22523 39973
rect 22465 39933 22477 39967
rect 22511 39964 22523 39967
rect 23198 39964 23204 39976
rect 22511 39936 23204 39964
rect 22511 39933 22523 39936
rect 22465 39927 22523 39933
rect 23198 39924 23204 39936
rect 23256 39924 23262 39976
rect 23400 39973 23428 40004
rect 23842 39992 23848 40004
rect 23900 39992 23906 40044
rect 24101 40035 24159 40041
rect 24101 40001 24113 40035
rect 24147 40032 24159 40035
rect 25222 40032 25228 40044
rect 24147 40004 25228 40032
rect 24147 40001 24159 40004
rect 24101 39995 24159 40001
rect 25222 39992 25228 40004
rect 25280 39992 25286 40044
rect 25314 39992 25320 40044
rect 25372 40032 25378 40044
rect 25869 40035 25927 40041
rect 25869 40032 25881 40035
rect 25372 40004 25881 40032
rect 25372 39992 25378 40004
rect 25869 40001 25881 40004
rect 25915 40001 25927 40035
rect 25869 39995 25927 40001
rect 23385 39967 23443 39973
rect 23385 39933 23397 39967
rect 23431 39933 23443 39967
rect 23385 39927 23443 39933
rect 23569 39967 23627 39973
rect 23569 39933 23581 39967
rect 23615 39964 23627 39967
rect 23658 39964 23664 39976
rect 23615 39936 23664 39964
rect 23615 39933 23627 39936
rect 23569 39927 23627 39933
rect 23658 39924 23664 39936
rect 23716 39924 23722 39976
rect 24210 39924 24216 39976
rect 24268 39964 24274 39976
rect 24305 39967 24363 39973
rect 24305 39964 24317 39967
rect 24268 39936 24317 39964
rect 24268 39924 24274 39936
rect 24305 39933 24317 39936
rect 24351 39933 24363 39967
rect 25406 39964 25412 39976
rect 25367 39936 25412 39964
rect 24305 39927 24363 39933
rect 25406 39924 25412 39936
rect 25464 39924 25470 39976
rect 25958 39924 25964 39976
rect 26016 39964 26022 39976
rect 26125 39967 26183 39973
rect 26125 39964 26137 39967
rect 26016 39936 26137 39964
rect 26016 39924 26022 39936
rect 26125 39933 26137 39936
rect 26171 39933 26183 39967
rect 27890 39964 27896 39976
rect 27851 39936 27896 39964
rect 26125 39927 26183 39933
rect 27890 39924 27896 39936
rect 27948 39924 27954 39976
rect 20732 39868 22094 39896
rect 23477 39899 23535 39905
rect 20732 39837 20760 39868
rect 23477 39865 23489 39899
rect 23523 39896 23535 39899
rect 24029 39899 24087 39905
rect 24029 39896 24041 39899
rect 23523 39868 24041 39896
rect 23523 39865 23535 39868
rect 23477 39859 23535 39865
rect 24029 39865 24041 39868
rect 24075 39865 24087 39899
rect 24029 39859 24087 39865
rect 24486 39856 24492 39908
rect 24544 39896 24550 39908
rect 24544 39868 27292 39896
rect 24544 39856 24550 39868
rect 18472 39800 19334 39828
rect 20717 39831 20775 39837
rect 18472 39788 18478 39800
rect 20717 39797 20729 39831
rect 20763 39797 20775 39831
rect 20717 39791 20775 39797
rect 21177 39831 21235 39837
rect 21177 39797 21189 39831
rect 21223 39828 21235 39831
rect 22646 39828 22652 39840
rect 21223 39800 22652 39828
rect 21223 39797 21235 39800
rect 21177 39791 21235 39797
rect 22646 39788 22652 39800
rect 22704 39788 22710 39840
rect 23566 39788 23572 39840
rect 23624 39828 23630 39840
rect 24213 39831 24271 39837
rect 24213 39828 24225 39831
rect 23624 39800 24225 39828
rect 23624 39788 23630 39800
rect 24213 39797 24225 39800
rect 24259 39828 24271 39831
rect 24394 39828 24400 39840
rect 24259 39800 24400 39828
rect 24259 39797 24271 39800
rect 24213 39791 24271 39797
rect 24394 39788 24400 39800
rect 24452 39788 24458 39840
rect 25222 39828 25228 39840
rect 25183 39800 25228 39828
rect 25222 39788 25228 39800
rect 25280 39788 25286 39840
rect 27264 39837 27292 39868
rect 27249 39831 27307 39837
rect 27249 39797 27261 39831
rect 27295 39797 27307 39831
rect 27249 39791 27307 39797
rect 27338 39788 27344 39840
rect 27396 39828 27402 39840
rect 27985 39831 28043 39837
rect 27985 39828 27997 39831
rect 27396 39800 27997 39828
rect 27396 39788 27402 39800
rect 27985 39797 27997 39800
rect 28031 39797 28043 39831
rect 27985 39791 28043 39797
rect 1104 39738 28888 39760
rect 1104 39686 10246 39738
rect 10298 39686 10310 39738
rect 10362 39686 10374 39738
rect 10426 39686 10438 39738
rect 10490 39686 19510 39738
rect 19562 39686 19574 39738
rect 19626 39686 19638 39738
rect 19690 39686 19702 39738
rect 19754 39686 28888 39738
rect 1104 39664 28888 39686
rect 3602 39584 3608 39636
rect 3660 39624 3666 39636
rect 4617 39627 4675 39633
rect 4617 39624 4629 39627
rect 3660 39596 4629 39624
rect 3660 39584 3666 39596
rect 4617 39593 4629 39596
rect 4663 39593 4675 39627
rect 11698 39624 11704 39636
rect 4617 39587 4675 39593
rect 5184 39596 11704 39624
rect 3697 39559 3755 39565
rect 3697 39525 3709 39559
rect 3743 39556 3755 39559
rect 4154 39556 4160 39568
rect 3743 39528 4160 39556
rect 3743 39525 3755 39528
rect 3697 39519 3755 39525
rect 4154 39516 4160 39528
rect 4212 39516 4218 39568
rect 4525 39559 4583 39565
rect 4525 39525 4537 39559
rect 4571 39556 4583 39559
rect 5184 39556 5212 39596
rect 11698 39584 11704 39596
rect 11756 39584 11762 39636
rect 11974 39584 11980 39636
rect 12032 39624 12038 39636
rect 12069 39627 12127 39633
rect 12069 39624 12081 39627
rect 12032 39596 12081 39624
rect 12032 39584 12038 39596
rect 12069 39593 12081 39596
rect 12115 39593 12127 39627
rect 12069 39587 12127 39593
rect 12710 39584 12716 39636
rect 12768 39584 12774 39636
rect 13909 39627 13967 39633
rect 13909 39593 13921 39627
rect 13955 39624 13967 39627
rect 14274 39624 14280 39636
rect 13955 39596 14280 39624
rect 13955 39593 13967 39596
rect 13909 39587 13967 39593
rect 14274 39584 14280 39596
rect 14332 39584 14338 39636
rect 15378 39624 15384 39636
rect 14389 39596 15384 39624
rect 4571 39528 5212 39556
rect 5261 39559 5319 39565
rect 4571 39525 4583 39528
rect 4525 39519 4583 39525
rect 5261 39525 5273 39559
rect 5307 39556 5319 39559
rect 10226 39556 10232 39568
rect 5307 39528 10232 39556
rect 5307 39525 5319 39528
rect 5261 39519 5319 39525
rect 10226 39516 10232 39528
rect 10284 39516 10290 39568
rect 10689 39559 10747 39565
rect 10689 39525 10701 39559
rect 10735 39556 10747 39559
rect 12728 39556 12756 39584
rect 10735 39528 10999 39556
rect 10735 39525 10747 39528
rect 10689 39519 10747 39525
rect 1857 39491 1915 39497
rect 1857 39457 1869 39491
rect 1903 39488 1915 39491
rect 2222 39488 2228 39500
rect 1903 39460 2228 39488
rect 1903 39457 1915 39460
rect 1857 39451 1915 39457
rect 2222 39448 2228 39460
rect 2280 39448 2286 39500
rect 2498 39448 2504 39500
rect 2556 39488 2562 39500
rect 2593 39491 2651 39497
rect 2593 39488 2605 39491
rect 2556 39460 2605 39488
rect 2556 39448 2562 39460
rect 2593 39457 2605 39460
rect 2639 39457 2651 39491
rect 3878 39488 3884 39500
rect 3839 39460 3884 39488
rect 2593 39451 2651 39457
rect 3878 39448 3884 39460
rect 3936 39448 3942 39500
rect 3970 39448 3976 39500
rect 4028 39488 4034 39500
rect 4028 39460 4073 39488
rect 4028 39448 4034 39460
rect 6914 39448 6920 39500
rect 6972 39488 6978 39500
rect 7009 39491 7067 39497
rect 7009 39488 7021 39491
rect 6972 39460 7021 39488
rect 6972 39448 6978 39460
rect 7009 39457 7021 39460
rect 7055 39457 7067 39491
rect 7009 39451 7067 39457
rect 8021 39491 8079 39497
rect 8021 39457 8033 39491
rect 8067 39457 8079 39491
rect 8021 39451 8079 39457
rect 8389 39491 8447 39497
rect 8389 39457 8401 39491
rect 8435 39488 8447 39491
rect 8478 39488 8484 39500
rect 8435 39460 8484 39488
rect 8435 39457 8447 39460
rect 8389 39451 8447 39457
rect 2682 39380 2688 39432
rect 2740 39420 2746 39432
rect 2740 39392 3740 39420
rect 2740 39380 2746 39392
rect 2777 39355 2835 39361
rect 2777 39321 2789 39355
rect 2823 39352 2835 39355
rect 2866 39352 2872 39364
rect 2823 39324 2872 39352
rect 2823 39321 2835 39324
rect 2777 39315 2835 39321
rect 2866 39312 2872 39324
rect 2924 39312 2930 39364
rect 1949 39287 2007 39293
rect 1949 39253 1961 39287
rect 1995 39284 2007 39287
rect 2958 39284 2964 39296
rect 1995 39256 2964 39284
rect 1995 39253 2007 39256
rect 1949 39247 2007 39253
rect 2958 39244 2964 39256
rect 3016 39244 3022 39296
rect 3712 39284 3740 39392
rect 3786 39380 3792 39432
rect 3844 39420 3850 39432
rect 5445 39423 5503 39429
rect 5445 39420 5457 39423
rect 3844 39392 5457 39420
rect 3844 39380 3850 39392
rect 5445 39389 5457 39392
rect 5491 39389 5503 39423
rect 5445 39383 5503 39389
rect 6362 39380 6368 39432
rect 6420 39420 6426 39432
rect 6825 39423 6883 39429
rect 6825 39420 6837 39423
rect 6420 39392 6837 39420
rect 6420 39380 6426 39392
rect 6825 39389 6837 39392
rect 6871 39420 6883 39423
rect 7098 39420 7104 39432
rect 6871 39392 7104 39420
rect 6871 39389 6883 39392
rect 6825 39383 6883 39389
rect 7098 39380 7104 39392
rect 7156 39380 7162 39432
rect 8036 39420 8064 39451
rect 8478 39448 8484 39460
rect 8536 39448 8542 39500
rect 8662 39488 8668 39500
rect 8623 39460 8668 39488
rect 8662 39448 8668 39460
rect 8720 39448 8726 39500
rect 9214 39448 9220 39500
rect 9272 39488 9278 39500
rect 9677 39491 9735 39497
rect 9677 39488 9689 39491
rect 9272 39460 9689 39488
rect 9272 39448 9278 39460
rect 9677 39457 9689 39460
rect 9723 39457 9735 39491
rect 9858 39488 9864 39500
rect 9819 39460 9864 39488
rect 9677 39451 9735 39457
rect 9858 39448 9864 39460
rect 9916 39448 9922 39500
rect 10318 39488 10324 39500
rect 10279 39460 10324 39488
rect 10318 39448 10324 39460
rect 10376 39448 10382 39500
rect 10502 39497 10508 39500
rect 10469 39491 10508 39497
rect 10469 39457 10481 39491
rect 10469 39451 10508 39457
rect 10502 39448 10508 39451
rect 10560 39448 10566 39500
rect 10870 39497 10876 39500
rect 10597 39491 10655 39497
rect 10597 39457 10609 39491
rect 10643 39457 10655 39491
rect 10597 39451 10655 39457
rect 10827 39491 10876 39497
rect 10827 39457 10839 39491
rect 10873 39457 10876 39491
rect 10827 39451 10876 39457
rect 8570 39420 8576 39432
rect 8036 39392 8576 39420
rect 8570 39380 8576 39392
rect 8628 39380 8634 39432
rect 8849 39423 8907 39429
rect 8849 39389 8861 39423
rect 8895 39389 8907 39423
rect 8849 39383 8907 39389
rect 3973 39355 4031 39361
rect 3973 39321 3985 39355
rect 4019 39352 4031 39355
rect 5258 39352 5264 39364
rect 4019 39324 5264 39352
rect 4019 39321 4031 39324
rect 3973 39315 4031 39321
rect 5258 39312 5264 39324
rect 5316 39312 5322 39364
rect 5368 39324 7880 39352
rect 5368 39284 5396 39324
rect 3712 39256 5396 39284
rect 7193 39287 7251 39293
rect 7193 39253 7205 39287
rect 7239 39284 7251 39287
rect 7742 39284 7748 39296
rect 7239 39256 7748 39284
rect 7239 39253 7251 39256
rect 7193 39247 7251 39253
rect 7742 39244 7748 39256
rect 7800 39244 7806 39296
rect 7852 39284 7880 39324
rect 8110 39312 8116 39364
rect 8168 39352 8174 39364
rect 8864 39352 8892 39383
rect 10226 39380 10232 39432
rect 10284 39420 10290 39432
rect 10612 39420 10640 39451
rect 10870 39448 10876 39451
rect 10928 39448 10934 39500
rect 10971 39488 10999 39528
rect 12544 39528 12756 39556
rect 11054 39488 11060 39500
rect 10971 39460 11060 39488
rect 11054 39448 11060 39460
rect 11112 39448 11118 39500
rect 11238 39448 11244 39500
rect 11296 39488 11302 39500
rect 11422 39488 11428 39500
rect 11296 39460 11428 39488
rect 11296 39448 11302 39460
rect 11422 39448 11428 39460
rect 11480 39448 11486 39500
rect 12066 39488 12072 39500
rect 11624 39460 12072 39488
rect 11624 39420 11652 39460
rect 12066 39448 12072 39460
rect 12124 39488 12130 39500
rect 12299 39491 12357 39497
rect 12299 39488 12311 39491
rect 12124 39460 12311 39488
rect 12124 39448 12130 39460
rect 12299 39457 12311 39460
rect 12345 39457 12357 39491
rect 12434 39488 12440 39500
rect 12395 39460 12440 39488
rect 12299 39451 12357 39457
rect 12434 39448 12440 39460
rect 12492 39448 12498 39500
rect 12544 39497 12572 39528
rect 12529 39491 12587 39497
rect 12529 39457 12541 39491
rect 12575 39457 12587 39491
rect 12529 39451 12587 39457
rect 12713 39491 12771 39497
rect 12713 39457 12725 39491
rect 12759 39488 12771 39491
rect 12802 39488 12808 39500
rect 12759 39460 12808 39488
rect 12759 39457 12771 39460
rect 12713 39451 12771 39457
rect 12802 39448 12808 39460
rect 12860 39448 12866 39500
rect 13814 39448 13820 39500
rect 13872 39488 13878 39500
rect 13998 39488 14004 39500
rect 13872 39460 14004 39488
rect 13872 39448 13878 39460
rect 13998 39448 14004 39460
rect 14056 39488 14062 39500
rect 14389 39497 14417 39596
rect 15378 39584 15384 39596
rect 15436 39584 15442 39636
rect 18049 39627 18107 39633
rect 18049 39593 18061 39627
rect 18095 39624 18107 39627
rect 20714 39624 20720 39636
rect 18095 39596 20720 39624
rect 18095 39593 18107 39596
rect 18049 39587 18107 39593
rect 20714 39584 20720 39596
rect 20772 39584 20778 39636
rect 22646 39624 22652 39636
rect 22607 39596 22652 39624
rect 22646 39584 22652 39596
rect 22704 39584 22710 39636
rect 27338 39624 27344 39636
rect 25056 39596 27344 39624
rect 14734 39516 14740 39568
rect 14792 39556 14798 39568
rect 14792 39528 15700 39556
rect 14792 39516 14798 39528
rect 14139 39491 14197 39497
rect 14139 39488 14151 39491
rect 14056 39460 14151 39488
rect 14056 39448 14062 39460
rect 14139 39457 14151 39460
rect 14185 39457 14197 39491
rect 14139 39451 14197 39457
rect 14277 39491 14335 39497
rect 14277 39457 14289 39491
rect 14323 39457 14335 39491
rect 14277 39451 14335 39457
rect 14374 39491 14432 39497
rect 14374 39457 14386 39491
rect 14420 39457 14432 39491
rect 14550 39488 14556 39500
rect 14511 39460 14556 39488
rect 14374 39451 14432 39457
rect 10284 39392 11652 39420
rect 10284 39380 10290 39392
rect 13722 39380 13728 39432
rect 13780 39420 13786 39432
rect 14292 39420 14320 39451
rect 13780 39392 14320 39420
rect 13780 39380 13786 39392
rect 8168 39324 8892 39352
rect 9125 39355 9183 39361
rect 8168 39312 8174 39324
rect 9125 39321 9137 39355
rect 9171 39352 9183 39355
rect 9306 39352 9312 39364
rect 9171 39324 9312 39352
rect 9171 39321 9183 39324
rect 9125 39315 9183 39321
rect 9306 39312 9312 39324
rect 9364 39312 9370 39364
rect 12526 39352 12532 39364
rect 9416 39324 12532 39352
rect 9416 39284 9444 39324
rect 12526 39312 12532 39324
rect 12584 39312 12590 39364
rect 7852 39256 9444 39284
rect 9674 39244 9680 39296
rect 9732 39284 9738 39296
rect 9769 39287 9827 39293
rect 9769 39284 9781 39287
rect 9732 39256 9781 39284
rect 9732 39244 9738 39256
rect 9769 39253 9781 39256
rect 9815 39253 9827 39287
rect 9769 39247 9827 39253
rect 9858 39244 9864 39296
rect 9916 39284 9922 39296
rect 10965 39287 11023 39293
rect 10965 39284 10977 39287
rect 9916 39256 10977 39284
rect 9916 39244 9922 39256
rect 10965 39253 10977 39256
rect 11011 39253 11023 39287
rect 10965 39247 11023 39253
rect 13630 39244 13636 39296
rect 13688 39284 13694 39296
rect 14389 39284 14417 39451
rect 14550 39448 14556 39460
rect 14608 39448 14614 39500
rect 14826 39448 14832 39500
rect 14884 39488 14890 39500
rect 15013 39491 15071 39497
rect 15013 39488 15025 39491
rect 14884 39460 15025 39488
rect 14884 39448 14890 39460
rect 15013 39457 15025 39460
rect 15059 39457 15071 39491
rect 15013 39451 15071 39457
rect 15102 39448 15108 39500
rect 15160 39488 15166 39500
rect 15286 39488 15292 39500
rect 15160 39460 15205 39488
rect 15247 39460 15292 39488
rect 15160 39448 15166 39460
rect 15286 39448 15292 39460
rect 15344 39448 15350 39500
rect 15378 39448 15384 39500
rect 15436 39488 15442 39500
rect 15519 39491 15577 39497
rect 15436 39460 15481 39488
rect 15436 39448 15442 39460
rect 15519 39457 15531 39491
rect 15565 39457 15577 39491
rect 15672 39488 15700 39528
rect 15838 39516 15844 39568
rect 15896 39556 15902 39568
rect 25056 39556 25084 39596
rect 27338 39584 27344 39596
rect 27396 39584 27402 39636
rect 15896 39528 25084 39556
rect 15896 39516 15902 39528
rect 25222 39516 25228 39568
rect 25280 39556 25286 39568
rect 27985 39559 28043 39565
rect 27985 39556 27997 39559
rect 25280 39528 27997 39556
rect 25280 39516 25286 39528
rect 27985 39525 27997 39528
rect 28031 39525 28043 39559
rect 27985 39519 28043 39525
rect 18233 39491 18291 39497
rect 18233 39488 18245 39491
rect 15672 39460 18245 39488
rect 15519 39451 15577 39457
rect 18233 39457 18245 39460
rect 18279 39457 18291 39491
rect 18233 39451 18291 39457
rect 14642 39380 14648 39432
rect 14700 39420 14706 39432
rect 15534 39420 15562 39451
rect 18598 39448 18604 39500
rect 18656 39488 18662 39500
rect 18949 39491 19007 39497
rect 18949 39488 18961 39491
rect 18656 39460 18961 39488
rect 18656 39448 18662 39460
rect 18949 39457 18961 39460
rect 18995 39457 19007 39491
rect 18949 39451 19007 39457
rect 22557 39491 22615 39497
rect 22557 39457 22569 39491
rect 22603 39488 22615 39491
rect 23658 39488 23664 39500
rect 22603 39460 23664 39488
rect 22603 39457 22615 39460
rect 22557 39451 22615 39457
rect 23658 39448 23664 39460
rect 23716 39448 23722 39500
rect 24210 39448 24216 39500
rect 24268 39488 24274 39500
rect 24489 39491 24547 39497
rect 24489 39488 24501 39491
rect 24268 39460 24501 39488
rect 24268 39448 24274 39460
rect 24489 39457 24501 39460
rect 24535 39457 24547 39491
rect 26878 39488 26884 39500
rect 26839 39460 26884 39488
rect 24489 39451 24547 39457
rect 26878 39448 26884 39460
rect 26936 39448 26942 39500
rect 14700 39392 15562 39420
rect 14700 39380 14706 39392
rect 15488 39364 15516 39392
rect 17218 39380 17224 39432
rect 17276 39420 17282 39432
rect 18693 39423 18751 39429
rect 18693 39420 18705 39423
rect 17276 39392 18705 39420
rect 17276 39380 17282 39392
rect 18693 39389 18705 39392
rect 18739 39389 18751 39423
rect 24394 39420 24400 39432
rect 24355 39392 24400 39420
rect 18693 39383 18751 39389
rect 24394 39380 24400 39392
rect 24452 39380 24458 39432
rect 24854 39420 24860 39432
rect 24815 39392 24860 39420
rect 24854 39380 24860 39392
rect 24912 39380 24918 39432
rect 15470 39312 15476 39364
rect 15528 39312 15534 39364
rect 28166 39352 28172 39364
rect 19628 39324 28172 39352
rect 15654 39284 15660 39296
rect 13688 39256 14417 39284
rect 15615 39256 15660 39284
rect 13688 39244 13694 39256
rect 15654 39244 15660 39256
rect 15712 39244 15718 39296
rect 15838 39244 15844 39296
rect 15896 39284 15902 39296
rect 19628 39284 19656 39324
rect 28166 39312 28172 39324
rect 28224 39312 28230 39364
rect 20070 39284 20076 39296
rect 15896 39256 19656 39284
rect 20031 39256 20076 39284
rect 15896 39244 15902 39256
rect 20070 39244 20076 39256
rect 20128 39244 20134 39296
rect 23658 39244 23664 39296
rect 23716 39284 23722 39296
rect 24486 39284 24492 39296
rect 23716 39256 24492 39284
rect 23716 39244 23722 39256
rect 24486 39244 24492 39256
rect 24544 39244 24550 39296
rect 26697 39287 26755 39293
rect 26697 39253 26709 39287
rect 26743 39284 26755 39287
rect 27890 39284 27896 39296
rect 26743 39256 27896 39284
rect 26743 39253 26755 39256
rect 26697 39247 26755 39253
rect 27890 39244 27896 39256
rect 27948 39244 27954 39296
rect 28074 39284 28080 39296
rect 28035 39256 28080 39284
rect 28074 39244 28080 39256
rect 28132 39244 28138 39296
rect 1104 39194 28888 39216
rect 1104 39142 5614 39194
rect 5666 39142 5678 39194
rect 5730 39142 5742 39194
rect 5794 39142 5806 39194
rect 5858 39142 14878 39194
rect 14930 39142 14942 39194
rect 14994 39142 15006 39194
rect 15058 39142 15070 39194
rect 15122 39142 24142 39194
rect 24194 39142 24206 39194
rect 24258 39142 24270 39194
rect 24322 39142 24334 39194
rect 24386 39142 28888 39194
rect 1104 39120 28888 39142
rect 2038 39040 2044 39092
rect 2096 39080 2102 39092
rect 2682 39080 2688 39092
rect 2096 39052 2688 39080
rect 2096 39040 2102 39052
rect 2682 39040 2688 39052
rect 2740 39040 2746 39092
rect 3237 39083 3295 39089
rect 3237 39049 3249 39083
rect 3283 39080 3295 39083
rect 3970 39080 3976 39092
rect 3283 39052 3976 39080
rect 3283 39049 3295 39052
rect 3237 39043 3295 39049
rect 3970 39040 3976 39052
rect 4028 39040 4034 39092
rect 5905 39083 5963 39089
rect 5905 39049 5917 39083
rect 5951 39080 5963 39083
rect 6178 39080 6184 39092
rect 5951 39052 6184 39080
rect 5951 39049 5963 39052
rect 5905 39043 5963 39049
rect 6178 39040 6184 39052
rect 6236 39040 6242 39092
rect 7745 39083 7803 39089
rect 7745 39049 7757 39083
rect 7791 39080 7803 39083
rect 8294 39080 8300 39092
rect 7791 39052 8300 39080
rect 7791 39049 7803 39052
rect 7745 39043 7803 39049
rect 8294 39040 8300 39052
rect 8352 39040 8358 39092
rect 8478 39080 8484 39092
rect 8439 39052 8484 39080
rect 8478 39040 8484 39052
rect 8536 39040 8542 39092
rect 9600 39052 12112 39080
rect 1854 39012 1860 39024
rect 1815 38984 1860 39012
rect 1854 38972 1860 38984
rect 1912 38972 1918 39024
rect 2590 38972 2596 39024
rect 2648 39012 2654 39024
rect 9600 39012 9628 39052
rect 11422 39012 11428 39024
rect 2648 38984 9628 39012
rect 10520 38984 11428 39012
rect 2648 38972 2654 38984
rect 1489 38947 1547 38953
rect 1489 38913 1501 38947
rect 1535 38944 1547 38947
rect 1578 38944 1584 38956
rect 1535 38916 1584 38944
rect 1535 38913 1547 38916
rect 1489 38907 1547 38913
rect 1578 38904 1584 38916
rect 1636 38904 1642 38956
rect 2038 38904 2044 38956
rect 2096 38944 2102 38956
rect 7285 38947 7343 38953
rect 2096 38916 5856 38944
rect 2096 38904 2102 38916
rect 3234 38876 3240 38888
rect 3195 38848 3240 38876
rect 3234 38836 3240 38848
rect 3292 38836 3298 38888
rect 3878 38836 3884 38888
rect 3936 38876 3942 38888
rect 4341 38879 4399 38885
rect 4341 38876 4353 38879
rect 3936 38848 4353 38876
rect 3936 38836 3942 38848
rect 4341 38845 4353 38848
rect 4387 38845 4399 38879
rect 4341 38839 4399 38845
rect 4433 38879 4491 38885
rect 4433 38845 4445 38879
rect 4479 38845 4491 38879
rect 4433 38839 4491 38845
rect 2961 38811 3019 38817
rect 2961 38777 2973 38811
rect 3007 38808 3019 38811
rect 3050 38808 3056 38820
rect 3007 38780 3056 38808
rect 3007 38777 3019 38780
rect 2961 38771 3019 38777
rect 3050 38768 3056 38780
rect 3108 38768 3114 38820
rect 3145 38811 3203 38817
rect 3145 38777 3157 38811
rect 3191 38808 3203 38811
rect 4448 38808 4476 38839
rect 4522 38836 4528 38888
rect 4580 38876 4586 38888
rect 4709 38879 4767 38885
rect 4580 38848 4625 38876
rect 4580 38836 4586 38848
rect 4709 38845 4721 38879
rect 4755 38876 4767 38879
rect 5169 38879 5227 38885
rect 5169 38876 5181 38879
rect 4755 38848 5181 38876
rect 4755 38845 4767 38848
rect 4709 38839 4767 38845
rect 5169 38845 5181 38848
rect 5215 38845 5227 38879
rect 5169 38839 5227 38845
rect 5258 38836 5264 38888
rect 5316 38876 5322 38888
rect 5828 38885 5856 38916
rect 7285 38913 7297 38947
rect 7331 38944 7343 38947
rect 8110 38944 8116 38956
rect 7331 38916 8116 38944
rect 7331 38913 7343 38916
rect 7285 38907 7343 38913
rect 5353 38879 5411 38885
rect 5353 38876 5365 38879
rect 5316 38848 5365 38876
rect 5316 38836 5322 38848
rect 5353 38845 5365 38848
rect 5399 38845 5411 38879
rect 5353 38839 5411 38845
rect 5813 38879 5871 38885
rect 5813 38845 5825 38879
rect 5859 38845 5871 38879
rect 5813 38839 5871 38845
rect 6825 38879 6883 38885
rect 6825 38845 6837 38879
rect 6871 38845 6883 38879
rect 6825 38839 6883 38845
rect 3191 38780 4476 38808
rect 6840 38808 6868 38839
rect 6914 38836 6920 38888
rect 6972 38876 6978 38888
rect 7009 38879 7067 38885
rect 7009 38876 7021 38879
rect 6972 38848 7021 38876
rect 6972 38836 6978 38848
rect 7009 38845 7021 38848
rect 7055 38845 7067 38879
rect 7742 38876 7748 38888
rect 7703 38848 7748 38876
rect 7009 38839 7067 38845
rect 7742 38836 7748 38848
rect 7800 38836 7806 38888
rect 7956 38885 7984 38916
rect 8110 38904 8116 38916
rect 8168 38904 8174 38956
rect 9674 38904 9680 38956
rect 9732 38944 9738 38956
rect 10520 38953 10548 38984
rect 11422 38972 11428 38984
rect 11480 38972 11486 39024
rect 11606 39012 11612 39024
rect 11567 38984 11612 39012
rect 11606 38972 11612 38984
rect 11664 38972 11670 39024
rect 12084 39012 12112 39052
rect 12158 39040 12164 39092
rect 12216 39080 12222 39092
rect 15654 39080 15660 39092
rect 12216 39052 15660 39080
rect 12216 39040 12222 39052
rect 15654 39040 15660 39052
rect 15712 39040 15718 39092
rect 22278 39080 22284 39092
rect 15764 39052 22284 39080
rect 15764 39012 15792 39052
rect 22278 39040 22284 39052
rect 22336 39040 22342 39092
rect 28074 39080 28080 39092
rect 22388 39052 28080 39080
rect 12084 38984 15792 39012
rect 16666 38972 16672 39024
rect 16724 38972 16730 39024
rect 18966 39012 18972 39024
rect 18927 38984 18972 39012
rect 18966 38972 18972 38984
rect 19024 38972 19030 39024
rect 9769 38947 9827 38953
rect 9769 38944 9781 38947
rect 9732 38916 9781 38944
rect 9732 38904 9738 38916
rect 9769 38913 9781 38916
rect 9815 38913 9827 38947
rect 10505 38947 10563 38953
rect 10505 38944 10517 38947
rect 9769 38907 9827 38913
rect 10428 38916 10517 38944
rect 7941 38879 7999 38885
rect 7941 38845 7953 38879
rect 7987 38845 7999 38879
rect 7941 38839 7999 38845
rect 8389 38879 8447 38885
rect 8389 38845 8401 38879
rect 8435 38845 8447 38879
rect 8389 38839 8447 38845
rect 7098 38808 7104 38820
rect 6840 38780 7104 38808
rect 3191 38777 3203 38780
rect 3145 38771 3203 38777
rect 4356 38752 4384 38780
rect 7098 38768 7104 38780
rect 7156 38768 7162 38820
rect 7760 38808 7788 38836
rect 8404 38808 8432 38839
rect 9858 38836 9864 38888
rect 9916 38876 9922 38888
rect 10045 38879 10103 38885
rect 9916 38848 9961 38876
rect 9916 38836 9922 38848
rect 10045 38845 10057 38879
rect 10091 38876 10103 38879
rect 10226 38876 10232 38888
rect 10091 38848 10232 38876
rect 10091 38845 10103 38848
rect 10045 38839 10103 38845
rect 10226 38836 10232 38848
rect 10284 38836 10290 38888
rect 7760 38780 8432 38808
rect 9582 38768 9588 38820
rect 9640 38808 9646 38820
rect 10428 38808 10456 38916
rect 10505 38913 10517 38916
rect 10551 38913 10563 38947
rect 10505 38907 10563 38913
rect 11238 38904 11244 38956
rect 11296 38904 11302 38956
rect 16684 38944 16712 38972
rect 16684 38916 16896 38944
rect 10965 38879 11023 38885
rect 10965 38876 10977 38879
rect 10796 38848 10977 38876
rect 9640 38780 10456 38808
rect 9640 38768 9646 38780
rect 10502 38768 10508 38820
rect 10560 38808 10566 38820
rect 10796 38808 10824 38848
rect 10965 38845 10977 38848
rect 11011 38845 11023 38879
rect 10965 38839 11023 38845
rect 11113 38879 11171 38885
rect 11113 38845 11125 38879
rect 11159 38876 11171 38879
rect 11256 38876 11284 38904
rect 11514 38885 11520 38888
rect 11159 38848 11284 38876
rect 11471 38879 11520 38885
rect 11159 38845 11171 38848
rect 11113 38839 11171 38845
rect 11471 38845 11483 38879
rect 11517 38845 11520 38879
rect 11471 38839 11520 38845
rect 11514 38836 11520 38839
rect 11572 38836 11578 38888
rect 12066 38876 12072 38888
rect 11624 38848 12072 38876
rect 10560 38780 10824 38808
rect 11241 38811 11299 38817
rect 10560 38768 10566 38780
rect 11241 38777 11253 38811
rect 11287 38777 11299 38811
rect 11241 38771 11299 38777
rect 11333 38811 11391 38817
rect 11333 38777 11345 38811
rect 11379 38808 11391 38811
rect 11624 38808 11652 38848
rect 12066 38836 12072 38848
rect 12124 38836 12130 38888
rect 14642 38836 14648 38888
rect 14700 38876 14706 38888
rect 14921 38879 14979 38885
rect 14921 38876 14933 38879
rect 14700 38848 14933 38876
rect 14700 38836 14706 38848
rect 14921 38845 14933 38848
rect 14967 38845 14979 38879
rect 14921 38839 14979 38845
rect 16574 38836 16580 38888
rect 16632 38885 16638 38888
rect 16632 38879 16681 38885
rect 16632 38845 16635 38879
rect 16669 38845 16681 38879
rect 16758 38876 16764 38888
rect 16719 38848 16764 38876
rect 16632 38839 16681 38845
rect 16632 38836 16638 38839
rect 16758 38836 16764 38848
rect 16816 38836 16822 38888
rect 16868 38885 16896 38916
rect 17144 38916 17724 38944
rect 16853 38879 16911 38885
rect 16853 38845 16865 38879
rect 16899 38845 16911 38879
rect 17034 38876 17040 38888
rect 16995 38848 17040 38876
rect 16853 38839 16911 38845
rect 17034 38836 17040 38848
rect 17092 38836 17098 38888
rect 11379 38780 11652 38808
rect 11379 38777 11391 38780
rect 11333 38771 11391 38777
rect 1949 38743 2007 38749
rect 1949 38709 1961 38743
rect 1995 38740 2007 38743
rect 3878 38740 3884 38752
rect 1995 38712 3884 38740
rect 1995 38709 2007 38712
rect 1949 38703 2007 38709
rect 3878 38700 3884 38712
rect 3936 38700 3942 38752
rect 4338 38700 4344 38752
rect 4396 38700 4402 38752
rect 4798 38700 4804 38752
rect 4856 38740 4862 38752
rect 5261 38743 5319 38749
rect 5261 38740 5273 38743
rect 4856 38712 5273 38740
rect 4856 38700 4862 38712
rect 5261 38709 5273 38712
rect 5307 38709 5319 38743
rect 11256 38740 11284 38771
rect 11698 38768 11704 38820
rect 11756 38808 11762 38820
rect 17144 38808 17172 38916
rect 17218 38836 17224 38888
rect 17276 38876 17282 38888
rect 17589 38879 17647 38885
rect 17589 38876 17601 38879
rect 17276 38848 17601 38876
rect 17276 38836 17282 38848
rect 17589 38845 17601 38848
rect 17635 38845 17647 38879
rect 17696 38876 17724 38916
rect 22388 38876 22416 39052
rect 28074 39040 28080 39052
rect 28132 39040 28138 39092
rect 25869 39015 25927 39021
rect 25869 38981 25881 39015
rect 25915 38981 25927 39015
rect 25869 38975 25927 38981
rect 26513 39015 26571 39021
rect 26513 38981 26525 39015
rect 26559 39012 26571 39015
rect 27798 39012 27804 39024
rect 26559 38984 27804 39012
rect 26559 38981 26571 38984
rect 26513 38975 26571 38981
rect 22462 38904 22468 38956
rect 22520 38944 22526 38956
rect 25884 38944 25912 38975
rect 27798 38972 27804 38984
rect 27856 38972 27862 39024
rect 28166 39012 28172 39024
rect 28127 38984 28172 39012
rect 28166 38972 28172 38984
rect 28224 38972 28230 39024
rect 22520 38916 25636 38944
rect 25884 38916 28028 38944
rect 22520 38904 22526 38916
rect 17696 38848 22416 38876
rect 22557 38879 22615 38885
rect 17589 38839 17647 38845
rect 22557 38845 22569 38879
rect 22603 38876 22615 38879
rect 22646 38876 22652 38888
rect 22603 38848 22652 38876
rect 22603 38845 22615 38848
rect 22557 38839 22615 38845
rect 22646 38836 22652 38848
rect 22704 38836 22710 38888
rect 22741 38879 22799 38885
rect 22741 38845 22753 38879
rect 22787 38876 22799 38879
rect 22787 38848 25544 38876
rect 22787 38845 22799 38848
rect 22741 38839 22799 38845
rect 11756 38780 17172 38808
rect 11756 38768 11762 38780
rect 17402 38768 17408 38820
rect 17460 38808 17466 38820
rect 17834 38811 17892 38817
rect 17834 38808 17846 38811
rect 17460 38780 17846 38808
rect 17460 38768 17466 38780
rect 17834 38777 17846 38780
rect 17880 38777 17892 38811
rect 22756 38808 22784 38839
rect 17834 38771 17892 38777
rect 22066 38780 22784 38808
rect 11606 38740 11612 38752
rect 11256 38712 11612 38740
rect 5261 38703 5319 38709
rect 11606 38700 11612 38712
rect 11664 38700 11670 38752
rect 11974 38700 11980 38752
rect 12032 38740 12038 38752
rect 12526 38740 12532 38752
rect 12032 38712 12532 38740
rect 12032 38700 12038 38712
rect 12526 38700 12532 38712
rect 12584 38700 12590 38752
rect 14734 38740 14740 38752
rect 14695 38712 14740 38740
rect 14734 38700 14740 38712
rect 14792 38700 14798 38752
rect 16390 38740 16396 38752
rect 16351 38712 16396 38740
rect 16390 38700 16396 38712
rect 16448 38700 16454 38752
rect 20162 38700 20168 38752
rect 20220 38740 20226 38752
rect 22066 38740 22094 38780
rect 25516 38752 25544 38848
rect 25608 38808 25636 38916
rect 26050 38876 26056 38888
rect 26011 38848 26056 38876
rect 26050 38836 26056 38848
rect 26108 38836 26114 38888
rect 26697 38879 26755 38885
rect 26697 38845 26709 38879
rect 26743 38876 26755 38879
rect 26786 38876 26792 38888
rect 26743 38848 26792 38876
rect 26743 38845 26755 38848
rect 26697 38839 26755 38845
rect 26786 38836 26792 38848
rect 26844 38836 26850 38888
rect 27246 38876 27252 38888
rect 27207 38848 27252 38876
rect 27246 38836 27252 38848
rect 27304 38836 27310 38888
rect 28000 38885 28028 38916
rect 27985 38879 28043 38885
rect 27985 38845 27997 38879
rect 28031 38845 28043 38879
rect 27985 38839 28043 38845
rect 27433 38811 27491 38817
rect 27433 38808 27445 38811
rect 25608 38780 27445 38808
rect 27433 38777 27445 38780
rect 27479 38777 27491 38811
rect 27433 38771 27491 38777
rect 22738 38740 22744 38752
rect 20220 38712 22094 38740
rect 22699 38712 22744 38740
rect 20220 38700 20226 38712
rect 22738 38700 22744 38712
rect 22796 38700 22802 38752
rect 25498 38700 25504 38752
rect 25556 38740 25562 38752
rect 25866 38740 25872 38752
rect 25556 38712 25872 38740
rect 25556 38700 25562 38712
rect 25866 38700 25872 38712
rect 25924 38700 25930 38752
rect 1104 38650 28888 38672
rect 1104 38598 10246 38650
rect 10298 38598 10310 38650
rect 10362 38598 10374 38650
rect 10426 38598 10438 38650
rect 10490 38598 19510 38650
rect 19562 38598 19574 38650
rect 19626 38598 19638 38650
rect 19690 38598 19702 38650
rect 19754 38598 28888 38650
rect 1104 38576 28888 38598
rect 19521 38539 19579 38545
rect 19521 38536 19533 38539
rect 2700 38508 19533 38536
rect 1673 38471 1731 38477
rect 1673 38437 1685 38471
rect 1719 38468 1731 38471
rect 1854 38468 1860 38480
rect 1719 38440 1860 38468
rect 1719 38437 1731 38440
rect 1673 38431 1731 38437
rect 1854 38428 1860 38440
rect 1912 38428 1918 38480
rect 2700 38477 2728 38508
rect 19521 38505 19533 38508
rect 19567 38505 19579 38539
rect 20070 38536 20076 38548
rect 20031 38508 20076 38536
rect 19521 38499 19579 38505
rect 20070 38496 20076 38508
rect 20128 38496 20134 38548
rect 28074 38536 28080 38548
rect 20180 38508 28080 38536
rect 2685 38471 2743 38477
rect 2685 38437 2697 38471
rect 2731 38437 2743 38471
rect 2685 38431 2743 38437
rect 3050 38428 3056 38480
rect 3108 38468 3114 38480
rect 4154 38468 4160 38480
rect 3108 38440 3832 38468
rect 3108 38428 3114 38440
rect 2590 38360 2596 38412
rect 2648 38400 2654 38412
rect 3068 38400 3096 38428
rect 2648 38372 3096 38400
rect 3605 38403 3663 38409
rect 2648 38360 2654 38372
rect 3605 38369 3617 38403
rect 3651 38400 3663 38403
rect 3651 38372 3740 38400
rect 3651 38369 3663 38372
rect 3605 38363 3663 38369
rect 1578 38224 1584 38276
rect 1636 38264 1642 38276
rect 1949 38267 2007 38273
rect 1949 38264 1961 38267
rect 1636 38236 1961 38264
rect 1636 38224 1642 38236
rect 1949 38233 1961 38236
rect 1995 38233 2007 38267
rect 1949 38227 2007 38233
rect 2133 38199 2191 38205
rect 2133 38165 2145 38199
rect 2179 38196 2191 38199
rect 2222 38196 2228 38208
rect 2179 38168 2228 38196
rect 2179 38165 2191 38168
rect 2133 38159 2191 38165
rect 2222 38156 2228 38168
rect 2280 38156 2286 38208
rect 2774 38156 2780 38208
rect 2832 38196 2838 38208
rect 3712 38196 3740 38372
rect 3804 38264 3832 38440
rect 3988 38440 4160 38468
rect 3988 38409 4016 38440
rect 4154 38428 4160 38440
rect 4212 38428 4218 38480
rect 4522 38468 4528 38480
rect 4483 38440 4528 38468
rect 4522 38428 4528 38440
rect 4580 38428 4586 38480
rect 5074 38428 5080 38480
rect 5132 38468 5138 38480
rect 5721 38471 5779 38477
rect 5721 38468 5733 38471
rect 5132 38440 5733 38468
rect 5132 38428 5138 38440
rect 5721 38437 5733 38440
rect 5767 38437 5779 38471
rect 5721 38431 5779 38437
rect 9490 38428 9496 38480
rect 9548 38468 9554 38480
rect 9674 38468 9680 38480
rect 9548 38440 9680 38468
rect 9548 38428 9554 38440
rect 9674 38428 9680 38440
rect 9732 38428 9738 38480
rect 10689 38471 10747 38477
rect 10689 38437 10701 38471
rect 10735 38468 10747 38471
rect 11514 38468 11520 38480
rect 10735 38440 11520 38468
rect 10735 38437 10747 38440
rect 10689 38431 10747 38437
rect 11514 38428 11520 38440
rect 11572 38428 11578 38480
rect 12406 38440 16344 38468
rect 3973 38403 4031 38409
rect 3973 38369 3985 38403
rect 4019 38369 4031 38403
rect 3973 38363 4031 38369
rect 4341 38403 4399 38409
rect 4341 38369 4353 38403
rect 4387 38400 4399 38403
rect 4614 38400 4620 38412
rect 4387 38372 4620 38400
rect 4387 38369 4399 38372
rect 4341 38363 4399 38369
rect 4614 38360 4620 38372
rect 4672 38360 4678 38412
rect 4985 38403 5043 38409
rect 4985 38369 4997 38403
rect 5031 38369 5043 38403
rect 4985 38363 5043 38369
rect 5629 38403 5687 38409
rect 5629 38369 5641 38403
rect 5675 38400 5687 38403
rect 5902 38400 5908 38412
rect 5675 38372 5908 38400
rect 5675 38369 5687 38372
rect 5629 38363 5687 38369
rect 3878 38292 3884 38344
rect 3936 38332 3942 38344
rect 5000 38332 5028 38363
rect 5902 38360 5908 38372
rect 5960 38360 5966 38412
rect 8846 38360 8852 38412
rect 8904 38400 8910 38412
rect 8941 38403 8999 38409
rect 8941 38400 8953 38403
rect 8904 38372 8953 38400
rect 8904 38360 8910 38372
rect 8941 38369 8953 38372
rect 8987 38369 8999 38403
rect 8941 38363 8999 38369
rect 10413 38403 10471 38409
rect 10413 38369 10425 38403
rect 10459 38369 10471 38403
rect 10413 38363 10471 38369
rect 9030 38332 9036 38344
rect 3936 38304 5028 38332
rect 8991 38304 9036 38332
rect 3936 38292 3942 38304
rect 9030 38292 9036 38304
rect 9088 38292 9094 38344
rect 9214 38332 9220 38344
rect 9175 38304 9220 38332
rect 9214 38292 9220 38304
rect 9272 38292 9278 38344
rect 9398 38292 9404 38344
rect 9456 38332 9462 38344
rect 10428 38332 10456 38363
rect 10502 38360 10508 38412
rect 10560 38400 10566 38412
rect 10778 38400 10784 38412
rect 10560 38372 10605 38400
rect 10739 38372 10784 38400
rect 10560 38360 10566 38372
rect 10778 38360 10784 38372
rect 10836 38360 10842 38412
rect 10870 38360 10876 38412
rect 10928 38409 10934 38412
rect 10928 38400 10936 38409
rect 12406 38400 12434 38440
rect 10928 38372 10973 38400
rect 11532 38372 12434 38400
rect 10928 38363 10936 38372
rect 10928 38360 10934 38363
rect 11422 38332 11428 38344
rect 9456 38304 9996 38332
rect 10428 38304 11428 38332
rect 9456 38292 9462 38304
rect 5077 38267 5135 38273
rect 5077 38264 5089 38267
rect 3804 38236 5089 38264
rect 5077 38233 5089 38236
rect 5123 38233 5135 38267
rect 5077 38227 5135 38233
rect 8573 38267 8631 38273
rect 8573 38233 8585 38267
rect 8619 38264 8631 38267
rect 9858 38264 9864 38276
rect 8619 38236 9864 38264
rect 8619 38233 8631 38236
rect 8573 38227 8631 38233
rect 9858 38224 9864 38236
rect 9916 38224 9922 38276
rect 9968 38264 9996 38304
rect 11422 38292 11428 38304
rect 11480 38292 11486 38344
rect 11532 38264 11560 38372
rect 13262 38360 13268 38412
rect 13320 38400 13326 38412
rect 13429 38403 13487 38409
rect 13429 38400 13441 38403
rect 13320 38372 13441 38400
rect 13320 38360 13326 38372
rect 13429 38369 13441 38372
rect 13475 38369 13487 38403
rect 13429 38363 13487 38369
rect 15105 38403 15163 38409
rect 15105 38369 15117 38403
rect 15151 38400 15163 38403
rect 15286 38400 15292 38412
rect 15151 38372 15292 38400
rect 15151 38369 15163 38372
rect 15105 38363 15163 38369
rect 15286 38360 15292 38372
rect 15344 38360 15350 38412
rect 16316 38400 16344 38440
rect 16390 38428 16396 38480
rect 16448 38468 16454 38480
rect 17558 38471 17616 38477
rect 17558 38468 17570 38471
rect 16448 38440 17570 38468
rect 16448 38428 16454 38440
rect 17558 38437 17570 38440
rect 17604 38437 17616 38471
rect 20180 38468 20208 38508
rect 28074 38496 28080 38508
rect 28132 38496 28138 38548
rect 27246 38468 27252 38480
rect 17558 38431 17616 38437
rect 18432 38440 20208 38468
rect 20272 38440 27252 38468
rect 18432 38400 18460 38440
rect 19981 38403 20039 38409
rect 19981 38400 19993 38403
rect 16316 38372 18460 38400
rect 18984 38372 19993 38400
rect 11974 38292 11980 38344
rect 12032 38332 12038 38344
rect 13173 38335 13231 38341
rect 13173 38332 13185 38335
rect 12032 38304 13185 38332
rect 12032 38292 12038 38304
rect 13173 38301 13185 38304
rect 13219 38301 13231 38335
rect 13173 38295 13231 38301
rect 17218 38292 17224 38344
rect 17276 38332 17282 38344
rect 17313 38335 17371 38341
rect 17313 38332 17325 38335
rect 17276 38304 17325 38332
rect 17276 38292 17282 38304
rect 17313 38301 17325 38304
rect 17359 38301 17371 38335
rect 17313 38295 17371 38301
rect 18414 38292 18420 38344
rect 18472 38332 18478 38344
rect 18984 38332 19012 38372
rect 19981 38369 19993 38372
rect 20027 38369 20039 38403
rect 20272 38400 20300 38440
rect 27246 38428 27252 38440
rect 27304 38428 27310 38480
rect 27890 38468 27896 38480
rect 27851 38440 27896 38468
rect 27890 38428 27896 38440
rect 27948 38428 27954 38480
rect 19981 38363 20039 38369
rect 20088 38372 20300 38400
rect 20809 38403 20867 38409
rect 18472 38304 19012 38332
rect 19521 38335 19579 38341
rect 18472 38292 18478 38304
rect 19521 38301 19533 38335
rect 19567 38332 19579 38335
rect 20088 38332 20116 38372
rect 20809 38369 20821 38403
rect 20855 38400 20867 38403
rect 20898 38400 20904 38412
rect 20855 38372 20904 38400
rect 20855 38369 20867 38372
rect 20809 38363 20867 38369
rect 20898 38360 20904 38372
rect 20956 38360 20962 38412
rect 20993 38403 21051 38409
rect 20993 38369 21005 38403
rect 21039 38369 21051 38403
rect 20993 38363 21051 38369
rect 19567 38304 20116 38332
rect 20257 38335 20315 38341
rect 19567 38301 19579 38304
rect 19521 38295 19579 38301
rect 20257 38301 20269 38335
rect 20303 38332 20315 38335
rect 20346 38332 20352 38344
rect 20303 38304 20352 38332
rect 20303 38301 20315 38304
rect 20257 38295 20315 38301
rect 20346 38292 20352 38304
rect 20404 38292 20410 38344
rect 21008 38332 21036 38363
rect 21266 38360 21272 38412
rect 21324 38400 21330 38412
rect 22925 38403 22983 38409
rect 22925 38400 22937 38403
rect 21324 38372 22937 38400
rect 21324 38360 21330 38372
rect 22925 38369 22937 38372
rect 22971 38369 22983 38403
rect 22925 38363 22983 38369
rect 24480 38403 24538 38409
rect 24480 38369 24492 38403
rect 24526 38400 24538 38403
rect 25038 38400 25044 38412
rect 24526 38372 25044 38400
rect 24526 38369 24538 38372
rect 24480 38363 24538 38369
rect 25038 38360 25044 38372
rect 25096 38360 25102 38412
rect 26142 38360 26148 38412
rect 26200 38400 26206 38412
rect 26237 38403 26295 38409
rect 26237 38400 26249 38403
rect 26200 38372 26249 38400
rect 26200 38360 26206 38372
rect 26237 38369 26249 38372
rect 26283 38369 26295 38403
rect 26878 38400 26884 38412
rect 26839 38372 26884 38400
rect 26237 38363 26295 38369
rect 26878 38360 26884 38372
rect 26936 38360 26942 38412
rect 20916 38304 21036 38332
rect 9968 38236 11560 38264
rect 18782 38224 18788 38276
rect 18840 38264 18846 38276
rect 20916 38264 20944 38304
rect 22186 38292 22192 38344
rect 22244 38332 22250 38344
rect 23017 38335 23075 38341
rect 23017 38332 23029 38335
rect 22244 38304 23029 38332
rect 22244 38292 22250 38304
rect 23017 38301 23029 38304
rect 23063 38301 23075 38335
rect 23017 38295 23075 38301
rect 23109 38335 23167 38341
rect 23109 38301 23121 38335
rect 23155 38301 23167 38335
rect 23109 38295 23167 38301
rect 24213 38335 24271 38341
rect 24213 38301 24225 38335
rect 24259 38301 24271 38335
rect 24213 38295 24271 38301
rect 21358 38264 21364 38276
rect 18840 38236 21364 38264
rect 18840 38224 18846 38236
rect 21358 38224 21364 38236
rect 21416 38224 21422 38276
rect 22646 38224 22652 38276
rect 22704 38264 22710 38276
rect 23124 38264 23152 38295
rect 22704 38236 23152 38264
rect 22704 38224 22710 38236
rect 4154 38196 4160 38208
rect 2832 38168 2877 38196
rect 3712 38168 4160 38196
rect 2832 38156 2838 38168
rect 4154 38156 4160 38168
rect 4212 38156 4218 38208
rect 4522 38156 4528 38208
rect 4580 38196 4586 38208
rect 5350 38196 5356 38208
rect 4580 38168 5356 38196
rect 4580 38156 4586 38168
rect 5350 38156 5356 38168
rect 5408 38156 5414 38208
rect 6178 38156 6184 38208
rect 6236 38196 6242 38208
rect 11057 38199 11115 38205
rect 11057 38196 11069 38199
rect 6236 38168 11069 38196
rect 6236 38156 6242 38168
rect 11057 38165 11069 38168
rect 11103 38165 11115 38199
rect 11057 38159 11115 38165
rect 11330 38156 11336 38208
rect 11388 38196 11394 38208
rect 12066 38196 12072 38208
rect 11388 38168 12072 38196
rect 11388 38156 11394 38168
rect 12066 38156 12072 38168
rect 12124 38156 12130 38208
rect 13538 38156 13544 38208
rect 13596 38196 13602 38208
rect 14366 38196 14372 38208
rect 13596 38168 14372 38196
rect 13596 38156 13602 38168
rect 14366 38156 14372 38168
rect 14424 38196 14430 38208
rect 14553 38199 14611 38205
rect 14553 38196 14565 38199
rect 14424 38168 14565 38196
rect 14424 38156 14430 38168
rect 14553 38165 14565 38168
rect 14599 38165 14611 38199
rect 15194 38196 15200 38208
rect 15155 38168 15200 38196
rect 14553 38159 14611 38165
rect 15194 38156 15200 38168
rect 15252 38156 15258 38208
rect 17954 38156 17960 38208
rect 18012 38196 18018 38208
rect 18693 38199 18751 38205
rect 18693 38196 18705 38199
rect 18012 38168 18705 38196
rect 18012 38156 18018 38168
rect 18693 38165 18705 38168
rect 18739 38165 18751 38199
rect 18693 38159 18751 38165
rect 19613 38199 19671 38205
rect 19613 38165 19625 38199
rect 19659 38196 19671 38199
rect 20438 38196 20444 38208
rect 19659 38168 20444 38196
rect 19659 38165 19671 38168
rect 19613 38159 19671 38165
rect 20438 38156 20444 38168
rect 20496 38156 20502 38208
rect 21082 38156 21088 38208
rect 21140 38196 21146 38208
rect 21177 38199 21235 38205
rect 21177 38196 21189 38199
rect 21140 38168 21189 38196
rect 21140 38156 21146 38168
rect 21177 38165 21189 38168
rect 21223 38165 21235 38199
rect 21177 38159 21235 38165
rect 22557 38199 22615 38205
rect 22557 38165 22569 38199
rect 22603 38196 22615 38199
rect 23106 38196 23112 38208
rect 22603 38168 23112 38196
rect 22603 38165 22615 38168
rect 22557 38159 22615 38165
rect 23106 38156 23112 38168
rect 23164 38156 23170 38208
rect 23198 38156 23204 38208
rect 23256 38196 23262 38208
rect 24228 38196 24256 38295
rect 24854 38196 24860 38208
rect 23256 38168 24860 38196
rect 23256 38156 23262 38168
rect 24854 38156 24860 38168
rect 24912 38196 24918 38208
rect 25314 38196 25320 38208
rect 24912 38168 25320 38196
rect 24912 38156 24918 38168
rect 25314 38156 25320 38168
rect 25372 38156 25378 38208
rect 25593 38199 25651 38205
rect 25593 38165 25605 38199
rect 25639 38196 25651 38199
rect 25866 38196 25872 38208
rect 25639 38168 25872 38196
rect 25639 38165 25651 38168
rect 25593 38159 25651 38165
rect 25866 38156 25872 38168
rect 25924 38156 25930 38208
rect 26050 38196 26056 38208
rect 26011 38168 26056 38196
rect 26050 38156 26056 38168
rect 26108 38156 26114 38208
rect 26694 38196 26700 38208
rect 26655 38168 26700 38196
rect 26694 38156 26700 38168
rect 26752 38156 26758 38208
rect 27982 38196 27988 38208
rect 27943 38168 27988 38196
rect 27982 38156 27988 38168
rect 28040 38156 28046 38208
rect 1104 38106 28888 38128
rect 1104 38054 5614 38106
rect 5666 38054 5678 38106
rect 5730 38054 5742 38106
rect 5794 38054 5806 38106
rect 5858 38054 14878 38106
rect 14930 38054 14942 38106
rect 14994 38054 15006 38106
rect 15058 38054 15070 38106
rect 15122 38054 24142 38106
rect 24194 38054 24206 38106
rect 24258 38054 24270 38106
rect 24322 38054 24334 38106
rect 24386 38054 28888 38106
rect 1104 38032 28888 38054
rect 2866 37952 2872 38004
rect 2924 37992 2930 38004
rect 2924 37964 3188 37992
rect 2924 37952 2930 37964
rect 2501 37927 2559 37933
rect 2501 37893 2513 37927
rect 2547 37924 2559 37927
rect 3160 37924 3188 37964
rect 3234 37952 3240 38004
rect 3292 37992 3298 38004
rect 4341 37995 4399 38001
rect 4341 37992 4353 37995
rect 3292 37964 4353 37992
rect 3292 37952 3298 37964
rect 4341 37961 4353 37964
rect 4387 37961 4399 37995
rect 22186 37992 22192 38004
rect 4341 37955 4399 37961
rect 4448 37964 22094 37992
rect 22147 37964 22192 37992
rect 4448 37924 4476 37964
rect 2547 37896 3096 37924
rect 3160 37896 4476 37924
rect 2547 37893 2559 37896
rect 2501 37887 2559 37893
rect 1394 37816 1400 37868
rect 1452 37856 1458 37868
rect 1578 37856 1584 37868
rect 1452 37828 1584 37856
rect 1452 37816 1458 37828
rect 1578 37816 1584 37828
rect 1636 37816 1642 37868
rect 3068 37856 3096 37896
rect 13354 37884 13360 37936
rect 13412 37924 13418 37936
rect 16117 37927 16175 37933
rect 16117 37924 16129 37927
rect 13412 37896 16129 37924
rect 13412 37884 13418 37896
rect 16117 37893 16129 37896
rect 16163 37893 16175 37927
rect 16117 37887 16175 37893
rect 16666 37884 16672 37936
rect 16724 37924 16730 37936
rect 16853 37927 16911 37933
rect 16853 37924 16865 37927
rect 16724 37896 16865 37924
rect 16724 37884 16730 37896
rect 16853 37893 16865 37896
rect 16899 37893 16911 37927
rect 16853 37887 16911 37893
rect 20070 37884 20076 37936
rect 20128 37924 20134 37936
rect 20346 37924 20352 37936
rect 20128 37896 20352 37924
rect 20128 37884 20134 37896
rect 20346 37884 20352 37896
rect 20404 37884 20410 37936
rect 22066 37924 22094 37964
rect 22186 37952 22192 37964
rect 22244 37952 22250 38004
rect 27246 37992 27252 38004
rect 27207 37964 27252 37992
rect 27246 37952 27252 37964
rect 27304 37952 27310 38004
rect 27982 37924 27988 37936
rect 22066 37896 27988 37924
rect 27982 37884 27988 37896
rect 28040 37884 28046 37936
rect 4154 37856 4160 37868
rect 3068 37828 4160 37856
rect 4154 37816 4160 37828
rect 4212 37816 4218 37868
rect 11606 37816 11612 37868
rect 11664 37856 11670 37868
rect 16022 37856 16028 37868
rect 11664 37828 12112 37856
rect 11664 37816 11670 37828
rect 2222 37748 2228 37800
rect 2280 37788 2286 37800
rect 2409 37791 2467 37797
rect 2409 37788 2421 37791
rect 2280 37760 2421 37788
rect 2280 37748 2286 37760
rect 2409 37757 2421 37760
rect 2455 37757 2467 37791
rect 2409 37751 2467 37757
rect 1578 37720 1584 37732
rect 1539 37692 1584 37720
rect 1578 37680 1584 37692
rect 1636 37680 1642 37732
rect 2424 37720 2452 37751
rect 2590 37748 2596 37800
rect 2648 37788 2654 37800
rect 2777 37791 2835 37797
rect 2777 37788 2789 37791
rect 2648 37760 2789 37788
rect 2648 37748 2654 37760
rect 2777 37757 2789 37760
rect 2823 37757 2835 37791
rect 2777 37751 2835 37757
rect 3142 37748 3148 37800
rect 3200 37788 3206 37800
rect 4246 37788 4252 37800
rect 3200 37760 3245 37788
rect 4207 37760 4252 37788
rect 3200 37748 3206 37760
rect 4246 37748 4252 37760
rect 4304 37748 4310 37800
rect 4433 37791 4491 37797
rect 4433 37757 4445 37791
rect 4479 37757 4491 37791
rect 4433 37751 4491 37757
rect 5077 37791 5135 37797
rect 5077 37757 5089 37791
rect 5123 37788 5135 37791
rect 5902 37788 5908 37800
rect 5123 37760 5908 37788
rect 5123 37757 5135 37760
rect 5077 37751 5135 37757
rect 3050 37720 3056 37732
rect 2424 37692 3056 37720
rect 3050 37680 3056 37692
rect 3108 37680 3114 37732
rect 1670 37652 1676 37664
rect 1631 37624 1676 37652
rect 1670 37612 1676 37624
rect 1728 37612 1734 37664
rect 2498 37612 2504 37664
rect 2556 37652 2562 37664
rect 2866 37652 2872 37664
rect 2556 37624 2872 37652
rect 2556 37612 2562 37624
rect 2866 37612 2872 37624
rect 2924 37612 2930 37664
rect 3418 37612 3424 37664
rect 3476 37652 3482 37664
rect 4448 37652 4476 37751
rect 5902 37748 5908 37760
rect 5960 37748 5966 37800
rect 10137 37791 10195 37797
rect 10137 37757 10149 37791
rect 10183 37788 10195 37791
rect 11146 37788 11152 37800
rect 10183 37760 11152 37788
rect 10183 37757 10195 37760
rect 10137 37751 10195 37757
rect 11146 37748 11152 37760
rect 11204 37788 11210 37800
rect 11974 37788 11980 37800
rect 11204 37760 11980 37788
rect 11204 37748 11210 37760
rect 11974 37748 11980 37760
rect 12032 37748 12038 37800
rect 12084 37788 12112 37828
rect 15856 37828 16028 37856
rect 12084 37760 12434 37788
rect 5350 37729 5356 37732
rect 5344 37683 5356 37729
rect 5408 37720 5414 37732
rect 5408 37692 5444 37720
rect 5350 37680 5356 37683
rect 5408 37680 5414 37692
rect 9950 37680 9956 37732
rect 10008 37720 10014 37732
rect 10226 37720 10232 37732
rect 10008 37692 10232 37720
rect 10008 37680 10014 37692
rect 10226 37680 10232 37692
rect 10284 37680 10290 37732
rect 10404 37723 10462 37729
rect 10404 37689 10416 37723
rect 10450 37720 10462 37723
rect 10962 37720 10968 37732
rect 10450 37692 10968 37720
rect 10450 37689 10462 37692
rect 10404 37683 10462 37689
rect 10962 37680 10968 37692
rect 11020 37680 11026 37732
rect 12066 37680 12072 37732
rect 12124 37720 12130 37732
rect 12222 37723 12280 37729
rect 12222 37720 12234 37723
rect 12124 37692 12234 37720
rect 12124 37680 12130 37692
rect 12222 37689 12234 37692
rect 12268 37689 12280 37723
rect 12222 37683 12280 37689
rect 12406 37664 12434 37760
rect 13354 37748 13360 37800
rect 13412 37788 13418 37800
rect 13722 37788 13728 37800
rect 13412 37760 13728 37788
rect 13412 37748 13418 37760
rect 13722 37748 13728 37760
rect 13780 37748 13786 37800
rect 13998 37748 14004 37800
rect 14056 37788 14062 37800
rect 14734 37788 14740 37800
rect 14056 37760 14740 37788
rect 14056 37748 14062 37760
rect 14734 37748 14740 37760
rect 14792 37748 14798 37800
rect 15378 37748 15384 37800
rect 15436 37788 15442 37800
rect 15654 37797 15660 37800
rect 15473 37791 15531 37797
rect 15473 37788 15485 37791
rect 15436 37760 15485 37788
rect 15436 37748 15442 37760
rect 15473 37757 15485 37760
rect 15519 37757 15531 37791
rect 15473 37751 15531 37757
rect 15621 37791 15660 37797
rect 15621 37757 15633 37791
rect 15621 37751 15660 37757
rect 15654 37748 15660 37751
rect 15712 37748 15718 37800
rect 15856 37797 15884 37828
rect 16022 37816 16028 37828
rect 16080 37816 16086 37868
rect 18598 37816 18604 37868
rect 18656 37856 18662 37868
rect 20806 37856 20812 37868
rect 18656 37828 20812 37856
rect 18656 37816 18662 37828
rect 20806 37816 20812 37828
rect 20864 37816 20870 37868
rect 22738 37816 22744 37868
rect 22796 37856 22802 37868
rect 23017 37859 23075 37865
rect 23017 37856 23029 37859
rect 22796 37828 23029 37856
rect 22796 37816 22802 37828
rect 23017 37825 23029 37828
rect 23063 37825 23075 37859
rect 25866 37856 25872 37868
rect 25827 37828 25872 37856
rect 23017 37819 23075 37825
rect 25866 37816 25872 37828
rect 25924 37816 25930 37868
rect 25958 37816 25964 37868
rect 26016 37856 26022 37868
rect 26016 37828 26061 37856
rect 26016 37816 26022 37828
rect 15841 37791 15899 37797
rect 15841 37757 15853 37791
rect 15887 37757 15899 37791
rect 15841 37751 15899 37757
rect 15930 37748 15936 37800
rect 15988 37797 15994 37800
rect 15988 37788 15996 37797
rect 16574 37788 16580 37800
rect 15988 37760 16033 37788
rect 16408 37760 16580 37788
rect 15988 37751 15996 37760
rect 15988 37748 15994 37751
rect 14826 37720 14832 37732
rect 14787 37692 14832 37720
rect 14826 37680 14832 37692
rect 14884 37680 14890 37732
rect 15749 37723 15807 37729
rect 15749 37689 15761 37723
rect 15795 37720 15807 37723
rect 16408 37720 16436 37760
rect 16574 37748 16580 37760
rect 16632 37748 16638 37800
rect 20070 37788 20076 37800
rect 20031 37760 20076 37788
rect 20070 37748 20076 37760
rect 20128 37748 20134 37800
rect 20162 37748 20168 37800
rect 20220 37788 20226 37800
rect 21082 37797 21088 37800
rect 20257 37791 20315 37797
rect 20257 37788 20269 37791
rect 20220 37760 20269 37788
rect 20220 37748 20226 37760
rect 20257 37757 20269 37760
rect 20303 37757 20315 37791
rect 21076 37788 21088 37797
rect 21043 37760 21088 37788
rect 20257 37751 20315 37757
rect 21076 37751 21088 37760
rect 21082 37748 21088 37751
rect 21140 37748 21146 37800
rect 23106 37748 23112 37800
rect 23164 37788 23170 37800
rect 23293 37791 23351 37797
rect 23164 37760 23209 37788
rect 23164 37748 23170 37760
rect 23293 37757 23305 37791
rect 23339 37788 23351 37791
rect 24026 37788 24032 37800
rect 23339 37760 24032 37788
rect 23339 37757 23351 37760
rect 23293 37751 23351 37757
rect 24026 37748 24032 37760
rect 24084 37748 24090 37800
rect 26050 37748 26056 37800
rect 26108 37788 26114 37800
rect 27157 37791 27215 37797
rect 27157 37788 27169 37791
rect 26108 37760 27169 37788
rect 26108 37748 26114 37760
rect 27157 37757 27169 37760
rect 27203 37757 27215 37791
rect 27157 37751 27215 37757
rect 27798 37748 27804 37800
rect 27856 37788 27862 37800
rect 27893 37791 27951 37797
rect 27893 37788 27905 37791
rect 27856 37760 27905 37788
rect 27856 37748 27862 37760
rect 27893 37757 27905 37760
rect 27939 37757 27951 37791
rect 27893 37751 27951 37757
rect 15795 37692 16436 37720
rect 15795 37689 15807 37692
rect 15749 37683 15807 37689
rect 16482 37680 16488 37732
rect 16540 37720 16546 37732
rect 16669 37723 16727 37729
rect 16669 37720 16681 37723
rect 16540 37692 16681 37720
rect 16540 37680 16546 37692
rect 16669 37689 16681 37692
rect 16715 37689 16727 37723
rect 16669 37683 16727 37689
rect 23753 37723 23811 37729
rect 23753 37689 23765 37723
rect 23799 37720 23811 37723
rect 25314 37720 25320 37732
rect 23799 37692 25320 37720
rect 23799 37689 23811 37692
rect 23753 37683 23811 37689
rect 25314 37680 25320 37692
rect 25372 37720 25378 37732
rect 25777 37723 25835 37729
rect 25777 37720 25789 37723
rect 25372 37692 25789 37720
rect 25372 37680 25378 37692
rect 25777 37689 25789 37692
rect 25823 37689 25835 37723
rect 25777 37683 25835 37689
rect 3476 37624 4476 37652
rect 6457 37655 6515 37661
rect 3476 37612 3482 37624
rect 6457 37621 6469 37655
rect 6503 37652 6515 37655
rect 6822 37652 6828 37664
rect 6503 37624 6828 37652
rect 6503 37621 6515 37624
rect 6457 37615 6515 37621
rect 6822 37612 6828 37624
rect 6880 37612 6886 37664
rect 11514 37652 11520 37664
rect 11427 37624 11520 37652
rect 11514 37612 11520 37624
rect 11572 37652 11578 37664
rect 11974 37652 11980 37664
rect 11572 37624 11980 37652
rect 11572 37612 11578 37624
rect 11974 37612 11980 37624
rect 12032 37612 12038 37664
rect 12342 37612 12348 37664
rect 12400 37652 12434 37664
rect 13357 37655 13415 37661
rect 13357 37652 13369 37655
rect 12400 37624 13369 37652
rect 12400 37612 12406 37624
rect 13357 37621 13369 37624
rect 13403 37621 13415 37655
rect 13357 37615 13415 37621
rect 13446 37612 13452 37664
rect 13504 37652 13510 37664
rect 13814 37652 13820 37664
rect 13504 37624 13820 37652
rect 13504 37612 13510 37624
rect 13814 37612 13820 37624
rect 13872 37612 13878 37664
rect 14921 37655 14979 37661
rect 14921 37621 14933 37655
rect 14967 37652 14979 37655
rect 15470 37652 15476 37664
rect 14967 37624 15476 37652
rect 14967 37621 14979 37624
rect 14921 37615 14979 37621
rect 15470 37612 15476 37624
rect 15528 37612 15534 37664
rect 15562 37612 15568 37664
rect 15620 37652 15626 37664
rect 15930 37652 15936 37664
rect 15620 37624 15936 37652
rect 15620 37612 15626 37624
rect 15930 37612 15936 37624
rect 15988 37612 15994 37664
rect 20257 37655 20315 37661
rect 20257 37621 20269 37655
rect 20303 37652 20315 37655
rect 20346 37652 20352 37664
rect 20303 37624 20352 37652
rect 20303 37621 20315 37624
rect 20257 37615 20315 37621
rect 20346 37612 20352 37624
rect 20404 37612 20410 37664
rect 25406 37652 25412 37664
rect 25367 37624 25412 37652
rect 25406 37612 25412 37624
rect 25464 37612 25470 37664
rect 27338 37612 27344 37664
rect 27396 37652 27402 37664
rect 27985 37655 28043 37661
rect 27985 37652 27997 37655
rect 27396 37624 27997 37652
rect 27396 37612 27402 37624
rect 27985 37621 27997 37624
rect 28031 37621 28043 37655
rect 27985 37615 28043 37621
rect 1104 37562 28888 37584
rect 1104 37510 10246 37562
rect 10298 37510 10310 37562
rect 10362 37510 10374 37562
rect 10426 37510 10438 37562
rect 10490 37510 19510 37562
rect 19562 37510 19574 37562
rect 19626 37510 19638 37562
rect 19690 37510 19702 37562
rect 19754 37510 28888 37562
rect 1104 37488 28888 37510
rect 2406 37408 2412 37460
rect 2464 37448 2470 37460
rect 13446 37448 13452 37460
rect 2464 37420 13452 37448
rect 2464 37408 2470 37420
rect 13446 37408 13452 37420
rect 13504 37408 13510 37460
rect 13814 37408 13820 37460
rect 13872 37448 13878 37460
rect 27338 37448 27344 37460
rect 13872 37420 27344 37448
rect 13872 37408 13878 37420
rect 27338 37408 27344 37420
rect 27396 37408 27402 37460
rect 28074 37448 28080 37460
rect 28035 37420 28080 37448
rect 28074 37408 28080 37420
rect 28132 37408 28138 37460
rect 2041 37383 2099 37389
rect 2041 37349 2053 37383
rect 2087 37380 2099 37383
rect 2866 37380 2872 37392
rect 2087 37352 2872 37380
rect 2087 37349 2099 37352
rect 2041 37343 2099 37349
rect 2866 37340 2872 37352
rect 2924 37340 2930 37392
rect 4709 37383 4767 37389
rect 4709 37349 4721 37383
rect 4755 37380 4767 37383
rect 5350 37380 5356 37392
rect 4755 37352 5120 37380
rect 5311 37352 5356 37380
rect 4755 37349 4767 37352
rect 4709 37343 4767 37349
rect 1857 37315 1915 37321
rect 1857 37281 1869 37315
rect 1903 37312 1915 37315
rect 2406 37312 2412 37324
rect 1903 37284 2412 37312
rect 1903 37281 1915 37284
rect 1857 37275 1915 37281
rect 2406 37272 2412 37284
rect 2464 37272 2470 37324
rect 2590 37312 2596 37324
rect 2551 37284 2596 37312
rect 2590 37272 2596 37284
rect 2648 37272 2654 37324
rect 3510 37312 3516 37324
rect 3471 37284 3516 37312
rect 3510 37272 3516 37284
rect 3568 37272 3574 37324
rect 4522 37272 4528 37324
rect 4580 37312 4586 37324
rect 4617 37315 4675 37321
rect 4617 37312 4629 37315
rect 4580 37284 4629 37312
rect 4580 37272 4586 37284
rect 4617 37281 4629 37284
rect 4663 37281 4675 37315
rect 4798 37312 4804 37324
rect 4759 37284 4804 37312
rect 4617 37275 4675 37281
rect 3602 37244 3608 37256
rect 3563 37216 3608 37244
rect 3602 37204 3608 37216
rect 3660 37204 3666 37256
rect 4632 37244 4660 37275
rect 4798 37272 4804 37284
rect 4856 37272 4862 37324
rect 4890 37244 4896 37256
rect 4632 37216 4896 37244
rect 4890 37204 4896 37216
rect 4948 37204 4954 37256
rect 5092 37244 5120 37352
rect 5350 37340 5356 37352
rect 5408 37340 5414 37392
rect 8754 37340 8760 37392
rect 8812 37380 8818 37392
rect 9217 37383 9275 37389
rect 9217 37380 9229 37383
rect 8812 37352 9229 37380
rect 8812 37340 8818 37352
rect 9217 37349 9229 37352
rect 9263 37349 9275 37383
rect 9953 37383 10011 37389
rect 9953 37380 9965 37383
rect 9217 37343 9275 37349
rect 9416 37352 9965 37380
rect 5258 37312 5264 37324
rect 5219 37284 5264 37312
rect 5258 37272 5264 37284
rect 5316 37272 5322 37324
rect 5445 37315 5503 37321
rect 5445 37312 5457 37315
rect 5368 37284 5457 37312
rect 5368 37244 5396 37284
rect 5445 37281 5457 37284
rect 5491 37281 5503 37315
rect 8846 37312 8852 37324
rect 5445 37275 5503 37281
rect 5552 37284 8852 37312
rect 5552 37244 5580 37284
rect 5092 37216 5396 37244
rect 5460 37216 5580 37244
rect 2774 37136 2780 37188
rect 2832 37176 2838 37188
rect 3881 37179 3939 37185
rect 2832 37148 2877 37176
rect 2832 37136 2838 37148
rect 3881 37145 3893 37179
rect 3927 37176 3939 37179
rect 3970 37176 3976 37188
rect 3927 37148 3976 37176
rect 3927 37145 3939 37148
rect 3881 37139 3939 37145
rect 3970 37136 3976 37148
rect 4028 37136 4034 37188
rect 4430 37136 4436 37188
rect 4488 37176 4494 37188
rect 5460 37176 5488 37216
rect 8772 37185 8800 37284
rect 8846 37272 8852 37284
rect 8904 37272 8910 37324
rect 9033 37315 9091 37321
rect 9033 37281 9045 37315
rect 9079 37312 9091 37315
rect 9416 37312 9444 37352
rect 9953 37349 9965 37352
rect 9999 37349 10011 37383
rect 10870 37380 10876 37392
rect 9953 37343 10011 37349
rect 10060 37352 10876 37380
rect 9858 37312 9864 37324
rect 9079 37284 9444 37312
rect 9819 37284 9864 37312
rect 9079 37281 9091 37284
rect 9033 37275 9091 37281
rect 9858 37272 9864 37284
rect 9916 37272 9922 37324
rect 10060 37321 10088 37352
rect 10870 37340 10876 37352
rect 10928 37340 10934 37392
rect 12066 37380 12072 37392
rect 12027 37352 12072 37380
rect 12066 37340 12072 37352
rect 12124 37340 12130 37392
rect 12158 37340 12164 37392
rect 12216 37380 12222 37392
rect 13173 37383 13231 37389
rect 12216 37352 12848 37380
rect 12216 37340 12222 37352
rect 10045 37315 10103 37321
rect 10045 37281 10057 37315
rect 10091 37281 10103 37315
rect 11514 37312 11520 37324
rect 10045 37275 10103 37281
rect 10152 37284 11520 37312
rect 9309 37247 9367 37253
rect 9309 37213 9321 37247
rect 9355 37244 9367 37247
rect 10152 37244 10180 37284
rect 11514 37272 11520 37284
rect 11572 37272 11578 37324
rect 12250 37272 12256 37324
rect 12308 37321 12314 37324
rect 12406 37321 12434 37352
rect 12308 37315 12357 37321
rect 12308 37281 12311 37315
rect 12345 37281 12357 37315
rect 12406 37315 12476 37321
rect 12406 37284 12430 37315
rect 12308 37275 12357 37281
rect 12418 37281 12430 37284
rect 12464 37281 12476 37315
rect 12418 37275 12476 37281
rect 12518 37315 12576 37321
rect 12518 37281 12530 37315
rect 12564 37281 12576 37315
rect 12710 37312 12716 37324
rect 12671 37284 12716 37312
rect 12518 37275 12576 37281
rect 12308 37272 12314 37275
rect 9355 37216 10180 37244
rect 9355 37213 9367 37216
rect 9309 37207 9367 37213
rect 12158 37204 12164 37256
rect 12216 37244 12222 37256
rect 12544 37244 12572 37275
rect 12710 37272 12716 37284
rect 12768 37272 12774 37324
rect 12216 37216 12572 37244
rect 12820 37244 12848 37352
rect 13173 37349 13185 37383
rect 13219 37380 13231 37383
rect 13262 37380 13268 37392
rect 13219 37352 13268 37380
rect 13219 37349 13231 37352
rect 13173 37343 13231 37349
rect 13262 37340 13268 37352
rect 13320 37340 13326 37392
rect 13722 37340 13728 37392
rect 13780 37340 13786 37392
rect 13998 37340 14004 37392
rect 14056 37380 14062 37392
rect 14553 37383 14611 37389
rect 14553 37380 14565 37383
rect 14056 37352 14565 37380
rect 14056 37340 14062 37352
rect 13446 37312 13452 37324
rect 13407 37284 13452 37312
rect 13446 37272 13452 37284
rect 13504 37272 13510 37324
rect 13538 37315 13596 37321
rect 13538 37281 13550 37315
rect 13584 37281 13596 37315
rect 13538 37275 13596 37281
rect 13633 37315 13691 37321
rect 13633 37281 13645 37315
rect 13679 37312 13691 37315
rect 13740 37312 13768 37340
rect 13679 37284 13768 37312
rect 13817 37315 13875 37321
rect 13817 37286 13829 37315
rect 13863 37286 13875 37315
rect 13679 37281 13691 37284
rect 13633 37275 13691 37281
rect 13556 37244 13584 37275
rect 12820 37216 13584 37244
rect 13814 37234 13820 37286
rect 13872 37234 13878 37286
rect 14292 37244 14320 37352
rect 14553 37349 14565 37352
rect 14599 37349 14611 37383
rect 14553 37343 14611 37349
rect 14645 37383 14703 37389
rect 14645 37349 14657 37383
rect 14691 37380 14703 37383
rect 14826 37380 14832 37392
rect 14691 37352 14832 37380
rect 14691 37349 14703 37352
rect 14645 37343 14703 37349
rect 14826 37340 14832 37352
rect 14884 37380 14890 37392
rect 15562 37380 15568 37392
rect 14884 37352 15568 37380
rect 14884 37340 14890 37352
rect 15562 37340 15568 37352
rect 15620 37340 15626 37392
rect 15654 37340 15660 37392
rect 15712 37380 15718 37392
rect 15933 37383 15991 37389
rect 15933 37380 15945 37383
rect 15712 37352 15945 37380
rect 15712 37340 15718 37352
rect 15933 37349 15945 37352
rect 15979 37380 15991 37383
rect 20346 37380 20352 37392
rect 15979 37352 19334 37380
rect 20307 37352 20352 37380
rect 15979 37349 15991 37352
rect 15933 37343 15991 37349
rect 14369 37315 14427 37321
rect 14369 37281 14381 37315
rect 14415 37312 14427 37315
rect 14734 37312 14740 37324
rect 14415 37284 14596 37312
rect 14695 37284 14740 37312
rect 14415 37281 14427 37284
rect 14369 37275 14427 37281
rect 14568 37244 14596 37284
rect 14734 37272 14740 37284
rect 14792 37272 14798 37324
rect 15286 37312 15292 37324
rect 14844 37284 15292 37312
rect 14844 37244 14872 37284
rect 15286 37272 15292 37284
rect 15344 37312 15350 37324
rect 15749 37315 15807 37321
rect 15749 37312 15761 37315
rect 15344 37284 15761 37312
rect 15344 37272 15350 37284
rect 15749 37281 15761 37284
rect 15795 37281 15807 37315
rect 15749 37275 15807 37281
rect 17954 37272 17960 37324
rect 18012 37312 18018 37324
rect 18305 37315 18363 37321
rect 18305 37312 18317 37315
rect 18012 37284 18317 37312
rect 18012 37272 18018 37284
rect 18305 37281 18317 37284
rect 18351 37281 18363 37315
rect 19306 37312 19334 37352
rect 20346 37340 20352 37352
rect 20404 37340 20410 37392
rect 20438 37340 20444 37392
rect 20496 37380 20502 37392
rect 20496 37352 20541 37380
rect 20496 37340 20502 37352
rect 20898 37340 20904 37392
rect 20956 37380 20962 37392
rect 21266 37380 21272 37392
rect 20956 37352 21272 37380
rect 20956 37340 20962 37352
rect 21266 37340 21272 37352
rect 21324 37340 21330 37392
rect 21358 37340 21364 37392
rect 21416 37380 21422 37392
rect 25038 37380 25044 37392
rect 21416 37352 24900 37380
rect 24999 37352 25044 37380
rect 21416 37340 21422 37352
rect 21082 37312 21088 37324
rect 19306 37284 21088 37312
rect 18305 37275 18363 37281
rect 21082 37272 21088 37284
rect 21140 37272 21146 37324
rect 22738 37272 22744 37324
rect 22796 37312 22802 37324
rect 24872 37321 24900 37352
rect 25038 37340 25044 37352
rect 25096 37340 25102 37392
rect 26694 37340 26700 37392
rect 26752 37380 26758 37392
rect 27985 37383 28043 37389
rect 27985 37380 27997 37383
rect 26752 37352 27997 37380
rect 26752 37340 26758 37352
rect 27985 37349 27997 37352
rect 28031 37349 28043 37383
rect 27985 37343 28043 37349
rect 23089 37315 23147 37321
rect 23089 37312 23101 37315
rect 22796 37284 23101 37312
rect 22796 37272 22802 37284
rect 23089 37281 23101 37284
rect 23135 37281 23147 37315
rect 23089 37275 23147 37281
rect 24673 37315 24731 37321
rect 24673 37281 24685 37315
rect 24719 37312 24731 37315
rect 24857 37315 24915 37321
rect 24719 37284 24808 37312
rect 24719 37281 24731 37284
rect 24673 37275 24731 37281
rect 14292 37216 14412 37244
rect 14568 37216 14872 37244
rect 12216 37204 12222 37216
rect 14384 37188 14412 37216
rect 15654 37204 15660 37256
rect 15712 37244 15718 37256
rect 17218 37244 17224 37256
rect 15712 37216 17224 37244
rect 15712 37204 15718 37216
rect 17218 37204 17224 37216
rect 17276 37244 17282 37256
rect 18046 37244 18052 37256
rect 17276 37216 18052 37244
rect 17276 37204 17282 37216
rect 18046 37204 18052 37216
rect 18104 37204 18110 37256
rect 20346 37204 20352 37256
rect 20404 37244 20410 37256
rect 20533 37247 20591 37253
rect 20533 37244 20545 37247
rect 20404 37216 20545 37244
rect 20404 37204 20410 37216
rect 20533 37213 20545 37216
rect 20579 37213 20591 37247
rect 20533 37207 20591 37213
rect 22833 37247 22891 37253
rect 22833 37213 22845 37247
rect 22879 37213 22891 37247
rect 24780 37244 24808 37284
rect 24857 37281 24869 37315
rect 24903 37281 24915 37315
rect 25314 37312 25320 37324
rect 24857 37275 24915 37281
rect 24964 37284 25320 37312
rect 24964 37244 24992 37284
rect 25314 37272 25320 37284
rect 25372 37272 25378 37324
rect 25406 37272 25412 37324
rect 25464 37312 25470 37324
rect 25869 37315 25927 37321
rect 25869 37312 25881 37315
rect 25464 37284 25881 37312
rect 25464 37272 25470 37284
rect 25869 37281 25881 37284
rect 25915 37281 25927 37315
rect 25869 37275 25927 37281
rect 26053 37315 26111 37321
rect 26053 37281 26065 37315
rect 26099 37281 26111 37315
rect 26053 37275 26111 37281
rect 26513 37315 26571 37321
rect 26513 37281 26525 37315
rect 26559 37312 26571 37315
rect 26970 37312 26976 37324
rect 26559 37284 26976 37312
rect 26559 37281 26571 37284
rect 26513 37275 26571 37281
rect 25774 37244 25780 37256
rect 24780 37216 24992 37244
rect 25735 37216 25780 37244
rect 22833 37207 22891 37213
rect 4488 37148 5488 37176
rect 8757 37179 8815 37185
rect 4488 37136 4494 37148
rect 8757 37145 8769 37179
rect 8803 37145 8815 37179
rect 8757 37139 8815 37145
rect 11146 37136 11152 37188
rect 11204 37176 11210 37188
rect 11514 37176 11520 37188
rect 11204 37148 11520 37176
rect 11204 37136 11210 37148
rect 11514 37136 11520 37148
rect 11572 37136 11578 37188
rect 14366 37136 14372 37188
rect 14424 37136 14430 37188
rect 15194 37176 15200 37188
rect 14660 37148 15200 37176
rect 7282 37068 7288 37120
rect 7340 37108 7346 37120
rect 14660 37108 14688 37148
rect 15194 37136 15200 37148
rect 15252 37176 15258 37188
rect 17862 37176 17868 37188
rect 15252 37148 17868 37176
rect 15252 37136 15258 37148
rect 17862 37136 17868 37148
rect 17920 37136 17926 37188
rect 7340 37080 14688 37108
rect 7340 37068 7346 37080
rect 14734 37068 14740 37120
rect 14792 37108 14798 37120
rect 14921 37111 14979 37117
rect 14921 37108 14933 37111
rect 14792 37080 14933 37108
rect 14792 37068 14798 37080
rect 14921 37077 14933 37080
rect 14967 37077 14979 37111
rect 14921 37071 14979 37077
rect 19334 37068 19340 37120
rect 19392 37108 19398 37120
rect 19429 37111 19487 37117
rect 19429 37108 19441 37111
rect 19392 37080 19441 37108
rect 19392 37068 19398 37080
rect 19429 37077 19441 37080
rect 19475 37077 19487 37111
rect 19429 37071 19487 37077
rect 19981 37111 20039 37117
rect 19981 37077 19993 37111
rect 20027 37108 20039 37111
rect 20898 37108 20904 37120
rect 20027 37080 20904 37108
rect 20027 37077 20039 37080
rect 19981 37071 20039 37077
rect 20898 37068 20904 37080
rect 20956 37068 20962 37120
rect 20990 37068 20996 37120
rect 21048 37108 21054 37120
rect 21361 37111 21419 37117
rect 21361 37108 21373 37111
rect 21048 37080 21373 37108
rect 21048 37068 21054 37080
rect 21361 37077 21373 37080
rect 21407 37077 21419 37111
rect 22848 37108 22876 37207
rect 25774 37204 25780 37216
rect 25832 37204 25838 37256
rect 26068 37244 26096 37275
rect 26970 37272 26976 37284
rect 27028 37272 27034 37324
rect 26602 37244 26608 37256
rect 26068 37216 26608 37244
rect 26602 37204 26608 37216
rect 26660 37204 26666 37256
rect 23014 37108 23020 37120
rect 22848 37080 23020 37108
rect 21361 37071 21419 37077
rect 23014 37068 23020 37080
rect 23072 37108 23078 37120
rect 23198 37108 23204 37120
rect 23072 37080 23204 37108
rect 23072 37068 23078 37080
rect 23198 37068 23204 37080
rect 23256 37068 23262 37120
rect 24026 37068 24032 37120
rect 24084 37108 24090 37120
rect 24213 37111 24271 37117
rect 24213 37108 24225 37111
rect 24084 37080 24225 37108
rect 24084 37068 24090 37080
rect 24213 37077 24225 37080
rect 24259 37077 24271 37111
rect 24213 37071 24271 37077
rect 1104 37018 28888 37040
rect 1104 36966 5614 37018
rect 5666 36966 5678 37018
rect 5730 36966 5742 37018
rect 5794 36966 5806 37018
rect 5858 36966 14878 37018
rect 14930 36966 14942 37018
rect 14994 36966 15006 37018
rect 15058 36966 15070 37018
rect 15122 36966 24142 37018
rect 24194 36966 24206 37018
rect 24258 36966 24270 37018
rect 24322 36966 24334 37018
rect 24386 36966 28888 37018
rect 1104 36944 28888 36966
rect 2746 36876 22094 36904
rect 2590 36796 2596 36848
rect 2648 36836 2654 36848
rect 2746 36836 2774 36876
rect 2648 36808 2774 36836
rect 2648 36796 2654 36808
rect 3602 36796 3608 36848
rect 3660 36836 3666 36848
rect 4341 36839 4399 36845
rect 4341 36836 4353 36839
rect 3660 36808 4353 36836
rect 3660 36796 3666 36808
rect 4341 36805 4353 36808
rect 4387 36805 4399 36839
rect 4341 36799 4399 36805
rect 7193 36839 7251 36845
rect 7193 36805 7205 36839
rect 7239 36836 7251 36839
rect 9030 36836 9036 36848
rect 7239 36808 9036 36836
rect 7239 36805 7251 36808
rect 7193 36799 7251 36805
rect 9030 36796 9036 36808
rect 9088 36796 9094 36848
rect 10962 36796 10968 36848
rect 11020 36836 11026 36848
rect 11701 36839 11759 36845
rect 11701 36836 11713 36839
rect 11020 36808 11713 36836
rect 11020 36796 11026 36808
rect 11701 36805 11713 36808
rect 11747 36805 11759 36839
rect 11701 36799 11759 36805
rect 13722 36796 13728 36848
rect 13780 36836 13786 36848
rect 15197 36839 15255 36845
rect 15197 36836 15209 36839
rect 13780 36808 15209 36836
rect 13780 36796 13786 36808
rect 15197 36805 15209 36808
rect 15243 36805 15255 36839
rect 15197 36799 15255 36805
rect 16758 36796 16764 36848
rect 16816 36836 16822 36848
rect 17494 36836 17500 36848
rect 16816 36808 17500 36836
rect 16816 36796 16822 36808
rect 17494 36796 17500 36808
rect 17552 36836 17558 36848
rect 18049 36839 18107 36845
rect 18049 36836 18061 36839
rect 17552 36808 18061 36836
rect 17552 36796 17558 36808
rect 18049 36805 18061 36808
rect 18095 36805 18107 36839
rect 22066 36836 22094 36876
rect 25774 36864 25780 36916
rect 25832 36904 25838 36916
rect 25961 36907 26019 36913
rect 25961 36904 25973 36907
rect 25832 36876 25973 36904
rect 25832 36864 25838 36876
rect 25961 36873 25973 36876
rect 26007 36873 26019 36907
rect 28077 36907 28135 36913
rect 28077 36904 28089 36907
rect 25961 36867 26019 36873
rect 26068 36876 28089 36904
rect 26068 36836 26096 36876
rect 28077 36873 28089 36876
rect 28123 36873 28135 36907
rect 28077 36867 28135 36873
rect 22066 36808 26096 36836
rect 26605 36839 26663 36845
rect 18049 36799 18107 36805
rect 26605 36805 26617 36839
rect 26651 36836 26663 36839
rect 27890 36836 27896 36848
rect 26651 36808 27896 36836
rect 26651 36805 26663 36808
rect 26605 36799 26663 36805
rect 27890 36796 27896 36808
rect 27948 36796 27954 36848
rect 2682 36728 2688 36780
rect 2740 36768 2746 36780
rect 12434 36768 12440 36780
rect 2740 36740 5212 36768
rect 2740 36728 2746 36740
rect 4154 36660 4160 36712
rect 4212 36700 4218 36712
rect 4249 36703 4307 36709
rect 4249 36700 4261 36703
rect 4212 36672 4261 36700
rect 4212 36660 4218 36672
rect 4249 36669 4261 36672
rect 4295 36669 4307 36703
rect 4249 36663 4307 36669
rect 4433 36703 4491 36709
rect 4433 36669 4445 36703
rect 4479 36700 4491 36703
rect 4614 36700 4620 36712
rect 4479 36672 4620 36700
rect 4479 36669 4491 36672
rect 4433 36663 4491 36669
rect 4614 36660 4620 36672
rect 4672 36660 4678 36712
rect 5184 36709 5212 36740
rect 12084 36740 12440 36768
rect 5169 36703 5227 36709
rect 5169 36669 5181 36703
rect 5215 36669 5227 36703
rect 5169 36663 5227 36669
rect 5813 36703 5871 36709
rect 5813 36669 5825 36703
rect 5859 36700 5871 36703
rect 5902 36700 5908 36712
rect 5859 36672 5908 36700
rect 5859 36669 5871 36672
rect 5813 36663 5871 36669
rect 1854 36632 1860 36644
rect 1815 36604 1860 36632
rect 1854 36592 1860 36604
rect 1912 36592 1918 36644
rect 2590 36632 2596 36644
rect 2551 36604 2596 36632
rect 2590 36592 2596 36604
rect 2648 36592 2654 36644
rect 2774 36592 2780 36644
rect 2832 36632 2838 36644
rect 2832 36604 2877 36632
rect 2832 36592 2838 36604
rect 4706 36592 4712 36644
rect 4764 36632 4770 36644
rect 4985 36635 5043 36641
rect 4985 36632 4997 36635
rect 4764 36604 4997 36632
rect 4764 36592 4770 36604
rect 4985 36601 4997 36604
rect 5031 36601 5043 36635
rect 4985 36595 5043 36601
rect 1946 36564 1952 36576
rect 1907 36536 1952 36564
rect 1946 36524 1952 36536
rect 2004 36524 2010 36576
rect 5184 36564 5212 36663
rect 5902 36660 5908 36672
rect 5960 36700 5966 36712
rect 6362 36700 6368 36712
rect 5960 36672 6368 36700
rect 5960 36660 5966 36672
rect 6362 36660 6368 36672
rect 6420 36660 6426 36712
rect 9674 36700 9680 36712
rect 9635 36672 9680 36700
rect 9674 36660 9680 36672
rect 9732 36660 9738 36712
rect 11974 36700 11980 36712
rect 11935 36672 11980 36700
rect 11974 36660 11980 36672
rect 12032 36660 12038 36712
rect 12084 36709 12112 36740
rect 12434 36728 12440 36740
rect 12492 36768 12498 36780
rect 13817 36771 13875 36777
rect 13817 36768 13829 36771
rect 12492 36740 13829 36768
rect 12492 36728 12498 36740
rect 13817 36737 13829 36740
rect 13863 36737 13875 36771
rect 13817 36731 13875 36737
rect 15470 36728 15476 36780
rect 15528 36768 15534 36780
rect 16022 36768 16028 36780
rect 15528 36740 16028 36768
rect 15528 36728 15534 36740
rect 16022 36728 16028 36740
rect 16080 36768 16086 36780
rect 17037 36771 17095 36777
rect 17037 36768 17049 36771
rect 16080 36740 17049 36768
rect 16080 36728 16086 36740
rect 17037 36737 17049 36740
rect 17083 36737 17095 36771
rect 17037 36731 17095 36737
rect 17218 36728 17224 36780
rect 17276 36768 17282 36780
rect 18966 36768 18972 36780
rect 17276 36740 18972 36768
rect 17276 36728 17282 36740
rect 18966 36728 18972 36740
rect 19024 36728 19030 36780
rect 25498 36728 25504 36780
rect 25556 36768 25562 36780
rect 25556 36740 26096 36768
rect 25556 36728 25562 36740
rect 12069 36703 12127 36709
rect 12069 36669 12081 36703
rect 12115 36669 12127 36703
rect 12069 36663 12127 36669
rect 12158 36660 12164 36712
rect 12216 36700 12222 36712
rect 12345 36703 12403 36709
rect 12216 36672 12261 36700
rect 12216 36660 12222 36672
rect 12345 36669 12357 36703
rect 12391 36700 12403 36703
rect 13262 36700 13268 36712
rect 12391 36672 13268 36700
rect 12391 36669 12403 36672
rect 12345 36663 12403 36669
rect 13262 36660 13268 36672
rect 13320 36660 13326 36712
rect 13633 36703 13691 36709
rect 13633 36669 13645 36703
rect 13679 36700 13691 36703
rect 13679 36672 15608 36700
rect 13679 36669 13691 36672
rect 13633 36663 13691 36669
rect 5353 36635 5411 36641
rect 5353 36601 5365 36635
rect 5399 36632 5411 36635
rect 6058 36635 6116 36641
rect 6058 36632 6070 36635
rect 5399 36604 6070 36632
rect 5399 36601 5411 36604
rect 5353 36595 5411 36601
rect 6058 36601 6070 36604
rect 6104 36601 6116 36635
rect 6058 36595 6116 36601
rect 14090 36592 14096 36644
rect 14148 36632 14154 36644
rect 14366 36632 14372 36644
rect 14148 36604 14372 36632
rect 14148 36592 14154 36604
rect 14366 36592 14372 36604
rect 14424 36592 14430 36644
rect 15013 36635 15071 36641
rect 15013 36601 15025 36635
rect 15059 36632 15071 36635
rect 15194 36632 15200 36644
rect 15059 36604 15200 36632
rect 15059 36601 15071 36604
rect 15013 36595 15071 36601
rect 15194 36592 15200 36604
rect 15252 36592 15258 36644
rect 7282 36564 7288 36576
rect 5184 36536 7288 36564
rect 7282 36524 7288 36536
rect 7340 36524 7346 36576
rect 9490 36564 9496 36576
rect 9451 36536 9496 36564
rect 9490 36524 9496 36536
rect 9548 36524 9554 36576
rect 10870 36524 10876 36576
rect 10928 36564 10934 36576
rect 13354 36564 13360 36576
rect 10928 36536 13360 36564
rect 10928 36524 10934 36536
rect 13354 36524 13360 36536
rect 13412 36524 13418 36576
rect 15580 36564 15608 36672
rect 15654 36660 15660 36712
rect 15712 36700 15718 36712
rect 15930 36700 15936 36712
rect 15712 36672 15757 36700
rect 15891 36672 15936 36700
rect 15712 36660 15718 36672
rect 15930 36660 15936 36672
rect 15988 36660 15994 36712
rect 16206 36660 16212 36712
rect 16264 36700 16270 36712
rect 16390 36700 16396 36712
rect 16264 36672 16396 36700
rect 16264 36660 16270 36672
rect 16390 36660 16396 36672
rect 16448 36660 16454 36712
rect 18693 36703 18751 36709
rect 18693 36669 18705 36703
rect 18739 36700 18751 36703
rect 20714 36700 20720 36712
rect 18739 36672 20576 36700
rect 20675 36672 20720 36700
rect 18739 36669 18751 36672
rect 18693 36663 18751 36669
rect 17865 36635 17923 36641
rect 17865 36601 17877 36635
rect 17911 36632 17923 36635
rect 17911 36604 18736 36632
rect 17911 36601 17923 36604
rect 17865 36595 17923 36601
rect 16574 36564 16580 36576
rect 15580 36536 16580 36564
rect 16574 36524 16580 36536
rect 16632 36564 16638 36576
rect 17880 36564 17908 36595
rect 18708 36576 18736 36604
rect 20548 36576 20576 36672
rect 20714 36660 20720 36672
rect 20772 36660 20778 36712
rect 21266 36660 21272 36712
rect 21324 36700 21330 36712
rect 21453 36703 21511 36709
rect 21453 36700 21465 36703
rect 21324 36672 21465 36700
rect 21324 36660 21330 36672
rect 21453 36669 21465 36672
rect 21499 36669 21511 36703
rect 25406 36700 25412 36712
rect 25367 36672 25412 36700
rect 21453 36663 21511 36669
rect 25406 36660 25412 36672
rect 25464 36660 25470 36712
rect 25774 36660 25780 36712
rect 25832 36700 25838 36712
rect 26068 36709 26096 36740
rect 25869 36703 25927 36709
rect 25869 36700 25881 36703
rect 25832 36672 25881 36700
rect 25832 36660 25838 36672
rect 25869 36669 25881 36672
rect 25915 36669 25927 36703
rect 25869 36663 25927 36669
rect 26053 36703 26111 36709
rect 26053 36669 26065 36703
rect 26099 36669 26111 36703
rect 26786 36700 26792 36712
rect 26747 36672 26792 36700
rect 26053 36663 26111 36669
rect 26786 36660 26792 36672
rect 26844 36660 26850 36712
rect 27430 36700 27436 36712
rect 27391 36672 27436 36700
rect 27430 36660 27436 36672
rect 27488 36660 27494 36712
rect 25498 36592 25504 36644
rect 25556 36632 25562 36644
rect 27985 36635 28043 36641
rect 27985 36632 27997 36635
rect 25556 36604 27997 36632
rect 25556 36592 25562 36604
rect 27985 36601 27997 36604
rect 28031 36601 28043 36635
rect 27985 36595 28043 36601
rect 16632 36536 17908 36564
rect 16632 36524 16638 36536
rect 18046 36524 18052 36576
rect 18104 36564 18110 36576
rect 18509 36567 18567 36573
rect 18509 36564 18521 36567
rect 18104 36536 18521 36564
rect 18104 36524 18110 36536
rect 18509 36533 18521 36536
rect 18555 36564 18567 36567
rect 18598 36564 18604 36576
rect 18555 36536 18604 36564
rect 18555 36533 18567 36536
rect 18509 36527 18567 36533
rect 18598 36524 18604 36536
rect 18656 36524 18662 36576
rect 18690 36524 18696 36576
rect 18748 36524 18754 36576
rect 20530 36564 20536 36576
rect 20491 36536 20536 36564
rect 20530 36524 20536 36536
rect 20588 36524 20594 36576
rect 21545 36567 21603 36573
rect 21545 36533 21557 36567
rect 21591 36564 21603 36567
rect 21910 36564 21916 36576
rect 21591 36536 21916 36564
rect 21591 36533 21603 36536
rect 21545 36527 21603 36533
rect 21910 36524 21916 36536
rect 21968 36524 21974 36576
rect 25222 36564 25228 36576
rect 25183 36536 25228 36564
rect 25222 36524 25228 36536
rect 25280 36524 25286 36576
rect 25774 36524 25780 36576
rect 25832 36564 25838 36576
rect 26050 36564 26056 36576
rect 25832 36536 26056 36564
rect 25832 36524 25838 36536
rect 26050 36524 26056 36536
rect 26108 36524 26114 36576
rect 27249 36567 27307 36573
rect 27249 36533 27261 36567
rect 27295 36564 27307 36567
rect 27798 36564 27804 36576
rect 27295 36536 27804 36564
rect 27295 36533 27307 36536
rect 27249 36527 27307 36533
rect 27798 36524 27804 36536
rect 27856 36524 27862 36576
rect 1104 36474 28888 36496
rect 1104 36422 10246 36474
rect 10298 36422 10310 36474
rect 10362 36422 10374 36474
rect 10426 36422 10438 36474
rect 10490 36422 19510 36474
rect 19562 36422 19574 36474
rect 19626 36422 19638 36474
rect 19690 36422 19702 36474
rect 19754 36422 28888 36474
rect 1104 36400 28888 36422
rect 3053 36363 3111 36369
rect 3053 36329 3065 36363
rect 3099 36360 3111 36363
rect 4246 36360 4252 36372
rect 3099 36332 4252 36360
rect 3099 36329 3111 36332
rect 3053 36323 3111 36329
rect 4246 36320 4252 36332
rect 4304 36320 4310 36372
rect 4893 36363 4951 36369
rect 4893 36329 4905 36363
rect 4939 36360 4951 36363
rect 5258 36360 5264 36372
rect 4939 36332 5264 36360
rect 4939 36329 4951 36332
rect 4893 36323 4951 36329
rect 5258 36320 5264 36332
rect 5316 36320 5322 36372
rect 5537 36363 5595 36369
rect 5537 36329 5549 36363
rect 5583 36360 5595 36363
rect 6086 36360 6092 36372
rect 5583 36332 6092 36360
rect 5583 36329 5595 36332
rect 5537 36323 5595 36329
rect 6086 36320 6092 36332
rect 6144 36320 6150 36372
rect 8297 36363 8355 36369
rect 8297 36329 8309 36363
rect 8343 36360 8355 36363
rect 9217 36363 9275 36369
rect 9217 36360 9229 36363
rect 8343 36332 9229 36360
rect 8343 36329 8355 36332
rect 8297 36323 8355 36329
rect 9217 36329 9229 36332
rect 9263 36329 9275 36363
rect 9217 36323 9275 36329
rect 9490 36320 9496 36372
rect 9548 36360 9554 36372
rect 11606 36360 11612 36372
rect 9548 36332 11612 36360
rect 9548 36320 9554 36332
rect 11606 36320 11612 36332
rect 11664 36320 11670 36372
rect 14093 36363 14151 36369
rect 14093 36329 14105 36363
rect 14139 36360 14151 36363
rect 14550 36360 14556 36372
rect 14139 36332 14556 36360
rect 14139 36329 14151 36332
rect 14093 36323 14151 36329
rect 14550 36320 14556 36332
rect 14608 36320 14614 36372
rect 15197 36363 15255 36369
rect 15197 36329 15209 36363
rect 15243 36360 15255 36363
rect 15930 36360 15936 36372
rect 15243 36332 15936 36360
rect 15243 36329 15255 36332
rect 15197 36323 15255 36329
rect 15930 36320 15936 36332
rect 15988 36320 15994 36372
rect 22738 36360 22744 36372
rect 17696 36332 22600 36360
rect 22699 36332 22744 36360
rect 17696 36292 17724 36332
rect 2746 36264 17724 36292
rect 1394 36184 1400 36236
rect 1452 36224 1458 36236
rect 1670 36224 1676 36236
rect 1452 36196 1676 36224
rect 1452 36184 1458 36196
rect 1670 36184 1676 36196
rect 1728 36184 1734 36236
rect 1762 36156 1768 36168
rect 1723 36128 1768 36156
rect 1762 36116 1768 36128
rect 1820 36116 1826 36168
rect 2222 36116 2228 36168
rect 2280 36156 2286 36168
rect 2409 36159 2467 36165
rect 2409 36156 2421 36159
rect 2280 36128 2421 36156
rect 2280 36116 2286 36128
rect 2409 36125 2421 36128
rect 2455 36125 2467 36159
rect 2409 36119 2467 36125
rect 1578 36048 1584 36100
rect 1636 36088 1642 36100
rect 2746 36088 2774 36264
rect 18506 36252 18512 36304
rect 18564 36292 18570 36304
rect 18874 36292 18880 36304
rect 18564 36264 18880 36292
rect 18564 36252 18570 36264
rect 18874 36252 18880 36264
rect 18932 36252 18938 36304
rect 2961 36227 3019 36233
rect 2961 36193 2973 36227
rect 3007 36224 3019 36227
rect 3050 36224 3056 36236
rect 3007 36196 3056 36224
rect 3007 36193 3019 36196
rect 2961 36187 3019 36193
rect 3050 36184 3056 36196
rect 3108 36184 3114 36236
rect 3142 36184 3148 36236
rect 3200 36224 3206 36236
rect 3789 36227 3847 36233
rect 3200 36196 3245 36224
rect 3200 36184 3206 36196
rect 3789 36193 3801 36227
rect 3835 36224 3847 36227
rect 4430 36224 4436 36236
rect 3835 36196 4436 36224
rect 3835 36193 3847 36196
rect 3789 36187 3847 36193
rect 4430 36184 4436 36196
rect 4488 36184 4494 36236
rect 4617 36227 4675 36233
rect 4617 36193 4629 36227
rect 4663 36224 4675 36227
rect 4709 36227 4767 36233
rect 4709 36224 4721 36227
rect 4663 36196 4721 36224
rect 4663 36193 4675 36196
rect 4617 36187 4675 36193
rect 4709 36193 4721 36196
rect 4755 36193 4767 36227
rect 4709 36187 4767 36193
rect 4901 36227 4959 36233
rect 4901 36193 4913 36227
rect 4947 36193 4959 36227
rect 4901 36187 4959 36193
rect 5445 36227 5503 36233
rect 5445 36193 5457 36227
rect 5491 36224 5503 36227
rect 6822 36224 6828 36236
rect 5491 36196 6828 36224
rect 5491 36193 5503 36196
rect 5445 36187 5503 36193
rect 4338 36116 4344 36168
rect 4396 36156 4402 36168
rect 4908 36156 4936 36187
rect 4396 36128 4936 36156
rect 4396 36116 4402 36128
rect 1636 36060 2774 36088
rect 4617 36091 4675 36097
rect 1636 36048 1642 36060
rect 4617 36057 4629 36091
rect 4663 36088 4675 36091
rect 5460 36088 5488 36187
rect 6822 36184 6828 36196
rect 6880 36184 6886 36236
rect 7190 36233 7196 36236
rect 7184 36187 7196 36233
rect 7248 36224 7254 36236
rect 9122 36224 9128 36236
rect 7248 36196 7284 36224
rect 9083 36196 9128 36224
rect 7190 36184 7196 36187
rect 7248 36184 7254 36196
rect 9122 36184 9128 36196
rect 9180 36184 9186 36236
rect 10410 36184 10416 36236
rect 10468 36224 10474 36236
rect 10735 36227 10793 36233
rect 10735 36224 10747 36227
rect 10468 36196 10747 36224
rect 10468 36184 10474 36196
rect 10735 36193 10747 36196
rect 10781 36193 10793 36227
rect 10870 36224 10876 36236
rect 10831 36196 10876 36224
rect 10735 36187 10793 36193
rect 10870 36184 10876 36196
rect 10928 36184 10934 36236
rect 10965 36227 11023 36233
rect 10965 36193 10977 36227
rect 11011 36193 11023 36227
rect 11146 36224 11152 36236
rect 11107 36196 11152 36224
rect 10965 36187 11023 36193
rect 6362 36116 6368 36168
rect 6420 36156 6426 36168
rect 6917 36159 6975 36165
rect 6917 36156 6929 36159
rect 6420 36128 6929 36156
rect 6420 36116 6426 36128
rect 6917 36125 6929 36128
rect 6963 36125 6975 36159
rect 6917 36119 6975 36125
rect 9401 36159 9459 36165
rect 9401 36125 9413 36159
rect 9447 36156 9459 36159
rect 9858 36156 9864 36168
rect 9447 36128 9864 36156
rect 9447 36125 9459 36128
rect 9401 36119 9459 36125
rect 9858 36116 9864 36128
rect 9916 36116 9922 36168
rect 10980 36156 11008 36187
rect 11146 36184 11152 36196
rect 11204 36184 11210 36236
rect 11606 36184 11612 36236
rect 11664 36224 11670 36236
rect 12253 36227 12311 36233
rect 12253 36224 12265 36227
rect 11664 36196 12265 36224
rect 11664 36184 11670 36196
rect 12253 36193 12265 36196
rect 12299 36193 12311 36227
rect 12253 36187 12311 36193
rect 13909 36227 13967 36233
rect 13909 36193 13921 36227
rect 13955 36224 13967 36227
rect 13998 36224 14004 36236
rect 13955 36196 14004 36224
rect 13955 36193 13967 36196
rect 13909 36187 13967 36193
rect 13998 36184 14004 36196
rect 14056 36184 14062 36236
rect 14093 36227 14151 36233
rect 14093 36193 14105 36227
rect 14139 36193 14151 36227
rect 15470 36224 15476 36236
rect 15431 36196 15476 36224
rect 14093 36187 14151 36193
rect 13722 36156 13728 36168
rect 10980 36128 13728 36156
rect 8754 36088 8760 36100
rect 4663 36060 5488 36088
rect 8715 36060 8760 36088
rect 4663 36057 4675 36060
rect 4617 36051 4675 36057
rect 8754 36048 8760 36060
rect 8812 36048 8818 36100
rect 9876 36088 9904 36116
rect 9876 36060 10824 36088
rect 3878 36020 3884 36032
rect 3839 35992 3884 36020
rect 3878 35980 3884 35992
rect 3936 35980 3942 36032
rect 9674 35980 9680 36032
rect 9732 36020 9738 36032
rect 9950 36020 9956 36032
rect 9732 35992 9956 36020
rect 9732 35980 9738 35992
rect 9950 35980 9956 35992
rect 10008 35980 10014 36032
rect 10502 36020 10508 36032
rect 10463 35992 10508 36020
rect 10502 35980 10508 35992
rect 10560 35980 10566 36032
rect 10796 36020 10824 36060
rect 10870 36048 10876 36100
rect 10928 36088 10934 36100
rect 10980 36088 11008 36128
rect 13722 36116 13728 36128
rect 13780 36116 13786 36168
rect 11974 36088 11980 36100
rect 10928 36060 11008 36088
rect 11440 36060 11980 36088
rect 10928 36048 10934 36060
rect 11440 36020 11468 36060
rect 11974 36048 11980 36060
rect 12032 36048 12038 36100
rect 13630 36048 13636 36100
rect 13688 36088 13694 36100
rect 14108 36088 14136 36187
rect 15470 36184 15476 36196
rect 15528 36184 15534 36236
rect 15565 36227 15623 36233
rect 15565 36193 15577 36227
rect 15611 36193 15623 36227
rect 15565 36187 15623 36193
rect 15657 36227 15715 36233
rect 15657 36193 15669 36227
rect 15703 36193 15715 36227
rect 15838 36224 15844 36236
rect 15799 36196 15844 36224
rect 15657 36187 15715 36193
rect 14550 36116 14556 36168
rect 14608 36156 14614 36168
rect 15102 36156 15108 36168
rect 14608 36128 15108 36156
rect 14608 36116 14614 36128
rect 15102 36116 15108 36128
rect 15160 36116 15166 36168
rect 15580 36088 15608 36187
rect 15672 36156 15700 36187
rect 15838 36184 15844 36196
rect 15896 36184 15902 36236
rect 17218 36184 17224 36236
rect 17276 36224 17282 36236
rect 17635 36227 17693 36233
rect 17635 36224 17647 36227
rect 17276 36196 17647 36224
rect 17276 36184 17282 36196
rect 17635 36193 17647 36196
rect 17681 36193 17693 36227
rect 17635 36187 17693 36193
rect 17754 36227 17812 36233
rect 17754 36193 17766 36227
rect 17800 36224 17812 36227
rect 17854 36227 17912 36233
rect 17800 36193 17813 36224
rect 17754 36187 17813 36193
rect 17854 36193 17866 36227
rect 17900 36193 17912 36227
rect 18046 36224 18052 36236
rect 18007 36196 18052 36224
rect 17854 36187 17912 36193
rect 16482 36156 16488 36168
rect 15672 36128 16488 36156
rect 16482 36116 16488 36128
rect 16540 36116 16546 36168
rect 16850 36116 16856 36168
rect 16908 36156 16914 36168
rect 17310 36156 17316 36168
rect 16908 36128 17316 36156
rect 16908 36116 16914 36128
rect 17310 36116 17316 36128
rect 17368 36116 17374 36168
rect 17402 36116 17408 36168
rect 17460 36156 17466 36168
rect 17460 36128 17505 36156
rect 17460 36116 17466 36128
rect 13688 36060 15608 36088
rect 13688 36048 13694 36060
rect 17494 36048 17500 36100
rect 17552 36088 17558 36100
rect 17785 36088 17813 36187
rect 17880 36100 17908 36187
rect 18046 36184 18052 36196
rect 18104 36184 18110 36236
rect 18598 36184 18604 36236
rect 18656 36224 18662 36236
rect 18966 36233 18972 36236
rect 18693 36227 18751 36233
rect 18693 36224 18705 36227
rect 18656 36196 18705 36224
rect 18656 36184 18662 36196
rect 18693 36193 18705 36196
rect 18739 36193 18751 36227
rect 18693 36187 18751 36193
rect 18960 36187 18972 36233
rect 19024 36224 19030 36236
rect 19024 36196 19060 36224
rect 18966 36184 18972 36187
rect 19024 36184 19030 36196
rect 17552 36060 17813 36088
rect 17552 36048 17558 36060
rect 17862 36048 17868 36100
rect 17920 36048 17926 36100
rect 22572 36088 22600 36332
rect 22738 36320 22744 36332
rect 22796 36320 22802 36372
rect 25409 36363 25467 36369
rect 25409 36329 25421 36363
rect 25455 36360 25467 36363
rect 25498 36360 25504 36372
rect 25455 36332 25504 36360
rect 25455 36329 25467 36332
rect 25409 36323 25467 36329
rect 25498 36320 25504 36332
rect 25556 36320 25562 36372
rect 25222 36252 25228 36304
rect 25280 36292 25286 36304
rect 27985 36295 28043 36301
rect 27985 36292 27997 36295
rect 25280 36264 27997 36292
rect 25280 36252 25286 36264
rect 27985 36261 27997 36264
rect 28031 36261 28043 36295
rect 27985 36255 28043 36261
rect 22971 36227 23029 36233
rect 22971 36224 22983 36227
rect 22848 36196 22983 36224
rect 22848 36156 22876 36196
rect 22971 36193 22983 36196
rect 23017 36193 23029 36227
rect 23106 36224 23112 36236
rect 23067 36196 23112 36224
rect 22971 36187 23029 36193
rect 23106 36184 23112 36196
rect 23164 36184 23170 36236
rect 23198 36184 23204 36236
rect 23256 36224 23262 36236
rect 23382 36224 23388 36236
rect 23256 36196 23301 36224
rect 23343 36196 23388 36224
rect 23256 36184 23262 36196
rect 23382 36184 23388 36196
rect 23440 36184 23446 36236
rect 25593 36227 25651 36233
rect 25593 36193 25605 36227
rect 25639 36224 25651 36227
rect 25866 36224 25872 36236
rect 25639 36196 25872 36224
rect 25639 36193 25651 36196
rect 25593 36187 25651 36193
rect 25866 36184 25872 36196
rect 25924 36184 25930 36236
rect 26142 36184 26148 36236
rect 26200 36224 26206 36236
rect 26237 36227 26295 36233
rect 26237 36224 26249 36227
rect 26200 36196 26249 36224
rect 26200 36184 26206 36196
rect 26237 36193 26249 36196
rect 26283 36193 26295 36227
rect 26878 36224 26884 36236
rect 26839 36196 26884 36224
rect 26237 36187 26295 36193
rect 26878 36184 26884 36196
rect 26936 36184 26942 36236
rect 23658 36156 23664 36168
rect 22848 36128 23664 36156
rect 23658 36116 23664 36128
rect 23716 36156 23722 36168
rect 24026 36156 24032 36168
rect 23716 36128 24032 36156
rect 23716 36116 23722 36128
rect 24026 36116 24032 36128
rect 24084 36116 24090 36168
rect 28169 36091 28227 36097
rect 28169 36088 28181 36091
rect 22572 36060 28181 36088
rect 28169 36057 28181 36060
rect 28215 36057 28227 36091
rect 28169 36051 28227 36057
rect 10796 35992 11468 36020
rect 11514 35980 11520 36032
rect 11572 36020 11578 36032
rect 12069 36023 12127 36029
rect 12069 36020 12081 36023
rect 11572 35992 12081 36020
rect 11572 35980 11578 35992
rect 12069 35989 12081 35992
rect 12115 35989 12127 36023
rect 12069 35983 12127 35989
rect 12158 35980 12164 36032
rect 12216 36020 12222 36032
rect 16206 36020 16212 36032
rect 12216 35992 16212 36020
rect 12216 35980 12222 35992
rect 16206 35980 16212 35992
rect 16264 35980 16270 36032
rect 16298 35980 16304 36032
rect 16356 36020 16362 36032
rect 18138 36020 18144 36032
rect 16356 35992 18144 36020
rect 16356 35980 16362 35992
rect 18138 35980 18144 35992
rect 18196 35980 18202 36032
rect 18230 35980 18236 36032
rect 18288 36020 18294 36032
rect 18966 36020 18972 36032
rect 18288 35992 18972 36020
rect 18288 35980 18294 35992
rect 18966 35980 18972 35992
rect 19024 35980 19030 36032
rect 19886 35980 19892 36032
rect 19944 36020 19950 36032
rect 20070 36020 20076 36032
rect 19944 35992 20076 36020
rect 19944 35980 19950 35992
rect 20070 35980 20076 35992
rect 20128 35980 20134 36032
rect 21174 35980 21180 36032
rect 21232 36020 21238 36032
rect 22646 36020 22652 36032
rect 21232 35992 22652 36020
rect 21232 35980 21238 35992
rect 22646 35980 22652 35992
rect 22704 35980 22710 36032
rect 22738 35980 22744 36032
rect 22796 36020 22802 36032
rect 23382 36020 23388 36032
rect 22796 35992 23388 36020
rect 22796 35980 22802 35992
rect 23382 35980 23388 35992
rect 23440 35980 23446 36032
rect 26050 36020 26056 36032
rect 26011 35992 26056 36020
rect 26050 35980 26056 35992
rect 26108 35980 26114 36032
rect 26697 36023 26755 36029
rect 26697 35989 26709 36023
rect 26743 36020 26755 36023
rect 27982 36020 27988 36032
rect 26743 35992 27988 36020
rect 26743 35989 26755 35992
rect 26697 35983 26755 35989
rect 27982 35980 27988 35992
rect 28040 35980 28046 36032
rect 1104 35930 28888 35952
rect 1104 35878 5614 35930
rect 5666 35878 5678 35930
rect 5730 35878 5742 35930
rect 5794 35878 5806 35930
rect 5858 35878 14878 35930
rect 14930 35878 14942 35930
rect 14994 35878 15006 35930
rect 15058 35878 15070 35930
rect 15122 35878 24142 35930
rect 24194 35878 24206 35930
rect 24258 35878 24270 35930
rect 24322 35878 24334 35930
rect 24386 35878 28888 35930
rect 1104 35856 28888 35878
rect 2406 35776 2412 35828
rect 2464 35816 2470 35828
rect 2464 35788 7144 35816
rect 2464 35776 2470 35788
rect 1762 35708 1768 35760
rect 1820 35748 1826 35760
rect 1857 35751 1915 35757
rect 1857 35748 1869 35751
rect 1820 35720 1869 35748
rect 1820 35708 1826 35720
rect 1857 35717 1869 35720
rect 1903 35717 1915 35751
rect 1857 35711 1915 35717
rect 2041 35751 2099 35757
rect 2041 35717 2053 35751
rect 2087 35748 2099 35751
rect 3142 35748 3148 35760
rect 2087 35720 3148 35748
rect 2087 35717 2099 35720
rect 2041 35711 2099 35717
rect 1872 35612 1900 35711
rect 3142 35708 3148 35720
rect 3200 35708 3206 35760
rect 3326 35708 3332 35760
rect 3384 35748 3390 35760
rect 3510 35748 3516 35760
rect 3384 35720 3516 35748
rect 3384 35708 3390 35720
rect 3510 35708 3516 35720
rect 3568 35748 3574 35760
rect 6638 35748 6644 35760
rect 3568 35720 6644 35748
rect 3568 35708 3574 35720
rect 6638 35708 6644 35720
rect 6696 35708 6702 35760
rect 3878 35680 3884 35692
rect 3068 35652 3884 35680
rect 2038 35612 2044 35624
rect 1872 35584 2044 35612
rect 2038 35572 2044 35584
rect 2096 35572 2102 35624
rect 3068 35621 3096 35652
rect 3878 35640 3884 35652
rect 3936 35680 3942 35692
rect 7116 35680 7144 35788
rect 7190 35776 7196 35828
rect 7248 35816 7254 35828
rect 7377 35819 7435 35825
rect 7377 35816 7389 35819
rect 7248 35788 7389 35816
rect 7248 35776 7254 35788
rect 7377 35785 7389 35788
rect 7423 35785 7435 35819
rect 7377 35779 7435 35785
rect 9950 35776 9956 35828
rect 10008 35816 10014 35828
rect 10410 35816 10416 35828
rect 10008 35788 10416 35816
rect 10008 35776 10014 35788
rect 10410 35776 10416 35788
rect 10468 35816 10474 35828
rect 11054 35816 11060 35828
rect 10468 35788 11060 35816
rect 10468 35776 10474 35788
rect 11054 35776 11060 35788
rect 11112 35776 11118 35828
rect 12069 35819 12127 35825
rect 12069 35785 12081 35819
rect 12115 35816 12127 35819
rect 12802 35816 12808 35828
rect 12115 35788 12808 35816
rect 12115 35785 12127 35788
rect 12069 35779 12127 35785
rect 12802 35776 12808 35788
rect 12860 35776 12866 35828
rect 13633 35819 13691 35825
rect 13633 35785 13645 35819
rect 13679 35816 13691 35819
rect 13814 35816 13820 35828
rect 13679 35788 13820 35816
rect 13679 35785 13691 35788
rect 13633 35779 13691 35785
rect 13814 35776 13820 35788
rect 13872 35776 13878 35828
rect 28077 35819 28135 35825
rect 28077 35816 28089 35819
rect 13924 35788 28089 35816
rect 13538 35748 13544 35760
rect 11900 35720 13544 35748
rect 9769 35683 9827 35689
rect 3936 35652 4292 35680
rect 7116 35652 9628 35680
rect 3936 35640 3942 35652
rect 3053 35615 3111 35621
rect 3053 35581 3065 35615
rect 3099 35581 3111 35615
rect 3053 35575 3111 35581
rect 3329 35615 3387 35621
rect 3329 35581 3341 35615
rect 3375 35612 3387 35615
rect 3602 35612 3608 35624
rect 3375 35584 3608 35612
rect 3375 35581 3387 35584
rect 3329 35575 3387 35581
rect 3602 35572 3608 35584
rect 3660 35572 3666 35624
rect 4264 35621 4292 35652
rect 4249 35615 4307 35621
rect 4249 35581 4261 35615
rect 4295 35581 4307 35615
rect 4249 35575 4307 35581
rect 7193 35615 7251 35621
rect 7193 35581 7205 35615
rect 7239 35612 7251 35615
rect 7282 35612 7288 35624
rect 7239 35584 7288 35612
rect 7239 35581 7251 35584
rect 7193 35575 7251 35581
rect 7282 35572 7288 35584
rect 7340 35572 7346 35624
rect 9398 35572 9404 35624
rect 9456 35612 9462 35624
rect 9493 35615 9551 35621
rect 9493 35612 9505 35615
rect 9456 35584 9505 35612
rect 9456 35572 9462 35584
rect 9493 35581 9505 35584
rect 9539 35581 9551 35615
rect 9600 35612 9628 35652
rect 9769 35649 9781 35683
rect 9815 35680 9827 35683
rect 10502 35680 10508 35692
rect 9815 35652 10508 35680
rect 9815 35649 9827 35652
rect 9769 35643 9827 35649
rect 10502 35640 10508 35652
rect 10560 35640 10566 35692
rect 11606 35640 11612 35692
rect 11664 35680 11670 35692
rect 11664 35652 11836 35680
rect 11664 35640 11670 35652
rect 11698 35612 11704 35624
rect 9600 35584 11560 35612
rect 11659 35584 11704 35612
rect 9493 35575 9551 35581
rect 1486 35504 1492 35556
rect 1544 35544 1550 35556
rect 1581 35547 1639 35553
rect 1581 35544 1593 35547
rect 1544 35516 1593 35544
rect 1544 35504 1550 35516
rect 1581 35513 1593 35516
rect 1627 35513 1639 35547
rect 1581 35507 1639 35513
rect 1854 35504 1860 35556
rect 1912 35544 1918 35556
rect 6914 35544 6920 35556
rect 1912 35516 6920 35544
rect 1912 35504 1918 35516
rect 6914 35504 6920 35516
rect 6972 35504 6978 35556
rect 7009 35547 7067 35553
rect 7009 35513 7021 35547
rect 7055 35544 7067 35547
rect 8018 35544 8024 35556
rect 7055 35516 8024 35544
rect 7055 35513 7067 35516
rect 7009 35507 7067 35513
rect 8018 35504 8024 35516
rect 8076 35544 8082 35556
rect 9122 35544 9128 35556
rect 8076 35516 9128 35544
rect 8076 35504 8082 35516
rect 9122 35504 9128 35516
rect 9180 35504 9186 35556
rect 11532 35544 11560 35584
rect 11698 35572 11704 35584
rect 11756 35572 11762 35624
rect 11808 35621 11836 35652
rect 11900 35621 11928 35720
rect 13538 35708 13544 35720
rect 13596 35708 13602 35760
rect 13924 35680 13952 35788
rect 28077 35785 28089 35788
rect 28123 35785 28135 35819
rect 28077 35779 28135 35785
rect 15562 35708 15568 35760
rect 15620 35748 15626 35760
rect 16114 35748 16120 35760
rect 15620 35720 16120 35748
rect 15620 35708 15626 35720
rect 16114 35708 16120 35720
rect 16172 35708 16178 35760
rect 18230 35748 18236 35760
rect 18191 35720 18236 35748
rect 18230 35708 18236 35720
rect 18288 35708 18294 35760
rect 18782 35708 18788 35760
rect 18840 35748 18846 35760
rect 19426 35748 19432 35760
rect 18840 35720 19432 35748
rect 18840 35708 18846 35720
rect 19426 35708 19432 35720
rect 19484 35708 19490 35760
rect 22557 35751 22615 35757
rect 22557 35717 22569 35751
rect 22603 35748 22615 35751
rect 22646 35748 22652 35760
rect 22603 35720 22652 35748
rect 22603 35717 22615 35720
rect 22557 35711 22615 35717
rect 22646 35708 22652 35720
rect 22704 35708 22710 35760
rect 23014 35748 23020 35760
rect 22975 35720 23020 35748
rect 23014 35708 23020 35720
rect 23072 35708 23078 35760
rect 23198 35708 23204 35760
rect 23256 35748 23262 35760
rect 23256 35720 24164 35748
rect 23256 35708 23262 35720
rect 12084 35652 13952 35680
rect 11793 35615 11851 35621
rect 11793 35581 11805 35615
rect 11839 35581 11851 35615
rect 11793 35575 11851 35581
rect 11885 35615 11943 35621
rect 11885 35581 11897 35615
rect 11931 35581 11943 35615
rect 12084 35612 12112 35652
rect 14182 35640 14188 35692
rect 14240 35680 14246 35692
rect 16666 35680 16672 35692
rect 14240 35652 16672 35680
rect 14240 35640 14246 35652
rect 16666 35640 16672 35652
rect 16724 35640 16730 35692
rect 17494 35640 17500 35692
rect 17552 35680 17558 35692
rect 17552 35652 18644 35680
rect 17552 35640 17558 35652
rect 11885 35575 11943 35581
rect 11992 35584 12112 35612
rect 13265 35615 13323 35621
rect 11992 35544 12020 35584
rect 13265 35581 13277 35615
rect 13311 35581 13323 35615
rect 13265 35575 13323 35581
rect 13357 35615 13415 35621
rect 13357 35581 13369 35615
rect 13403 35581 13415 35615
rect 13357 35575 13415 35581
rect 13449 35615 13507 35621
rect 13449 35581 13461 35615
rect 13495 35612 13507 35615
rect 13538 35612 13544 35624
rect 13495 35584 13544 35612
rect 13495 35581 13507 35584
rect 13449 35575 13507 35581
rect 11532 35516 12020 35544
rect 2866 35476 2872 35488
rect 2827 35448 2872 35476
rect 2866 35436 2872 35448
rect 2924 35436 2930 35488
rect 3234 35476 3240 35488
rect 3195 35448 3240 35476
rect 3234 35436 3240 35448
rect 3292 35436 3298 35488
rect 4338 35436 4344 35488
rect 4396 35476 4402 35488
rect 4433 35479 4491 35485
rect 4433 35476 4445 35479
rect 4396 35448 4445 35476
rect 4396 35436 4402 35448
rect 4433 35445 4445 35448
rect 4479 35445 4491 35479
rect 4433 35439 4491 35445
rect 9858 35436 9864 35488
rect 9916 35476 9922 35488
rect 11606 35476 11612 35488
rect 9916 35448 11612 35476
rect 9916 35436 9922 35448
rect 11606 35436 11612 35448
rect 11664 35436 11670 35488
rect 11698 35436 11704 35488
rect 11756 35476 11762 35488
rect 12342 35476 12348 35488
rect 11756 35448 12348 35476
rect 11756 35436 11762 35448
rect 12342 35436 12348 35448
rect 12400 35476 12406 35488
rect 13280 35476 13308 35575
rect 13372 35544 13400 35575
rect 13538 35572 13544 35584
rect 13596 35572 13602 35624
rect 14550 35572 14556 35624
rect 14608 35612 14614 35624
rect 14737 35615 14795 35621
rect 14737 35612 14749 35615
rect 14608 35584 14749 35612
rect 14608 35572 14614 35584
rect 14737 35581 14749 35584
rect 14783 35581 14795 35615
rect 14737 35575 14795 35581
rect 15194 35572 15200 35624
rect 15252 35612 15258 35624
rect 15933 35615 15991 35621
rect 15933 35612 15945 35615
rect 15252 35584 15945 35612
rect 15252 35572 15258 35584
rect 15933 35581 15945 35584
rect 15979 35612 15991 35615
rect 16114 35612 16120 35624
rect 15979 35584 16120 35612
rect 15979 35581 15991 35584
rect 15933 35575 15991 35581
rect 16114 35572 16120 35584
rect 16172 35612 16178 35624
rect 16482 35612 16488 35624
rect 16172 35584 16488 35612
rect 16172 35572 16178 35584
rect 16482 35572 16488 35584
rect 16540 35612 16546 35624
rect 16761 35615 16819 35621
rect 16761 35612 16773 35615
rect 16540 35584 16773 35612
rect 16540 35572 16546 35584
rect 16761 35581 16773 35584
rect 16807 35581 16819 35615
rect 18506 35612 18512 35624
rect 18467 35584 18512 35612
rect 16761 35575 16819 35581
rect 18506 35572 18512 35584
rect 18564 35572 18570 35624
rect 18616 35621 18644 35652
rect 20530 35640 20536 35692
rect 20588 35680 20594 35692
rect 20588 35652 21312 35680
rect 20588 35640 20594 35652
rect 18601 35615 18659 35621
rect 18601 35581 18613 35615
rect 18647 35581 18659 35615
rect 18601 35575 18659 35581
rect 18693 35615 18751 35621
rect 18693 35581 18705 35615
rect 18739 35581 18751 35615
rect 18693 35575 18751 35581
rect 18889 35615 18947 35621
rect 18889 35581 18901 35615
rect 18935 35612 18947 35615
rect 19150 35612 19156 35624
rect 18935 35584 19156 35612
rect 18935 35581 18947 35584
rect 18889 35575 18947 35581
rect 13630 35544 13636 35556
rect 13372 35516 13636 35544
rect 13630 35504 13636 35516
rect 13688 35544 13694 35556
rect 13998 35544 14004 35556
rect 13688 35516 14004 35544
rect 13688 35504 13694 35516
rect 13998 35504 14004 35516
rect 14056 35504 14062 35556
rect 16945 35547 17003 35553
rect 16945 35513 16957 35547
rect 16991 35544 17003 35547
rect 17862 35544 17868 35556
rect 16991 35516 17868 35544
rect 16991 35513 17003 35516
rect 16945 35507 17003 35513
rect 17862 35504 17868 35516
rect 17920 35544 17926 35556
rect 18230 35544 18236 35556
rect 17920 35516 18236 35544
rect 17920 35504 17926 35516
rect 18230 35504 18236 35516
rect 18288 35544 18294 35556
rect 18708 35544 18736 35575
rect 19150 35572 19156 35584
rect 19208 35572 19214 35624
rect 20806 35572 20812 35624
rect 20864 35612 20870 35624
rect 21177 35615 21235 35621
rect 21177 35612 21189 35615
rect 20864 35584 21189 35612
rect 20864 35572 20870 35584
rect 21177 35581 21189 35584
rect 21223 35581 21235 35615
rect 21284 35612 21312 35652
rect 23106 35640 23112 35692
rect 23164 35680 23170 35692
rect 24136 35680 24164 35720
rect 24394 35680 24400 35692
rect 23164 35652 24072 35680
rect 23164 35640 23170 35652
rect 23201 35615 23259 35621
rect 23201 35612 23213 35615
rect 21284 35584 23213 35612
rect 21177 35575 21235 35581
rect 23201 35581 23213 35584
rect 23247 35581 23259 35615
rect 23201 35575 23259 35581
rect 23842 35572 23848 35624
rect 23900 35621 23906 35624
rect 24044 35621 24072 35652
rect 24136 35652 24400 35680
rect 24136 35621 24164 35652
rect 24394 35640 24400 35652
rect 24452 35640 24458 35692
rect 24854 35640 24860 35692
rect 24912 35680 24918 35692
rect 25225 35683 25283 35689
rect 25225 35680 25237 35683
rect 24912 35652 25237 35680
rect 24912 35640 24918 35652
rect 25225 35649 25237 35652
rect 25271 35649 25283 35683
rect 25225 35643 25283 35649
rect 23900 35615 23949 35621
rect 23900 35581 23903 35615
rect 23937 35581 23949 35615
rect 23900 35575 23949 35581
rect 24029 35615 24087 35621
rect 24029 35581 24041 35615
rect 24075 35581 24087 35615
rect 24029 35575 24087 35581
rect 24121 35615 24179 35621
rect 24121 35581 24133 35615
rect 24167 35581 24179 35615
rect 24121 35575 24179 35581
rect 24305 35615 24363 35621
rect 24305 35581 24317 35615
rect 24351 35612 24363 35615
rect 24578 35612 24584 35624
rect 24351 35584 24584 35612
rect 24351 35581 24363 35584
rect 24305 35575 24363 35581
rect 23900 35572 23906 35575
rect 24578 35572 24584 35584
rect 24636 35572 24642 35624
rect 26050 35572 26056 35624
rect 26108 35612 26114 35624
rect 27249 35615 27307 35621
rect 27249 35612 27261 35615
rect 26108 35584 27261 35612
rect 26108 35572 26114 35584
rect 27249 35581 27261 35584
rect 27295 35581 27307 35615
rect 27249 35575 27307 35581
rect 27890 35572 27896 35624
rect 27948 35612 27954 35624
rect 27985 35615 28043 35621
rect 27985 35612 27997 35615
rect 27948 35584 27997 35612
rect 27948 35572 27954 35584
rect 27985 35581 27997 35584
rect 28031 35581 28043 35615
rect 27985 35575 28043 35581
rect 20070 35544 20076 35556
rect 18288 35516 20076 35544
rect 18288 35504 18294 35516
rect 20070 35504 20076 35516
rect 20128 35504 20134 35556
rect 20714 35504 20720 35556
rect 20772 35544 20778 35556
rect 21422 35547 21480 35553
rect 21422 35544 21434 35547
rect 20772 35516 21434 35544
rect 20772 35504 20778 35516
rect 21422 35513 21434 35516
rect 21468 35513 21480 35547
rect 21422 35507 21480 35513
rect 23661 35547 23719 35553
rect 23661 35513 23673 35547
rect 23707 35544 23719 35547
rect 25470 35547 25528 35553
rect 25470 35544 25482 35547
rect 23707 35516 25482 35544
rect 23707 35513 23719 35516
rect 23661 35507 23719 35513
rect 25470 35513 25482 35516
rect 25516 35513 25528 35547
rect 27433 35547 27491 35553
rect 27433 35544 27445 35547
rect 25470 35507 25528 35513
rect 25608 35516 27445 35544
rect 13722 35476 13728 35488
rect 12400 35448 13728 35476
rect 12400 35436 12406 35448
rect 13722 35436 13728 35448
rect 13780 35436 13786 35488
rect 14550 35436 14556 35488
rect 14608 35476 14614 35488
rect 14829 35479 14887 35485
rect 14829 35476 14841 35479
rect 14608 35448 14841 35476
rect 14608 35436 14614 35448
rect 14829 35445 14841 35448
rect 14875 35445 14887 35479
rect 16022 35476 16028 35488
rect 15983 35448 16028 35476
rect 14829 35439 14887 35445
rect 16022 35436 16028 35448
rect 16080 35436 16086 35488
rect 16206 35436 16212 35488
rect 16264 35476 16270 35488
rect 25608 35476 25636 35516
rect 27433 35513 27445 35516
rect 27479 35513 27491 35547
rect 27433 35507 27491 35513
rect 26602 35476 26608 35488
rect 16264 35448 25636 35476
rect 26563 35448 26608 35476
rect 16264 35436 16270 35448
rect 26602 35436 26608 35448
rect 26660 35436 26666 35488
rect 1104 35386 28888 35408
rect 1104 35334 10246 35386
rect 10298 35334 10310 35386
rect 10362 35334 10374 35386
rect 10426 35334 10438 35386
rect 10490 35334 19510 35386
rect 19562 35334 19574 35386
rect 19626 35334 19638 35386
rect 19690 35334 19702 35386
rect 19754 35334 28888 35386
rect 1104 35312 28888 35334
rect 2409 35275 2467 35281
rect 2409 35241 2421 35275
rect 2455 35272 2467 35275
rect 3234 35272 3240 35284
rect 2455 35244 3240 35272
rect 2455 35241 2467 35244
rect 2409 35235 2467 35241
rect 3234 35232 3240 35244
rect 3292 35232 3298 35284
rect 3602 35272 3608 35284
rect 3563 35244 3608 35272
rect 3602 35232 3608 35244
rect 3660 35232 3666 35284
rect 9953 35275 10011 35281
rect 9953 35241 9965 35275
rect 9999 35272 10011 35275
rect 11146 35272 11152 35284
rect 9999 35244 11152 35272
rect 9999 35241 10011 35244
rect 9953 35235 10011 35241
rect 11146 35232 11152 35244
rect 11204 35232 11210 35284
rect 12805 35275 12863 35281
rect 12805 35241 12817 35275
rect 12851 35272 12863 35275
rect 13078 35272 13084 35284
rect 12851 35244 13084 35272
rect 12851 35241 12863 35244
rect 12805 35235 12863 35241
rect 13078 35232 13084 35244
rect 13136 35232 13142 35284
rect 13449 35275 13507 35281
rect 13449 35241 13461 35275
rect 13495 35272 13507 35275
rect 13906 35272 13912 35284
rect 13495 35244 13912 35272
rect 13495 35241 13507 35244
rect 13449 35235 13507 35241
rect 13906 35232 13912 35244
rect 13964 35232 13970 35284
rect 14550 35232 14556 35284
rect 14608 35272 14614 35284
rect 14737 35275 14795 35281
rect 14608 35244 14688 35272
rect 14608 35232 14614 35244
rect 1581 35207 1639 35213
rect 1581 35173 1593 35207
rect 1627 35204 1639 35207
rect 10318 35204 10324 35216
rect 1627 35176 10324 35204
rect 1627 35173 1639 35176
rect 1581 35167 1639 35173
rect 10318 35164 10324 35176
rect 10376 35164 10382 35216
rect 10962 35204 10968 35216
rect 10796 35176 10968 35204
rect 2501 35139 2559 35145
rect 2501 35105 2513 35139
rect 2547 35105 2559 35139
rect 2501 35099 2559 35105
rect 2685 35139 2743 35145
rect 2685 35105 2697 35139
rect 2731 35136 2743 35139
rect 3234 35136 3240 35148
rect 2731 35108 3240 35136
rect 2731 35105 2743 35108
rect 2685 35099 2743 35105
rect 2516 35068 2544 35099
rect 3234 35096 3240 35108
rect 3292 35096 3298 35148
rect 3329 35139 3387 35145
rect 3329 35105 3341 35139
rect 3375 35105 3387 35139
rect 3329 35099 3387 35105
rect 3142 35068 3148 35080
rect 2516 35040 3148 35068
rect 3142 35028 3148 35040
rect 3200 35028 3206 35080
rect 3344 35068 3372 35099
rect 3418 35096 3424 35148
rect 3476 35136 3482 35148
rect 4433 35139 4491 35145
rect 3476 35108 3521 35136
rect 3476 35096 3482 35108
rect 4433 35105 4445 35139
rect 4479 35136 4491 35139
rect 4522 35136 4528 35148
rect 4479 35108 4528 35136
rect 4479 35105 4491 35108
rect 4433 35099 4491 35105
rect 4522 35096 4528 35108
rect 4580 35096 4586 35148
rect 4700 35139 4758 35145
rect 4700 35105 4712 35139
rect 4746 35136 4758 35139
rect 4982 35136 4988 35148
rect 4746 35108 4988 35136
rect 4746 35105 4758 35108
rect 4700 35099 4758 35105
rect 4982 35096 4988 35108
rect 5040 35096 5046 35148
rect 7929 35139 7987 35145
rect 7929 35105 7941 35139
rect 7975 35136 7987 35139
rect 9490 35136 9496 35148
rect 7975 35108 9496 35136
rect 7975 35105 7987 35108
rect 7929 35099 7987 35105
rect 9490 35096 9496 35108
rect 9548 35096 9554 35148
rect 9769 35139 9827 35145
rect 9769 35105 9781 35139
rect 9815 35136 9827 35139
rect 9858 35136 9864 35148
rect 9815 35108 9864 35136
rect 9815 35105 9827 35108
rect 9769 35099 9827 35105
rect 9858 35096 9864 35108
rect 9916 35096 9922 35148
rect 9953 35139 10011 35145
rect 9953 35105 9965 35139
rect 9999 35136 10011 35139
rect 10502 35136 10508 35148
rect 9999 35108 10508 35136
rect 9999 35105 10011 35108
rect 9953 35099 10011 35105
rect 10502 35096 10508 35108
rect 10560 35096 10566 35148
rect 10796 35145 10824 35176
rect 10962 35164 10968 35176
rect 11020 35164 11026 35216
rect 14660 35204 14688 35244
rect 14737 35241 14749 35275
rect 14783 35272 14795 35275
rect 15562 35272 15568 35284
rect 14783 35244 15568 35272
rect 14783 35241 14795 35244
rect 14737 35235 14795 35241
rect 15562 35232 15568 35244
rect 15620 35232 15626 35284
rect 16114 35272 16120 35284
rect 16075 35244 16120 35272
rect 16114 35232 16120 35244
rect 16172 35232 16178 35284
rect 17681 35275 17739 35281
rect 17681 35241 17693 35275
rect 17727 35272 17739 35275
rect 17954 35272 17960 35284
rect 17727 35244 17960 35272
rect 17727 35241 17739 35244
rect 17681 35235 17739 35241
rect 17954 35232 17960 35244
rect 18012 35232 18018 35284
rect 18506 35232 18512 35284
rect 18564 35272 18570 35284
rect 19886 35272 19892 35284
rect 18564 35244 19892 35272
rect 18564 35232 18570 35244
rect 19886 35232 19892 35244
rect 19944 35232 19950 35284
rect 23106 35272 23112 35284
rect 19996 35244 23112 35272
rect 12544 35176 13308 35204
rect 14660 35176 15976 35204
rect 12544 35148 12572 35176
rect 10689 35139 10747 35145
rect 10689 35105 10701 35139
rect 10735 35105 10747 35139
rect 10689 35099 10747 35105
rect 10781 35139 10839 35145
rect 10781 35105 10793 35139
rect 10827 35105 10839 35139
rect 10781 35099 10839 35105
rect 10410 35068 10416 35080
rect 3252 35040 3372 35068
rect 5736 35040 10416 35068
rect 3252 35000 3280 35040
rect 2240 34972 3280 35000
rect 2240 34944 2268 34972
rect 1670 34932 1676 34944
rect 1631 34904 1676 34932
rect 1670 34892 1676 34904
rect 1728 34892 1734 34944
rect 2222 34932 2228 34944
rect 2183 34904 2228 34932
rect 2222 34892 2228 34904
rect 2280 34892 2286 34944
rect 2406 34892 2412 34944
rect 2464 34932 2470 34944
rect 5736 34932 5764 35040
rect 10410 35028 10416 35040
rect 10468 35028 10474 35080
rect 10704 35068 10732 35099
rect 10870 35096 10876 35148
rect 10928 35136 10934 35148
rect 11054 35136 11060 35148
rect 10928 35108 10973 35136
rect 11015 35108 11060 35136
rect 10928 35096 10934 35108
rect 11054 35096 11060 35108
rect 11112 35096 11118 35148
rect 12342 35096 12348 35148
rect 12400 35145 12406 35148
rect 12400 35139 12459 35145
rect 12400 35105 12413 35139
rect 12447 35105 12459 35139
rect 12526 35136 12532 35148
rect 12487 35108 12532 35136
rect 12400 35099 12459 35105
rect 12400 35096 12406 35099
rect 12526 35096 12532 35108
rect 12584 35096 12590 35148
rect 12621 35139 12679 35145
rect 12621 35105 12633 35139
rect 12667 35136 12679 35139
rect 12802 35136 12808 35148
rect 12667 35108 12808 35136
rect 12667 35105 12679 35108
rect 12621 35099 12679 35105
rect 12802 35096 12808 35108
rect 12860 35096 12866 35148
rect 13280 35145 13308 35176
rect 13265 35139 13323 35145
rect 13265 35105 13277 35139
rect 13311 35105 13323 35139
rect 13446 35136 13452 35148
rect 13407 35108 13452 35136
rect 13265 35099 13323 35105
rect 13446 35096 13452 35108
rect 13504 35096 13510 35148
rect 13998 35096 14004 35148
rect 14056 35136 14062 35148
rect 14553 35139 14611 35145
rect 14553 35136 14565 35139
rect 14056 35108 14565 35136
rect 14056 35096 14062 35108
rect 14553 35105 14565 35108
rect 14599 35105 14611 35139
rect 14553 35099 14611 35105
rect 14737 35139 14795 35145
rect 14737 35105 14749 35139
rect 14783 35136 14795 35139
rect 14826 35136 14832 35148
rect 14783 35108 14832 35136
rect 14783 35105 14795 35108
rect 14737 35099 14795 35105
rect 14826 35096 14832 35108
rect 14884 35096 14890 35148
rect 15286 35096 15292 35148
rect 15344 35136 15350 35148
rect 15948 35145 15976 35176
rect 17494 35164 17500 35216
rect 17552 35204 17558 35216
rect 19153 35207 19211 35213
rect 17552 35176 18092 35204
rect 17552 35164 17558 35176
rect 15933 35139 15991 35145
rect 15344 35108 15389 35136
rect 15344 35096 15350 35108
rect 15933 35105 15945 35139
rect 15979 35105 15991 35139
rect 15933 35099 15991 35105
rect 17402 35096 17408 35148
rect 17460 35136 17466 35148
rect 18064 35145 18092 35176
rect 19153 35173 19165 35207
rect 19199 35204 19211 35207
rect 19996 35204 20024 35244
rect 19199 35176 20024 35204
rect 19199 35173 19211 35176
rect 19153 35167 19211 35173
rect 17911 35139 17969 35145
rect 17911 35136 17923 35139
rect 17460 35108 17923 35136
rect 17460 35096 17466 35108
rect 17911 35105 17923 35108
rect 17957 35105 17969 35139
rect 17911 35099 17969 35105
rect 18049 35139 18107 35145
rect 18049 35105 18061 35139
rect 18095 35105 18107 35139
rect 18049 35099 18107 35105
rect 18141 35139 18199 35145
rect 18141 35105 18153 35139
rect 18187 35136 18199 35139
rect 18230 35136 18236 35148
rect 18187 35108 18236 35136
rect 18187 35105 18199 35108
rect 18141 35099 18199 35105
rect 18230 35096 18236 35108
rect 18288 35096 18294 35148
rect 18325 35139 18383 35145
rect 18325 35105 18337 35139
rect 18371 35136 18383 35139
rect 18598 35136 18604 35148
rect 18371 35108 18604 35136
rect 18371 35105 18383 35108
rect 18325 35099 18383 35105
rect 18598 35096 18604 35108
rect 18656 35096 18662 35148
rect 18690 35096 18696 35148
rect 18748 35136 18754 35148
rect 18969 35139 19027 35145
rect 18969 35136 18981 35139
rect 18748 35108 18981 35136
rect 18748 35096 18754 35108
rect 18969 35105 18981 35108
rect 19015 35105 19027 35139
rect 18969 35099 19027 35105
rect 19702 35096 19708 35148
rect 19760 35136 19766 35148
rect 19996 35145 20024 35176
rect 20180 35176 20576 35204
rect 19843 35139 19901 35145
rect 19843 35136 19855 35139
rect 19760 35108 19855 35136
rect 19760 35096 19766 35108
rect 19843 35105 19855 35108
rect 19889 35105 19901 35139
rect 19843 35099 19901 35105
rect 19981 35139 20039 35145
rect 19981 35105 19993 35139
rect 20027 35105 20039 35139
rect 19981 35099 20039 35105
rect 20070 35096 20076 35148
rect 20128 35136 20134 35148
rect 20180 35136 20208 35176
rect 20257 35139 20315 35145
rect 20128 35108 20221 35136
rect 20128 35096 20134 35108
rect 20257 35105 20269 35139
rect 20303 35136 20315 35139
rect 20438 35136 20444 35148
rect 20303 35108 20444 35136
rect 20303 35105 20315 35108
rect 20257 35099 20315 35105
rect 20438 35096 20444 35108
rect 20496 35096 20502 35148
rect 20548 35136 20576 35176
rect 20714 35164 20720 35216
rect 20772 35204 20778 35216
rect 20901 35207 20959 35213
rect 20901 35204 20913 35207
rect 20772 35176 20913 35204
rect 20772 35164 20778 35176
rect 20901 35173 20913 35176
rect 20947 35173 20959 35207
rect 20901 35167 20959 35173
rect 21174 35145 21180 35148
rect 21157 35139 21180 35145
rect 20548 35108 21128 35136
rect 11330 35068 11336 35080
rect 10704 35040 11336 35068
rect 11330 35028 11336 35040
rect 11388 35028 11394 35080
rect 12066 35028 12072 35080
rect 12124 35068 12130 35080
rect 20990 35068 20996 35080
rect 12124 35040 20996 35068
rect 12124 35028 12130 35040
rect 20990 35028 20996 35040
rect 21048 35028 21054 35080
rect 21100 35068 21128 35108
rect 21157 35105 21169 35139
rect 21157 35099 21180 35105
rect 21174 35096 21180 35099
rect 21232 35096 21238 35148
rect 21284 35145 21312 35244
rect 23106 35232 23112 35244
rect 23164 35232 23170 35284
rect 23477 35275 23535 35281
rect 23477 35241 23489 35275
rect 23523 35272 23535 35275
rect 24578 35272 24584 35284
rect 23523 35244 24584 35272
rect 23523 35241 23535 35244
rect 23477 35235 23535 35241
rect 24578 35232 24584 35244
rect 24636 35232 24642 35284
rect 24854 35232 24860 35284
rect 24912 35272 24918 35284
rect 25774 35272 25780 35284
rect 24912 35244 25780 35272
rect 24912 35232 24918 35244
rect 25774 35232 25780 35244
rect 25832 35272 25838 35284
rect 26421 35275 26479 35281
rect 26421 35272 26433 35275
rect 25832 35244 26433 35272
rect 25832 35232 25838 35244
rect 26421 35241 26433 35244
rect 26467 35241 26479 35275
rect 26421 35235 26479 35241
rect 23124 35204 23152 35232
rect 23937 35207 23995 35213
rect 23124 35176 23888 35204
rect 21269 35139 21327 35145
rect 21269 35105 21281 35139
rect 21315 35105 21327 35139
rect 21269 35099 21327 35105
rect 21361 35139 21419 35145
rect 21361 35105 21373 35139
rect 21407 35105 21419 35139
rect 21542 35136 21548 35148
rect 21503 35108 21548 35136
rect 21361 35099 21419 35105
rect 21376 35068 21404 35099
rect 21542 35096 21548 35108
rect 21600 35096 21606 35148
rect 22462 35096 22468 35148
rect 22520 35136 22526 35148
rect 23198 35145 23204 35148
rect 23073 35139 23131 35145
rect 23073 35136 23085 35139
rect 22520 35108 23085 35136
rect 22520 35096 22526 35108
rect 23073 35105 23085 35108
rect 23119 35105 23131 35139
rect 23191 35139 23204 35145
rect 23191 35136 23203 35139
rect 23159 35108 23203 35136
rect 23073 35099 23131 35105
rect 23191 35105 23203 35108
rect 23191 35099 23204 35105
rect 23198 35096 23204 35099
rect 23256 35096 23262 35148
rect 23293 35139 23351 35145
rect 23293 35105 23305 35139
rect 23339 35136 23351 35139
rect 23382 35136 23388 35148
rect 23339 35108 23388 35136
rect 23339 35105 23351 35108
rect 23293 35099 23351 35105
rect 23382 35096 23388 35108
rect 23440 35096 23446 35148
rect 21100 35040 21404 35068
rect 23860 35068 23888 35176
rect 23937 35173 23949 35207
rect 23983 35204 23995 35207
rect 25286 35207 25344 35213
rect 25286 35204 25298 35207
rect 23983 35176 25298 35204
rect 23983 35173 23995 35176
rect 23937 35167 23995 35173
rect 25286 35173 25298 35176
rect 25332 35173 25344 35207
rect 27982 35204 27988 35216
rect 27943 35176 27988 35204
rect 25286 35167 25344 35173
rect 27982 35164 27988 35176
rect 28040 35164 28046 35216
rect 24210 35136 24216 35148
rect 24171 35108 24216 35136
rect 24210 35096 24216 35108
rect 24268 35096 24274 35148
rect 24305 35139 24363 35145
rect 24305 35105 24317 35139
rect 24351 35105 24363 35139
rect 24305 35099 24363 35105
rect 24320 35068 24348 35099
rect 24394 35096 24400 35148
rect 24452 35136 24458 35148
rect 24578 35136 24584 35148
rect 24452 35108 24497 35136
rect 24539 35108 24584 35136
rect 24452 35096 24458 35108
rect 24578 35096 24584 35108
rect 24636 35096 24642 35148
rect 24762 35096 24768 35148
rect 24820 35136 24826 35148
rect 25041 35139 25099 35145
rect 25041 35136 25053 35139
rect 24820 35108 25053 35136
rect 24820 35096 24826 35108
rect 25041 35105 25053 35108
rect 25087 35105 25099 35139
rect 25041 35099 25099 35105
rect 23860 35040 24348 35068
rect 6914 34960 6920 35012
rect 6972 35000 6978 35012
rect 6972 34972 10640 35000
rect 6972 34960 6978 34972
rect 2464 34904 5764 34932
rect 5813 34935 5871 34941
rect 2464 34892 2470 34904
rect 5813 34901 5825 34935
rect 5859 34932 5871 34935
rect 5902 34932 5908 34944
rect 5859 34904 5908 34932
rect 5859 34901 5871 34904
rect 5813 34895 5871 34901
rect 5902 34892 5908 34904
rect 5960 34892 5966 34944
rect 7742 34932 7748 34944
rect 7703 34904 7748 34932
rect 7742 34892 7748 34904
rect 7800 34892 7806 34944
rect 10410 34932 10416 34944
rect 10371 34904 10416 34932
rect 10410 34892 10416 34904
rect 10468 34892 10474 34944
rect 10612 34932 10640 34972
rect 11440 34972 19932 35000
rect 11440 34932 11468 34972
rect 10612 34904 11468 34932
rect 12802 34892 12808 34944
rect 12860 34932 12866 34944
rect 13538 34932 13544 34944
rect 12860 34904 13544 34932
rect 12860 34892 12866 34904
rect 13538 34892 13544 34904
rect 13596 34932 13602 34944
rect 15381 34935 15439 34941
rect 15381 34932 15393 34935
rect 13596 34904 15393 34932
rect 13596 34892 13602 34904
rect 15381 34901 15393 34904
rect 15427 34932 15439 34935
rect 16022 34932 16028 34944
rect 15427 34904 16028 34932
rect 15427 34901 15439 34904
rect 15381 34895 15439 34901
rect 16022 34892 16028 34904
rect 16080 34892 16086 34944
rect 17218 34892 17224 34944
rect 17276 34932 17282 34944
rect 17494 34932 17500 34944
rect 17276 34904 17500 34932
rect 17276 34892 17282 34904
rect 17494 34892 17500 34904
rect 17552 34892 17558 34944
rect 19610 34932 19616 34944
rect 19571 34904 19616 34932
rect 19610 34892 19616 34904
rect 19668 34892 19674 34944
rect 19904 34932 19932 34972
rect 19978 34960 19984 35012
rect 20036 35000 20042 35012
rect 22370 35000 22376 35012
rect 20036 34972 22376 35000
rect 20036 34960 20042 34972
rect 22370 34960 22376 34972
rect 22428 35000 22434 35012
rect 23014 35000 23020 35012
rect 22428 34972 23020 35000
rect 22428 34960 22434 34972
rect 23014 34960 23020 34972
rect 23072 34960 23078 35012
rect 24210 34960 24216 35012
rect 24268 35000 24274 35012
rect 24854 35000 24860 35012
rect 24268 34972 24860 35000
rect 24268 34960 24274 34972
rect 24854 34960 24860 34972
rect 24912 34960 24918 35012
rect 28077 34935 28135 34941
rect 28077 34932 28089 34935
rect 19904 34904 28089 34932
rect 28077 34901 28089 34904
rect 28123 34901 28135 34935
rect 28077 34895 28135 34901
rect 1104 34842 28888 34864
rect 1104 34790 5614 34842
rect 5666 34790 5678 34842
rect 5730 34790 5742 34842
rect 5794 34790 5806 34842
rect 5858 34790 14878 34842
rect 14930 34790 14942 34842
rect 14994 34790 15006 34842
rect 15058 34790 15070 34842
rect 15122 34790 24142 34842
rect 24194 34790 24206 34842
rect 24258 34790 24270 34842
rect 24322 34790 24334 34842
rect 24386 34790 28888 34842
rect 1104 34768 28888 34790
rect 1673 34731 1731 34737
rect 1673 34697 1685 34731
rect 1719 34728 1731 34731
rect 2406 34728 2412 34740
rect 1719 34700 2412 34728
rect 1719 34697 1731 34700
rect 1673 34691 1731 34697
rect 1872 34533 1900 34700
rect 2406 34688 2412 34700
rect 2464 34688 2470 34740
rect 4982 34728 4988 34740
rect 4943 34700 4988 34728
rect 4982 34688 4988 34700
rect 5040 34688 5046 34740
rect 16114 34728 16120 34740
rect 5920 34700 16120 34728
rect 2590 34620 2596 34672
rect 2648 34660 2654 34672
rect 5920 34660 5948 34700
rect 16114 34688 16120 34700
rect 16172 34688 16178 34740
rect 16209 34731 16267 34737
rect 16209 34697 16221 34731
rect 16255 34728 16267 34731
rect 16942 34728 16948 34740
rect 16255 34700 16948 34728
rect 16255 34697 16267 34700
rect 16209 34691 16267 34697
rect 16942 34688 16948 34700
rect 17000 34688 17006 34740
rect 17313 34731 17371 34737
rect 17313 34697 17325 34731
rect 17359 34728 17371 34731
rect 18046 34728 18052 34740
rect 17359 34700 18052 34728
rect 17359 34697 17371 34700
rect 17313 34691 17371 34697
rect 18046 34688 18052 34700
rect 18104 34688 18110 34740
rect 18233 34731 18291 34737
rect 18233 34697 18245 34731
rect 18279 34728 18291 34731
rect 18598 34728 18604 34740
rect 18279 34700 18604 34728
rect 18279 34697 18291 34700
rect 18233 34691 18291 34697
rect 18598 34688 18604 34700
rect 18656 34688 18662 34740
rect 19702 34688 19708 34740
rect 19760 34728 19766 34740
rect 20346 34728 20352 34740
rect 19760 34700 20352 34728
rect 19760 34688 19766 34700
rect 20346 34688 20352 34700
rect 20404 34688 20410 34740
rect 22738 34688 22744 34740
rect 22796 34728 22802 34740
rect 22833 34731 22891 34737
rect 22833 34728 22845 34731
rect 22796 34700 22845 34728
rect 22796 34688 22802 34700
rect 22833 34697 22845 34700
rect 22879 34697 22891 34731
rect 22833 34691 22891 34697
rect 23845 34731 23903 34737
rect 23845 34697 23857 34731
rect 23891 34728 23903 34731
rect 24578 34728 24584 34740
rect 23891 34700 24584 34728
rect 23891 34697 23903 34700
rect 23845 34691 23903 34697
rect 24578 34688 24584 34700
rect 24636 34688 24642 34740
rect 25225 34731 25283 34737
rect 25225 34697 25237 34731
rect 25271 34728 25283 34731
rect 25958 34728 25964 34740
rect 25271 34700 25964 34728
rect 25271 34697 25283 34700
rect 25225 34691 25283 34697
rect 25958 34688 25964 34700
rect 26016 34688 26022 34740
rect 27338 34728 27344 34740
rect 27299 34700 27344 34728
rect 27338 34688 27344 34700
rect 27396 34688 27402 34740
rect 2648 34632 5948 34660
rect 2648 34620 2654 34632
rect 9398 34620 9404 34672
rect 9456 34660 9462 34672
rect 9456 34632 9536 34660
rect 9456 34620 9462 34632
rect 3970 34552 3976 34604
rect 4028 34592 4034 34604
rect 4028 34564 5212 34592
rect 4028 34552 4034 34564
rect 1857 34527 1915 34533
rect 1857 34493 1869 34527
rect 1903 34493 1915 34527
rect 2038 34524 2044 34536
rect 1999 34496 2044 34524
rect 1857 34487 1915 34493
rect 2038 34484 2044 34496
rect 2096 34484 2102 34536
rect 2774 34484 2780 34536
rect 2832 34524 2838 34536
rect 4522 34524 4528 34536
rect 2832 34496 2877 34524
rect 4483 34496 4528 34524
rect 2832 34484 2838 34496
rect 4522 34484 4528 34496
rect 4580 34484 4586 34536
rect 4706 34484 4712 34536
rect 4764 34524 4770 34536
rect 5184 34533 5212 34564
rect 5534 34552 5540 34604
rect 5592 34592 5598 34604
rect 5905 34595 5963 34601
rect 5905 34592 5917 34595
rect 5592 34564 5917 34592
rect 5592 34552 5598 34564
rect 5905 34561 5917 34564
rect 5951 34592 5963 34595
rect 6362 34592 6368 34604
rect 5951 34564 6368 34592
rect 5951 34561 5963 34564
rect 5905 34555 5963 34561
rect 6362 34552 6368 34564
rect 6420 34552 6426 34604
rect 6638 34552 6644 34604
rect 6696 34592 6702 34604
rect 7285 34595 7343 34601
rect 7285 34592 7297 34595
rect 6696 34564 7297 34592
rect 6696 34552 6702 34564
rect 7285 34561 7297 34564
rect 7331 34561 7343 34595
rect 7285 34555 7343 34561
rect 5169 34527 5227 34533
rect 4764 34496 5120 34524
rect 4764 34484 4770 34496
rect 2590 34456 2596 34468
rect 2551 34428 2596 34456
rect 2590 34416 2596 34428
rect 2648 34416 2654 34468
rect 4341 34459 4399 34465
rect 4341 34425 4353 34459
rect 4387 34456 4399 34459
rect 4430 34456 4436 34468
rect 4387 34428 4436 34456
rect 4387 34425 4399 34428
rect 4341 34419 4399 34425
rect 4430 34416 4436 34428
rect 4488 34416 4494 34468
rect 4982 34456 4988 34468
rect 4943 34428 4988 34456
rect 4982 34416 4988 34428
rect 5040 34416 5046 34468
rect 5092 34456 5120 34496
rect 5169 34493 5181 34527
rect 5215 34493 5227 34527
rect 5169 34487 5227 34493
rect 5261 34527 5319 34533
rect 5261 34493 5273 34527
rect 5307 34493 5319 34527
rect 5261 34487 5319 34493
rect 6181 34527 6239 34533
rect 6181 34493 6193 34527
rect 6227 34524 6239 34527
rect 9398 34524 9404 34536
rect 6227 34496 9404 34524
rect 6227 34493 6239 34496
rect 6181 34487 6239 34493
rect 5276 34456 5304 34487
rect 9398 34484 9404 34496
rect 9456 34484 9462 34536
rect 9508 34533 9536 34632
rect 10502 34620 10508 34672
rect 10560 34660 10566 34672
rect 11146 34660 11152 34672
rect 10560 34632 11152 34660
rect 10560 34620 10566 34632
rect 11146 34620 11152 34632
rect 11204 34620 11210 34672
rect 12161 34663 12219 34669
rect 12161 34629 12173 34663
rect 12207 34660 12219 34663
rect 12710 34660 12716 34672
rect 12207 34632 12716 34660
rect 12207 34629 12219 34632
rect 12161 34623 12219 34629
rect 12710 34620 12716 34632
rect 12768 34620 12774 34672
rect 13354 34620 13360 34672
rect 13412 34660 13418 34672
rect 13541 34663 13599 34669
rect 13541 34660 13553 34663
rect 13412 34632 13553 34660
rect 13412 34620 13418 34632
rect 13541 34629 13553 34632
rect 13587 34629 13599 34663
rect 13541 34623 13599 34629
rect 19610 34620 19616 34672
rect 19668 34660 19674 34672
rect 28169 34663 28227 34669
rect 28169 34660 28181 34663
rect 19668 34632 20024 34660
rect 19668 34620 19674 34632
rect 9769 34595 9827 34601
rect 9769 34561 9781 34595
rect 9815 34592 9827 34595
rect 10410 34592 10416 34604
rect 9815 34564 10416 34592
rect 9815 34561 9827 34564
rect 9769 34555 9827 34561
rect 10410 34552 10416 34564
rect 10468 34552 10474 34604
rect 12342 34592 12348 34604
rect 11808 34564 12348 34592
rect 9493 34527 9551 34533
rect 9493 34493 9505 34527
rect 9539 34524 9551 34527
rect 11514 34524 11520 34536
rect 9539 34496 11520 34524
rect 9539 34493 9551 34496
rect 9493 34487 9551 34493
rect 11514 34484 11520 34496
rect 11572 34484 11578 34536
rect 11808 34533 11836 34564
rect 12342 34552 12348 34564
rect 12400 34552 12406 34604
rect 13722 34552 13728 34604
rect 13780 34552 13786 34604
rect 13998 34552 14004 34604
rect 14056 34592 14062 34604
rect 15194 34592 15200 34604
rect 14056 34564 15200 34592
rect 14056 34552 14062 34564
rect 15194 34552 15200 34564
rect 15252 34592 15258 34604
rect 17218 34592 17224 34604
rect 15252 34564 15976 34592
rect 15252 34552 15258 34564
rect 11793 34527 11851 34533
rect 11793 34493 11805 34527
rect 11839 34493 11851 34527
rect 11793 34487 11851 34493
rect 11885 34527 11943 34533
rect 11885 34493 11897 34527
rect 11931 34493 11943 34527
rect 11885 34487 11943 34493
rect 11977 34527 12035 34533
rect 11977 34493 11989 34527
rect 12023 34524 12035 34527
rect 12802 34524 12808 34536
rect 12023 34496 12808 34524
rect 12023 34493 12035 34496
rect 11977 34487 12035 34493
rect 5092 34428 5304 34456
rect 10962 34416 10968 34468
rect 11020 34456 11026 34468
rect 11900 34456 11928 34487
rect 12802 34484 12808 34496
rect 12860 34484 12866 34536
rect 13538 34484 13544 34536
rect 13596 34524 13602 34536
rect 13740 34524 13768 34552
rect 15948 34533 15976 34564
rect 17052 34564 17224 34592
rect 13596 34496 13768 34524
rect 15841 34527 15899 34533
rect 13596 34484 13602 34496
rect 15841 34493 15853 34527
rect 15887 34493 15899 34527
rect 15841 34487 15899 34493
rect 15933 34527 15991 34533
rect 15933 34493 15945 34527
rect 15979 34493 15991 34527
rect 15933 34487 15991 34493
rect 11020 34428 11928 34456
rect 11020 34416 11026 34428
rect 13078 34416 13084 34468
rect 13136 34456 13142 34468
rect 13357 34459 13415 34465
rect 13357 34456 13369 34459
rect 13136 34428 13369 34456
rect 13136 34416 13142 34428
rect 13357 34425 13369 34428
rect 13403 34425 13415 34459
rect 13357 34419 13415 34425
rect 15856 34456 15884 34487
rect 16022 34484 16028 34536
rect 16080 34524 16086 34536
rect 17052 34533 17080 34564
rect 17218 34552 17224 34564
rect 17276 34552 17282 34604
rect 18230 34592 18236 34604
rect 17972 34564 18236 34592
rect 16945 34527 17003 34533
rect 16080 34496 16125 34524
rect 16080 34484 16086 34496
rect 16945 34493 16957 34527
rect 16991 34493 17003 34527
rect 16945 34487 17003 34493
rect 17037 34527 17095 34533
rect 17037 34493 17049 34527
rect 17083 34493 17095 34527
rect 17037 34487 17095 34493
rect 17129 34527 17187 34533
rect 17129 34493 17141 34527
rect 17175 34493 17187 34527
rect 17129 34487 17187 34493
rect 16482 34456 16488 34468
rect 15856 34428 16488 34456
rect 4890 34348 4896 34400
rect 4948 34388 4954 34400
rect 5258 34388 5264 34400
rect 4948 34360 5264 34388
rect 4948 34348 4954 34360
rect 5258 34348 5264 34360
rect 5316 34348 5322 34400
rect 10870 34388 10876 34400
rect 10831 34360 10876 34388
rect 10870 34348 10876 34360
rect 10928 34348 10934 34400
rect 11882 34348 11888 34400
rect 11940 34388 11946 34400
rect 13814 34388 13820 34400
rect 11940 34360 13820 34388
rect 11940 34348 11946 34360
rect 13814 34348 13820 34360
rect 13872 34348 13878 34400
rect 15856 34388 15884 34428
rect 16482 34416 16488 34428
rect 16540 34456 16546 34468
rect 16960 34456 16988 34487
rect 17144 34456 17172 34487
rect 17678 34484 17684 34536
rect 17736 34524 17742 34536
rect 17972 34533 18000 34564
rect 18230 34552 18236 34564
rect 18288 34552 18294 34604
rect 19886 34552 19892 34604
rect 19944 34552 19950 34604
rect 19996 34592 20024 34632
rect 22572 34632 28181 34660
rect 22572 34592 22600 34632
rect 28169 34629 28181 34632
rect 28215 34629 28227 34663
rect 28169 34623 28227 34629
rect 23382 34592 23388 34604
rect 19996 34564 20116 34592
rect 17865 34527 17923 34533
rect 17865 34524 17877 34527
rect 17736 34496 17877 34524
rect 17736 34484 17742 34496
rect 17865 34493 17877 34496
rect 17911 34493 17923 34527
rect 17865 34487 17923 34493
rect 17957 34527 18015 34533
rect 17957 34493 17969 34527
rect 18003 34493 18015 34527
rect 17957 34487 18015 34493
rect 18049 34527 18107 34533
rect 18049 34493 18061 34527
rect 18095 34524 18107 34527
rect 19150 34524 19156 34536
rect 18095 34496 19156 34524
rect 18095 34493 18107 34496
rect 18049 34487 18107 34493
rect 18064 34456 18092 34487
rect 19150 34484 19156 34496
rect 19208 34484 19214 34536
rect 19904 34524 19932 34552
rect 19981 34527 20039 34533
rect 19981 34524 19993 34527
rect 19904 34496 19993 34524
rect 19981 34493 19993 34496
rect 20027 34493 20039 34527
rect 20088 34524 20116 34564
rect 21008 34564 22600 34592
rect 22756 34564 23388 34592
rect 20237 34527 20295 34533
rect 20237 34524 20249 34527
rect 20088 34496 20249 34524
rect 19981 34487 20039 34493
rect 20237 34493 20249 34496
rect 20283 34493 20295 34527
rect 20237 34487 20295 34493
rect 21008 34456 21036 34564
rect 22462 34524 22468 34536
rect 22423 34496 22468 34524
rect 22462 34484 22468 34496
rect 22520 34484 22526 34536
rect 22557 34527 22615 34533
rect 22557 34493 22569 34527
rect 22603 34493 22615 34527
rect 22557 34487 22615 34493
rect 22661 34527 22719 34533
rect 22661 34493 22673 34527
rect 22707 34524 22719 34527
rect 22756 34524 22784 34564
rect 23382 34552 23388 34564
rect 23440 34592 23446 34604
rect 23440 34564 23704 34592
rect 23440 34552 23446 34564
rect 23676 34533 23704 34564
rect 23842 34552 23848 34604
rect 23900 34592 23906 34604
rect 25222 34592 25228 34604
rect 23900 34564 25228 34592
rect 23900 34552 23906 34564
rect 25222 34552 25228 34564
rect 25280 34592 25286 34604
rect 26602 34592 26608 34604
rect 25280 34564 26608 34592
rect 25280 34552 25286 34564
rect 26602 34552 26608 34564
rect 26660 34552 26666 34604
rect 23477 34527 23535 34533
rect 23477 34524 23489 34527
rect 22707 34496 22784 34524
rect 22848 34496 23489 34524
rect 22707 34493 22719 34496
rect 22661 34487 22719 34493
rect 16540 34428 16988 34456
rect 17052 34428 18092 34456
rect 19306 34428 21036 34456
rect 16540 34416 16546 34428
rect 16022 34388 16028 34400
rect 15856 34360 16028 34388
rect 16022 34348 16028 34360
rect 16080 34348 16086 34400
rect 16206 34348 16212 34400
rect 16264 34388 16270 34400
rect 17052 34388 17080 34428
rect 17880 34400 17908 34428
rect 16264 34360 17080 34388
rect 16264 34348 16270 34360
rect 17862 34348 17868 34400
rect 17920 34348 17926 34400
rect 17954 34348 17960 34400
rect 18012 34388 18018 34400
rect 19306 34388 19334 34428
rect 22186 34416 22192 34468
rect 22244 34456 22250 34468
rect 22572 34456 22600 34487
rect 22244 34428 22600 34456
rect 22244 34416 22250 34428
rect 18012 34360 19334 34388
rect 18012 34348 18018 34360
rect 20346 34348 20352 34400
rect 20404 34388 20410 34400
rect 21361 34391 21419 34397
rect 21361 34388 21373 34391
rect 20404 34360 21373 34388
rect 20404 34348 20410 34360
rect 21361 34357 21373 34360
rect 21407 34357 21419 34391
rect 21361 34351 21419 34357
rect 22462 34348 22468 34400
rect 22520 34388 22526 34400
rect 22848 34388 22876 34496
rect 23477 34493 23489 34496
rect 23523 34493 23535 34527
rect 23477 34487 23535 34493
rect 23569 34527 23627 34533
rect 23569 34493 23581 34527
rect 23615 34493 23627 34527
rect 23569 34487 23627 34493
rect 23661 34527 23719 34533
rect 23661 34493 23673 34527
rect 23707 34493 23719 34527
rect 25406 34524 25412 34536
rect 25367 34496 25412 34524
rect 23661 34487 23719 34493
rect 23584 34400 23612 34487
rect 25406 34484 25412 34496
rect 25464 34484 25470 34536
rect 26050 34524 26056 34536
rect 26011 34496 26056 34524
rect 26050 34484 26056 34496
rect 26108 34484 26114 34536
rect 26694 34524 26700 34536
rect 26655 34496 26700 34524
rect 26694 34484 26700 34496
rect 26752 34484 26758 34536
rect 27249 34459 27307 34465
rect 27249 34456 27261 34459
rect 25884 34428 27261 34456
rect 22520 34360 22876 34388
rect 22520 34348 22526 34360
rect 23566 34348 23572 34400
rect 23624 34348 23630 34400
rect 25884 34397 25912 34428
rect 27249 34425 27261 34428
rect 27295 34425 27307 34459
rect 27249 34419 27307 34425
rect 27798 34416 27804 34468
rect 27856 34456 27862 34468
rect 27985 34459 28043 34465
rect 27985 34456 27997 34459
rect 27856 34428 27997 34456
rect 27856 34416 27862 34428
rect 27985 34425 27997 34428
rect 28031 34425 28043 34459
rect 27985 34419 28043 34425
rect 25869 34391 25927 34397
rect 25869 34357 25881 34391
rect 25915 34357 25927 34391
rect 26510 34388 26516 34400
rect 26471 34360 26516 34388
rect 25869 34351 25927 34357
rect 26510 34348 26516 34360
rect 26568 34348 26574 34400
rect 1104 34298 28888 34320
rect 1104 34246 10246 34298
rect 10298 34246 10310 34298
rect 10362 34246 10374 34298
rect 10426 34246 10438 34298
rect 10490 34246 19510 34298
rect 19562 34246 19574 34298
rect 19626 34246 19638 34298
rect 19690 34246 19702 34298
rect 19754 34246 28888 34298
rect 1104 34224 28888 34246
rect 3878 34184 3884 34196
rect 3791 34156 3884 34184
rect 3878 34144 3884 34156
rect 3936 34184 3942 34196
rect 4890 34184 4896 34196
rect 3936 34156 4896 34184
rect 3936 34144 3942 34156
rect 4890 34144 4896 34156
rect 4948 34144 4954 34196
rect 4982 34144 4988 34196
rect 5040 34184 5046 34196
rect 5261 34187 5319 34193
rect 5261 34184 5273 34187
rect 5040 34156 5273 34184
rect 5040 34144 5046 34156
rect 5261 34153 5273 34156
rect 5307 34153 5319 34187
rect 5261 34147 5319 34153
rect 7285 34187 7343 34193
rect 7285 34153 7297 34187
rect 7331 34184 7343 34187
rect 11054 34184 11060 34196
rect 7331 34156 8616 34184
rect 11015 34156 11060 34184
rect 7331 34153 7343 34156
rect 7285 34147 7343 34153
rect 4525 34119 4583 34125
rect 4525 34085 4537 34119
rect 4571 34116 4583 34119
rect 8588 34116 8616 34156
rect 11054 34144 11060 34156
rect 11112 34144 11118 34196
rect 24673 34187 24731 34193
rect 11164 34156 22094 34184
rect 11164 34116 11192 34156
rect 12805 34119 12863 34125
rect 12805 34116 12817 34119
rect 4571 34088 8524 34116
rect 8588 34088 11192 34116
rect 12406 34088 12817 34116
rect 4571 34085 4583 34088
rect 4525 34079 4583 34085
rect 1857 34051 1915 34057
rect 1857 34017 1869 34051
rect 1903 34017 1915 34051
rect 2038 34048 2044 34060
rect 1999 34020 2044 34048
rect 1857 34011 1915 34017
rect 1872 33980 1900 34011
rect 2038 34008 2044 34020
rect 2096 34008 2102 34060
rect 2406 34008 2412 34060
rect 2464 34048 2470 34060
rect 2593 34051 2651 34057
rect 2593 34048 2605 34051
rect 2464 34020 2605 34048
rect 2464 34008 2470 34020
rect 2593 34017 2605 34020
rect 2639 34017 2651 34051
rect 2593 34011 2651 34017
rect 3789 34051 3847 34057
rect 3789 34017 3801 34051
rect 3835 34048 3847 34051
rect 4430 34048 4436 34060
rect 3835 34020 4436 34048
rect 3835 34017 3847 34020
rect 3789 34011 3847 34017
rect 4430 34008 4436 34020
rect 4488 34008 4494 34060
rect 5166 34048 5172 34060
rect 5127 34020 5172 34048
rect 5166 34008 5172 34020
rect 5224 34008 5230 34060
rect 5258 34008 5264 34060
rect 5316 34048 5322 34060
rect 7650 34057 7656 34060
rect 5353 34051 5411 34057
rect 5353 34048 5365 34051
rect 5316 34020 5365 34048
rect 5316 34008 5322 34020
rect 5353 34017 5365 34020
rect 5399 34017 5411 34051
rect 5353 34011 5411 34017
rect 7644 34011 7656 34057
rect 7708 34048 7714 34060
rect 7708 34020 7744 34048
rect 7650 34008 7656 34011
rect 7708 34008 7714 34020
rect 7285 33983 7343 33989
rect 7285 33980 7297 33983
rect 1872 33952 7297 33980
rect 7285 33949 7297 33952
rect 7331 33949 7343 33983
rect 7285 33943 7343 33949
rect 7377 33983 7435 33989
rect 7377 33949 7389 33983
rect 7423 33949 7435 33983
rect 7377 33943 7435 33949
rect 2777 33915 2835 33921
rect 2777 33881 2789 33915
rect 2823 33912 2835 33915
rect 3050 33912 3056 33924
rect 2823 33884 3056 33912
rect 2823 33881 2835 33884
rect 2777 33875 2835 33881
rect 3050 33872 3056 33884
rect 3108 33872 3114 33924
rect 6362 33872 6368 33924
rect 6420 33912 6426 33924
rect 7392 33912 7420 33943
rect 6420 33884 7420 33912
rect 8496 33912 8524 34088
rect 10962 34048 10968 34060
rect 10923 34020 10968 34048
rect 10962 34008 10968 34020
rect 11020 34008 11026 34060
rect 11146 34048 11152 34060
rect 11107 34020 11152 34048
rect 11146 34008 11152 34020
rect 11204 34048 11210 34060
rect 12406 34048 12434 34088
rect 12805 34085 12817 34088
rect 12851 34116 12863 34119
rect 13446 34116 13452 34128
rect 12851 34088 13452 34116
rect 12851 34085 12863 34088
rect 12805 34079 12863 34085
rect 13446 34076 13452 34088
rect 13504 34076 13510 34128
rect 14182 34076 14188 34128
rect 14240 34116 14246 34128
rect 15105 34119 15163 34125
rect 14240 34088 14964 34116
rect 14240 34076 14246 34088
rect 11204 34020 12434 34048
rect 12621 34051 12679 34057
rect 11204 34008 11210 34020
rect 12621 34017 12633 34051
rect 12667 34048 12679 34051
rect 13078 34048 13084 34060
rect 12667 34020 13084 34048
rect 12667 34017 12679 34020
rect 12621 34011 12679 34017
rect 12636 33980 12664 34011
rect 13078 34008 13084 34020
rect 13136 34048 13142 34060
rect 13357 34051 13415 34057
rect 13357 34048 13369 34051
rect 13136 34020 13369 34048
rect 13136 34008 13142 34020
rect 13357 34017 13369 34020
rect 13403 34017 13415 34051
rect 13998 34048 14004 34060
rect 13959 34020 14004 34048
rect 13357 34011 13415 34017
rect 13998 34008 14004 34020
rect 14056 34008 14062 34060
rect 14274 34008 14280 34060
rect 14332 34048 14338 34060
rect 14936 34057 14964 34088
rect 15105 34085 15117 34119
rect 15151 34116 15163 34119
rect 15838 34116 15844 34128
rect 15151 34088 15844 34116
rect 15151 34085 15163 34088
rect 15105 34079 15163 34085
rect 15838 34076 15844 34088
rect 15896 34076 15902 34128
rect 16393 34119 16451 34125
rect 16393 34085 16405 34119
rect 16439 34116 16451 34119
rect 17034 34116 17040 34128
rect 16439 34088 17040 34116
rect 16439 34085 16451 34088
rect 16393 34079 16451 34085
rect 17034 34076 17040 34088
rect 17092 34076 17098 34128
rect 18046 34116 18052 34128
rect 18007 34088 18052 34116
rect 18046 34076 18052 34088
rect 18104 34076 18110 34128
rect 18690 34076 18696 34128
rect 18748 34116 18754 34128
rect 19245 34119 19303 34125
rect 18748 34088 19012 34116
rect 18748 34076 18754 34088
rect 14737 34051 14795 34057
rect 14737 34048 14749 34051
rect 14332 34020 14749 34048
rect 14332 34008 14338 34020
rect 14737 34017 14749 34020
rect 14783 34017 14795 34051
rect 14737 34011 14795 34017
rect 14829 34051 14887 34057
rect 14829 34017 14841 34051
rect 14875 34017 14887 34051
rect 14829 34011 14887 34017
rect 14921 34051 14979 34057
rect 14921 34017 14933 34051
rect 14967 34048 14979 34051
rect 15654 34048 15660 34060
rect 14967 34020 15660 34048
rect 14967 34017 14979 34020
rect 14921 34011 14979 34017
rect 12802 33980 12808 33992
rect 12636 33952 12808 33980
rect 12802 33940 12808 33952
rect 12860 33940 12866 33992
rect 13446 33940 13452 33992
rect 13504 33980 13510 33992
rect 13541 33983 13599 33989
rect 13541 33980 13553 33983
rect 13504 33952 13553 33980
rect 13504 33940 13510 33952
rect 13541 33949 13553 33952
rect 13587 33980 13599 33983
rect 13906 33980 13912 33992
rect 13587 33952 13912 33980
rect 13587 33949 13599 33952
rect 13541 33943 13599 33949
rect 13906 33940 13912 33952
rect 13964 33940 13970 33992
rect 14844 33980 14872 34011
rect 15654 34008 15660 34020
rect 15712 34008 15718 34060
rect 16022 34048 16028 34060
rect 15983 34020 16028 34048
rect 16022 34008 16028 34020
rect 16080 34008 16086 34060
rect 16117 34051 16175 34057
rect 16117 34017 16129 34051
rect 16163 34017 16175 34051
rect 16117 34011 16175 34017
rect 15562 33980 15568 33992
rect 14844 33952 15568 33980
rect 15562 33940 15568 33952
rect 15620 33980 15626 33992
rect 16132 33980 16160 34011
rect 16206 34008 16212 34060
rect 16264 34048 16270 34060
rect 16264 34020 16309 34048
rect 16264 34008 16270 34020
rect 16482 34008 16488 34060
rect 16540 34048 16546 34060
rect 17678 34048 17684 34060
rect 16540 34020 17684 34048
rect 16540 34008 16546 34020
rect 17678 34008 17684 34020
rect 17736 34008 17742 34060
rect 17773 34051 17831 34057
rect 17773 34017 17785 34051
rect 17819 34017 17831 34051
rect 17773 34011 17831 34017
rect 15620 33952 16160 33980
rect 15620 33940 15626 33952
rect 17310 33940 17316 33992
rect 17368 33980 17374 33992
rect 17788 33980 17816 34011
rect 17862 34008 17868 34060
rect 17920 34048 17926 34060
rect 17920 34020 17965 34048
rect 17920 34008 17926 34020
rect 18782 34008 18788 34060
rect 18840 34048 18846 34060
rect 18984 34057 19012 34088
rect 19245 34085 19257 34119
rect 19291 34116 19303 34119
rect 20438 34116 20444 34128
rect 19291 34088 20444 34116
rect 19291 34085 19303 34088
rect 19245 34079 19303 34085
rect 20438 34076 20444 34088
rect 20496 34076 20502 34128
rect 21269 34119 21327 34125
rect 21269 34085 21281 34119
rect 21315 34116 21327 34119
rect 21542 34116 21548 34128
rect 21315 34088 21548 34116
rect 21315 34085 21327 34088
rect 21269 34079 21327 34085
rect 21542 34076 21548 34088
rect 21600 34076 21606 34128
rect 22066 34116 22094 34156
rect 24673 34153 24685 34187
rect 24719 34184 24731 34187
rect 25774 34184 25780 34196
rect 24719 34156 25780 34184
rect 24719 34153 24731 34156
rect 24673 34147 24731 34153
rect 25774 34144 25780 34156
rect 25832 34144 25838 34196
rect 25961 34187 26019 34193
rect 25961 34153 25973 34187
rect 26007 34184 26019 34187
rect 26007 34156 27936 34184
rect 26007 34153 26019 34156
rect 25961 34147 26019 34153
rect 22066 34088 26280 34116
rect 18877 34051 18935 34057
rect 18877 34048 18889 34051
rect 18840 34020 18889 34048
rect 18840 34008 18846 34020
rect 18877 34017 18889 34020
rect 18923 34017 18935 34051
rect 18877 34011 18935 34017
rect 18969 34051 19027 34057
rect 18969 34017 18981 34051
rect 19015 34017 19027 34051
rect 18969 34011 19027 34017
rect 19061 34051 19119 34057
rect 19061 34017 19073 34051
rect 19107 34048 19119 34051
rect 19150 34048 19156 34060
rect 19107 34020 19156 34048
rect 19107 34017 19119 34020
rect 19061 34011 19119 34017
rect 17368 33952 17816 33980
rect 18892 33980 18920 34011
rect 19150 34008 19156 34020
rect 19208 34008 19214 34060
rect 20865 34051 20923 34057
rect 20865 34017 20877 34051
rect 20911 34017 20923 34051
rect 20990 34048 20996 34060
rect 20951 34020 20996 34048
rect 20865 34011 20923 34017
rect 20880 33980 20908 34011
rect 20990 34008 20996 34020
rect 21048 34008 21054 34060
rect 21082 34008 21088 34060
rect 21140 34048 21146 34060
rect 23382 34048 23388 34060
rect 21140 34020 23388 34048
rect 21140 34008 21146 34020
rect 23382 34008 23388 34020
rect 23440 34008 23446 34060
rect 24854 34048 24860 34060
rect 24815 34020 24860 34048
rect 24854 34008 24860 34020
rect 24912 34008 24918 34060
rect 25498 34048 25504 34060
rect 25459 34020 25504 34048
rect 25498 34008 25504 34020
rect 25556 34008 25562 34060
rect 26142 34048 26148 34060
rect 26103 34020 26148 34048
rect 26142 34008 26148 34020
rect 26200 34008 26206 34060
rect 26252 34048 26280 34088
rect 26510 34076 26516 34128
rect 26568 34116 26574 34128
rect 27908 34125 27936 34156
rect 26697 34119 26755 34125
rect 26697 34116 26709 34119
rect 26568 34088 26709 34116
rect 26568 34076 26574 34088
rect 26697 34085 26709 34088
rect 26743 34085 26755 34119
rect 26697 34079 26755 34085
rect 27893 34119 27951 34125
rect 27893 34085 27905 34119
rect 27939 34085 27951 34119
rect 27893 34079 27951 34085
rect 28077 34051 28135 34057
rect 28077 34048 28089 34051
rect 26252 34020 28089 34048
rect 28077 34017 28089 34020
rect 28123 34017 28135 34051
rect 28077 34011 28135 34017
rect 22462 33980 22468 33992
rect 18892 33952 22468 33980
rect 17368 33940 17374 33952
rect 22462 33940 22468 33952
rect 22520 33940 22526 33992
rect 23106 33940 23112 33992
rect 23164 33980 23170 33992
rect 23290 33980 23296 33992
rect 23164 33952 23296 33980
rect 23164 33940 23170 33952
rect 23290 33940 23296 33952
rect 23348 33940 23354 33992
rect 24486 33940 24492 33992
rect 24544 33980 24550 33992
rect 24670 33980 24676 33992
rect 24544 33952 24676 33980
rect 24544 33940 24550 33952
rect 24670 33940 24676 33952
rect 24728 33940 24734 33992
rect 27246 33912 27252 33924
rect 8496 33884 27252 33912
rect 6420 33872 6426 33884
rect 4154 33804 4160 33856
rect 4212 33844 4218 33856
rect 4617 33847 4675 33853
rect 4617 33844 4629 33847
rect 4212 33816 4629 33844
rect 4212 33804 4218 33816
rect 4617 33813 4629 33816
rect 4663 33813 4675 33847
rect 7392 33844 7420 33884
rect 27246 33872 27252 33884
rect 27304 33872 27310 33924
rect 7742 33844 7748 33856
rect 7392 33816 7748 33844
rect 4617 33807 4675 33813
rect 7742 33804 7748 33816
rect 7800 33804 7806 33856
rect 8757 33847 8815 33853
rect 8757 33813 8769 33847
rect 8803 33844 8815 33847
rect 9490 33844 9496 33856
rect 8803 33816 9496 33844
rect 8803 33813 8815 33816
rect 8757 33807 8815 33813
rect 9490 33804 9496 33816
rect 9548 33804 9554 33856
rect 13538 33804 13544 33856
rect 13596 33844 13602 33856
rect 14185 33847 14243 33853
rect 14185 33844 14197 33847
rect 13596 33816 14197 33844
rect 13596 33804 13602 33816
rect 14185 33813 14197 33816
rect 14231 33813 14243 33847
rect 14185 33807 14243 33813
rect 15470 33804 15476 33856
rect 15528 33844 15534 33856
rect 15838 33844 15844 33856
rect 15528 33816 15844 33844
rect 15528 33804 15534 33816
rect 15838 33804 15844 33816
rect 15896 33804 15902 33856
rect 17954 33804 17960 33856
rect 18012 33844 18018 33856
rect 18414 33844 18420 33856
rect 18012 33816 18420 33844
rect 18012 33804 18018 33816
rect 18414 33804 18420 33816
rect 18472 33804 18478 33856
rect 22002 33804 22008 33856
rect 22060 33844 22066 33856
rect 24486 33844 24492 33856
rect 22060 33816 24492 33844
rect 22060 33804 22066 33816
rect 24486 33804 24492 33816
rect 24544 33804 24550 33856
rect 25317 33847 25375 33853
rect 25317 33813 25329 33847
rect 25363 33844 25375 33847
rect 26510 33844 26516 33856
rect 25363 33816 26516 33844
rect 25363 33813 25375 33816
rect 25317 33807 25375 33813
rect 26510 33804 26516 33816
rect 26568 33804 26574 33856
rect 26786 33844 26792 33856
rect 26747 33816 26792 33844
rect 26786 33804 26792 33816
rect 26844 33804 26850 33856
rect 1104 33754 28888 33776
rect 1104 33702 5614 33754
rect 5666 33702 5678 33754
rect 5730 33702 5742 33754
rect 5794 33702 5806 33754
rect 5858 33702 14878 33754
rect 14930 33702 14942 33754
rect 14994 33702 15006 33754
rect 15058 33702 15070 33754
rect 15122 33702 24142 33754
rect 24194 33702 24206 33754
rect 24258 33702 24270 33754
rect 24322 33702 24334 33754
rect 24386 33702 28888 33754
rect 1104 33680 28888 33702
rect 1394 33600 1400 33652
rect 1452 33640 1458 33652
rect 1581 33643 1639 33649
rect 1581 33640 1593 33643
rect 1452 33612 1593 33640
rect 1452 33600 1458 33612
rect 1581 33609 1593 33612
rect 1627 33609 1639 33643
rect 1581 33603 1639 33609
rect 3142 33600 3148 33652
rect 3200 33640 3206 33652
rect 5077 33643 5135 33649
rect 5077 33640 5089 33643
rect 3200 33612 5089 33640
rect 3200 33600 3206 33612
rect 5077 33609 5089 33612
rect 5123 33609 5135 33643
rect 5077 33603 5135 33609
rect 7650 33600 7656 33652
rect 7708 33640 7714 33652
rect 7837 33643 7895 33649
rect 7837 33640 7849 33643
rect 7708 33612 7849 33640
rect 7708 33600 7714 33612
rect 7837 33609 7849 33612
rect 7883 33609 7895 33643
rect 26786 33640 26792 33652
rect 7837 33603 7895 33609
rect 7944 33612 26792 33640
rect 4798 33532 4804 33584
rect 4856 33572 4862 33584
rect 5258 33572 5264 33584
rect 4856 33544 5264 33572
rect 4856 33532 4862 33544
rect 5258 33532 5264 33544
rect 5316 33572 5322 33584
rect 5721 33575 5779 33581
rect 5721 33572 5733 33575
rect 5316 33544 5733 33572
rect 5316 33532 5322 33544
rect 5721 33541 5733 33544
rect 5767 33541 5779 33575
rect 5721 33535 5779 33541
rect 7944 33504 7972 33612
rect 26786 33600 26792 33612
rect 26844 33600 26850 33652
rect 27246 33640 27252 33652
rect 27207 33612 27252 33640
rect 27246 33600 27252 33612
rect 27304 33600 27310 33652
rect 27982 33640 27988 33652
rect 27943 33612 27988 33640
rect 27982 33600 27988 33612
rect 28040 33600 28046 33652
rect 23842 33572 23848 33584
rect 1504 33476 7972 33504
rect 8128 33544 23848 33572
rect 1504 33445 1532 33476
rect 1489 33439 1547 33445
rect 1489 33405 1501 33439
rect 1535 33405 1547 33439
rect 1489 33399 1547 33405
rect 2409 33439 2467 33445
rect 2409 33405 2421 33439
rect 2455 33436 2467 33439
rect 2498 33436 2504 33448
rect 2455 33408 2504 33436
rect 2455 33405 2467 33408
rect 2409 33399 2467 33405
rect 2498 33396 2504 33408
rect 2556 33396 2562 33448
rect 2682 33436 2688 33448
rect 2643 33408 2688 33436
rect 2682 33396 2688 33408
rect 2740 33396 2746 33448
rect 3142 33436 3148 33448
rect 3103 33408 3148 33436
rect 3142 33396 3148 33408
rect 3200 33396 3206 33448
rect 3329 33439 3387 33445
rect 3329 33405 3341 33439
rect 3375 33436 3387 33439
rect 3418 33436 3424 33448
rect 3375 33408 3424 33436
rect 3375 33405 3387 33408
rect 3329 33399 3387 33405
rect 3418 33396 3424 33408
rect 3476 33436 3482 33448
rect 4985 33439 5043 33445
rect 4985 33436 4997 33439
rect 3476 33408 4997 33436
rect 3476 33396 3482 33408
rect 4985 33405 4997 33408
rect 5031 33405 5043 33439
rect 4985 33399 5043 33405
rect 5166 33396 5172 33448
rect 5224 33436 5230 33448
rect 5629 33439 5687 33445
rect 5629 33436 5641 33439
rect 5224 33408 5641 33436
rect 5224 33396 5230 33408
rect 5629 33405 5641 33408
rect 5675 33436 5687 33439
rect 5902 33436 5908 33448
rect 5675 33408 5908 33436
rect 5675 33405 5687 33408
rect 5629 33399 5687 33405
rect 5902 33396 5908 33408
rect 5960 33436 5966 33448
rect 6638 33436 6644 33448
rect 5960 33408 6644 33436
rect 5960 33396 5966 33408
rect 6638 33396 6644 33408
rect 6696 33396 6702 33448
rect 4341 33371 4399 33377
rect 4341 33337 4353 33371
rect 4387 33368 4399 33371
rect 8128 33368 8156 33544
rect 23842 33532 23848 33544
rect 23900 33532 23906 33584
rect 24394 33532 24400 33584
rect 24452 33572 24458 33584
rect 24670 33572 24676 33584
rect 24452 33544 24676 33572
rect 24452 33532 24458 33544
rect 24670 33532 24676 33544
rect 24728 33532 24734 33584
rect 25774 33532 25780 33584
rect 25832 33572 25838 33584
rect 25832 33544 27936 33572
rect 25832 33532 25838 33544
rect 8481 33507 8539 33513
rect 8481 33473 8493 33507
rect 8527 33504 8539 33507
rect 9122 33504 9128 33516
rect 8527 33476 9128 33504
rect 8527 33473 8539 33476
rect 8481 33467 8539 33473
rect 9122 33464 9128 33476
rect 9180 33464 9186 33516
rect 12802 33504 12808 33516
rect 12763 33476 12808 33504
rect 12802 33464 12808 33476
rect 12860 33464 12866 33516
rect 13725 33507 13783 33513
rect 13725 33473 13737 33507
rect 13771 33504 13783 33507
rect 14182 33504 14188 33516
rect 13771 33476 14188 33504
rect 13771 33473 13783 33476
rect 13725 33467 13783 33473
rect 14182 33464 14188 33476
rect 14240 33464 14246 33516
rect 14550 33464 14556 33516
rect 14608 33504 14614 33516
rect 14826 33504 14832 33516
rect 14608 33476 14832 33504
rect 14608 33464 14614 33476
rect 14826 33464 14832 33476
rect 14884 33464 14890 33516
rect 15764 33476 16804 33504
rect 9677 33439 9735 33445
rect 9677 33405 9689 33439
rect 9723 33436 9735 33439
rect 9950 33436 9956 33448
rect 9723 33408 9956 33436
rect 9723 33405 9735 33408
rect 9677 33399 9735 33405
rect 9950 33396 9956 33408
rect 10008 33436 10014 33448
rect 10870 33436 10876 33448
rect 10008 33408 10876 33436
rect 10008 33396 10014 33408
rect 10870 33396 10876 33408
rect 10928 33396 10934 33448
rect 12713 33439 12771 33445
rect 12713 33405 12725 33439
rect 12759 33405 12771 33439
rect 12713 33399 12771 33405
rect 12897 33439 12955 33445
rect 12897 33405 12909 33439
rect 12943 33436 12955 33439
rect 13078 33436 13084 33448
rect 12943 33408 13084 33436
rect 12943 33405 12955 33408
rect 12897 33399 12955 33405
rect 4387 33340 8156 33368
rect 8205 33371 8263 33377
rect 4387 33337 4399 33340
rect 4341 33331 4399 33337
rect 8205 33337 8217 33371
rect 8251 33368 8263 33371
rect 9490 33368 9496 33380
rect 8251 33340 9496 33368
rect 8251 33337 8263 33340
rect 8205 33331 8263 33337
rect 9490 33328 9496 33340
rect 9548 33328 9554 33380
rect 3602 33260 3608 33312
rect 3660 33300 3666 33312
rect 4433 33303 4491 33309
rect 4433 33300 4445 33303
rect 3660 33272 4445 33300
rect 3660 33260 3666 33272
rect 4433 33269 4445 33272
rect 4479 33269 4491 33303
rect 4433 33263 4491 33269
rect 5166 33260 5172 33312
rect 5224 33300 5230 33312
rect 5442 33300 5448 33312
rect 5224 33272 5448 33300
rect 5224 33260 5230 33272
rect 5442 33260 5448 33272
rect 5500 33260 5506 33312
rect 8110 33260 8116 33312
rect 8168 33300 8174 33312
rect 8297 33303 8355 33309
rect 8297 33300 8309 33303
rect 8168 33272 8309 33300
rect 8168 33260 8174 33272
rect 8297 33269 8309 33272
rect 8343 33269 8355 33303
rect 8297 33263 8355 33269
rect 9861 33303 9919 33309
rect 9861 33269 9873 33303
rect 9907 33300 9919 33303
rect 11054 33300 11060 33312
rect 9907 33272 11060 33300
rect 9907 33269 9919 33272
rect 9861 33263 9919 33269
rect 11054 33260 11060 33272
rect 11112 33300 11118 33312
rect 11330 33300 11336 33312
rect 11112 33272 11336 33300
rect 11112 33260 11118 33272
rect 11330 33260 11336 33272
rect 11388 33260 11394 33312
rect 12728 33300 12756 33399
rect 13078 33396 13084 33408
rect 13136 33396 13142 33448
rect 13354 33436 13360 33448
rect 13315 33408 13360 33436
rect 13354 33396 13360 33408
rect 13412 33396 13418 33448
rect 13541 33439 13599 33445
rect 13541 33405 13553 33439
rect 13587 33405 13599 33439
rect 13541 33399 13599 33405
rect 12802 33328 12808 33380
rect 12860 33368 12866 33380
rect 13556 33368 13584 33399
rect 13906 33396 13912 33448
rect 13964 33436 13970 33448
rect 15010 33436 15016 33448
rect 13964 33408 15016 33436
rect 13964 33396 13970 33408
rect 15010 33396 15016 33408
rect 15068 33396 15074 33448
rect 15764 33368 15792 33476
rect 16776 33445 16804 33476
rect 20714 33464 20720 33516
rect 20772 33504 20778 33516
rect 20772 33476 24072 33504
rect 20772 33464 20778 33476
rect 16025 33439 16083 33445
rect 16025 33405 16037 33439
rect 16071 33405 16083 33439
rect 16025 33399 16083 33405
rect 16761 33439 16819 33445
rect 16761 33405 16773 33439
rect 16807 33436 16819 33439
rect 16942 33436 16948 33448
rect 16807 33408 16948 33436
rect 16807 33405 16819 33408
rect 16761 33399 16819 33405
rect 12860 33340 13584 33368
rect 14016 33340 15792 33368
rect 12860 33328 12866 33340
rect 14016 33312 14044 33340
rect 13998 33300 14004 33312
rect 12728 33272 14004 33300
rect 13998 33260 14004 33272
rect 14056 33260 14062 33312
rect 15197 33303 15255 33309
rect 15197 33269 15209 33303
rect 15243 33300 15255 33303
rect 15286 33300 15292 33312
rect 15243 33272 15292 33300
rect 15243 33269 15255 33272
rect 15197 33263 15255 33269
rect 15286 33260 15292 33272
rect 15344 33300 15350 33312
rect 16040 33300 16068 33399
rect 16942 33396 16948 33408
rect 17000 33436 17006 33448
rect 18141 33439 18199 33445
rect 18141 33436 18153 33439
rect 17000 33408 18153 33436
rect 17000 33396 17006 33408
rect 18141 33405 18153 33408
rect 18187 33405 18199 33439
rect 18141 33399 18199 33405
rect 21174 33396 21180 33448
rect 21232 33436 21238 33448
rect 21453 33439 21511 33445
rect 21453 33436 21465 33439
rect 21232 33408 21465 33436
rect 21232 33396 21238 33408
rect 21453 33405 21465 33408
rect 21499 33405 21511 33439
rect 21453 33399 21511 33405
rect 21542 33396 21548 33448
rect 21600 33436 21606 33448
rect 21836 33445 21864 33476
rect 21729 33439 21787 33445
rect 21729 33436 21741 33439
rect 21600 33408 21741 33436
rect 21600 33396 21606 33408
rect 21729 33405 21741 33408
rect 21775 33405 21787 33439
rect 21729 33399 21787 33405
rect 21821 33439 21879 33445
rect 21821 33405 21833 33439
rect 21867 33405 21879 33439
rect 23658 33436 23664 33448
rect 23619 33408 23664 33436
rect 21821 33399 21879 33405
rect 23658 33396 23664 33408
rect 23716 33396 23722 33448
rect 24044 33445 24072 33476
rect 24486 33464 24492 33516
rect 24544 33504 24550 33516
rect 25593 33507 25651 33513
rect 25593 33504 25605 33507
rect 24544 33476 25605 33504
rect 24544 33464 24550 33476
rect 25593 33473 25605 33476
rect 25639 33473 25651 33507
rect 25593 33467 25651 33473
rect 25961 33507 26019 33513
rect 25961 33473 25973 33507
rect 26007 33504 26019 33507
rect 26326 33504 26332 33516
rect 26007 33476 26332 33504
rect 26007 33473 26019 33476
rect 25961 33467 26019 33473
rect 26326 33464 26332 33476
rect 26384 33464 26390 33516
rect 24029 33439 24087 33445
rect 24029 33405 24041 33439
rect 24075 33436 24087 33439
rect 24302 33436 24308 33448
rect 24075 33408 24308 33436
rect 24075 33405 24087 33408
rect 24029 33399 24087 33405
rect 24302 33396 24308 33408
rect 24360 33396 24366 33448
rect 25777 33439 25835 33445
rect 25777 33405 25789 33439
rect 25823 33405 25835 33439
rect 25777 33399 25835 33405
rect 25869 33439 25927 33445
rect 25869 33405 25881 33439
rect 25915 33405 25927 33439
rect 25869 33399 25927 33405
rect 18414 33328 18420 33380
rect 18472 33368 18478 33380
rect 20073 33371 20131 33377
rect 20073 33368 20085 33371
rect 18472 33340 20085 33368
rect 18472 33328 18478 33340
rect 20073 33337 20085 33340
rect 20119 33337 20131 33371
rect 20073 33331 20131 33337
rect 20257 33371 20315 33377
rect 20257 33337 20269 33371
rect 20303 33368 20315 33371
rect 20438 33368 20444 33380
rect 20303 33340 20444 33368
rect 20303 33337 20315 33340
rect 20257 33331 20315 33337
rect 20438 33328 20444 33340
rect 20496 33368 20502 33380
rect 21637 33371 21695 33377
rect 21637 33368 21649 33371
rect 20496 33340 21649 33368
rect 20496 33328 20502 33340
rect 21637 33337 21649 33340
rect 21683 33368 21695 33371
rect 23842 33368 23848 33380
rect 21683 33340 23848 33368
rect 21683 33337 21695 33340
rect 21637 33331 21695 33337
rect 23842 33328 23848 33340
rect 23900 33328 23906 33380
rect 23934 33328 23940 33380
rect 23992 33368 23998 33380
rect 23992 33340 24037 33368
rect 23992 33328 23998 33340
rect 16206 33300 16212 33312
rect 15344 33272 16068 33300
rect 16167 33272 16212 33300
rect 15344 33260 15350 33272
rect 16206 33260 16212 33272
rect 16264 33260 16270 33312
rect 16482 33260 16488 33312
rect 16540 33300 16546 33312
rect 16945 33303 17003 33309
rect 16945 33300 16957 33303
rect 16540 33272 16957 33300
rect 16540 33260 16546 33272
rect 16945 33269 16957 33272
rect 16991 33269 17003 33303
rect 16945 33263 17003 33269
rect 18325 33303 18383 33309
rect 18325 33269 18337 33303
rect 18371 33300 18383 33303
rect 18782 33300 18788 33312
rect 18371 33272 18788 33300
rect 18371 33269 18383 33272
rect 18325 33263 18383 33269
rect 18782 33260 18788 33272
rect 18840 33260 18846 33312
rect 22002 33300 22008 33312
rect 21963 33272 22008 33300
rect 22002 33260 22008 33272
rect 22060 33260 22066 33312
rect 24026 33260 24032 33312
rect 24084 33300 24090 33312
rect 24213 33303 24271 33309
rect 24213 33300 24225 33303
rect 24084 33272 24225 33300
rect 24084 33260 24090 33272
rect 24213 33269 24225 33272
rect 24259 33269 24271 33303
rect 25792 33300 25820 33399
rect 25884 33368 25912 33399
rect 26050 33396 26056 33448
rect 26108 33436 26114 33448
rect 26108 33408 26153 33436
rect 26108 33396 26114 33408
rect 26234 33396 26240 33448
rect 26292 33436 26298 33448
rect 27908 33445 27936 33544
rect 27157 33439 27215 33445
rect 27157 33436 27169 33439
rect 26292 33408 27169 33436
rect 26292 33396 26298 33408
rect 27157 33405 27169 33408
rect 27203 33405 27215 33439
rect 27157 33399 27215 33405
rect 27893 33439 27951 33445
rect 27893 33405 27905 33439
rect 27939 33405 27951 33439
rect 27893 33399 27951 33405
rect 26418 33368 26424 33380
rect 25884 33340 26424 33368
rect 26418 33328 26424 33340
rect 26476 33328 26482 33380
rect 26234 33300 26240 33312
rect 25792 33272 26240 33300
rect 24213 33263 24271 33269
rect 26234 33260 26240 33272
rect 26292 33260 26298 33312
rect 1104 33210 28888 33232
rect 1104 33158 10246 33210
rect 10298 33158 10310 33210
rect 10362 33158 10374 33210
rect 10426 33158 10438 33210
rect 10490 33158 19510 33210
rect 19562 33158 19574 33210
rect 19626 33158 19638 33210
rect 19690 33158 19702 33210
rect 19754 33158 28888 33210
rect 1104 33136 28888 33158
rect 27985 33099 28043 33105
rect 27985 33096 27997 33099
rect 2746 33068 27997 33096
rect 2590 32988 2596 33040
rect 2648 33028 2654 33040
rect 2746 33028 2774 33068
rect 27985 33065 27997 33068
rect 28031 33065 28043 33099
rect 27985 33059 28043 33065
rect 2648 33000 2774 33028
rect 2648 32988 2654 33000
rect 4246 32988 4252 33040
rect 4304 33028 4310 33040
rect 4430 33028 4436 33040
rect 4304 33000 4436 33028
rect 4304 32988 4310 33000
rect 4430 32988 4436 33000
rect 4488 33028 4494 33040
rect 4893 33031 4951 33037
rect 4893 33028 4905 33031
rect 4488 33000 4905 33028
rect 4488 32988 4494 33000
rect 4893 32997 4905 33000
rect 4939 32997 4951 33031
rect 13078 33028 13084 33040
rect 13039 33000 13084 33028
rect 4893 32991 4951 32997
rect 13078 32988 13084 33000
rect 13136 32988 13142 33040
rect 13998 32988 14004 33040
rect 14056 33028 14062 33040
rect 14461 33031 14519 33037
rect 14461 33028 14473 33031
rect 14056 33000 14473 33028
rect 14056 32988 14062 33000
rect 14461 32997 14473 33000
rect 14507 32997 14519 33031
rect 14461 32991 14519 32997
rect 15010 32988 15016 33040
rect 15068 33028 15074 33040
rect 18141 33031 18199 33037
rect 18141 33028 18153 33031
rect 15068 33000 18153 33028
rect 15068 32988 15074 33000
rect 18141 32997 18153 33000
rect 18187 33028 18199 33031
rect 18414 33028 18420 33040
rect 18187 33000 18420 33028
rect 18187 32997 18199 33000
rect 18141 32991 18199 32997
rect 18414 32988 18420 33000
rect 18472 32988 18478 33040
rect 18690 32988 18696 33040
rect 18748 33028 18754 33040
rect 18969 33031 19027 33037
rect 18969 33028 18981 33031
rect 18748 33000 18981 33028
rect 18748 32988 18754 33000
rect 18969 32997 18981 33000
rect 19015 32997 19027 33031
rect 18969 32991 19027 32997
rect 19061 33031 19119 33037
rect 19061 32997 19073 33031
rect 19107 33028 19119 33031
rect 19978 33028 19984 33040
rect 19107 33000 19984 33028
rect 19107 32997 19119 33000
rect 19061 32991 19119 32997
rect 19978 32988 19984 33000
rect 20036 32988 20042 33040
rect 24762 32988 24768 33040
rect 24820 33028 24826 33040
rect 27893 33031 27951 33037
rect 27893 33028 27905 33031
rect 24820 33000 25452 33028
rect 24820 32988 24826 33000
rect 1486 32960 1492 32972
rect 1447 32932 1492 32960
rect 1486 32920 1492 32932
rect 1544 32920 1550 32972
rect 1762 32920 1768 32972
rect 1820 32960 1826 32972
rect 1857 32963 1915 32969
rect 1857 32960 1869 32963
rect 1820 32932 1869 32960
rect 1820 32920 1826 32932
rect 1857 32929 1869 32932
rect 1903 32929 1915 32963
rect 1857 32923 1915 32929
rect 2038 32920 2044 32972
rect 2096 32960 2102 32972
rect 4157 32963 4215 32969
rect 4157 32960 4169 32963
rect 2096 32932 4169 32960
rect 2096 32920 2102 32932
rect 4157 32929 4169 32932
rect 4203 32929 4215 32963
rect 4157 32923 4215 32929
rect 4801 32963 4859 32969
rect 4801 32929 4813 32963
rect 4847 32960 4859 32963
rect 4982 32960 4988 32972
rect 4847 32932 4988 32960
rect 4847 32929 4859 32932
rect 4801 32923 4859 32929
rect 4982 32920 4988 32932
rect 5040 32920 5046 32972
rect 8662 32960 8668 32972
rect 8623 32932 8668 32960
rect 8662 32920 8668 32932
rect 8720 32920 8726 32972
rect 9490 32960 9496 32972
rect 9451 32932 9496 32960
rect 9490 32920 9496 32932
rect 9548 32920 9554 32972
rect 10689 32963 10747 32969
rect 10689 32929 10701 32963
rect 10735 32929 10747 32963
rect 10689 32923 10747 32929
rect 10873 32963 10931 32969
rect 10873 32929 10885 32963
rect 10919 32960 10931 32963
rect 11146 32960 11152 32972
rect 10919 32932 11152 32960
rect 10919 32929 10931 32932
rect 10873 32923 10931 32929
rect 3418 32852 3424 32904
rect 3476 32892 3482 32904
rect 3973 32895 4031 32901
rect 3973 32892 3985 32895
rect 3476 32864 3985 32892
rect 3476 32852 3482 32864
rect 3973 32861 3985 32864
rect 4019 32861 4031 32895
rect 3973 32855 4031 32861
rect 4065 32895 4123 32901
rect 4065 32861 4077 32895
rect 4111 32861 4123 32895
rect 4246 32892 4252 32904
rect 4207 32864 4252 32892
rect 4065 32855 4123 32861
rect 2682 32824 2688 32836
rect 2643 32796 2688 32824
rect 2682 32784 2688 32796
rect 2740 32784 2746 32836
rect 3878 32784 3884 32836
rect 3936 32824 3942 32836
rect 4080 32824 4108 32855
rect 4246 32852 4252 32864
rect 4304 32852 4310 32904
rect 8754 32892 8760 32904
rect 8715 32864 8760 32892
rect 8754 32852 8760 32864
rect 8812 32852 8818 32904
rect 8849 32895 8907 32901
rect 8849 32861 8861 32895
rect 8895 32892 8907 32895
rect 9858 32892 9864 32904
rect 8895 32864 9864 32892
rect 8895 32861 8907 32864
rect 8849 32855 8907 32861
rect 3936 32796 4108 32824
rect 3936 32784 3942 32796
rect 8478 32784 8484 32836
rect 8536 32824 8542 32836
rect 8864 32824 8892 32855
rect 9858 32852 9864 32864
rect 9916 32852 9922 32904
rect 10704 32892 10732 32923
rect 11146 32920 11152 32932
rect 11204 32920 11210 32972
rect 12158 32960 12164 32972
rect 12119 32932 12164 32960
rect 12158 32920 12164 32932
rect 12216 32920 12222 32972
rect 12253 32963 12311 32969
rect 12253 32929 12265 32963
rect 12299 32929 12311 32963
rect 12253 32923 12311 32929
rect 12066 32892 12072 32904
rect 10704 32864 12072 32892
rect 12066 32852 12072 32864
rect 12124 32892 12130 32904
rect 12268 32892 12296 32923
rect 12342 32920 12348 32972
rect 12400 32960 12406 32972
rect 12400 32932 12445 32960
rect 12400 32920 12406 32932
rect 12802 32920 12808 32972
rect 12860 32960 12866 32972
rect 12989 32963 13047 32969
rect 12989 32960 13001 32963
rect 12860 32932 13001 32960
rect 12860 32920 12866 32932
rect 12989 32929 13001 32932
rect 13035 32929 13047 32963
rect 12989 32923 13047 32929
rect 13173 32963 13231 32969
rect 13173 32929 13185 32963
rect 13219 32960 13231 32963
rect 13354 32960 13360 32972
rect 13219 32932 13360 32960
rect 13219 32929 13231 32932
rect 13173 32923 13231 32929
rect 12124 32864 12296 32892
rect 12124 32852 12130 32864
rect 8536 32796 8892 32824
rect 8536 32784 8542 32796
rect 12710 32784 12716 32836
rect 12768 32824 12774 32836
rect 13188 32824 13216 32923
rect 13354 32920 13360 32932
rect 13412 32920 13418 32972
rect 13814 32920 13820 32972
rect 13872 32960 13878 32972
rect 14093 32963 14151 32969
rect 14093 32960 14105 32963
rect 13872 32932 14105 32960
rect 13872 32920 13878 32932
rect 14093 32929 14105 32932
rect 14139 32929 14151 32963
rect 14093 32923 14151 32929
rect 14277 32963 14335 32969
rect 14277 32929 14289 32963
rect 14323 32929 14335 32963
rect 14277 32923 14335 32929
rect 14369 32963 14427 32969
rect 14369 32929 14381 32963
rect 14415 32929 14427 32963
rect 14369 32923 14427 32929
rect 12768 32796 13216 32824
rect 12768 32784 12774 32796
rect 14182 32784 14188 32836
rect 14240 32824 14246 32836
rect 14292 32824 14320 32923
rect 14384 32892 14412 32923
rect 14550 32920 14556 32972
rect 14608 32960 14614 32972
rect 14734 32960 14740 32972
rect 14608 32932 14653 32960
rect 14695 32932 14740 32960
rect 14608 32920 14614 32932
rect 14734 32920 14740 32932
rect 14792 32920 14798 32972
rect 18506 32920 18512 32972
rect 18564 32960 18570 32972
rect 18785 32963 18843 32969
rect 18785 32960 18797 32963
rect 18564 32932 18797 32960
rect 18564 32920 18570 32932
rect 18785 32929 18797 32932
rect 18831 32929 18843 32963
rect 18785 32923 18843 32929
rect 19153 32963 19211 32969
rect 19153 32929 19165 32963
rect 19199 32960 19211 32963
rect 19199 32932 19840 32960
rect 19199 32929 19211 32932
rect 19153 32923 19211 32929
rect 16114 32892 16120 32904
rect 14384 32864 16120 32892
rect 16114 32852 16120 32864
rect 16172 32852 16178 32904
rect 16482 32852 16488 32904
rect 16540 32892 16546 32904
rect 16540 32864 18368 32892
rect 16540 32852 16546 32864
rect 16500 32824 16528 32852
rect 14240 32796 16528 32824
rect 18340 32824 18368 32864
rect 19150 32824 19156 32836
rect 18340 32796 19156 32824
rect 14240 32784 14246 32796
rect 19150 32784 19156 32796
rect 19208 32784 19214 32836
rect 3786 32756 3792 32768
rect 3747 32728 3792 32756
rect 3786 32716 3792 32728
rect 3844 32716 3850 32768
rect 7834 32716 7840 32768
rect 7892 32756 7898 32768
rect 8297 32759 8355 32765
rect 8297 32756 8309 32759
rect 7892 32728 8309 32756
rect 7892 32716 7898 32728
rect 8297 32725 8309 32728
rect 8343 32725 8355 32759
rect 8297 32719 8355 32725
rect 9585 32759 9643 32765
rect 9585 32725 9597 32759
rect 9631 32756 9643 32759
rect 9858 32756 9864 32768
rect 9631 32728 9864 32756
rect 9631 32725 9643 32728
rect 9585 32719 9643 32725
rect 9858 32716 9864 32728
rect 9916 32716 9922 32768
rect 10781 32759 10839 32765
rect 10781 32725 10793 32759
rect 10827 32756 10839 32759
rect 11330 32756 11336 32768
rect 10827 32728 11336 32756
rect 10827 32725 10839 32728
rect 10781 32719 10839 32725
rect 11330 32716 11336 32728
rect 11388 32716 11394 32768
rect 11974 32716 11980 32768
rect 12032 32756 12038 32768
rect 12158 32756 12164 32768
rect 12032 32728 12164 32756
rect 12032 32716 12038 32728
rect 12158 32716 12164 32728
rect 12216 32716 12222 32768
rect 12529 32759 12587 32765
rect 12529 32725 12541 32759
rect 12575 32756 12587 32759
rect 13262 32756 13268 32768
rect 12575 32728 13268 32756
rect 12575 32725 12587 32728
rect 12529 32719 12587 32725
rect 13262 32716 13268 32728
rect 13320 32716 13326 32768
rect 17862 32716 17868 32768
rect 17920 32756 17926 32768
rect 18233 32759 18291 32765
rect 18233 32756 18245 32759
rect 17920 32728 18245 32756
rect 17920 32716 17926 32728
rect 18233 32725 18245 32728
rect 18279 32756 18291 32759
rect 18690 32756 18696 32768
rect 18279 32728 18696 32756
rect 18279 32725 18291 32728
rect 18233 32719 18291 32725
rect 18690 32716 18696 32728
rect 18748 32716 18754 32768
rect 18966 32716 18972 32768
rect 19024 32756 19030 32768
rect 19337 32759 19395 32765
rect 19337 32756 19349 32759
rect 19024 32728 19349 32756
rect 19024 32716 19030 32728
rect 19337 32725 19349 32728
rect 19383 32725 19395 32759
rect 19812 32756 19840 32932
rect 19886 32920 19892 32972
rect 19944 32960 19950 32972
rect 20625 32963 20683 32969
rect 20625 32960 20637 32963
rect 19944 32932 20637 32960
rect 19944 32920 19950 32932
rect 20625 32929 20637 32932
rect 20671 32929 20683 32963
rect 20625 32923 20683 32929
rect 22094 32920 22100 32972
rect 22152 32960 22158 32972
rect 24486 32960 24492 32972
rect 22152 32932 24492 32960
rect 22152 32920 22158 32932
rect 24486 32920 24492 32932
rect 24544 32920 24550 32972
rect 24854 32920 24860 32972
rect 24912 32960 24918 32972
rect 25424 32969 25452 33000
rect 25516 33000 27905 33028
rect 25041 32963 25099 32969
rect 25041 32960 25053 32963
rect 24912 32932 25053 32960
rect 24912 32920 24918 32932
rect 25041 32929 25053 32932
rect 25087 32929 25099 32963
rect 25041 32923 25099 32929
rect 25225 32963 25283 32969
rect 25225 32929 25237 32963
rect 25271 32929 25283 32963
rect 25225 32923 25283 32929
rect 25317 32963 25375 32969
rect 25317 32929 25329 32963
rect 25363 32929 25375 32963
rect 25317 32923 25375 32929
rect 25409 32963 25467 32969
rect 25409 32929 25421 32963
rect 25455 32929 25467 32963
rect 25409 32923 25467 32929
rect 20254 32892 20260 32904
rect 20215 32864 20260 32892
rect 20254 32852 20260 32864
rect 20312 32852 20318 32904
rect 20441 32895 20499 32901
rect 20441 32861 20453 32895
rect 20487 32861 20499 32895
rect 20441 32855 20499 32861
rect 20456 32824 20484 32855
rect 20530 32852 20536 32904
rect 20588 32892 20594 32904
rect 20717 32895 20775 32901
rect 20588 32864 20633 32892
rect 20588 32852 20594 32864
rect 20717 32861 20729 32895
rect 20763 32892 20775 32895
rect 20806 32892 20812 32904
rect 20763 32864 20812 32892
rect 20763 32861 20775 32864
rect 20717 32855 20775 32861
rect 20806 32852 20812 32864
rect 20864 32852 20870 32904
rect 22370 32852 22376 32904
rect 22428 32892 22434 32904
rect 22557 32895 22615 32901
rect 22557 32892 22569 32895
rect 22428 32864 22569 32892
rect 22428 32852 22434 32864
rect 22557 32861 22569 32864
rect 22603 32861 22615 32895
rect 22830 32892 22836 32904
rect 22791 32864 22836 32892
rect 22557 32855 22615 32861
rect 22830 32852 22836 32864
rect 22888 32852 22894 32904
rect 23842 32852 23848 32904
rect 23900 32892 23906 32904
rect 25240 32892 25268 32923
rect 23900 32864 25268 32892
rect 23900 32852 23906 32864
rect 21082 32824 21088 32836
rect 20456 32796 21088 32824
rect 21082 32784 21088 32796
rect 21140 32784 21146 32836
rect 23492 32796 24072 32824
rect 20714 32756 20720 32768
rect 19812 32728 20720 32756
rect 19337 32719 19395 32725
rect 20714 32716 20720 32728
rect 20772 32716 20778 32768
rect 23014 32716 23020 32768
rect 23072 32756 23078 32768
rect 23492 32756 23520 32796
rect 23934 32756 23940 32768
rect 23072 32728 23520 32756
rect 23895 32728 23940 32756
rect 23072 32716 23078 32728
rect 23934 32716 23940 32728
rect 23992 32716 23998 32768
rect 24044 32756 24072 32796
rect 24302 32784 24308 32836
rect 24360 32824 24366 32836
rect 24762 32824 24768 32836
rect 24360 32796 24768 32824
rect 24360 32784 24366 32796
rect 24762 32784 24768 32796
rect 24820 32784 24826 32836
rect 24854 32784 24860 32836
rect 24912 32824 24918 32836
rect 24964 32824 24992 32864
rect 24912 32796 24992 32824
rect 24912 32784 24918 32796
rect 25130 32784 25136 32836
rect 25188 32824 25194 32836
rect 25332 32824 25360 32923
rect 25188 32796 25360 32824
rect 25188 32784 25194 32796
rect 25516 32756 25544 33000
rect 27893 32997 27905 33000
rect 27939 32997 27951 33031
rect 27893 32991 27951 32997
rect 26421 32963 26479 32969
rect 26421 32929 26433 32963
rect 26467 32960 26479 32963
rect 27246 32960 27252 32972
rect 26467 32932 27252 32960
rect 26467 32929 26479 32932
rect 26421 32923 26479 32929
rect 27246 32920 27252 32932
rect 27304 32920 27310 32972
rect 26234 32892 26240 32904
rect 26195 32864 26240 32892
rect 26234 32852 26240 32864
rect 26292 32852 26298 32904
rect 26326 32852 26332 32904
rect 26384 32892 26390 32904
rect 26513 32895 26571 32901
rect 26384 32864 26429 32892
rect 26384 32852 26390 32864
rect 26513 32861 26525 32895
rect 26559 32861 26571 32895
rect 26513 32855 26571 32861
rect 25593 32827 25651 32833
rect 25593 32793 25605 32827
rect 25639 32824 25651 32827
rect 26528 32824 26556 32855
rect 25639 32796 26556 32824
rect 25639 32793 25651 32796
rect 25593 32787 25651 32793
rect 24044 32728 25544 32756
rect 25774 32716 25780 32768
rect 25832 32756 25838 32768
rect 26053 32759 26111 32765
rect 26053 32756 26065 32759
rect 25832 32728 26065 32756
rect 25832 32716 25838 32728
rect 26053 32725 26065 32728
rect 26099 32725 26111 32759
rect 26053 32719 26111 32725
rect 1104 32666 28888 32688
rect 1104 32614 5614 32666
rect 5666 32614 5678 32666
rect 5730 32614 5742 32666
rect 5794 32614 5806 32666
rect 5858 32614 14878 32666
rect 14930 32614 14942 32666
rect 14994 32614 15006 32666
rect 15058 32614 15070 32666
rect 15122 32614 24142 32666
rect 24194 32614 24206 32666
rect 24258 32614 24270 32666
rect 24322 32614 24334 32666
rect 24386 32614 28888 32666
rect 1104 32592 28888 32614
rect 1489 32555 1547 32561
rect 1489 32521 1501 32555
rect 1535 32552 1547 32555
rect 4614 32552 4620 32564
rect 1535 32524 4620 32552
rect 1535 32521 1547 32524
rect 1489 32515 1547 32521
rect 4614 32512 4620 32524
rect 4672 32512 4678 32564
rect 4724 32524 7420 32552
rect 2406 32444 2412 32496
rect 2464 32484 2470 32496
rect 4724 32484 4752 32524
rect 2464 32456 4752 32484
rect 4801 32487 4859 32493
rect 2464 32444 2470 32456
rect 4801 32453 4813 32487
rect 4847 32484 4859 32487
rect 6270 32484 6276 32496
rect 4847 32456 6276 32484
rect 4847 32453 4859 32456
rect 4801 32447 4859 32453
rect 6270 32444 6276 32456
rect 6328 32444 6334 32496
rect 7098 32444 7104 32496
rect 7156 32484 7162 32496
rect 7193 32487 7251 32493
rect 7193 32484 7205 32487
rect 7156 32456 7205 32484
rect 7156 32444 7162 32456
rect 7193 32453 7205 32456
rect 7239 32453 7251 32487
rect 7392 32484 7420 32524
rect 8110 32512 8116 32564
rect 8168 32552 8174 32564
rect 8389 32555 8447 32561
rect 8389 32552 8401 32555
rect 8168 32524 8401 32552
rect 8168 32512 8174 32524
rect 8389 32521 8401 32524
rect 8435 32521 8447 32555
rect 18509 32555 18567 32561
rect 8389 32515 8447 32521
rect 9508 32524 17264 32552
rect 9508 32484 9536 32524
rect 7392 32456 9536 32484
rect 9600 32456 13492 32484
rect 7193 32447 7251 32453
rect 1780 32388 2774 32416
rect 1780 32357 1808 32388
rect 2746 32360 2774 32388
rect 4430 32376 4436 32428
rect 4488 32416 4494 32428
rect 4614 32416 4620 32428
rect 4488 32388 4620 32416
rect 4488 32376 4494 32388
rect 4614 32376 4620 32388
rect 4672 32376 4678 32428
rect 5626 32376 5632 32428
rect 5684 32416 5690 32428
rect 6457 32419 6515 32425
rect 6457 32416 6469 32419
rect 5684 32388 6469 32416
rect 5684 32376 5690 32388
rect 6457 32385 6469 32388
rect 6503 32385 6515 32419
rect 6457 32379 6515 32385
rect 7745 32419 7803 32425
rect 7745 32385 7757 32419
rect 7791 32416 7803 32419
rect 9600 32416 9628 32456
rect 7791 32388 9628 32416
rect 7791 32385 7803 32388
rect 7745 32379 7803 32385
rect 1765 32351 1823 32357
rect 1765 32317 1777 32351
rect 1811 32317 1823 32351
rect 1765 32311 1823 32317
rect 2041 32351 2099 32357
rect 2041 32317 2053 32351
rect 2087 32348 2099 32351
rect 2222 32348 2228 32360
rect 2087 32320 2228 32348
rect 2087 32317 2099 32320
rect 2041 32311 2099 32317
rect 2222 32308 2228 32320
rect 2280 32308 2286 32360
rect 2501 32351 2559 32357
rect 2501 32317 2513 32351
rect 2547 32348 2559 32351
rect 2590 32348 2596 32360
rect 2547 32320 2596 32348
rect 2547 32317 2559 32320
rect 2501 32311 2559 32317
rect 2590 32308 2596 32320
rect 2648 32308 2654 32360
rect 2746 32320 2780 32360
rect 2774 32308 2780 32320
rect 2832 32308 2838 32360
rect 2869 32351 2927 32357
rect 2869 32317 2881 32351
rect 2915 32348 2927 32351
rect 2958 32348 2964 32360
rect 2915 32320 2964 32348
rect 2915 32317 2927 32320
rect 2869 32311 2927 32317
rect 2958 32308 2964 32320
rect 3016 32308 3022 32360
rect 3053 32351 3111 32357
rect 3053 32317 3065 32351
rect 3099 32317 3111 32351
rect 3053 32311 3111 32317
rect 5077 32351 5135 32357
rect 5077 32317 5089 32351
rect 5123 32348 5135 32351
rect 6086 32348 6092 32360
rect 5123 32320 6092 32348
rect 5123 32317 5135 32320
rect 5077 32311 5135 32317
rect 2130 32240 2136 32292
rect 2188 32280 2194 32292
rect 3068 32280 3096 32311
rect 6086 32308 6092 32320
rect 6144 32308 6150 32360
rect 6178 32308 6184 32360
rect 6236 32348 6242 32360
rect 6273 32351 6331 32357
rect 6273 32348 6285 32351
rect 6236 32320 6285 32348
rect 6236 32308 6242 32320
rect 6273 32317 6285 32320
rect 6319 32317 6331 32351
rect 6273 32311 6331 32317
rect 6362 32308 6368 32360
rect 6420 32348 6426 32360
rect 7760 32348 7788 32379
rect 9674 32376 9680 32428
rect 9732 32416 9738 32428
rect 9950 32416 9956 32428
rect 9732 32388 9956 32416
rect 9732 32376 9738 32388
rect 9950 32376 9956 32388
rect 10008 32416 10014 32428
rect 10045 32419 10103 32425
rect 10045 32416 10057 32419
rect 10008 32388 10057 32416
rect 10008 32376 10014 32388
rect 10045 32385 10057 32388
rect 10091 32385 10103 32419
rect 10045 32379 10103 32385
rect 10778 32376 10784 32428
rect 10836 32376 10842 32428
rect 11164 32388 12664 32416
rect 8294 32348 8300 32360
rect 6420 32320 7788 32348
rect 8255 32320 8300 32348
rect 6420 32308 6426 32320
rect 8294 32308 8300 32320
rect 8352 32308 8358 32360
rect 9858 32348 9864 32360
rect 9819 32320 9864 32348
rect 9858 32308 9864 32320
rect 9916 32308 9922 32360
rect 10796 32348 10824 32376
rect 11164 32357 11192 32388
rect 10965 32351 11023 32357
rect 10965 32348 10977 32351
rect 10796 32320 10977 32348
rect 10965 32317 10977 32320
rect 11011 32317 11023 32351
rect 10965 32311 11023 32317
rect 11057 32351 11115 32357
rect 11057 32317 11069 32351
rect 11103 32317 11115 32351
rect 11057 32311 11115 32317
rect 11149 32351 11207 32357
rect 11149 32317 11161 32351
rect 11195 32317 11207 32351
rect 11330 32348 11336 32360
rect 11291 32320 11336 32348
rect 11149 32311 11207 32317
rect 2188 32252 3096 32280
rect 5353 32283 5411 32289
rect 2188 32240 2194 32252
rect 5353 32249 5365 32283
rect 5399 32280 5411 32283
rect 5534 32280 5540 32292
rect 5399 32252 5540 32280
rect 5399 32249 5411 32252
rect 5353 32243 5411 32249
rect 5534 32240 5540 32252
rect 5592 32240 5598 32292
rect 5920 32252 7052 32280
rect 4890 32172 4896 32224
rect 4948 32212 4954 32224
rect 5920 32221 5948 32252
rect 5261 32215 5319 32221
rect 5261 32212 5273 32215
rect 4948 32184 5273 32212
rect 4948 32172 4954 32184
rect 5261 32181 5273 32184
rect 5307 32181 5319 32215
rect 5261 32175 5319 32181
rect 5905 32215 5963 32221
rect 5905 32181 5917 32215
rect 5951 32181 5963 32215
rect 5905 32175 5963 32181
rect 6362 32172 6368 32224
rect 6420 32212 6426 32224
rect 7024 32212 7052 32252
rect 7098 32240 7104 32292
rect 7156 32280 7162 32292
rect 7469 32283 7527 32289
rect 7469 32280 7481 32283
rect 7156 32252 7481 32280
rect 7156 32240 7162 32252
rect 7469 32249 7481 32252
rect 7515 32249 7527 32283
rect 7469 32243 7527 32249
rect 9398 32240 9404 32292
rect 9456 32280 9462 32292
rect 11072 32280 11100 32311
rect 11330 32308 11336 32320
rect 11388 32308 11394 32360
rect 11882 32308 11888 32360
rect 11940 32348 11946 32360
rect 12268 32357 12296 32388
rect 12069 32351 12127 32357
rect 12069 32348 12081 32351
rect 11940 32320 12081 32348
rect 11940 32308 11946 32320
rect 12069 32317 12081 32320
rect 12115 32317 12127 32351
rect 12069 32311 12127 32317
rect 12161 32351 12219 32357
rect 12161 32317 12173 32351
rect 12207 32317 12219 32351
rect 12161 32311 12219 32317
rect 12253 32351 12311 32357
rect 12253 32317 12265 32351
rect 12299 32317 12311 32351
rect 12253 32311 12311 32317
rect 12176 32280 12204 32311
rect 12434 32308 12440 32360
rect 12492 32348 12498 32360
rect 12636 32348 12664 32388
rect 12802 32376 12808 32428
rect 12860 32416 12866 32428
rect 13262 32416 13268 32428
rect 12860 32388 13268 32416
rect 12860 32376 12866 32388
rect 13262 32376 13268 32388
rect 13320 32416 13326 32428
rect 13357 32419 13415 32425
rect 13357 32416 13369 32419
rect 13320 32388 13369 32416
rect 13320 32376 13326 32388
rect 13357 32385 13369 32388
rect 13403 32385 13415 32419
rect 13464 32416 13492 32456
rect 13538 32444 13544 32496
rect 13596 32484 13602 32496
rect 13633 32487 13691 32493
rect 13633 32484 13645 32487
rect 13596 32456 13645 32484
rect 13596 32444 13602 32456
rect 13633 32453 13645 32456
rect 13679 32453 13691 32487
rect 13633 32447 13691 32453
rect 13817 32487 13875 32493
rect 13817 32453 13829 32487
rect 13863 32484 13875 32487
rect 13906 32484 13912 32496
rect 13863 32456 13912 32484
rect 13863 32453 13875 32456
rect 13817 32447 13875 32453
rect 13906 32444 13912 32456
rect 13964 32444 13970 32496
rect 15930 32444 15936 32496
rect 15988 32444 15994 32496
rect 16117 32487 16175 32493
rect 16117 32453 16129 32487
rect 16163 32484 16175 32487
rect 16482 32484 16488 32496
rect 16163 32456 16488 32484
rect 16163 32453 16175 32456
rect 16117 32447 16175 32453
rect 16482 32444 16488 32456
rect 16540 32444 16546 32496
rect 17236 32484 17264 32524
rect 18509 32521 18521 32555
rect 18555 32552 18567 32555
rect 18598 32552 18604 32564
rect 18555 32524 18604 32552
rect 18555 32521 18567 32524
rect 18509 32515 18567 32521
rect 18598 32512 18604 32524
rect 18656 32512 18662 32564
rect 18782 32512 18788 32564
rect 18840 32552 18846 32564
rect 20530 32552 20536 32564
rect 18840 32524 20536 32552
rect 18840 32512 18846 32524
rect 20530 32512 20536 32524
rect 20588 32512 20594 32564
rect 20806 32552 20812 32564
rect 20767 32524 20812 32552
rect 20806 32512 20812 32524
rect 20864 32512 20870 32564
rect 21269 32555 21327 32561
rect 21269 32521 21281 32555
rect 21315 32552 21327 32555
rect 21726 32552 21732 32564
rect 21315 32524 21732 32552
rect 21315 32521 21327 32524
rect 21269 32515 21327 32521
rect 21726 32512 21732 32524
rect 21784 32512 21790 32564
rect 22370 32512 22376 32564
rect 22428 32552 22434 32564
rect 22646 32552 22652 32564
rect 22428 32524 22652 32552
rect 22428 32512 22434 32524
rect 22646 32512 22652 32524
rect 22704 32512 22710 32564
rect 23014 32552 23020 32564
rect 22975 32524 23020 32552
rect 23014 32512 23020 32524
rect 23072 32512 23078 32564
rect 23661 32555 23719 32561
rect 23661 32521 23673 32555
rect 23707 32552 23719 32555
rect 23750 32552 23756 32564
rect 23707 32524 23756 32552
rect 23707 32521 23719 32524
rect 23661 32515 23719 32521
rect 23750 32512 23756 32524
rect 23808 32512 23814 32564
rect 25777 32555 25835 32561
rect 25777 32521 25789 32555
rect 25823 32552 25835 32555
rect 26050 32552 26056 32564
rect 25823 32524 26056 32552
rect 25823 32521 25835 32524
rect 25777 32515 25835 32521
rect 26050 32512 26056 32524
rect 26108 32512 26114 32564
rect 17236 32456 19104 32484
rect 15102 32416 15108 32428
rect 13464 32388 15108 32416
rect 13357 32379 13415 32385
rect 15102 32376 15108 32388
rect 15160 32376 15166 32428
rect 15948 32416 15976 32444
rect 17494 32416 17500 32428
rect 15212 32388 15976 32416
rect 17420 32388 17500 32416
rect 15212 32348 15240 32388
rect 12492 32320 12537 32348
rect 12636 32320 15240 32348
rect 12492 32308 12498 32320
rect 15286 32308 15292 32360
rect 15344 32348 15350 32360
rect 15933 32351 15991 32357
rect 15933 32348 15945 32351
rect 15344 32320 15945 32348
rect 15344 32308 15350 32320
rect 15933 32317 15945 32320
rect 15979 32348 15991 32351
rect 16022 32348 16028 32360
rect 15979 32320 16028 32348
rect 15979 32317 15991 32320
rect 15933 32311 15991 32317
rect 16022 32308 16028 32320
rect 16080 32308 16086 32360
rect 17420 32357 17448 32388
rect 17494 32376 17500 32388
rect 17552 32376 17558 32428
rect 18506 32376 18512 32428
rect 18564 32416 18570 32428
rect 18693 32419 18751 32425
rect 18693 32416 18705 32419
rect 18564 32388 18705 32416
rect 18564 32376 18570 32388
rect 18693 32385 18705 32388
rect 18739 32385 18751 32419
rect 18966 32416 18972 32428
rect 18927 32388 18972 32416
rect 18693 32379 18751 32385
rect 18966 32376 18972 32388
rect 19024 32376 19030 32428
rect 19076 32416 19104 32456
rect 19150 32444 19156 32496
rect 19208 32484 19214 32496
rect 24118 32484 24124 32496
rect 19208 32456 23612 32484
rect 19208 32444 19214 32456
rect 20346 32416 20352 32428
rect 19076 32388 19288 32416
rect 17405 32351 17463 32357
rect 17405 32317 17417 32351
rect 17451 32317 17463 32351
rect 17770 32348 17776 32360
rect 17405 32311 17463 32317
rect 17512 32320 17776 32348
rect 13446 32280 13452 32292
rect 9456 32252 10824 32280
rect 11072 32252 13452 32280
rect 9456 32240 9462 32252
rect 7653 32215 7711 32221
rect 7653 32212 7665 32215
rect 6420 32184 6465 32212
rect 7024 32184 7665 32212
rect 6420 32172 6426 32184
rect 7653 32181 7665 32184
rect 7699 32181 7711 32215
rect 7653 32175 7711 32181
rect 8754 32172 8760 32224
rect 8812 32212 8818 32224
rect 9493 32215 9551 32221
rect 9493 32212 9505 32215
rect 8812 32184 9505 32212
rect 8812 32172 8818 32184
rect 9493 32181 9505 32184
rect 9539 32181 9551 32215
rect 9493 32175 9551 32181
rect 9582 32172 9588 32224
rect 9640 32212 9646 32224
rect 9858 32212 9864 32224
rect 9640 32184 9864 32212
rect 9640 32172 9646 32184
rect 9858 32172 9864 32184
rect 9916 32172 9922 32224
rect 9950 32172 9956 32224
rect 10008 32212 10014 32224
rect 10686 32212 10692 32224
rect 10008 32184 10053 32212
rect 10647 32184 10692 32212
rect 10008 32172 10014 32184
rect 10686 32172 10692 32184
rect 10744 32172 10750 32224
rect 10796 32212 10824 32252
rect 13446 32240 13452 32252
rect 13504 32240 13510 32292
rect 14918 32240 14924 32292
rect 14976 32280 14982 32292
rect 17512 32280 17540 32320
rect 17770 32308 17776 32320
rect 17828 32308 17834 32360
rect 18782 32348 18788 32360
rect 18743 32320 18788 32348
rect 18782 32308 18788 32320
rect 18840 32308 18846 32360
rect 18877 32351 18935 32357
rect 18877 32317 18889 32351
rect 18923 32317 18935 32351
rect 18877 32311 18935 32317
rect 14976 32252 17540 32280
rect 17589 32283 17647 32289
rect 14976 32240 14982 32252
rect 17589 32249 17601 32283
rect 17635 32249 17647 32283
rect 17589 32243 17647 32249
rect 11793 32215 11851 32221
rect 11793 32212 11805 32215
rect 10796 32184 11805 32212
rect 11793 32181 11805 32184
rect 11839 32181 11851 32215
rect 11793 32175 11851 32181
rect 15930 32172 15936 32224
rect 15988 32212 15994 32224
rect 16574 32212 16580 32224
rect 15988 32184 16580 32212
rect 15988 32172 15994 32184
rect 16574 32172 16580 32184
rect 16632 32172 16638 32224
rect 17034 32172 17040 32224
rect 17092 32212 17098 32224
rect 17604 32212 17632 32243
rect 17678 32240 17684 32292
rect 17736 32280 17742 32292
rect 17736 32252 17781 32280
rect 17736 32240 17742 32252
rect 18046 32240 18052 32292
rect 18104 32280 18110 32292
rect 18892 32280 18920 32311
rect 19150 32280 19156 32292
rect 18104 32252 18920 32280
rect 18984 32252 19156 32280
rect 18104 32240 18110 32252
rect 17862 32212 17868 32224
rect 17092 32184 17868 32212
rect 17092 32172 17098 32184
rect 17862 32172 17868 32184
rect 17920 32172 17926 32224
rect 17957 32215 18015 32221
rect 17957 32181 17969 32215
rect 18003 32212 18015 32215
rect 18984 32212 19012 32252
rect 19150 32240 19156 32252
rect 19208 32240 19214 32292
rect 18003 32184 19012 32212
rect 19260 32212 19288 32388
rect 20272 32388 20352 32416
rect 20272 32357 20300 32388
rect 20346 32376 20352 32388
rect 20404 32376 20410 32428
rect 20530 32376 20536 32428
rect 20588 32416 20594 32428
rect 21545 32419 21603 32425
rect 21545 32416 21557 32419
rect 20588 32388 21557 32416
rect 20588 32376 20594 32388
rect 21545 32385 21557 32388
rect 21591 32385 21603 32419
rect 21545 32379 21603 32385
rect 21729 32419 21787 32425
rect 21729 32385 21741 32419
rect 21775 32416 21787 32419
rect 22002 32416 22008 32428
rect 21775 32388 22008 32416
rect 21775 32385 21787 32388
rect 21729 32379 21787 32385
rect 22002 32376 22008 32388
rect 22060 32376 22066 32428
rect 23584 32416 23612 32456
rect 23952 32456 24124 32484
rect 23952 32425 23980 32456
rect 24118 32444 24124 32456
rect 24176 32484 24182 32496
rect 26326 32484 26332 32496
rect 24176 32456 26332 32484
rect 24176 32444 24182 32456
rect 26326 32444 26332 32456
rect 26384 32444 26390 32496
rect 23845 32419 23903 32425
rect 23845 32416 23857 32419
rect 23584 32388 23857 32416
rect 20257 32351 20315 32357
rect 20257 32317 20269 32351
rect 20303 32317 20315 32351
rect 20438 32348 20444 32360
rect 20399 32320 20444 32348
rect 20257 32311 20315 32317
rect 20438 32308 20444 32320
rect 20496 32308 20502 32360
rect 20625 32351 20683 32357
rect 20625 32317 20637 32351
rect 20671 32348 20683 32351
rect 20714 32348 20720 32360
rect 20671 32320 20720 32348
rect 20671 32317 20683 32320
rect 20625 32311 20683 32317
rect 20714 32308 20720 32320
rect 20772 32308 20778 32360
rect 21082 32308 21088 32360
rect 21140 32348 21146 32360
rect 21453 32351 21511 32357
rect 21453 32348 21465 32351
rect 21140 32320 21465 32348
rect 21140 32308 21146 32320
rect 21453 32317 21465 32320
rect 21499 32317 21511 32351
rect 21453 32311 21511 32317
rect 21628 32351 21686 32357
rect 21628 32317 21640 32351
rect 21674 32348 21686 32351
rect 22094 32348 22100 32360
rect 21674 32320 22100 32348
rect 21674 32317 21686 32320
rect 21628 32311 21686 32317
rect 22094 32308 22100 32320
rect 22152 32308 22158 32360
rect 23201 32351 23259 32357
rect 23201 32317 23213 32351
rect 23247 32317 23259 32351
rect 23201 32311 23259 32317
rect 20530 32240 20536 32292
rect 20588 32280 20594 32292
rect 23216 32280 23244 32311
rect 23290 32280 23296 32292
rect 20588 32252 20633 32280
rect 23216 32252 23296 32280
rect 20588 32240 20594 32252
rect 23290 32240 23296 32252
rect 23348 32240 23354 32292
rect 23584 32280 23612 32388
rect 23845 32385 23857 32388
rect 23891 32385 23903 32419
rect 23845 32379 23903 32385
rect 23937 32419 23995 32425
rect 23937 32385 23949 32419
rect 23983 32385 23995 32419
rect 23937 32379 23995 32385
rect 24029 32419 24087 32425
rect 24029 32385 24041 32419
rect 24075 32385 24087 32419
rect 24029 32379 24087 32385
rect 23658 32308 23664 32360
rect 23716 32348 23722 32360
rect 24044 32348 24072 32379
rect 24394 32376 24400 32428
rect 24452 32416 24458 32428
rect 24452 32388 25636 32416
rect 24452 32376 24458 32388
rect 23716 32320 24072 32348
rect 24121 32351 24179 32357
rect 23716 32308 23722 32320
rect 24121 32317 24133 32351
rect 24167 32317 24179 32351
rect 25222 32348 25228 32360
rect 25183 32320 25228 32348
rect 24121 32311 24179 32317
rect 23584 32252 23980 32280
rect 23842 32212 23848 32224
rect 19260 32184 23848 32212
rect 18003 32181 18015 32184
rect 17957 32175 18015 32181
rect 23842 32172 23848 32184
rect 23900 32172 23906 32224
rect 23952 32212 23980 32252
rect 24026 32240 24032 32292
rect 24084 32280 24090 32292
rect 24136 32280 24164 32311
rect 25222 32308 25228 32320
rect 25280 32308 25286 32360
rect 25608 32357 25636 32388
rect 25593 32351 25651 32357
rect 25593 32317 25605 32351
rect 25639 32317 25651 32351
rect 25593 32311 25651 32317
rect 25774 32308 25780 32360
rect 25832 32348 25838 32360
rect 26789 32351 26847 32357
rect 26789 32348 26801 32351
rect 25832 32320 26801 32348
rect 25832 32308 25838 32320
rect 26789 32317 26801 32320
rect 26835 32317 26847 32351
rect 26789 32311 26847 32317
rect 24084 32252 24164 32280
rect 24084 32240 24090 32252
rect 24854 32240 24860 32292
rect 24912 32280 24918 32292
rect 25409 32283 25467 32289
rect 25409 32280 25421 32283
rect 24912 32252 25421 32280
rect 24912 32240 24918 32252
rect 25409 32249 25421 32252
rect 25455 32249 25467 32283
rect 25409 32243 25467 32249
rect 25501 32283 25559 32289
rect 25501 32249 25513 32283
rect 25547 32280 25559 32283
rect 25866 32280 25872 32292
rect 25547 32252 25872 32280
rect 25547 32249 25559 32252
rect 25501 32243 25559 32249
rect 25866 32240 25872 32252
rect 25924 32240 25930 32292
rect 27056 32283 27114 32289
rect 27056 32249 27068 32283
rect 27102 32280 27114 32283
rect 27430 32280 27436 32292
rect 27102 32252 27436 32280
rect 27102 32249 27114 32252
rect 27056 32243 27114 32249
rect 27430 32240 27436 32252
rect 27488 32240 27494 32292
rect 26234 32212 26240 32224
rect 23952 32184 26240 32212
rect 26234 32172 26240 32184
rect 26292 32172 26298 32224
rect 27614 32172 27620 32224
rect 27672 32212 27678 32224
rect 28169 32215 28227 32221
rect 28169 32212 28181 32215
rect 27672 32184 28181 32212
rect 27672 32172 27678 32184
rect 28169 32181 28181 32184
rect 28215 32181 28227 32215
rect 28169 32175 28227 32181
rect 1104 32122 28888 32144
rect 1104 32070 10246 32122
rect 10298 32070 10310 32122
rect 10362 32070 10374 32122
rect 10426 32070 10438 32122
rect 10490 32070 19510 32122
rect 19562 32070 19574 32122
rect 19626 32070 19638 32122
rect 19690 32070 19702 32122
rect 19754 32070 28888 32122
rect 1104 32048 28888 32070
rect 2038 32008 2044 32020
rect 1999 31980 2044 32008
rect 2038 31968 2044 31980
rect 2096 31968 2102 32020
rect 2409 32011 2467 32017
rect 2409 31977 2421 32011
rect 2455 32008 2467 32011
rect 2774 32008 2780 32020
rect 2455 31980 2780 32008
rect 2455 31977 2467 31980
rect 2409 31971 2467 31977
rect 2774 31968 2780 31980
rect 2832 32008 2838 32020
rect 3142 32008 3148 32020
rect 2832 31980 3148 32008
rect 2832 31968 2838 31980
rect 3142 31968 3148 31980
rect 3200 32008 3206 32020
rect 3602 32008 3608 32020
rect 3200 31980 3608 32008
rect 3200 31968 3206 31980
rect 3602 31968 3608 31980
rect 3660 31968 3666 32020
rect 4890 32008 4896 32020
rect 4851 31980 4896 32008
rect 4890 31968 4896 31980
rect 4948 31968 4954 32020
rect 5258 32008 5264 32020
rect 5219 31980 5264 32008
rect 5258 31968 5264 31980
rect 5316 31968 5322 32020
rect 5534 31968 5540 32020
rect 5592 32008 5598 32020
rect 6270 32008 6276 32020
rect 5592 31980 6276 32008
rect 5592 31968 5598 31980
rect 6270 31968 6276 31980
rect 6328 31968 6334 32020
rect 8662 31968 8668 32020
rect 8720 32008 8726 32020
rect 8849 32011 8907 32017
rect 8849 32008 8861 32011
rect 8720 31980 8861 32008
rect 8720 31968 8726 31980
rect 8849 31977 8861 31980
rect 8895 31977 8907 32011
rect 8849 31971 8907 31977
rect 10689 32011 10747 32017
rect 10689 31977 10701 32011
rect 10735 32008 10747 32011
rect 12434 32008 12440 32020
rect 10735 31980 12440 32008
rect 10735 31977 10747 31980
rect 10689 31971 10747 31977
rect 12434 31968 12440 31980
rect 12492 31968 12498 32020
rect 13262 32008 13268 32020
rect 12912 31980 13268 32008
rect 2590 31940 2596 31952
rect 2240 31912 2596 31940
rect 1394 31872 1400 31884
rect 1355 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 2240 31881 2268 31912
rect 2590 31900 2596 31912
rect 2648 31900 2654 31952
rect 3228 31943 3286 31949
rect 3228 31909 3240 31943
rect 3274 31940 3286 31943
rect 3786 31940 3792 31952
rect 3274 31912 3792 31940
rect 3274 31909 3286 31912
rect 3228 31903 3286 31909
rect 3786 31900 3792 31912
rect 3844 31900 3850 31952
rect 7282 31940 7288 31952
rect 6932 31912 7288 31940
rect 2225 31875 2283 31881
rect 2225 31841 2237 31875
rect 2271 31841 2283 31875
rect 2225 31835 2283 31841
rect 2498 31832 2504 31884
rect 2556 31872 2562 31884
rect 2961 31875 3019 31881
rect 2556 31844 2601 31872
rect 2556 31832 2562 31844
rect 2961 31841 2973 31875
rect 3007 31872 3019 31875
rect 3050 31872 3056 31884
rect 3007 31844 3056 31872
rect 3007 31841 3019 31844
rect 2961 31835 3019 31841
rect 3050 31832 3056 31844
rect 3108 31832 3114 31884
rect 5353 31875 5411 31881
rect 5353 31841 5365 31875
rect 5399 31872 5411 31875
rect 6730 31872 6736 31884
rect 5399 31844 6736 31872
rect 5399 31841 5411 31844
rect 5353 31835 5411 31841
rect 6730 31832 6736 31844
rect 6788 31832 6794 31884
rect 1489 31807 1547 31813
rect 1489 31773 1501 31807
rect 1535 31804 1547 31807
rect 2516 31804 2544 31832
rect 1535 31776 2544 31804
rect 1535 31773 1547 31776
rect 1489 31767 1547 31773
rect 5442 31764 5448 31816
rect 5500 31804 5506 31816
rect 5537 31807 5595 31813
rect 5537 31804 5549 31807
rect 5500 31776 5549 31804
rect 5500 31764 5506 31776
rect 5537 31773 5549 31776
rect 5583 31804 5595 31807
rect 5626 31804 5632 31816
rect 5583 31776 5632 31804
rect 5583 31773 5595 31776
rect 5537 31767 5595 31773
rect 5626 31764 5632 31776
rect 5684 31764 5690 31816
rect 6932 31813 6960 31912
rect 7282 31900 7288 31912
rect 7340 31940 7346 31952
rect 7834 31940 7840 31952
rect 7340 31912 7840 31940
rect 7340 31900 7346 31912
rect 7834 31900 7840 31912
rect 7892 31900 7898 31952
rect 8110 31900 8116 31952
rect 8168 31940 8174 31952
rect 8168 31912 8984 31940
rect 8168 31900 8174 31912
rect 7006 31832 7012 31884
rect 7064 31881 7070 31884
rect 7064 31875 7113 31881
rect 7064 31841 7067 31875
rect 7101 31872 7113 31875
rect 8294 31872 8300 31884
rect 7101 31844 8300 31872
rect 7101 31841 7113 31844
rect 7064 31835 7113 31841
rect 7064 31832 7070 31835
rect 6917 31807 6975 31813
rect 6917 31773 6929 31807
rect 6963 31773 6975 31807
rect 6917 31767 6975 31773
rect 8128 31745 8156 31844
rect 8294 31832 8300 31844
rect 8352 31832 8358 31884
rect 8754 31872 8760 31884
rect 8715 31844 8760 31872
rect 8754 31832 8760 31844
rect 8812 31832 8818 31884
rect 8956 31881 8984 31912
rect 10042 31900 10048 31952
rect 10100 31940 10106 31952
rect 10318 31940 10324 31952
rect 10100 31912 10324 31940
rect 10100 31900 10106 31912
rect 10318 31900 10324 31912
rect 10376 31900 10382 31952
rect 12912 31949 12940 31980
rect 13262 31968 13268 31980
rect 13320 31968 13326 32020
rect 14550 32008 14556 32020
rect 14511 31980 14556 32008
rect 14550 31968 14556 31980
rect 14608 31968 14614 32020
rect 18138 31968 18144 32020
rect 18196 32008 18202 32020
rect 18325 32011 18383 32017
rect 18325 32008 18337 32011
rect 18196 31980 18337 32008
rect 18196 31968 18202 31980
rect 18325 31977 18337 31980
rect 18371 31977 18383 32011
rect 18325 31971 18383 31977
rect 18506 31968 18512 32020
rect 18564 32008 18570 32020
rect 21082 32008 21088 32020
rect 18564 31980 21088 32008
rect 18564 31968 18570 31980
rect 21082 31968 21088 31980
rect 21140 31968 21146 32020
rect 21174 31968 21180 32020
rect 21232 32008 21238 32020
rect 22741 32011 22799 32017
rect 22741 32008 22753 32011
rect 21232 31980 22753 32008
rect 21232 31968 21238 31980
rect 22741 31977 22753 31980
rect 22787 32008 22799 32011
rect 22787 31980 22968 32008
rect 22787 31977 22799 31980
rect 22741 31971 22799 31977
rect 12897 31943 12955 31949
rect 12897 31909 12909 31943
rect 12943 31909 12955 31943
rect 12897 31903 12955 31909
rect 13722 31900 13728 31952
rect 13780 31940 13786 31952
rect 14918 31940 14924 31952
rect 13780 31912 14924 31940
rect 13780 31900 13786 31912
rect 14918 31900 14924 31912
rect 14976 31900 14982 31952
rect 15286 31940 15292 31952
rect 15028 31912 15292 31940
rect 8941 31875 8999 31881
rect 8941 31841 8953 31875
rect 8987 31841 8999 31875
rect 8941 31835 8999 31841
rect 9214 31832 9220 31884
rect 9272 31872 9278 31884
rect 9766 31872 9772 31884
rect 9272 31844 9772 31872
rect 9272 31832 9278 31844
rect 9766 31832 9772 31844
rect 9824 31832 9830 31884
rect 10505 31875 10563 31881
rect 10505 31841 10517 31875
rect 10551 31841 10563 31875
rect 10505 31835 10563 31841
rect 10689 31875 10747 31881
rect 10689 31841 10701 31875
rect 10735 31872 10747 31875
rect 11146 31872 11152 31884
rect 10735 31844 11152 31872
rect 10735 31841 10747 31844
rect 10689 31835 10747 31841
rect 10520 31804 10548 31835
rect 11146 31832 11152 31844
rect 11204 31832 11210 31884
rect 12161 31875 12219 31881
rect 12161 31841 12173 31875
rect 12207 31872 12219 31875
rect 13538 31872 13544 31884
rect 12207 31844 13544 31872
rect 12207 31841 12219 31844
rect 12161 31835 12219 31841
rect 13538 31832 13544 31844
rect 13596 31832 13602 31884
rect 13814 31832 13820 31884
rect 13872 31872 13878 31884
rect 14277 31875 14335 31881
rect 14277 31872 14289 31875
rect 13872 31844 14289 31872
rect 13872 31832 13878 31844
rect 14277 31841 14289 31844
rect 14323 31841 14335 31875
rect 14277 31835 14335 31841
rect 14553 31875 14611 31881
rect 14553 31841 14565 31875
rect 14599 31872 14611 31875
rect 15028 31872 15056 31912
rect 15286 31900 15292 31912
rect 15344 31900 15350 31952
rect 15470 31900 15476 31952
rect 15528 31940 15534 31952
rect 16298 31940 16304 31952
rect 15528 31912 15976 31940
rect 15528 31900 15534 31912
rect 15948 31884 15976 31912
rect 16040 31912 16304 31940
rect 14599 31844 15056 31872
rect 14599 31841 14611 31844
rect 14553 31835 14611 31841
rect 11330 31804 11336 31816
rect 10520 31776 11336 31804
rect 11330 31764 11336 31776
rect 11388 31764 11394 31816
rect 12250 31764 12256 31816
rect 12308 31804 12314 31816
rect 13081 31807 13139 31813
rect 13081 31804 13093 31807
rect 12308 31776 13093 31804
rect 12308 31764 12314 31776
rect 13081 31773 13093 31776
rect 13127 31773 13139 31807
rect 13081 31767 13139 31773
rect 13633 31807 13691 31813
rect 13633 31773 13645 31807
rect 13679 31804 13691 31807
rect 13906 31804 13912 31816
rect 13679 31776 13912 31804
rect 13679 31773 13691 31776
rect 13633 31767 13691 31773
rect 8113 31739 8171 31745
rect 8113 31705 8125 31739
rect 8159 31705 8171 31739
rect 8113 31699 8171 31705
rect 8570 31696 8576 31748
rect 8628 31736 8634 31748
rect 12802 31736 12808 31748
rect 8628 31708 12808 31736
rect 8628 31696 8634 31708
rect 12802 31696 12808 31708
rect 12860 31696 12866 31748
rect 4341 31671 4399 31677
rect 4341 31637 4353 31671
rect 4387 31668 4399 31671
rect 4982 31668 4988 31680
rect 4387 31640 4988 31668
rect 4387 31637 4399 31640
rect 4341 31631 4399 31637
rect 4982 31628 4988 31640
rect 5040 31628 5046 31680
rect 7098 31628 7104 31680
rect 7156 31668 7162 31680
rect 7285 31671 7343 31677
rect 7285 31668 7297 31671
rect 7156 31640 7297 31668
rect 7156 31628 7162 31640
rect 7285 31637 7297 31640
rect 7331 31637 7343 31671
rect 8294 31668 8300 31680
rect 8255 31640 8300 31668
rect 7285 31631 7343 31637
rect 8294 31628 8300 31640
rect 8352 31628 8358 31680
rect 10318 31628 10324 31680
rect 10376 31668 10382 31680
rect 11146 31668 11152 31680
rect 10376 31640 11152 31668
rect 10376 31628 10382 31640
rect 11146 31628 11152 31640
rect 11204 31628 11210 31680
rect 12345 31671 12403 31677
rect 12345 31637 12357 31671
rect 12391 31668 12403 31671
rect 12710 31668 12716 31680
rect 12391 31640 12716 31668
rect 12391 31637 12403 31640
rect 12345 31631 12403 31637
rect 12710 31628 12716 31640
rect 12768 31628 12774 31680
rect 13096 31668 13124 31767
rect 13906 31764 13912 31776
rect 13964 31764 13970 31816
rect 14185 31807 14243 31813
rect 14185 31773 14197 31807
rect 14231 31804 14243 31807
rect 14568 31804 14596 31835
rect 15102 31832 15108 31884
rect 15160 31872 15166 31884
rect 15795 31875 15853 31881
rect 15795 31872 15807 31875
rect 15160 31844 15205 31872
rect 15304 31844 15807 31872
rect 15160 31832 15166 31844
rect 14231 31776 14596 31804
rect 14231 31773 14243 31776
rect 14185 31767 14243 31773
rect 14185 31671 14243 31677
rect 14185 31668 14197 31671
rect 13096 31640 14197 31668
rect 14185 31637 14197 31640
rect 14231 31637 14243 31671
rect 14185 31631 14243 31637
rect 14550 31628 14556 31680
rect 14608 31668 14614 31680
rect 15304 31668 15332 31844
rect 15795 31841 15807 31844
rect 15841 31841 15853 31875
rect 15930 31872 15936 31884
rect 15891 31844 15936 31872
rect 15795 31835 15853 31841
rect 15810 31804 15838 31835
rect 15930 31832 15936 31844
rect 15988 31832 15994 31884
rect 16040 31881 16068 31912
rect 16298 31900 16304 31912
rect 16356 31900 16362 31952
rect 18782 31900 18788 31952
rect 18840 31940 18846 31952
rect 22554 31940 22560 31952
rect 18840 31912 22560 31940
rect 18840 31900 18846 31912
rect 22554 31900 22560 31912
rect 22612 31900 22618 31952
rect 16025 31875 16083 31881
rect 16025 31841 16037 31875
rect 16071 31841 16083 31875
rect 16025 31835 16083 31841
rect 16209 31875 16267 31881
rect 16209 31841 16221 31875
rect 16255 31872 16267 31875
rect 16482 31872 16488 31884
rect 16255 31844 16488 31872
rect 16255 31841 16267 31844
rect 16209 31835 16267 31841
rect 16482 31832 16488 31844
rect 16540 31832 16546 31884
rect 17313 31875 17371 31881
rect 17313 31841 17325 31875
rect 17359 31872 17371 31875
rect 17402 31872 17408 31884
rect 17359 31844 17408 31872
rect 17359 31841 17371 31844
rect 17313 31835 17371 31841
rect 17402 31832 17408 31844
rect 17460 31832 17466 31884
rect 17497 31875 17555 31881
rect 17497 31841 17509 31875
rect 17543 31841 17555 31875
rect 17497 31835 17555 31841
rect 17589 31875 17647 31881
rect 17589 31841 17601 31875
rect 17635 31841 17647 31875
rect 17589 31835 17647 31841
rect 17681 31875 17739 31881
rect 17681 31841 17693 31875
rect 17727 31872 17739 31875
rect 17770 31872 17776 31884
rect 17727 31844 17776 31872
rect 17727 31841 17739 31844
rect 17681 31835 17739 31841
rect 16574 31804 16580 31816
rect 15810 31776 16580 31804
rect 16574 31764 16580 31776
rect 16632 31764 16638 31816
rect 17034 31764 17040 31816
rect 17092 31804 17098 31816
rect 17512 31804 17540 31835
rect 17092 31776 17540 31804
rect 17092 31764 17098 31776
rect 17494 31696 17500 31748
rect 17552 31736 17558 31748
rect 17604 31736 17632 31835
rect 17770 31832 17776 31844
rect 17828 31832 17834 31884
rect 18506 31872 18512 31884
rect 18467 31844 18512 31872
rect 18506 31832 18512 31844
rect 18564 31832 18570 31884
rect 19150 31872 19156 31884
rect 18892 31844 19156 31872
rect 18598 31804 18604 31816
rect 18559 31776 18604 31804
rect 18598 31764 18604 31776
rect 18656 31764 18662 31816
rect 18693 31807 18751 31813
rect 18693 31773 18705 31807
rect 18739 31773 18751 31807
rect 18693 31767 18751 31773
rect 18785 31807 18843 31813
rect 18785 31773 18797 31807
rect 18831 31804 18843 31807
rect 18892 31804 18920 31844
rect 19150 31832 19156 31844
rect 19208 31832 19214 31884
rect 20438 31832 20444 31884
rect 20496 31872 20502 31884
rect 21174 31872 21180 31884
rect 20496 31844 21180 31872
rect 20496 31832 20502 31844
rect 21174 31832 21180 31844
rect 21232 31881 21238 31884
rect 21232 31875 21291 31881
rect 21232 31841 21245 31875
rect 21279 31841 21291 31875
rect 21358 31872 21364 31884
rect 21319 31844 21364 31872
rect 21232 31835 21291 31841
rect 21232 31832 21238 31835
rect 21358 31832 21364 31844
rect 21416 31832 21422 31884
rect 21453 31875 21511 31881
rect 21453 31841 21465 31875
rect 21499 31872 21511 31875
rect 22186 31872 22192 31884
rect 21499 31844 22192 31872
rect 21499 31841 21511 31844
rect 21453 31835 21511 31841
rect 22186 31832 22192 31844
rect 22244 31872 22250 31884
rect 22738 31872 22744 31884
rect 22244 31844 22744 31872
rect 22244 31832 22250 31844
rect 22738 31832 22744 31844
rect 22796 31832 22802 31884
rect 22940 31881 22968 31980
rect 23106 31968 23112 32020
rect 23164 32008 23170 32020
rect 24026 32008 24032 32020
rect 23164 31980 24032 32008
rect 23164 31968 23170 31980
rect 24026 31968 24032 31980
rect 24084 31968 24090 32020
rect 24121 32011 24179 32017
rect 24121 31977 24133 32011
rect 24167 31977 24179 32011
rect 24121 31971 24179 31977
rect 24136 31940 24164 31971
rect 24762 31968 24768 32020
rect 24820 32008 24826 32020
rect 24949 32011 25007 32017
rect 24949 32008 24961 32011
rect 24820 31980 24961 32008
rect 24820 31968 24826 31980
rect 24949 31977 24961 31980
rect 24995 31977 25007 32011
rect 24949 31971 25007 31977
rect 25961 32011 26019 32017
rect 25961 31977 25973 32011
rect 26007 32008 26019 32011
rect 26602 32008 26608 32020
rect 26007 31980 26608 32008
rect 26007 31977 26019 31980
rect 25961 31971 26019 31977
rect 26602 31968 26608 31980
rect 26660 31968 26666 32020
rect 27893 31943 27951 31949
rect 27893 31940 27905 31943
rect 24136 31912 27905 31940
rect 27893 31909 27905 31912
rect 27939 31909 27951 31943
rect 27893 31903 27951 31909
rect 22925 31875 22983 31881
rect 22925 31841 22937 31875
rect 22971 31841 22983 31875
rect 22925 31835 22983 31841
rect 23017 31875 23075 31881
rect 23017 31841 23029 31875
rect 23063 31841 23075 31875
rect 23017 31835 23075 31841
rect 23109 31875 23167 31881
rect 23109 31841 23121 31875
rect 23155 31872 23167 31875
rect 23566 31872 23572 31884
rect 23155 31844 23572 31872
rect 23155 31841 23167 31844
rect 23109 31835 23167 31841
rect 18831 31776 18920 31804
rect 18831 31773 18843 31776
rect 18785 31767 18843 31773
rect 17552 31708 17632 31736
rect 17552 31696 17558 31708
rect 15562 31668 15568 31680
rect 14608 31640 15332 31668
rect 15523 31640 15568 31668
rect 14608 31628 14614 31640
rect 15562 31628 15568 31640
rect 15620 31628 15626 31680
rect 17862 31668 17868 31680
rect 17823 31640 17868 31668
rect 17862 31628 17868 31640
rect 17920 31628 17926 31680
rect 18598 31628 18604 31680
rect 18656 31668 18662 31680
rect 18708 31668 18736 31767
rect 18966 31764 18972 31816
rect 19024 31804 19030 31816
rect 21082 31804 21088 31816
rect 19024 31776 21088 31804
rect 19024 31764 19030 31776
rect 21082 31764 21088 31776
rect 21140 31764 21146 31816
rect 21376 31804 21404 31832
rect 23032 31804 23060 31835
rect 23566 31832 23572 31844
rect 23624 31872 23630 31884
rect 23750 31872 23756 31884
rect 23624 31844 23756 31872
rect 23624 31832 23630 31844
rect 23750 31832 23756 31844
rect 23808 31832 23814 31884
rect 24305 31875 24363 31881
rect 24305 31841 24317 31875
rect 24351 31841 24363 31875
rect 24305 31835 24363 31841
rect 23290 31804 23296 31816
rect 21376 31776 23296 31804
rect 23290 31764 23296 31776
rect 23348 31764 23354 31816
rect 24320 31804 24348 31835
rect 24394 31832 24400 31884
rect 24452 31872 24458 31884
rect 24857 31875 24915 31881
rect 24857 31872 24869 31875
rect 24452 31844 24869 31872
rect 24452 31832 24458 31844
rect 24857 31841 24869 31844
rect 24903 31841 24915 31875
rect 25222 31872 25228 31884
rect 24857 31835 24915 31841
rect 24964 31844 25228 31872
rect 24964 31804 24992 31844
rect 25222 31832 25228 31844
rect 25280 31832 25286 31884
rect 26142 31872 26148 31884
rect 26103 31844 26148 31872
rect 26142 31832 26148 31844
rect 26200 31832 26206 31884
rect 26510 31832 26516 31884
rect 26568 31872 26574 31884
rect 26697 31875 26755 31881
rect 26697 31872 26709 31875
rect 26568 31844 26709 31872
rect 26568 31832 26574 31844
rect 26697 31841 26709 31844
rect 26743 31841 26755 31875
rect 26697 31835 26755 31841
rect 24320 31776 24992 31804
rect 22462 31696 22468 31748
rect 22520 31736 22526 31748
rect 23934 31736 23940 31748
rect 22520 31708 23940 31736
rect 22520 31696 22526 31708
rect 23934 31696 23940 31708
rect 23992 31696 23998 31748
rect 18656 31640 18736 31668
rect 18656 31628 18662 31640
rect 18874 31628 18880 31680
rect 18932 31668 18938 31680
rect 21266 31668 21272 31680
rect 18932 31640 21272 31668
rect 18932 31628 18938 31640
rect 21266 31628 21272 31640
rect 21324 31628 21330 31680
rect 21634 31668 21640 31680
rect 21595 31640 21640 31668
rect 21634 31628 21640 31640
rect 21692 31628 21698 31680
rect 21726 31628 21732 31680
rect 21784 31668 21790 31680
rect 22094 31668 22100 31680
rect 21784 31640 22100 31668
rect 21784 31628 21790 31640
rect 22094 31628 22100 31640
rect 22152 31668 22158 31680
rect 22646 31668 22652 31680
rect 22152 31640 22652 31668
rect 22152 31628 22158 31640
rect 22646 31628 22652 31640
rect 22704 31628 22710 31680
rect 22741 31671 22799 31677
rect 22741 31637 22753 31671
rect 22787 31668 22799 31671
rect 22922 31668 22928 31680
rect 22787 31640 22928 31668
rect 22787 31637 22799 31640
rect 22741 31631 22799 31637
rect 22922 31628 22928 31640
rect 22980 31628 22986 31680
rect 23293 31671 23351 31677
rect 23293 31637 23305 31671
rect 23339 31668 23351 31671
rect 23382 31668 23388 31680
rect 23339 31640 23388 31668
rect 23339 31637 23351 31640
rect 23293 31631 23351 31637
rect 23382 31628 23388 31640
rect 23440 31628 23446 31680
rect 23842 31628 23848 31680
rect 23900 31668 23906 31680
rect 26789 31671 26847 31677
rect 26789 31668 26801 31671
rect 23900 31640 26801 31668
rect 23900 31628 23906 31640
rect 26789 31637 26801 31640
rect 26835 31637 26847 31671
rect 27982 31668 27988 31680
rect 27943 31640 27988 31668
rect 26789 31631 26847 31637
rect 27982 31628 27988 31640
rect 28040 31628 28046 31680
rect 1104 31578 28888 31600
rect 1104 31526 5614 31578
rect 5666 31526 5678 31578
rect 5730 31526 5742 31578
rect 5794 31526 5806 31578
rect 5858 31526 14878 31578
rect 14930 31526 14942 31578
rect 14994 31526 15006 31578
rect 15058 31526 15070 31578
rect 15122 31526 24142 31578
rect 24194 31526 24206 31578
rect 24258 31526 24270 31578
rect 24322 31526 24334 31578
rect 24386 31526 28888 31578
rect 1104 31504 28888 31526
rect 1394 31424 1400 31476
rect 1452 31464 1458 31476
rect 2593 31467 2651 31473
rect 2593 31464 2605 31467
rect 1452 31436 2605 31464
rect 1452 31424 1458 31436
rect 2593 31433 2605 31436
rect 2639 31433 2651 31467
rect 2593 31427 2651 31433
rect 4246 31424 4252 31476
rect 4304 31464 4310 31476
rect 4709 31467 4767 31473
rect 4709 31464 4721 31467
rect 4304 31436 4721 31464
rect 4304 31424 4310 31436
rect 4709 31433 4721 31436
rect 4755 31433 4767 31467
rect 6362 31464 6368 31476
rect 6323 31436 6368 31464
rect 4709 31427 4767 31433
rect 6362 31424 6368 31436
rect 6420 31424 6426 31476
rect 8570 31464 8576 31476
rect 7116 31436 8576 31464
rect 2498 31396 2504 31408
rect 2459 31368 2504 31396
rect 2498 31356 2504 31368
rect 2556 31356 2562 31408
rect 4617 31399 4675 31405
rect 4617 31365 4629 31399
rect 4663 31396 4675 31399
rect 4982 31396 4988 31408
rect 4663 31368 4988 31396
rect 4663 31365 4675 31368
rect 4617 31359 4675 31365
rect 4982 31356 4988 31368
rect 5040 31356 5046 31408
rect 7116 31396 7144 31436
rect 8570 31424 8576 31436
rect 8628 31424 8634 31476
rect 8662 31424 8668 31476
rect 8720 31464 8726 31476
rect 22189 31467 22247 31473
rect 8720 31436 22094 31464
rect 8720 31424 8726 31436
rect 7282 31396 7288 31408
rect 5644 31368 7144 31396
rect 7243 31368 7288 31396
rect 5644 31328 5672 31368
rect 7282 31356 7288 31368
rect 7340 31356 7346 31408
rect 10870 31356 10876 31408
rect 10928 31396 10934 31408
rect 11149 31399 11207 31405
rect 11149 31396 11161 31399
rect 10928 31368 11161 31396
rect 10928 31356 10934 31368
rect 11149 31365 11161 31368
rect 11195 31365 11207 31399
rect 11149 31359 11207 31365
rect 12434 31356 12440 31408
rect 12492 31396 12498 31408
rect 14550 31396 14556 31408
rect 12492 31368 14556 31396
rect 12492 31356 12498 31368
rect 14550 31356 14556 31368
rect 14608 31356 14614 31408
rect 16574 31356 16580 31408
rect 16632 31396 16638 31408
rect 16761 31399 16819 31405
rect 16761 31396 16773 31399
rect 16632 31368 16773 31396
rect 16632 31356 16638 31368
rect 16761 31365 16773 31368
rect 16807 31365 16819 31399
rect 21726 31396 21732 31408
rect 16761 31359 16819 31365
rect 21008 31368 21732 31396
rect 3160 31300 5672 31328
rect 5721 31331 5779 31337
rect 1489 31263 1547 31269
rect 1489 31229 1501 31263
rect 1535 31260 1547 31263
rect 2682 31260 2688 31272
rect 1535 31232 2688 31260
rect 1535 31229 1547 31232
rect 1489 31223 1547 31229
rect 2682 31220 2688 31232
rect 2740 31220 2746 31272
rect 3160 31269 3188 31300
rect 5721 31297 5733 31331
rect 5767 31328 5779 31331
rect 7190 31328 7196 31340
rect 5767 31300 7196 31328
rect 5767 31297 5779 31300
rect 5721 31291 5779 31297
rect 7190 31288 7196 31300
rect 7248 31288 7254 31340
rect 7377 31331 7435 31337
rect 7377 31297 7389 31331
rect 7423 31328 7435 31331
rect 10045 31331 10103 31337
rect 7423 31300 7880 31328
rect 7423 31297 7435 31300
rect 7377 31291 7435 31297
rect 3145 31263 3203 31269
rect 3145 31229 3157 31263
rect 3191 31229 3203 31263
rect 3145 31223 3203 31229
rect 4154 31220 4160 31272
rect 4212 31260 4218 31272
rect 4249 31263 4307 31269
rect 4249 31260 4261 31263
rect 4212 31232 4261 31260
rect 4212 31220 4218 31232
rect 4249 31229 4261 31232
rect 4295 31260 4307 31263
rect 4522 31260 4528 31272
rect 4295 31232 4528 31260
rect 4295 31229 4307 31232
rect 4249 31223 4307 31229
rect 4522 31220 4528 31232
rect 4580 31220 4586 31272
rect 5629 31263 5687 31269
rect 5629 31229 5641 31263
rect 5675 31260 5687 31263
rect 5902 31260 5908 31272
rect 5675 31232 5908 31260
rect 5675 31229 5687 31232
rect 5629 31223 5687 31229
rect 5902 31220 5908 31232
rect 5960 31220 5966 31272
rect 6273 31263 6331 31269
rect 6273 31229 6285 31263
rect 6319 31260 6331 31263
rect 6362 31260 6368 31272
rect 6319 31232 6368 31260
rect 6319 31229 6331 31232
rect 6273 31223 6331 31229
rect 6362 31220 6368 31232
rect 6420 31220 6426 31272
rect 7852 31269 7880 31300
rect 10045 31297 10057 31331
rect 10091 31328 10103 31331
rect 10686 31328 10692 31340
rect 10091 31300 10692 31328
rect 10091 31297 10103 31300
rect 10045 31291 10103 31297
rect 10686 31288 10692 31300
rect 10744 31288 10750 31340
rect 14182 31328 14188 31340
rect 12544 31300 14188 31328
rect 7837 31263 7895 31269
rect 7837 31229 7849 31263
rect 7883 31229 7895 31263
rect 7837 31223 7895 31229
rect 9769 31263 9827 31269
rect 9769 31229 9781 31263
rect 9815 31260 9827 31263
rect 11514 31260 11520 31272
rect 9815 31232 11520 31260
rect 9815 31229 9827 31232
rect 9769 31223 9827 31229
rect 11514 31220 11520 31232
rect 11572 31220 11578 31272
rect 11882 31260 11888 31272
rect 11843 31232 11888 31260
rect 11882 31220 11888 31232
rect 11940 31220 11946 31272
rect 12544 31269 12572 31300
rect 14182 31288 14188 31300
rect 14240 31288 14246 31340
rect 18506 31328 18512 31340
rect 17604 31300 18512 31328
rect 12253 31263 12311 31269
rect 12253 31229 12265 31263
rect 12299 31229 12311 31263
rect 12253 31223 12311 31229
rect 12529 31263 12587 31269
rect 12529 31229 12541 31263
rect 12575 31229 12587 31263
rect 12529 31223 12587 31229
rect 2130 31192 2136 31204
rect 2091 31164 2136 31192
rect 2130 31152 2136 31164
rect 2188 31152 2194 31204
rect 6917 31195 6975 31201
rect 6917 31161 6929 31195
rect 6963 31192 6975 31195
rect 7006 31192 7012 31204
rect 6963 31164 7012 31192
rect 6963 31161 6975 31164
rect 6917 31155 6975 31161
rect 7006 31152 7012 31164
rect 7064 31192 7070 31204
rect 7282 31192 7288 31204
rect 7064 31164 7288 31192
rect 7064 31152 7070 31164
rect 7282 31152 7288 31164
rect 7340 31152 7346 31204
rect 11974 31192 11980 31204
rect 7392 31164 8064 31192
rect 11935 31164 11980 31192
rect 1394 31084 1400 31136
rect 1452 31124 1458 31136
rect 1581 31127 1639 31133
rect 1581 31124 1593 31127
rect 1452 31096 1593 31124
rect 1452 31084 1458 31096
rect 1581 31093 1593 31096
rect 1627 31093 1639 31127
rect 3234 31124 3240 31136
rect 3195 31096 3240 31124
rect 1581 31087 1639 31093
rect 3234 31084 3240 31096
rect 3292 31084 3298 31136
rect 3326 31084 3332 31136
rect 3384 31124 3390 31136
rect 7392 31124 7420 31164
rect 7926 31124 7932 31136
rect 3384 31096 7420 31124
rect 7887 31096 7932 31124
rect 3384 31084 3390 31096
rect 7926 31084 7932 31096
rect 7984 31084 7990 31136
rect 8036 31124 8064 31164
rect 11974 31152 11980 31164
rect 12032 31152 12038 31204
rect 12268 31192 12296 31223
rect 12710 31220 12716 31272
rect 12768 31260 12774 31272
rect 12989 31263 13047 31269
rect 12989 31260 13001 31263
rect 12768 31232 13001 31260
rect 12768 31220 12774 31232
rect 12989 31229 13001 31232
rect 13035 31260 13047 31263
rect 13170 31260 13176 31272
rect 13035 31232 13176 31260
rect 13035 31229 13047 31232
rect 12989 31223 13047 31229
rect 13170 31220 13176 31232
rect 13228 31220 13234 31272
rect 15381 31263 15439 31269
rect 15381 31229 15393 31263
rect 15427 31229 15439 31263
rect 15381 31223 15439 31229
rect 15396 31192 15424 31223
rect 15470 31220 15476 31272
rect 15528 31260 15534 31272
rect 15637 31263 15695 31269
rect 15637 31260 15649 31263
rect 15528 31232 15649 31260
rect 15528 31220 15534 31232
rect 15637 31229 15649 31232
rect 15683 31229 15695 31263
rect 15637 31223 15695 31229
rect 16022 31220 16028 31272
rect 16080 31260 16086 31272
rect 17313 31263 17371 31269
rect 17313 31260 17325 31263
rect 16080 31232 17325 31260
rect 16080 31220 16086 31232
rect 17313 31229 17325 31232
rect 17359 31229 17371 31263
rect 17313 31223 17371 31229
rect 17402 31220 17408 31272
rect 17460 31260 17466 31272
rect 17604 31269 17632 31300
rect 18506 31288 18512 31300
rect 18564 31288 18570 31340
rect 19981 31331 20039 31337
rect 19981 31297 19993 31331
rect 20027 31328 20039 31331
rect 21008 31328 21036 31368
rect 21726 31356 21732 31368
rect 21784 31356 21790 31408
rect 22066 31396 22094 31436
rect 22189 31433 22201 31467
rect 22235 31464 22247 31467
rect 22830 31464 22836 31476
rect 22235 31436 22836 31464
rect 22235 31433 22247 31436
rect 22189 31427 22247 31433
rect 22830 31424 22836 31436
rect 22888 31424 22894 31476
rect 27525 31467 27583 31473
rect 27525 31464 27537 31467
rect 22940 31436 27537 31464
rect 22940 31396 22968 31436
rect 27525 31433 27537 31436
rect 27571 31433 27583 31467
rect 27525 31427 27583 31433
rect 22066 31368 22968 31396
rect 24118 31356 24124 31408
rect 24176 31396 24182 31408
rect 24762 31396 24768 31408
rect 24176 31368 24768 31396
rect 24176 31356 24182 31368
rect 24762 31356 24768 31368
rect 24820 31356 24826 31408
rect 20027 31300 21036 31328
rect 21361 31331 21419 31337
rect 20027 31297 20039 31300
rect 19981 31291 20039 31297
rect 21361 31297 21373 31331
rect 21407 31297 21419 31331
rect 21361 31291 21419 31297
rect 17589 31263 17647 31269
rect 17589 31260 17601 31263
rect 17460 31232 17601 31260
rect 17460 31220 17466 31232
rect 17589 31229 17601 31232
rect 17635 31229 17647 31263
rect 17589 31223 17647 31229
rect 18322 31220 18328 31272
rect 18380 31260 18386 31272
rect 18877 31263 18935 31269
rect 18877 31260 18889 31263
rect 18380 31232 18889 31260
rect 18380 31220 18386 31232
rect 18877 31229 18889 31232
rect 18923 31260 18935 31263
rect 18966 31260 18972 31272
rect 18923 31232 18972 31260
rect 18923 31229 18935 31232
rect 18877 31223 18935 31229
rect 18966 31220 18972 31232
rect 19024 31220 19030 31272
rect 20254 31260 20260 31272
rect 20215 31232 20260 31260
rect 20254 31220 20260 31232
rect 20312 31220 20318 31272
rect 20530 31220 20536 31272
rect 20588 31260 20594 31272
rect 21376 31260 21404 31291
rect 21634 31288 21640 31340
rect 21692 31328 21698 31340
rect 23661 31331 23719 31337
rect 21692 31300 22876 31328
rect 21692 31288 21698 31300
rect 22462 31260 22468 31272
rect 20588 31232 21404 31260
rect 22423 31232 22468 31260
rect 20588 31220 20594 31232
rect 22462 31220 22468 31232
rect 22520 31220 22526 31272
rect 22557 31263 22615 31269
rect 22557 31229 22569 31263
rect 22603 31229 22615 31263
rect 22557 31223 22615 31229
rect 15838 31192 15844 31204
rect 12268 31164 12756 31192
rect 15396 31164 15844 31192
rect 12728 31136 12756 31164
rect 15838 31152 15844 31164
rect 15896 31152 15902 31204
rect 21910 31152 21916 31204
rect 21968 31192 21974 31204
rect 22572 31192 22600 31223
rect 22646 31220 22652 31272
rect 22704 31260 22710 31272
rect 22848 31269 22876 31300
rect 23661 31297 23673 31331
rect 23707 31328 23719 31331
rect 25501 31331 25559 31337
rect 25501 31328 25513 31331
rect 23707 31300 25513 31328
rect 23707 31297 23719 31300
rect 23661 31291 23719 31297
rect 25501 31297 25513 31300
rect 25547 31297 25559 31331
rect 25501 31291 25559 31297
rect 22833 31263 22891 31269
rect 22704 31232 22749 31260
rect 22704 31220 22710 31232
rect 22833 31229 22845 31263
rect 22879 31229 22891 31263
rect 23934 31260 23940 31272
rect 23895 31232 23940 31260
rect 22833 31223 22891 31229
rect 23934 31220 23940 31232
rect 23992 31220 23998 31272
rect 24029 31263 24087 31269
rect 24029 31229 24041 31263
rect 24075 31229 24087 31263
rect 24029 31223 24087 31229
rect 24044 31192 24072 31223
rect 24118 31220 24124 31272
rect 24176 31260 24182 31272
rect 24305 31263 24363 31269
rect 24176 31232 24221 31260
rect 24176 31220 24182 31232
rect 24305 31229 24317 31263
rect 24351 31229 24363 31263
rect 25222 31260 25228 31272
rect 25183 31232 25228 31260
rect 24305 31223 24363 31229
rect 21968 31164 24072 31192
rect 21968 31152 21974 31164
rect 10870 31124 10876 31136
rect 8036 31096 10876 31124
rect 10870 31084 10876 31096
rect 10928 31084 10934 31136
rect 12158 31084 12164 31136
rect 12216 31124 12222 31136
rect 12434 31124 12440 31136
rect 12216 31096 12440 31124
rect 12216 31084 12222 31096
rect 12434 31084 12440 31096
rect 12492 31084 12498 31136
rect 12710 31084 12716 31136
rect 12768 31124 12774 31136
rect 13173 31127 13231 31133
rect 13173 31124 13185 31127
rect 12768 31096 13185 31124
rect 12768 31084 12774 31096
rect 13173 31093 13185 31096
rect 13219 31124 13231 31127
rect 13814 31124 13820 31136
rect 13219 31096 13820 31124
rect 13219 31093 13231 31096
rect 13173 31087 13231 31093
rect 13814 31084 13820 31096
rect 13872 31084 13878 31136
rect 14182 31084 14188 31136
rect 14240 31124 14246 31136
rect 18506 31124 18512 31136
rect 14240 31096 18512 31124
rect 14240 31084 14246 31096
rect 18506 31084 18512 31096
rect 18564 31084 18570 31136
rect 18966 31124 18972 31136
rect 18879 31096 18972 31124
rect 18966 31084 18972 31096
rect 19024 31124 19030 31136
rect 21358 31124 21364 31136
rect 19024 31096 21364 31124
rect 19024 31084 19030 31096
rect 21358 31084 21364 31096
rect 21416 31084 21422 31136
rect 24026 31084 24032 31136
rect 24084 31124 24090 31136
rect 24320 31124 24348 31223
rect 25222 31220 25228 31232
rect 25280 31260 25286 31272
rect 25774 31260 25780 31272
rect 25280 31232 25780 31260
rect 25280 31220 25286 31232
rect 25774 31220 25780 31232
rect 25832 31220 25838 31272
rect 26326 31152 26332 31204
rect 26384 31192 26390 31204
rect 27433 31195 27491 31201
rect 27433 31192 27445 31195
rect 26384 31164 27445 31192
rect 26384 31152 26390 31164
rect 27433 31161 27445 31164
rect 27479 31161 27491 31195
rect 27433 31155 27491 31161
rect 24084 31096 24348 31124
rect 24084 31084 24090 31096
rect 25866 31084 25872 31136
rect 25924 31124 25930 31136
rect 26605 31127 26663 31133
rect 26605 31124 26617 31127
rect 25924 31096 26617 31124
rect 25924 31084 25930 31096
rect 26605 31093 26617 31096
rect 26651 31093 26663 31127
rect 26605 31087 26663 31093
rect 1104 31034 28888 31056
rect 1104 30982 10246 31034
rect 10298 30982 10310 31034
rect 10362 30982 10374 31034
rect 10426 30982 10438 31034
rect 10490 30982 19510 31034
rect 19562 30982 19574 31034
rect 19626 30982 19638 31034
rect 19690 30982 19702 31034
rect 19754 30982 28888 31034
rect 1104 30960 28888 30982
rect 3786 30880 3792 30932
rect 3844 30920 3850 30932
rect 4709 30923 4767 30929
rect 4709 30920 4721 30923
rect 3844 30892 4721 30920
rect 3844 30880 3850 30892
rect 4709 30889 4721 30892
rect 4755 30889 4767 30923
rect 27982 30920 27988 30932
rect 4709 30883 4767 30889
rect 5368 30892 27988 30920
rect 5368 30861 5396 30892
rect 27982 30880 27988 30892
rect 28040 30880 28046 30932
rect 5353 30855 5411 30861
rect 5353 30821 5365 30855
rect 5399 30821 5411 30855
rect 8662 30852 8668 30864
rect 5353 30815 5411 30821
rect 7208 30824 8668 30852
rect 1854 30784 1860 30796
rect 1815 30756 1860 30784
rect 1854 30744 1860 30756
rect 1912 30744 1918 30796
rect 2590 30784 2596 30796
rect 2551 30756 2596 30784
rect 2590 30744 2596 30756
rect 2648 30744 2654 30796
rect 3510 30744 3516 30796
rect 3568 30784 3574 30796
rect 3789 30787 3847 30793
rect 3789 30784 3801 30787
rect 3568 30756 3801 30784
rect 3568 30744 3574 30756
rect 3789 30753 3801 30756
rect 3835 30753 3847 30787
rect 3789 30747 3847 30753
rect 4617 30787 4675 30793
rect 4617 30753 4629 30787
rect 4663 30784 4675 30787
rect 7208 30784 7236 30824
rect 8662 30812 8668 30824
rect 8720 30812 8726 30864
rect 10042 30812 10048 30864
rect 10100 30852 10106 30864
rect 11054 30852 11060 30864
rect 10100 30824 11060 30852
rect 10100 30812 10106 30824
rect 11054 30812 11060 30824
rect 11112 30812 11118 30864
rect 11330 30812 11336 30864
rect 11388 30852 11394 30864
rect 15565 30855 15623 30861
rect 11388 30824 15332 30852
rect 11388 30812 11394 30824
rect 7558 30784 7564 30796
rect 4663 30756 7236 30784
rect 7519 30756 7564 30784
rect 4663 30753 4675 30756
rect 4617 30747 4675 30753
rect 7558 30744 7564 30756
rect 7616 30744 7622 30796
rect 7926 30784 7932 30796
rect 7887 30756 7932 30784
rect 7926 30744 7932 30756
rect 7984 30744 7990 30796
rect 8021 30787 8079 30793
rect 8021 30753 8033 30787
rect 8067 30753 8079 30787
rect 8021 30747 8079 30753
rect 1946 30676 1952 30728
rect 2004 30716 2010 30728
rect 3234 30716 3240 30728
rect 2004 30688 3240 30716
rect 2004 30676 2010 30688
rect 3234 30676 3240 30688
rect 3292 30676 3298 30728
rect 4062 30676 4068 30728
rect 4120 30716 4126 30728
rect 5537 30719 5595 30725
rect 5537 30716 5549 30719
rect 4120 30688 5549 30716
rect 4120 30676 4126 30688
rect 5537 30685 5549 30688
rect 5583 30685 5595 30719
rect 5537 30679 5595 30685
rect 7466 30676 7472 30728
rect 7524 30716 7530 30728
rect 8036 30716 8064 30747
rect 8294 30744 8300 30796
rect 8352 30784 8358 30796
rect 8389 30787 8447 30793
rect 8389 30784 8401 30787
rect 8352 30756 8401 30784
rect 8352 30744 8358 30756
rect 8389 30753 8401 30756
rect 8435 30753 8447 30787
rect 8389 30747 8447 30753
rect 12161 30787 12219 30793
rect 12161 30753 12173 30787
rect 12207 30784 12219 30787
rect 12250 30784 12256 30796
rect 12207 30756 12256 30784
rect 12207 30753 12219 30756
rect 12161 30747 12219 30753
rect 12250 30744 12256 30756
rect 12308 30744 12314 30796
rect 12345 30787 12403 30793
rect 12345 30753 12357 30787
rect 12391 30753 12403 30787
rect 12345 30747 12403 30753
rect 7524 30688 8064 30716
rect 12360 30716 12388 30747
rect 12434 30744 12440 30796
rect 12492 30784 12498 30796
rect 13725 30787 13783 30793
rect 12492 30756 12537 30784
rect 12492 30744 12498 30756
rect 13725 30753 13737 30787
rect 13771 30753 13783 30787
rect 13906 30784 13912 30796
rect 13867 30756 13912 30784
rect 13725 30747 13783 30753
rect 12710 30716 12716 30728
rect 12360 30688 12716 30716
rect 7524 30676 7530 30688
rect 12710 30676 12716 30688
rect 12768 30676 12774 30728
rect 2774 30608 2780 30660
rect 2832 30648 2838 30660
rect 8665 30651 8723 30657
rect 2832 30620 2877 30648
rect 2832 30608 2838 30620
rect 8665 30617 8677 30651
rect 8711 30648 8723 30651
rect 8938 30648 8944 30660
rect 8711 30620 8944 30648
rect 8711 30617 8723 30620
rect 8665 30611 8723 30617
rect 8938 30608 8944 30620
rect 8996 30608 9002 30660
rect 9950 30608 9956 30660
rect 10008 30648 10014 30660
rect 10686 30648 10692 30660
rect 10008 30620 10692 30648
rect 10008 30608 10014 30620
rect 10686 30608 10692 30620
rect 10744 30608 10750 30660
rect 11330 30608 11336 30660
rect 11388 30648 11394 30660
rect 11514 30648 11520 30660
rect 11388 30620 11520 30648
rect 11388 30608 11394 30620
rect 11514 30608 11520 30620
rect 11572 30608 11578 30660
rect 1946 30580 1952 30592
rect 1907 30552 1952 30580
rect 1946 30540 1952 30552
rect 2004 30540 2010 30592
rect 3878 30540 3884 30592
rect 3936 30580 3942 30592
rect 3973 30583 4031 30589
rect 3973 30580 3985 30583
rect 3936 30552 3985 30580
rect 3936 30540 3942 30552
rect 3973 30549 3985 30552
rect 4019 30580 4031 30583
rect 11882 30580 11888 30592
rect 4019 30552 11888 30580
rect 4019 30549 4031 30552
rect 3973 30543 4031 30549
rect 11882 30540 11888 30552
rect 11940 30540 11946 30592
rect 12434 30540 12440 30592
rect 12492 30580 12498 30592
rect 13740 30580 13768 30747
rect 13906 30744 13912 30756
rect 13964 30744 13970 30796
rect 14274 30784 14280 30796
rect 14235 30756 14280 30784
rect 14274 30744 14280 30756
rect 14332 30744 14338 30796
rect 14553 30787 14611 30793
rect 14553 30753 14565 30787
rect 14599 30784 14611 30787
rect 15102 30784 15108 30796
rect 14599 30756 15108 30784
rect 14599 30753 14611 30756
rect 14553 30747 14611 30753
rect 15102 30744 15108 30756
rect 15160 30744 15166 30796
rect 15304 30793 15332 30824
rect 15565 30821 15577 30855
rect 15611 30852 15623 30855
rect 16206 30852 16212 30864
rect 15611 30824 16212 30852
rect 15611 30821 15623 30824
rect 15565 30815 15623 30821
rect 16206 30812 16212 30824
rect 16264 30812 16270 30864
rect 18506 30852 18512 30864
rect 18467 30824 18512 30852
rect 18506 30812 18512 30824
rect 18564 30812 18570 30864
rect 19153 30855 19211 30861
rect 19153 30821 19165 30855
rect 19199 30852 19211 30855
rect 20254 30852 20260 30864
rect 19199 30824 20260 30852
rect 19199 30821 19211 30824
rect 19153 30815 19211 30821
rect 20254 30812 20260 30824
rect 20312 30812 20318 30864
rect 21358 30852 21364 30864
rect 20916 30824 21364 30852
rect 15197 30787 15255 30793
rect 15197 30753 15209 30787
rect 15243 30753 15255 30787
rect 15197 30747 15255 30753
rect 15289 30787 15347 30793
rect 15289 30753 15301 30787
rect 15335 30753 15347 30787
rect 15289 30747 15347 30753
rect 15381 30787 15439 30793
rect 15381 30753 15393 30787
rect 15427 30784 15439 30787
rect 15470 30784 15476 30796
rect 15427 30756 15476 30784
rect 15427 30753 15439 30756
rect 15381 30747 15439 30753
rect 15212 30648 15240 30747
rect 15470 30744 15476 30756
rect 15528 30744 15534 30796
rect 16114 30784 16120 30796
rect 16075 30756 16120 30784
rect 16114 30744 16120 30756
rect 16172 30744 16178 30796
rect 17402 30744 17408 30796
rect 17460 30784 17466 30796
rect 17497 30787 17555 30793
rect 17497 30784 17509 30787
rect 17460 30756 17509 30784
rect 17460 30744 17466 30756
rect 17497 30753 17509 30756
rect 17543 30753 17555 30787
rect 17497 30747 17555 30753
rect 17773 30787 17831 30793
rect 17773 30753 17785 30787
rect 17819 30784 17831 30787
rect 17862 30784 17868 30796
rect 17819 30756 17868 30784
rect 17819 30753 17831 30756
rect 17773 30747 17831 30753
rect 17862 30744 17868 30756
rect 17920 30744 17926 30796
rect 19426 30784 19432 30796
rect 19387 30756 19432 30784
rect 19426 30744 19432 30756
rect 19484 30744 19490 30796
rect 19521 30787 19579 30793
rect 19521 30753 19533 30787
rect 19567 30753 19579 30787
rect 19521 30747 19579 30753
rect 19613 30787 19671 30793
rect 19613 30753 19625 30787
rect 19659 30753 19671 30787
rect 19613 30747 19671 30753
rect 16666 30676 16672 30728
rect 16724 30716 16730 30728
rect 17313 30719 17371 30725
rect 17313 30716 17325 30719
rect 16724 30688 17325 30716
rect 16724 30676 16730 30688
rect 17313 30685 17325 30688
rect 17359 30685 17371 30719
rect 17313 30679 17371 30685
rect 17589 30719 17647 30725
rect 17589 30685 17601 30719
rect 17635 30685 17647 30719
rect 17589 30679 17647 30685
rect 17681 30719 17739 30725
rect 17681 30685 17693 30719
rect 17727 30716 17739 30719
rect 18693 30719 18751 30725
rect 17727 30688 17816 30716
rect 17727 30685 17739 30688
rect 17681 30679 17739 30685
rect 17402 30648 17408 30660
rect 15212 30620 17408 30648
rect 17402 30608 17408 30620
rect 17460 30608 17466 30660
rect 13814 30580 13820 30592
rect 12492 30552 12537 30580
rect 13740 30552 13820 30580
rect 12492 30540 12498 30552
rect 13814 30540 13820 30552
rect 13872 30540 13878 30592
rect 16022 30540 16028 30592
rect 16080 30580 16086 30592
rect 16209 30583 16267 30589
rect 16209 30580 16221 30583
rect 16080 30552 16221 30580
rect 16080 30540 16086 30552
rect 16209 30549 16221 30552
rect 16255 30549 16267 30583
rect 16209 30543 16267 30549
rect 16574 30540 16580 30592
rect 16632 30580 16638 30592
rect 17604 30580 17632 30679
rect 17788 30660 17816 30688
rect 18693 30685 18705 30719
rect 18739 30716 18751 30719
rect 19536 30716 19564 30747
rect 18739 30688 19564 30716
rect 19628 30716 19656 30747
rect 19702 30744 19708 30796
rect 19760 30784 19766 30796
rect 19797 30787 19855 30793
rect 19797 30784 19809 30787
rect 19760 30756 19809 30784
rect 19760 30744 19766 30756
rect 19797 30753 19809 30756
rect 19843 30753 19855 30787
rect 19797 30747 19855 30753
rect 20438 30744 20444 30796
rect 20496 30784 20502 30796
rect 20916 30793 20944 30824
rect 21358 30812 21364 30824
rect 21416 30812 21422 30864
rect 22833 30855 22891 30861
rect 22833 30821 22845 30855
rect 22879 30852 22891 30855
rect 22879 30824 23612 30852
rect 22879 30821 22891 30824
rect 22833 30815 22891 30821
rect 20809 30787 20867 30793
rect 20809 30784 20821 30787
rect 20496 30756 20821 30784
rect 20496 30744 20502 30756
rect 20809 30753 20821 30756
rect 20855 30753 20867 30787
rect 20809 30747 20867 30753
rect 20901 30787 20959 30793
rect 20901 30753 20913 30787
rect 20947 30753 20959 30787
rect 20901 30747 20959 30753
rect 20990 30744 20996 30796
rect 21048 30784 21054 30796
rect 21174 30784 21180 30796
rect 21048 30756 21180 30784
rect 21048 30744 21054 30756
rect 21174 30744 21180 30756
rect 21232 30744 21238 30796
rect 23014 30744 23020 30796
rect 23072 30784 23078 30796
rect 23109 30787 23167 30793
rect 23109 30784 23121 30787
rect 23072 30756 23121 30784
rect 23072 30744 23078 30756
rect 23109 30753 23121 30756
rect 23155 30753 23167 30787
rect 23109 30747 23167 30753
rect 23201 30787 23259 30793
rect 23201 30753 23213 30787
rect 23247 30753 23259 30787
rect 23201 30747 23259 30753
rect 23293 30787 23351 30793
rect 23293 30753 23305 30787
rect 23339 30753 23351 30787
rect 23293 30747 23351 30753
rect 20070 30716 20076 30728
rect 19628 30688 20076 30716
rect 18739 30685 18751 30688
rect 18693 30679 18751 30685
rect 17770 30608 17776 30660
rect 17828 30608 17834 30660
rect 19536 30648 19564 30688
rect 20070 30676 20076 30688
rect 20128 30676 20134 30728
rect 21910 30716 21916 30728
rect 20824 30688 21916 30716
rect 20824 30660 20852 30688
rect 21910 30676 21916 30688
rect 21968 30716 21974 30728
rect 23216 30716 23244 30747
rect 21968 30688 23244 30716
rect 21968 30676 21974 30688
rect 20806 30648 20812 30660
rect 19536 30620 20812 30648
rect 20806 30608 20812 30620
rect 20864 30608 20870 30660
rect 20898 30608 20904 30660
rect 20956 30648 20962 30660
rect 22646 30648 22652 30660
rect 20956 30620 22652 30648
rect 20956 30608 20962 30620
rect 22646 30608 22652 30620
rect 22704 30648 22710 30660
rect 23308 30648 23336 30747
rect 23382 30744 23388 30796
rect 23440 30784 23446 30796
rect 23477 30787 23535 30793
rect 23477 30784 23489 30787
rect 23440 30756 23489 30784
rect 23440 30744 23446 30756
rect 23477 30753 23489 30756
rect 23523 30753 23535 30787
rect 23584 30784 23612 30824
rect 26602 30812 26608 30864
rect 26660 30852 26666 30864
rect 26697 30855 26755 30861
rect 26697 30852 26709 30855
rect 26660 30824 26709 30852
rect 26660 30812 26666 30824
rect 26697 30821 26709 30824
rect 26743 30821 26755 30855
rect 26697 30815 26755 30821
rect 24213 30787 24271 30793
rect 24213 30784 24225 30787
rect 23584 30756 24225 30784
rect 23477 30747 23535 30753
rect 24213 30753 24225 30756
rect 24259 30753 24271 30787
rect 24213 30747 24271 30753
rect 25406 30744 25412 30796
rect 25464 30784 25470 30796
rect 25774 30784 25780 30796
rect 25464 30756 25780 30784
rect 25464 30744 25470 30756
rect 25774 30744 25780 30756
rect 25832 30744 25838 30796
rect 27522 30744 27528 30796
rect 27580 30784 27586 30796
rect 28169 30787 28227 30793
rect 28169 30784 28181 30787
rect 27580 30756 28181 30784
rect 27580 30744 27586 30756
rect 28169 30753 28181 30756
rect 28215 30753 28227 30787
rect 28169 30747 28227 30753
rect 23937 30719 23995 30725
rect 23937 30685 23949 30719
rect 23983 30716 23995 30719
rect 25222 30716 25228 30728
rect 23983 30688 25228 30716
rect 23983 30685 23995 30688
rect 23937 30679 23995 30685
rect 25222 30676 25228 30688
rect 25280 30676 25286 30728
rect 26881 30651 26939 30657
rect 26881 30648 26893 30651
rect 22704 30620 23336 30648
rect 24872 30620 26893 30648
rect 22704 30608 22710 30620
rect 18690 30580 18696 30592
rect 16632 30552 18696 30580
rect 16632 30540 16638 30552
rect 18690 30540 18696 30552
rect 18748 30540 18754 30592
rect 19426 30540 19432 30592
rect 19484 30580 19490 30592
rect 20530 30580 20536 30592
rect 19484 30552 20536 30580
rect 19484 30540 19490 30552
rect 20530 30540 20536 30552
rect 20588 30540 20594 30592
rect 20990 30540 20996 30592
rect 21048 30580 21054 30592
rect 21177 30583 21235 30589
rect 21177 30580 21189 30583
rect 21048 30552 21189 30580
rect 21048 30540 21054 30552
rect 21177 30549 21189 30552
rect 21223 30549 21235 30583
rect 21177 30543 21235 30549
rect 21266 30540 21272 30592
rect 21324 30580 21330 30592
rect 24872 30580 24900 30620
rect 26881 30617 26893 30620
rect 26927 30617 26939 30651
rect 26881 30611 26939 30617
rect 21324 30552 24900 30580
rect 21324 30540 21330 30552
rect 25222 30540 25228 30592
rect 25280 30580 25286 30592
rect 25317 30583 25375 30589
rect 25317 30580 25329 30583
rect 25280 30552 25329 30580
rect 25280 30540 25286 30552
rect 25317 30549 25329 30552
rect 25363 30549 25375 30583
rect 27982 30580 27988 30592
rect 27943 30552 27988 30580
rect 25317 30543 25375 30549
rect 27982 30540 27988 30552
rect 28040 30540 28046 30592
rect 1104 30490 28888 30512
rect 1104 30438 5614 30490
rect 5666 30438 5678 30490
rect 5730 30438 5742 30490
rect 5794 30438 5806 30490
rect 5858 30438 14878 30490
rect 14930 30438 14942 30490
rect 14994 30438 15006 30490
rect 15058 30438 15070 30490
rect 15122 30438 24142 30490
rect 24194 30438 24206 30490
rect 24258 30438 24270 30490
rect 24322 30438 24334 30490
rect 24386 30438 28888 30490
rect 1104 30416 28888 30438
rect 4982 30336 4988 30388
rect 5040 30376 5046 30388
rect 5258 30376 5264 30388
rect 5040 30348 5264 30376
rect 5040 30336 5046 30348
rect 5258 30336 5264 30348
rect 5316 30336 5322 30388
rect 6638 30336 6644 30388
rect 6696 30376 6702 30388
rect 6914 30376 6920 30388
rect 6696 30348 6920 30376
rect 6696 30336 6702 30348
rect 6914 30336 6920 30348
rect 6972 30336 6978 30388
rect 12342 30336 12348 30388
rect 12400 30376 12406 30388
rect 13722 30376 13728 30388
rect 12400 30348 13728 30376
rect 12400 30336 12406 30348
rect 13722 30336 13728 30348
rect 13780 30336 13786 30388
rect 17402 30336 17408 30388
rect 17460 30376 17466 30388
rect 17681 30379 17739 30385
rect 17681 30376 17693 30379
rect 17460 30348 17693 30376
rect 17460 30336 17466 30348
rect 17681 30345 17693 30348
rect 17727 30345 17739 30379
rect 22094 30376 22100 30388
rect 17681 30339 17739 30345
rect 21468 30348 22100 30376
rect 1854 30268 1860 30320
rect 1912 30308 1918 30320
rect 6086 30308 6092 30320
rect 1912 30280 5948 30308
rect 6047 30280 6092 30308
rect 1912 30268 1918 30280
rect 2866 30200 2872 30252
rect 2924 30240 2930 30252
rect 3329 30243 3387 30249
rect 3329 30240 3341 30243
rect 2924 30212 3341 30240
rect 2924 30200 2930 30212
rect 3329 30209 3341 30212
rect 3375 30209 3387 30243
rect 5920 30240 5948 30280
rect 6086 30268 6092 30280
rect 6144 30268 6150 30320
rect 6730 30308 6736 30320
rect 6691 30280 6736 30308
rect 6730 30268 6736 30280
rect 6788 30268 6794 30320
rect 14829 30311 14887 30317
rect 12406 30280 13216 30308
rect 12406 30240 12434 30280
rect 5920 30212 12434 30240
rect 3329 30203 3387 30209
rect 3053 30175 3111 30181
rect 3053 30141 3065 30175
rect 3099 30141 3111 30175
rect 3053 30135 3111 30141
rect 3145 30175 3203 30181
rect 3145 30141 3157 30175
rect 3191 30172 3203 30175
rect 4338 30172 4344 30184
rect 3191 30144 4344 30172
rect 3191 30141 3203 30144
rect 3145 30135 3203 30141
rect 1854 30104 1860 30116
rect 1815 30076 1860 30104
rect 1854 30064 1860 30076
rect 1912 30064 1918 30116
rect 3068 30104 3096 30135
rect 4338 30132 4344 30144
rect 4396 30132 4402 30184
rect 4798 30172 4804 30184
rect 4759 30144 4804 30172
rect 4798 30132 4804 30144
rect 4856 30132 4862 30184
rect 4890 30132 4896 30184
rect 4948 30172 4954 30184
rect 5077 30175 5135 30181
rect 4948 30144 4993 30172
rect 4948 30132 4954 30144
rect 5077 30141 5089 30175
rect 5123 30141 5135 30175
rect 5077 30135 5135 30141
rect 5537 30175 5595 30181
rect 5537 30141 5549 30175
rect 5583 30172 5595 30175
rect 5902 30172 5908 30184
rect 5583 30144 5908 30172
rect 5583 30141 5595 30144
rect 5537 30135 5595 30141
rect 4062 30104 4068 30116
rect 3068 30076 4068 30104
rect 4062 30064 4068 30076
rect 4120 30104 4126 30116
rect 4706 30104 4712 30116
rect 4120 30076 4712 30104
rect 4120 30064 4126 30076
rect 4706 30064 4712 30076
rect 4764 30064 4770 30116
rect 5092 30104 5120 30135
rect 5902 30132 5908 30144
rect 5960 30132 5966 30184
rect 5997 30175 6055 30181
rect 5997 30141 6009 30175
rect 6043 30172 6055 30175
rect 6086 30172 6092 30184
rect 6043 30144 6092 30172
rect 6043 30141 6055 30144
rect 5997 30135 6055 30141
rect 6086 30132 6092 30144
rect 6144 30132 6150 30184
rect 6638 30172 6644 30184
rect 6599 30144 6644 30172
rect 6638 30132 6644 30144
rect 6696 30132 6702 30184
rect 9582 30172 9588 30184
rect 9543 30144 9588 30172
rect 9582 30132 9588 30144
rect 9640 30132 9646 30184
rect 11974 30172 11980 30184
rect 11935 30144 11980 30172
rect 11974 30132 11980 30144
rect 12032 30132 12038 30184
rect 12345 30175 12403 30181
rect 12345 30141 12357 30175
rect 12391 30172 12403 30175
rect 12434 30172 12440 30184
rect 12391 30144 12440 30172
rect 12391 30141 12403 30144
rect 12345 30135 12403 30141
rect 12434 30132 12440 30144
rect 12492 30132 12498 30184
rect 12802 30172 12808 30184
rect 12763 30144 12808 30172
rect 12802 30132 12808 30144
rect 12860 30132 12866 30184
rect 6178 30104 6184 30116
rect 5092 30076 6184 30104
rect 6178 30064 6184 30076
rect 6236 30064 6242 30116
rect 11885 30107 11943 30113
rect 11885 30104 11897 30107
rect 8036 30076 11897 30104
rect 1949 30039 2007 30045
rect 1949 30005 1961 30039
rect 1995 30036 2007 30039
rect 2406 30036 2412 30048
rect 1995 30008 2412 30036
rect 1995 30005 2007 30008
rect 1949 29999 2007 30005
rect 2406 29996 2412 30008
rect 2464 29996 2470 30048
rect 3326 30036 3332 30048
rect 3287 30008 3332 30036
rect 3326 29996 3332 30008
rect 3384 29996 3390 30048
rect 3970 29996 3976 30048
rect 4028 30036 4034 30048
rect 8036 30036 8064 30076
rect 11885 30073 11897 30076
rect 11931 30073 11943 30107
rect 11885 30067 11943 30073
rect 9674 30036 9680 30048
rect 4028 30008 8064 30036
rect 9635 30008 9680 30036
rect 4028 29996 4034 30008
rect 9674 29996 9680 30008
rect 9732 29996 9738 30048
rect 13188 30036 13216 30280
rect 14829 30277 14841 30311
rect 14875 30277 14887 30311
rect 16574 30308 16580 30320
rect 16535 30280 16580 30308
rect 14829 30271 14887 30277
rect 13722 30240 13728 30252
rect 13280 30212 13728 30240
rect 13280 30181 13308 30212
rect 13722 30200 13728 30212
rect 13780 30240 13786 30252
rect 14844 30240 14872 30271
rect 16574 30268 16580 30280
rect 16632 30268 16638 30320
rect 13780 30212 14872 30240
rect 13780 30200 13786 30212
rect 15102 30200 15108 30252
rect 15160 30240 15166 30252
rect 16942 30240 16948 30252
rect 15160 30212 16948 30240
rect 15160 30200 15166 30212
rect 16942 30200 16948 30212
rect 17000 30240 17006 30252
rect 17696 30240 17724 30339
rect 18969 30311 19027 30317
rect 18969 30277 18981 30311
rect 19015 30308 19027 30311
rect 19702 30308 19708 30320
rect 19015 30280 19708 30308
rect 19015 30277 19027 30280
rect 18969 30271 19027 30277
rect 19702 30268 19708 30280
rect 19760 30268 19766 30320
rect 20806 30268 20812 30320
rect 20864 30268 20870 30320
rect 20438 30240 20444 30252
rect 17000 30212 17540 30240
rect 17696 30212 20444 30240
rect 17000 30200 17006 30212
rect 13265 30175 13323 30181
rect 13265 30141 13277 30175
rect 13311 30141 13323 30175
rect 13446 30172 13452 30184
rect 13407 30144 13452 30172
rect 13265 30135 13323 30141
rect 13446 30132 13452 30144
rect 13504 30132 13510 30184
rect 13814 30132 13820 30184
rect 13872 30172 13878 30184
rect 14550 30172 14556 30184
rect 13872 30144 14556 30172
rect 13872 30132 13878 30144
rect 14550 30132 14556 30144
rect 14608 30172 14614 30184
rect 14737 30175 14795 30181
rect 14737 30172 14749 30175
rect 14608 30144 14749 30172
rect 14608 30132 14614 30144
rect 14737 30141 14749 30144
rect 14783 30141 14795 30175
rect 14737 30135 14795 30141
rect 14921 30175 14979 30181
rect 14921 30141 14933 30175
rect 14967 30172 14979 30175
rect 15657 30175 15715 30181
rect 15657 30172 15669 30175
rect 14967 30144 15669 30172
rect 14967 30141 14979 30144
rect 14921 30135 14979 30141
rect 15657 30141 15669 30144
rect 15703 30172 15715 30175
rect 16114 30172 16120 30184
rect 15703 30144 16120 30172
rect 15703 30141 15715 30144
rect 15657 30135 15715 30141
rect 13906 30064 13912 30116
rect 13964 30104 13970 30116
rect 14936 30104 14964 30135
rect 16114 30132 16120 30144
rect 16172 30132 16178 30184
rect 17512 30181 17540 30212
rect 20438 30200 20444 30212
rect 20496 30200 20502 30252
rect 20824 30240 20852 30268
rect 21468 30249 21496 30348
rect 22094 30336 22100 30348
rect 22152 30336 22158 30388
rect 23014 30336 23020 30388
rect 23072 30376 23078 30388
rect 24026 30376 24032 30388
rect 23072 30348 23888 30376
rect 23987 30348 24032 30376
rect 23072 30336 23078 30348
rect 23290 30268 23296 30320
rect 23348 30308 23354 30320
rect 23860 30308 23888 30348
rect 24026 30336 24032 30348
rect 24084 30336 24090 30388
rect 25222 30308 25228 30320
rect 23348 30280 23796 30308
rect 23860 30280 25228 30308
rect 23348 30268 23354 30280
rect 20732 30212 20852 30240
rect 21453 30243 21511 30249
rect 17497 30175 17555 30181
rect 17497 30141 17509 30175
rect 17543 30141 17555 30175
rect 17497 30135 17555 30141
rect 18601 30175 18659 30181
rect 18601 30141 18613 30175
rect 18647 30141 18659 30175
rect 18601 30135 18659 30141
rect 18693 30175 18751 30181
rect 18693 30141 18705 30175
rect 18739 30141 18751 30175
rect 18693 30135 18751 30141
rect 15838 30104 15844 30116
rect 13964 30076 14964 30104
rect 15751 30076 15844 30104
rect 13964 30064 13970 30076
rect 15838 30064 15844 30076
rect 15896 30104 15902 30116
rect 16393 30107 16451 30113
rect 16393 30104 16405 30107
rect 15896 30076 16405 30104
rect 15896 30064 15902 30076
rect 16393 30073 16405 30076
rect 16439 30073 16451 30107
rect 16393 30067 16451 30073
rect 16666 30064 16672 30116
rect 16724 30104 16730 30116
rect 18616 30104 18644 30135
rect 16724 30076 18644 30104
rect 18708 30104 18736 30135
rect 18782 30132 18788 30184
rect 18840 30172 18846 30184
rect 20732 30181 20760 30212
rect 21453 30209 21465 30243
rect 21499 30209 21511 30243
rect 21453 30203 21511 30209
rect 20625 30175 20683 30181
rect 18840 30144 18885 30172
rect 18840 30132 18846 30144
rect 20625 30141 20637 30175
rect 20671 30141 20683 30175
rect 20625 30135 20683 30141
rect 20717 30175 20775 30181
rect 20717 30141 20729 30175
rect 20763 30141 20775 30175
rect 20717 30135 20775 30141
rect 18966 30104 18972 30116
rect 18708 30076 18972 30104
rect 16724 30064 16730 30076
rect 18966 30064 18972 30076
rect 19024 30064 19030 30116
rect 20346 30104 20352 30116
rect 20307 30076 20352 30104
rect 20346 30064 20352 30076
rect 20404 30064 20410 30116
rect 20640 30104 20668 30135
rect 20806 30132 20812 30184
rect 20864 30172 20870 30184
rect 20990 30172 20996 30184
rect 20864 30144 20909 30172
rect 20951 30144 20996 30172
rect 20864 30132 20870 30144
rect 20990 30132 20996 30144
rect 21048 30132 21054 30184
rect 21726 30172 21732 30184
rect 21687 30144 21732 30172
rect 21726 30132 21732 30144
rect 21784 30132 21790 30184
rect 22922 30132 22928 30184
rect 22980 30172 22986 30184
rect 23768 30181 23796 30280
rect 25222 30268 25228 30280
rect 25280 30268 25286 30320
rect 26145 30311 26203 30317
rect 26145 30277 26157 30311
rect 26191 30277 26203 30311
rect 26145 30271 26203 30277
rect 26160 30240 26188 30271
rect 26160 30212 28028 30240
rect 23661 30175 23719 30181
rect 23661 30172 23673 30175
rect 22980 30144 23673 30172
rect 22980 30132 22986 30144
rect 23661 30141 23673 30144
rect 23707 30141 23719 30175
rect 23661 30135 23719 30141
rect 23753 30175 23811 30181
rect 23753 30141 23765 30175
rect 23799 30141 23811 30175
rect 23753 30135 23811 30141
rect 23845 30175 23903 30181
rect 23845 30141 23857 30175
rect 23891 30141 23903 30175
rect 25682 30172 25688 30184
rect 25643 30144 25688 30172
rect 23845 30135 23903 30141
rect 20640 30076 20760 30104
rect 17034 30036 17040 30048
rect 13188 30008 17040 30036
rect 17034 29996 17040 30008
rect 17092 29996 17098 30048
rect 20732 30036 20760 30076
rect 23198 30064 23204 30116
rect 23256 30104 23262 30116
rect 23860 30104 23888 30135
rect 25682 30132 25688 30144
rect 25740 30132 25746 30184
rect 26142 30132 26148 30184
rect 26200 30172 26206 30184
rect 28000 30181 28028 30212
rect 26329 30175 26387 30181
rect 26329 30172 26341 30175
rect 26200 30144 26341 30172
rect 26200 30132 26206 30144
rect 26329 30141 26341 30144
rect 26375 30141 26387 30175
rect 26329 30135 26387 30141
rect 27985 30175 28043 30181
rect 27985 30141 27997 30175
rect 28031 30141 28043 30175
rect 27985 30135 28043 30141
rect 26881 30107 26939 30113
rect 26881 30104 26893 30107
rect 23256 30076 23888 30104
rect 25516 30076 26893 30104
rect 23256 30064 23262 30076
rect 21450 30036 21456 30048
rect 20732 30008 21456 30036
rect 21450 29996 21456 30008
rect 21508 30036 21514 30048
rect 22462 30036 22468 30048
rect 21508 30008 22468 30036
rect 21508 29996 21514 30008
rect 22462 29996 22468 30008
rect 22520 30036 22526 30048
rect 25516 30045 25544 30076
rect 26881 30073 26893 30076
rect 26927 30073 26939 30107
rect 26881 30067 26939 30073
rect 22833 30039 22891 30045
rect 22833 30036 22845 30039
rect 22520 30008 22845 30036
rect 22520 29996 22526 30008
rect 22833 30005 22845 30008
rect 22879 30005 22891 30039
rect 22833 29999 22891 30005
rect 25501 30039 25559 30045
rect 25501 30005 25513 30039
rect 25547 30005 25559 30039
rect 25501 29999 25559 30005
rect 25590 29996 25596 30048
rect 25648 30036 25654 30048
rect 26973 30039 27031 30045
rect 26973 30036 26985 30039
rect 25648 30008 26985 30036
rect 25648 29996 25654 30008
rect 26973 30005 26985 30008
rect 27019 30005 27031 30039
rect 26973 29999 27031 30005
rect 27062 29996 27068 30048
rect 27120 30036 27126 30048
rect 28077 30039 28135 30045
rect 28077 30036 28089 30039
rect 27120 30008 28089 30036
rect 27120 29996 27126 30008
rect 28077 30005 28089 30008
rect 28123 30005 28135 30039
rect 28077 29999 28135 30005
rect 1104 29946 28888 29968
rect 1104 29894 10246 29946
rect 10298 29894 10310 29946
rect 10362 29894 10374 29946
rect 10426 29894 10438 29946
rect 10490 29894 19510 29946
rect 19562 29894 19574 29946
rect 19626 29894 19638 29946
rect 19690 29894 19702 29946
rect 19754 29894 28888 29946
rect 1104 29872 28888 29894
rect 2590 29792 2596 29844
rect 2648 29832 2654 29844
rect 13814 29832 13820 29844
rect 2648 29804 13820 29832
rect 2648 29792 2654 29804
rect 13814 29792 13820 29804
rect 13872 29792 13878 29844
rect 13906 29792 13912 29844
rect 13964 29832 13970 29844
rect 14182 29832 14188 29844
rect 13964 29804 14188 29832
rect 13964 29792 13970 29804
rect 14182 29792 14188 29804
rect 14240 29832 14246 29844
rect 14369 29835 14427 29841
rect 14369 29832 14381 29835
rect 14240 29804 14381 29832
rect 14240 29792 14246 29804
rect 14369 29801 14381 29804
rect 14415 29801 14427 29835
rect 15286 29832 15292 29844
rect 14369 29795 14427 29801
rect 15212 29804 15292 29832
rect 3326 29724 3332 29776
rect 3384 29773 3390 29776
rect 3384 29767 3448 29773
rect 3384 29733 3402 29767
rect 3436 29733 3448 29767
rect 3384 29727 3448 29733
rect 5629 29767 5687 29773
rect 5629 29733 5641 29767
rect 5675 29764 5687 29767
rect 5675 29736 6040 29764
rect 5675 29733 5687 29736
rect 5629 29727 5687 29733
rect 3384 29724 3390 29727
rect 2133 29699 2191 29705
rect 2133 29665 2145 29699
rect 2179 29696 2191 29699
rect 2774 29696 2780 29708
rect 2179 29668 2780 29696
rect 2179 29665 2191 29668
rect 2133 29659 2191 29665
rect 2774 29656 2780 29668
rect 2832 29656 2838 29708
rect 5442 29696 5448 29708
rect 3160 29668 5448 29696
rect 2222 29628 2228 29640
rect 2183 29600 2228 29628
rect 2222 29588 2228 29600
rect 2280 29588 2286 29640
rect 2314 29588 2320 29640
rect 2372 29628 2378 29640
rect 3160 29637 3188 29668
rect 5442 29656 5448 29668
rect 5500 29656 5506 29708
rect 5537 29699 5595 29705
rect 5537 29665 5549 29699
rect 5583 29696 5595 29699
rect 5902 29696 5908 29708
rect 5583 29668 5908 29696
rect 5583 29665 5595 29668
rect 5537 29659 5595 29665
rect 5902 29656 5908 29668
rect 5960 29656 5966 29708
rect 3145 29631 3203 29637
rect 2372 29600 2417 29628
rect 2372 29588 2378 29600
rect 3145 29597 3157 29631
rect 3191 29597 3203 29631
rect 3145 29591 3203 29597
rect 1394 29520 1400 29572
rect 1452 29560 1458 29572
rect 3050 29560 3056 29572
rect 1452 29532 3056 29560
rect 1452 29520 1458 29532
rect 3050 29520 3056 29532
rect 3108 29560 3114 29572
rect 3160 29560 3188 29591
rect 4982 29588 4988 29640
rect 5040 29628 5046 29640
rect 5718 29628 5724 29640
rect 5040 29600 5724 29628
rect 5040 29588 5046 29600
rect 5718 29588 5724 29600
rect 5776 29588 5782 29640
rect 3108 29532 3188 29560
rect 5169 29563 5227 29569
rect 3108 29520 3114 29532
rect 5169 29529 5181 29563
rect 5215 29560 5227 29563
rect 5534 29560 5540 29572
rect 5215 29532 5540 29560
rect 5215 29529 5227 29532
rect 5169 29523 5227 29529
rect 5534 29520 5540 29532
rect 5592 29520 5598 29572
rect 1670 29452 1676 29504
rect 1728 29492 1734 29504
rect 1765 29495 1823 29501
rect 1765 29492 1777 29495
rect 1728 29464 1777 29492
rect 1728 29452 1734 29464
rect 1765 29461 1777 29464
rect 1811 29461 1823 29495
rect 4522 29492 4528 29504
rect 4483 29464 4528 29492
rect 1765 29455 1823 29461
rect 4522 29452 4528 29464
rect 4580 29452 4586 29504
rect 6012 29492 6040 29736
rect 9122 29724 9128 29776
rect 9180 29764 9186 29776
rect 9180 29736 9904 29764
rect 9180 29724 9186 29736
rect 6638 29696 6644 29708
rect 6104 29668 6644 29696
rect 6104 29560 6132 29668
rect 6638 29656 6644 29668
rect 6696 29656 6702 29708
rect 8472 29699 8530 29705
rect 8472 29665 8484 29699
rect 8518 29696 8530 29699
rect 9876 29696 9904 29736
rect 9950 29724 9956 29776
rect 10008 29764 10014 29776
rect 10413 29767 10471 29773
rect 10413 29764 10425 29767
rect 10008 29736 10425 29764
rect 10008 29724 10014 29736
rect 10413 29733 10425 29736
rect 10459 29733 10471 29767
rect 10413 29727 10471 29733
rect 12158 29724 12164 29776
rect 12216 29764 12222 29776
rect 12216 29736 14320 29764
rect 12216 29724 12222 29736
rect 14292 29708 14320 29736
rect 8518 29668 9536 29696
rect 8518 29665 8530 29668
rect 8472 29659 8530 29665
rect 7742 29588 7748 29640
rect 7800 29628 7806 29640
rect 8205 29631 8263 29637
rect 8205 29628 8217 29631
rect 7800 29600 8217 29628
rect 7800 29588 7806 29600
rect 8205 29597 8217 29600
rect 8251 29597 8263 29631
rect 9508 29628 9536 29668
rect 9600 29668 9812 29696
rect 9876 29668 10640 29696
rect 9600 29628 9628 29668
rect 9508 29600 9628 29628
rect 9784 29628 9812 29668
rect 10612 29637 10640 29668
rect 12710 29656 12716 29708
rect 12768 29696 12774 29708
rect 13725 29699 13783 29705
rect 13725 29696 13737 29699
rect 12768 29668 13737 29696
rect 12768 29656 12774 29668
rect 13725 29665 13737 29668
rect 13771 29665 13783 29699
rect 14274 29696 14280 29708
rect 14235 29668 14280 29696
rect 13725 29659 13783 29665
rect 10505 29631 10563 29637
rect 9784 29600 10088 29628
rect 8205 29591 8263 29597
rect 6270 29560 6276 29572
rect 6104 29532 6276 29560
rect 6270 29520 6276 29532
rect 6328 29520 6334 29572
rect 9582 29560 9588 29572
rect 9543 29532 9588 29560
rect 9582 29520 9588 29532
rect 9640 29560 9646 29572
rect 9950 29560 9956 29572
rect 9640 29532 9956 29560
rect 9640 29520 9646 29532
rect 9950 29520 9956 29532
rect 10008 29520 10014 29572
rect 10060 29569 10088 29600
rect 10505 29597 10517 29631
rect 10551 29597 10563 29631
rect 10505 29591 10563 29597
rect 10597 29631 10655 29637
rect 10597 29597 10609 29631
rect 10643 29597 10655 29631
rect 13740 29628 13768 29659
rect 14274 29656 14280 29668
rect 14332 29656 14338 29708
rect 14461 29699 14519 29705
rect 14461 29665 14473 29699
rect 14507 29696 14519 29699
rect 14550 29696 14556 29708
rect 14507 29668 14556 29696
rect 14507 29665 14519 29668
rect 14461 29659 14519 29665
rect 14550 29656 14556 29668
rect 14608 29656 14614 29708
rect 15212 29705 15240 29804
rect 15286 29792 15292 29804
rect 15344 29792 15350 29844
rect 15378 29792 15384 29844
rect 15436 29832 15442 29844
rect 16025 29835 16083 29841
rect 16025 29832 16037 29835
rect 15436 29804 16037 29832
rect 15436 29792 15442 29804
rect 16025 29801 16037 29804
rect 16071 29801 16083 29835
rect 16025 29795 16083 29801
rect 20070 29792 20076 29844
rect 20128 29832 20134 29844
rect 20806 29832 20812 29844
rect 20128 29804 20812 29832
rect 20128 29792 20134 29804
rect 20806 29792 20812 29804
rect 20864 29792 20870 29844
rect 25961 29835 26019 29841
rect 25961 29801 25973 29835
rect 26007 29832 26019 29835
rect 26326 29832 26332 29844
rect 26007 29804 26332 29832
rect 26007 29801 26019 29804
rect 25961 29795 26019 29801
rect 26326 29792 26332 29804
rect 26384 29792 26390 29844
rect 15562 29724 15568 29776
rect 15620 29764 15626 29776
rect 27062 29764 27068 29776
rect 15620 29736 27068 29764
rect 15620 29724 15626 29736
rect 27062 29724 27068 29736
rect 27120 29724 27126 29776
rect 27982 29764 27988 29776
rect 27943 29736 27988 29764
rect 27982 29724 27988 29736
rect 28040 29724 28046 29776
rect 15105 29699 15163 29705
rect 15105 29665 15117 29699
rect 15151 29665 15163 29699
rect 15105 29659 15163 29665
rect 15197 29699 15255 29705
rect 15197 29665 15209 29699
rect 15243 29665 15255 29699
rect 15197 29659 15255 29665
rect 15289 29699 15347 29705
rect 15289 29665 15301 29699
rect 15335 29665 15347 29699
rect 15289 29659 15347 29665
rect 15473 29699 15531 29705
rect 15473 29665 15485 29699
rect 15519 29696 15531 29699
rect 15933 29699 15991 29705
rect 15933 29696 15945 29699
rect 15519 29668 15945 29696
rect 15519 29665 15531 29668
rect 15473 29659 15531 29665
rect 15933 29665 15945 29668
rect 15979 29665 15991 29699
rect 16114 29696 16120 29708
rect 16075 29668 16120 29696
rect 15933 29659 15991 29665
rect 15120 29628 15148 29659
rect 13740 29600 15148 29628
rect 10597 29591 10655 29597
rect 10045 29563 10103 29569
rect 10045 29529 10057 29563
rect 10091 29529 10103 29563
rect 10045 29523 10103 29529
rect 6822 29492 6828 29504
rect 6012 29464 6828 29492
rect 6822 29452 6828 29464
rect 6880 29452 6886 29504
rect 8386 29452 8392 29504
rect 8444 29492 8450 29504
rect 10520 29492 10548 29591
rect 15304 29572 15332 29659
rect 16114 29656 16120 29668
rect 16172 29656 16178 29708
rect 16942 29656 16948 29708
rect 17000 29696 17006 29708
rect 17218 29696 17224 29708
rect 17000 29668 17224 29696
rect 17000 29656 17006 29668
rect 17218 29656 17224 29668
rect 17276 29656 17282 29708
rect 26050 29656 26056 29708
rect 26108 29696 26114 29708
rect 26145 29699 26203 29705
rect 26145 29696 26157 29699
rect 26108 29668 26157 29696
rect 26108 29656 26114 29668
rect 26145 29665 26157 29668
rect 26191 29665 26203 29699
rect 26694 29696 26700 29708
rect 26655 29668 26700 29696
rect 26145 29659 26203 29665
rect 26694 29656 26700 29668
rect 26752 29656 26758 29708
rect 17034 29588 17040 29640
rect 17092 29628 17098 29640
rect 28169 29631 28227 29637
rect 28169 29628 28181 29631
rect 17092 29600 28181 29628
rect 17092 29588 17098 29600
rect 28169 29597 28181 29600
rect 28215 29597 28227 29631
rect 28169 29591 28227 29597
rect 15286 29520 15292 29572
rect 15344 29520 15350 29572
rect 15562 29520 15568 29572
rect 15620 29560 15626 29572
rect 26234 29560 26240 29572
rect 15620 29532 26240 29560
rect 15620 29520 15626 29532
rect 26234 29520 26240 29532
rect 26292 29520 26298 29572
rect 26878 29560 26884 29572
rect 26839 29532 26884 29560
rect 26878 29520 26884 29532
rect 26936 29520 26942 29572
rect 8444 29464 10548 29492
rect 8444 29452 8450 29464
rect 12434 29452 12440 29504
rect 12492 29492 12498 29504
rect 13446 29492 13452 29504
rect 12492 29464 13452 29492
rect 12492 29452 12498 29464
rect 13446 29452 13452 29464
rect 13504 29452 13510 29504
rect 15470 29452 15476 29504
rect 15528 29492 15534 29504
rect 20438 29492 20444 29504
rect 15528 29464 20444 29492
rect 15528 29452 15534 29464
rect 20438 29452 20444 29464
rect 20496 29452 20502 29504
rect 1104 29402 28888 29424
rect 1104 29350 5614 29402
rect 5666 29350 5678 29402
rect 5730 29350 5742 29402
rect 5794 29350 5806 29402
rect 5858 29350 14878 29402
rect 14930 29350 14942 29402
rect 14994 29350 15006 29402
rect 15058 29350 15070 29402
rect 15122 29350 24142 29402
rect 24194 29350 24206 29402
rect 24258 29350 24270 29402
rect 24322 29350 24334 29402
rect 24386 29350 28888 29402
rect 1104 29328 28888 29350
rect 25590 29288 25596 29300
rect 2746 29260 25596 29288
rect 2746 29164 2774 29260
rect 25590 29248 25596 29260
rect 25648 29248 25654 29300
rect 27430 29248 27436 29300
rect 27488 29288 27494 29300
rect 27985 29291 28043 29297
rect 27985 29288 27997 29291
rect 27488 29260 27997 29288
rect 27488 29248 27494 29260
rect 27985 29257 27997 29260
rect 28031 29257 28043 29291
rect 27985 29251 28043 29257
rect 4249 29223 4307 29229
rect 4249 29189 4261 29223
rect 4295 29220 4307 29223
rect 4890 29220 4896 29232
rect 4295 29192 4896 29220
rect 4295 29189 4307 29192
rect 4249 29183 4307 29189
rect 4890 29180 4896 29192
rect 4948 29180 4954 29232
rect 6822 29220 6828 29232
rect 6735 29192 6828 29220
rect 6822 29180 6828 29192
rect 6880 29180 6886 29232
rect 7558 29180 7564 29232
rect 7616 29220 7622 29232
rect 8021 29223 8079 29229
rect 8021 29220 8033 29223
rect 7616 29192 8033 29220
rect 7616 29180 7622 29192
rect 8021 29189 8033 29192
rect 8067 29189 8079 29223
rect 10502 29220 10508 29232
rect 8021 29183 8079 29189
rect 8588 29192 10508 29220
rect 1394 29152 1400 29164
rect 1355 29124 1400 29152
rect 1394 29112 1400 29124
rect 1452 29112 1458 29164
rect 2682 29112 2688 29164
rect 2740 29124 2774 29164
rect 4801 29155 4859 29161
rect 2740 29112 2746 29124
rect 4801 29121 4813 29155
rect 4847 29152 4859 29155
rect 4982 29152 4988 29164
rect 4847 29124 4988 29152
rect 4847 29121 4859 29124
rect 4801 29115 4859 29121
rect 4982 29112 4988 29124
rect 5040 29112 5046 29164
rect 5442 29152 5448 29164
rect 5403 29124 5448 29152
rect 5442 29112 5448 29124
rect 5500 29112 5506 29164
rect 6840 29152 6868 29180
rect 8588 29152 8616 29192
rect 10502 29180 10508 29192
rect 10560 29180 10566 29232
rect 11698 29180 11704 29232
rect 11756 29220 11762 29232
rect 22370 29220 22376 29232
rect 11756 29192 22376 29220
rect 11756 29180 11762 29192
rect 22370 29180 22376 29192
rect 22428 29180 22434 29232
rect 22922 29180 22928 29232
rect 22980 29220 22986 29232
rect 26510 29220 26516 29232
rect 22980 29192 26516 29220
rect 22980 29180 22986 29192
rect 26510 29180 26516 29192
rect 26568 29180 26574 29232
rect 6840 29124 8616 29152
rect 9122 29112 9128 29164
rect 9180 29152 9186 29164
rect 9398 29152 9404 29164
rect 9180 29124 9404 29152
rect 9180 29112 9186 29124
rect 9398 29112 9404 29124
rect 9456 29112 9462 29164
rect 10689 29155 10747 29161
rect 10689 29121 10701 29155
rect 10735 29152 10747 29155
rect 11054 29152 11060 29164
rect 10735 29124 11060 29152
rect 10735 29121 10747 29124
rect 10689 29115 10747 29121
rect 11054 29112 11060 29124
rect 11112 29112 11118 29164
rect 12250 29152 12256 29164
rect 11164 29124 12256 29152
rect 1670 29093 1676 29096
rect 1664 29084 1676 29093
rect 1631 29056 1676 29084
rect 1664 29047 1676 29056
rect 1670 29044 1676 29047
rect 1728 29044 1734 29096
rect 2774 29044 2780 29096
rect 2832 29044 2838 29096
rect 4338 29044 4344 29096
rect 4396 29084 4402 29096
rect 4617 29087 4675 29093
rect 4617 29084 4629 29087
rect 4396 29056 4629 29084
rect 4396 29044 4402 29056
rect 4617 29053 4629 29056
rect 4663 29084 4675 29087
rect 5350 29084 5356 29096
rect 4663 29056 5356 29084
rect 4663 29053 4675 29056
rect 4617 29047 4675 29053
rect 5350 29044 5356 29056
rect 5408 29044 5414 29096
rect 5460 29084 5488 29112
rect 7742 29084 7748 29096
rect 5460 29056 7748 29084
rect 7742 29044 7748 29056
rect 7800 29044 7806 29096
rect 7926 29084 7932 29096
rect 7887 29056 7932 29084
rect 7926 29044 7932 29056
rect 7984 29044 7990 29096
rect 8205 29087 8263 29093
rect 8205 29053 8217 29087
rect 8251 29084 8263 29087
rect 8386 29084 8392 29096
rect 8251 29056 8392 29084
rect 8251 29053 8263 29056
rect 8205 29047 8263 29053
rect 8386 29044 8392 29056
rect 8444 29044 8450 29096
rect 9769 29087 9827 29093
rect 9769 29053 9781 29087
rect 9815 29084 9827 29087
rect 9815 29056 9849 29084
rect 9815 29053 9827 29056
rect 9769 29047 9827 29053
rect 2792 29016 2820 29044
rect 4246 29016 4252 29028
rect 2792 28988 4252 29016
rect 2792 28957 2820 28988
rect 4246 28976 4252 28988
rect 4304 28976 4310 29028
rect 4706 29016 4712 29028
rect 4667 28988 4712 29016
rect 4706 28976 4712 28988
rect 4764 28976 4770 29028
rect 5712 29019 5770 29025
rect 5712 28985 5724 29019
rect 5758 29016 5770 29019
rect 5810 29016 5816 29028
rect 5758 28988 5816 29016
rect 5758 28985 5770 28988
rect 5712 28979 5770 28985
rect 5810 28976 5816 28988
rect 5868 28976 5874 29028
rect 9784 29016 9812 29047
rect 10778 29044 10784 29096
rect 10836 29084 10842 29096
rect 10965 29087 11023 29093
rect 10836 29056 10881 29084
rect 10836 29044 10842 29056
rect 10965 29053 10977 29087
rect 11011 29084 11023 29087
rect 11164 29084 11192 29124
rect 12250 29112 12256 29124
rect 12308 29152 12314 29164
rect 25682 29152 25688 29164
rect 12308 29124 15056 29152
rect 25643 29124 25688 29152
rect 12308 29112 12314 29124
rect 11011 29056 11192 29084
rect 11425 29087 11483 29093
rect 11011 29053 11023 29056
rect 10965 29047 11023 29053
rect 11425 29053 11437 29087
rect 11471 29084 11483 29087
rect 11698 29084 11704 29096
rect 11471 29056 11704 29084
rect 11471 29053 11483 29056
rect 11425 29047 11483 29053
rect 11698 29044 11704 29056
rect 11756 29044 11762 29096
rect 11882 29084 11888 29096
rect 11843 29056 11888 29084
rect 11882 29044 11888 29056
rect 11940 29044 11946 29096
rect 13446 29044 13452 29096
rect 13504 29084 13510 29096
rect 14550 29084 14556 29096
rect 13504 29056 14556 29084
rect 13504 29044 13510 29056
rect 14550 29044 14556 29056
rect 14608 29044 14614 29096
rect 15028 29093 15056 29124
rect 25682 29112 25688 29124
rect 25740 29112 25746 29164
rect 26436 29124 27660 29152
rect 15013 29087 15071 29093
rect 15013 29053 15025 29087
rect 15059 29053 15071 29087
rect 15013 29047 15071 29053
rect 15289 29087 15347 29093
rect 15289 29053 15301 29087
rect 15335 29084 15347 29087
rect 15838 29084 15844 29096
rect 15335 29056 15844 29084
rect 15335 29053 15347 29056
rect 15289 29047 15347 29053
rect 15838 29044 15844 29056
rect 15896 29044 15902 29096
rect 25501 29087 25559 29093
rect 25501 29053 25513 29087
rect 25547 29084 25559 29087
rect 26436 29084 26464 29124
rect 27632 29096 27660 29124
rect 25547 29056 26464 29084
rect 25547 29053 25559 29056
rect 25501 29047 25559 29053
rect 26510 29044 26516 29096
rect 26568 29084 26574 29096
rect 26973 29087 27031 29093
rect 26973 29084 26985 29087
rect 26568 29056 26985 29084
rect 26568 29044 26574 29056
rect 26973 29053 26985 29056
rect 27019 29053 27031 29087
rect 27614 29084 27620 29096
rect 27575 29056 27620 29084
rect 26973 29047 27031 29053
rect 27614 29044 27620 29056
rect 27672 29044 27678 29096
rect 27706 29044 27712 29096
rect 27764 29084 27770 29096
rect 27985 29087 28043 29093
rect 27985 29084 27997 29087
rect 27764 29056 27997 29084
rect 27764 29044 27770 29056
rect 27985 29053 27997 29056
rect 28031 29053 28043 29087
rect 27985 29047 28043 29053
rect 28169 29087 28227 29093
rect 28169 29053 28181 29087
rect 28215 29084 28227 29087
rect 28258 29084 28264 29096
rect 28215 29056 28264 29084
rect 28215 29053 28227 29056
rect 28169 29047 28227 29053
rect 28258 29044 28264 29056
rect 28316 29044 28322 29096
rect 10226 29016 10232 29028
rect 5920 28988 10232 29016
rect 2777 28951 2835 28957
rect 2777 28917 2789 28951
rect 2823 28948 2835 28951
rect 2823 28920 2857 28948
rect 2823 28917 2835 28920
rect 2777 28911 2835 28917
rect 3970 28908 3976 28960
rect 4028 28948 4034 28960
rect 5920 28948 5948 28988
rect 10226 28976 10232 28988
rect 10284 28976 10290 29028
rect 11977 29019 12035 29025
rect 11977 29016 11989 29019
rect 11256 28988 11989 29016
rect 9858 28948 9864 28960
rect 4028 28920 5948 28948
rect 9819 28920 9864 28948
rect 4028 28908 4034 28920
rect 9858 28908 9864 28920
rect 9916 28908 9922 28960
rect 11256 28948 11284 28988
rect 11977 28985 11989 28988
rect 12023 28985 12035 29019
rect 15197 29019 15255 29025
rect 15197 29016 15209 29019
rect 11977 28979 12035 28985
rect 15120 28988 15209 29016
rect 11330 28948 11336 28960
rect 11256 28920 11336 28948
rect 11330 28908 11336 28920
rect 11388 28908 11394 28960
rect 14274 28908 14280 28960
rect 14332 28948 14338 28960
rect 15120 28948 15148 28988
rect 15197 28985 15209 28988
rect 15243 28985 15255 29019
rect 15197 28979 15255 28985
rect 25590 28976 25596 29028
rect 25648 29016 25654 29028
rect 26237 29019 26295 29025
rect 26237 29016 26249 29019
rect 25648 28988 26249 29016
rect 25648 28976 25654 28988
rect 26237 28985 26249 28988
rect 26283 28985 26295 29019
rect 26418 29016 26424 29028
rect 26379 28988 26424 29016
rect 26237 28979 26295 28985
rect 26418 28976 26424 28988
rect 26476 28976 26482 29028
rect 27154 29016 27160 29028
rect 27115 28988 27160 29016
rect 27154 28976 27160 28988
rect 27212 28976 27218 29028
rect 14332 28920 15148 28948
rect 15289 28951 15347 28957
rect 14332 28908 14338 28920
rect 15289 28917 15301 28951
rect 15335 28948 15347 28951
rect 16114 28948 16120 28960
rect 15335 28920 16120 28948
rect 15335 28917 15347 28920
rect 15289 28911 15347 28917
rect 16114 28908 16120 28920
rect 16172 28908 16178 28960
rect 20162 28908 20168 28960
rect 20220 28948 20226 28960
rect 24854 28948 24860 28960
rect 20220 28920 24860 28948
rect 20220 28908 20226 28920
rect 24854 28908 24860 28920
rect 24912 28908 24918 28960
rect 25130 28908 25136 28960
rect 25188 28948 25194 28960
rect 26694 28948 26700 28960
rect 25188 28920 26700 28948
rect 25188 28908 25194 28920
rect 26694 28908 26700 28920
rect 26752 28908 26758 28960
rect 27709 28951 27767 28957
rect 27709 28917 27721 28951
rect 27755 28948 27767 28951
rect 27890 28948 27896 28960
rect 27755 28920 27896 28948
rect 27755 28917 27767 28920
rect 27709 28911 27767 28917
rect 27890 28908 27896 28920
rect 27948 28908 27954 28960
rect 1104 28858 28888 28880
rect 1104 28806 10246 28858
rect 10298 28806 10310 28858
rect 10362 28806 10374 28858
rect 10426 28806 10438 28858
rect 10490 28806 19510 28858
rect 19562 28806 19574 28858
rect 19626 28806 19638 28858
rect 19690 28806 19702 28858
rect 19754 28806 28888 28858
rect 1104 28784 28888 28806
rect 2222 28704 2228 28756
rect 2280 28744 2286 28756
rect 2593 28747 2651 28753
rect 2593 28744 2605 28747
rect 2280 28716 2605 28744
rect 2280 28704 2286 28716
rect 2593 28713 2605 28716
rect 2639 28713 2651 28747
rect 2593 28707 2651 28713
rect 1854 28676 1860 28688
rect 1815 28648 1860 28676
rect 1854 28636 1860 28648
rect 1912 28636 1918 28688
rect 2608 28676 2636 28707
rect 4338 28704 4344 28756
rect 4396 28744 4402 28756
rect 4433 28747 4491 28753
rect 4433 28744 4445 28747
rect 4396 28716 4445 28744
rect 4396 28704 4402 28716
rect 4433 28713 4445 28716
rect 4479 28713 4491 28747
rect 4433 28707 4491 28713
rect 4798 28704 4804 28756
rect 4856 28744 4862 28756
rect 5077 28747 5135 28753
rect 5077 28744 5089 28747
rect 4856 28716 5089 28744
rect 4856 28704 4862 28716
rect 5077 28713 5089 28716
rect 5123 28713 5135 28747
rect 5810 28744 5816 28756
rect 5771 28716 5816 28744
rect 5077 28707 5135 28713
rect 5810 28704 5816 28716
rect 5868 28704 5874 28756
rect 7926 28744 7932 28756
rect 5920 28716 7696 28744
rect 7887 28716 7932 28744
rect 4522 28676 4528 28688
rect 2608 28648 3372 28676
rect 2130 28568 2136 28620
rect 2188 28608 2194 28620
rect 3344 28617 3372 28648
rect 4356 28648 4528 28676
rect 4356 28617 4384 28648
rect 4522 28636 4528 28648
rect 4580 28676 4586 28688
rect 5258 28676 5264 28688
rect 4580 28648 5264 28676
rect 4580 28636 4586 28648
rect 5258 28636 5264 28648
rect 5316 28636 5322 28688
rect 5920 28676 5948 28716
rect 7558 28676 7564 28688
rect 5460 28648 5948 28676
rect 7208 28648 7564 28676
rect 2501 28611 2559 28617
rect 2501 28608 2513 28611
rect 2188 28580 2513 28608
rect 2188 28568 2194 28580
rect 2501 28577 2513 28580
rect 2547 28577 2559 28611
rect 2501 28571 2559 28577
rect 3145 28611 3203 28617
rect 3145 28577 3157 28611
rect 3191 28577 3203 28611
rect 3145 28571 3203 28577
rect 3329 28611 3387 28617
rect 3329 28577 3341 28611
rect 3375 28577 3387 28611
rect 3329 28571 3387 28577
rect 4341 28611 4399 28617
rect 4341 28577 4353 28611
rect 4387 28577 4399 28611
rect 4982 28608 4988 28620
rect 4943 28580 4988 28608
rect 4341 28571 4399 28577
rect 3160 28540 3188 28571
rect 4982 28568 4988 28580
rect 5040 28568 5046 28620
rect 5460 28552 5488 28648
rect 5721 28611 5779 28617
rect 5721 28577 5733 28611
rect 5767 28577 5779 28611
rect 5721 28571 5779 28577
rect 5905 28611 5963 28617
rect 5905 28577 5917 28611
rect 5951 28608 5963 28611
rect 7098 28608 7104 28620
rect 5951 28580 6960 28608
rect 7059 28580 7104 28608
rect 5951 28577 5963 28580
rect 5905 28571 5963 28577
rect 5166 28540 5172 28552
rect 3160 28512 5172 28540
rect 5166 28500 5172 28512
rect 5224 28500 5230 28552
rect 5442 28500 5448 28552
rect 5500 28500 5506 28552
rect 5736 28540 5764 28571
rect 6178 28540 6184 28552
rect 5736 28512 6184 28540
rect 6178 28500 6184 28512
rect 6236 28500 6242 28552
rect 6932 28540 6960 28580
rect 7098 28568 7104 28580
rect 7156 28568 7162 28620
rect 7208 28617 7236 28648
rect 7558 28636 7564 28648
rect 7616 28636 7622 28688
rect 7668 28676 7696 28716
rect 7926 28704 7932 28716
rect 7984 28704 7990 28756
rect 8389 28747 8447 28753
rect 8389 28713 8401 28747
rect 8435 28744 8447 28747
rect 9125 28747 9183 28753
rect 9125 28744 9137 28747
rect 8435 28716 9137 28744
rect 8435 28713 8447 28716
rect 8389 28707 8447 28713
rect 9125 28713 9137 28716
rect 9171 28713 9183 28747
rect 9125 28707 9183 28713
rect 9493 28747 9551 28753
rect 9493 28713 9505 28747
rect 9539 28744 9551 28747
rect 9674 28744 9680 28756
rect 9539 28716 9680 28744
rect 9539 28713 9551 28716
rect 9493 28707 9551 28713
rect 9674 28704 9680 28716
rect 9732 28704 9738 28756
rect 9858 28704 9864 28756
rect 9916 28744 9922 28756
rect 10781 28747 10839 28753
rect 10781 28744 10793 28747
rect 9916 28716 10793 28744
rect 9916 28704 9922 28716
rect 10781 28713 10793 28716
rect 10827 28713 10839 28747
rect 10781 28707 10839 28713
rect 11054 28704 11060 28756
rect 11112 28744 11118 28756
rect 12161 28747 12219 28753
rect 12161 28744 12173 28747
rect 11112 28716 12173 28744
rect 11112 28704 11118 28716
rect 12161 28713 12173 28716
rect 12207 28713 12219 28747
rect 21266 28744 21272 28756
rect 12161 28707 12219 28713
rect 12406 28716 21272 28744
rect 10686 28676 10692 28688
rect 7668 28648 8432 28676
rect 10647 28648 10692 28676
rect 7193 28611 7251 28617
rect 7193 28577 7205 28611
rect 7239 28577 7251 28611
rect 7193 28571 7251 28577
rect 7285 28611 7343 28617
rect 7285 28577 7297 28611
rect 7331 28608 7343 28611
rect 7466 28608 7472 28620
rect 7331 28580 7472 28608
rect 7331 28577 7343 28580
rect 7285 28571 7343 28577
rect 7466 28568 7472 28580
rect 7524 28568 7530 28620
rect 8294 28608 8300 28620
rect 8255 28580 8300 28608
rect 8294 28568 8300 28580
rect 8352 28568 8358 28620
rect 8404 28608 8432 28648
rect 10686 28636 10692 28648
rect 10744 28636 10750 28688
rect 12406 28676 12434 28716
rect 21266 28704 21272 28716
rect 21324 28704 21330 28756
rect 25130 28704 25136 28756
rect 25188 28704 25194 28756
rect 26694 28704 26700 28756
rect 26752 28744 26758 28756
rect 26789 28747 26847 28753
rect 26789 28744 26801 28747
rect 26752 28716 26801 28744
rect 26752 28704 26758 28716
rect 26789 28713 26801 28716
rect 26835 28713 26847 28747
rect 26789 28707 26847 28713
rect 10796 28648 12434 28676
rect 10796 28608 10824 28648
rect 12802 28636 12808 28688
rect 12860 28676 12866 28688
rect 13817 28679 13875 28685
rect 13817 28676 13829 28679
rect 12860 28648 13829 28676
rect 12860 28636 12866 28648
rect 13817 28645 13829 28648
rect 13863 28645 13875 28679
rect 13817 28639 13875 28645
rect 14090 28636 14096 28688
rect 14148 28676 14154 28688
rect 15473 28679 15531 28685
rect 15473 28676 15485 28679
rect 14148 28648 15485 28676
rect 14148 28636 14154 28648
rect 15473 28645 15485 28648
rect 15519 28645 15531 28679
rect 25148 28676 25176 28704
rect 25654 28679 25712 28685
rect 25654 28676 25666 28679
rect 15473 28639 15531 28645
rect 24780 28648 25176 28676
rect 25424 28648 25666 28676
rect 8404 28580 10824 28608
rect 11330 28568 11336 28620
rect 11388 28608 11394 28620
rect 12069 28611 12127 28617
rect 12069 28608 12081 28611
rect 11388 28580 12081 28608
rect 11388 28568 11394 28580
rect 12069 28577 12081 28580
rect 12115 28577 12127 28611
rect 12069 28571 12127 28577
rect 13725 28611 13783 28617
rect 13725 28577 13737 28611
rect 13771 28577 13783 28611
rect 13725 28571 13783 28577
rect 14001 28611 14059 28617
rect 14001 28577 14013 28611
rect 14047 28577 14059 28611
rect 14182 28608 14188 28620
rect 14143 28580 14188 28608
rect 14001 28571 14059 28577
rect 7374 28540 7380 28552
rect 6932 28512 7380 28540
rect 7374 28500 7380 28512
rect 7432 28500 7438 28552
rect 8570 28540 8576 28552
rect 8531 28512 8576 28540
rect 8570 28500 8576 28512
rect 8628 28500 8634 28552
rect 9585 28543 9643 28549
rect 9585 28509 9597 28543
rect 9631 28509 9643 28543
rect 9766 28540 9772 28552
rect 9727 28512 9772 28540
rect 9585 28503 9643 28509
rect 2038 28472 2044 28484
rect 1951 28444 2044 28472
rect 2038 28432 2044 28444
rect 2096 28472 2102 28484
rect 2096 28444 4016 28472
rect 2096 28432 2102 28444
rect 3142 28364 3148 28416
rect 3200 28404 3206 28416
rect 3237 28407 3295 28413
rect 3237 28404 3249 28407
rect 3200 28376 3249 28404
rect 3200 28364 3206 28376
rect 3237 28373 3249 28376
rect 3283 28373 3295 28407
rect 3988 28404 4016 28444
rect 4062 28432 4068 28484
rect 4120 28472 4126 28484
rect 4522 28472 4528 28484
rect 4120 28444 4528 28472
rect 4120 28432 4126 28444
rect 4522 28432 4528 28444
rect 4580 28432 4586 28484
rect 4632 28444 5396 28472
rect 4632 28404 4660 28444
rect 3988 28376 4660 28404
rect 5368 28404 5396 28444
rect 6638 28432 6644 28484
rect 6696 28472 6702 28484
rect 9600 28472 9628 28503
rect 9766 28500 9772 28512
rect 9824 28500 9830 28552
rect 10965 28543 11023 28549
rect 10965 28509 10977 28543
rect 11011 28540 11023 28543
rect 11054 28540 11060 28552
rect 11011 28512 11060 28540
rect 11011 28509 11023 28512
rect 10965 28503 11023 28509
rect 11054 28500 11060 28512
rect 11112 28500 11118 28552
rect 13740 28540 13768 28571
rect 13648 28512 13768 28540
rect 14016 28540 14044 28571
rect 14182 28568 14188 28580
rect 14240 28568 14246 28620
rect 15197 28611 15255 28617
rect 15197 28577 15209 28611
rect 15243 28608 15255 28611
rect 15243 28580 15700 28608
rect 15243 28577 15255 28580
rect 15197 28571 15255 28577
rect 14274 28540 14280 28552
rect 14016 28512 14280 28540
rect 9858 28472 9864 28484
rect 6696 28444 9536 28472
rect 9600 28444 9864 28472
rect 6696 28432 6702 28444
rect 6362 28404 6368 28416
rect 5368 28376 6368 28404
rect 3237 28367 3295 28373
rect 6362 28364 6368 28376
rect 6420 28364 6426 28416
rect 7098 28364 7104 28416
rect 7156 28404 7162 28416
rect 7469 28407 7527 28413
rect 7469 28404 7481 28407
rect 7156 28376 7481 28404
rect 7156 28364 7162 28376
rect 7469 28373 7481 28376
rect 7515 28373 7527 28407
rect 9508 28404 9536 28444
rect 9858 28432 9864 28444
rect 9916 28432 9922 28484
rect 10321 28475 10379 28481
rect 10321 28441 10333 28475
rect 10367 28472 10379 28475
rect 10778 28472 10784 28484
rect 10367 28444 10784 28472
rect 10367 28441 10379 28444
rect 10321 28435 10379 28441
rect 10778 28432 10784 28444
rect 10836 28432 10842 28484
rect 12802 28404 12808 28416
rect 9508 28376 12808 28404
rect 7469 28367 7527 28373
rect 12802 28364 12808 28376
rect 12860 28364 12866 28416
rect 13648 28404 13676 28512
rect 14274 28500 14280 28512
rect 14332 28500 14338 28552
rect 15470 28540 15476 28552
rect 15431 28512 15476 28540
rect 15470 28500 15476 28512
rect 15528 28500 15534 28552
rect 15672 28540 15700 28580
rect 16022 28568 16028 28620
rect 16080 28608 16086 28620
rect 16390 28608 16396 28620
rect 16080 28580 16396 28608
rect 16080 28568 16086 28580
rect 16390 28568 16396 28580
rect 16448 28568 16454 28620
rect 18966 28608 18972 28620
rect 18927 28580 18972 28608
rect 18966 28568 18972 28580
rect 19024 28568 19030 28620
rect 20254 28617 20260 28620
rect 20248 28571 20260 28617
rect 20312 28608 20318 28620
rect 24780 28617 24808 28648
rect 24765 28611 24823 28617
rect 20312 28580 20348 28608
rect 20254 28568 20260 28571
rect 20312 28568 20318 28580
rect 24765 28577 24777 28611
rect 24811 28577 24823 28611
rect 24765 28571 24823 28577
rect 24949 28611 25007 28617
rect 24949 28577 24961 28611
rect 24995 28577 25007 28611
rect 24949 28571 25007 28577
rect 16206 28540 16212 28552
rect 15672 28512 16212 28540
rect 16206 28500 16212 28512
rect 16264 28500 16270 28552
rect 19334 28500 19340 28552
rect 19392 28540 19398 28552
rect 19981 28543 20039 28549
rect 19981 28540 19993 28543
rect 19392 28512 19993 28540
rect 19392 28500 19398 28512
rect 19981 28509 19993 28512
rect 20027 28509 20039 28543
rect 19981 28503 20039 28509
rect 24854 28500 24860 28552
rect 24912 28500 24918 28552
rect 24964 28540 24992 28571
rect 25130 28568 25136 28620
rect 25188 28608 25194 28620
rect 25424 28608 25452 28648
rect 25654 28645 25666 28648
rect 25700 28645 25712 28679
rect 25654 28639 25712 28645
rect 26142 28608 26148 28620
rect 25188 28580 25452 28608
rect 25516 28580 26148 28608
rect 25188 28568 25194 28580
rect 25222 28540 25228 28552
rect 24964 28512 25228 28540
rect 25222 28500 25228 28512
rect 25280 28500 25286 28552
rect 25409 28543 25467 28549
rect 25409 28509 25421 28543
rect 25455 28540 25467 28543
rect 25516 28540 25544 28580
rect 26142 28568 26148 28580
rect 26200 28568 26206 28620
rect 27982 28608 27988 28620
rect 27943 28580 27988 28608
rect 27982 28568 27988 28580
rect 28040 28568 28046 28620
rect 25455 28512 25544 28540
rect 25455 28509 25467 28512
rect 25409 28503 25467 28509
rect 13722 28432 13728 28484
rect 13780 28472 13786 28484
rect 15289 28475 15347 28481
rect 15289 28472 15301 28475
rect 13780 28444 15301 28472
rect 13780 28432 13786 28444
rect 15289 28441 15301 28444
rect 15335 28441 15347 28475
rect 15289 28435 15347 28441
rect 19153 28475 19211 28481
rect 19153 28441 19165 28475
rect 19199 28472 19211 28475
rect 19242 28472 19248 28484
rect 19199 28444 19248 28472
rect 19199 28441 19211 28444
rect 19153 28435 19211 28441
rect 19242 28432 19248 28444
rect 19300 28432 19306 28484
rect 24872 28472 24900 28500
rect 28169 28475 28227 28481
rect 24872 28444 24992 28472
rect 15930 28404 15936 28416
rect 13648 28376 15936 28404
rect 15930 28364 15936 28376
rect 15988 28364 15994 28416
rect 21358 28404 21364 28416
rect 21319 28376 21364 28404
rect 21358 28364 21364 28376
rect 21416 28404 21422 28416
rect 22922 28404 22928 28416
rect 21416 28376 22928 28404
rect 21416 28364 21422 28376
rect 22922 28364 22928 28376
rect 22980 28364 22986 28416
rect 24854 28404 24860 28416
rect 24815 28376 24860 28404
rect 24854 28364 24860 28376
rect 24912 28364 24918 28416
rect 24964 28404 24992 28444
rect 28169 28441 28181 28475
rect 28215 28472 28227 28475
rect 28258 28472 28264 28484
rect 28215 28444 28264 28472
rect 28215 28441 28227 28444
rect 28169 28435 28227 28441
rect 28258 28432 28264 28444
rect 28316 28432 28322 28484
rect 26050 28404 26056 28416
rect 24964 28376 26056 28404
rect 26050 28364 26056 28376
rect 26108 28364 26114 28416
rect 1104 28314 28888 28336
rect 1104 28262 5614 28314
rect 5666 28262 5678 28314
rect 5730 28262 5742 28314
rect 5794 28262 5806 28314
rect 5858 28262 14878 28314
rect 14930 28262 14942 28314
rect 14994 28262 15006 28314
rect 15058 28262 15070 28314
rect 15122 28262 24142 28314
rect 24194 28262 24206 28314
rect 24258 28262 24270 28314
rect 24322 28262 24334 28314
rect 24386 28262 28888 28314
rect 1104 28240 28888 28262
rect 2498 28160 2504 28212
rect 2556 28200 2562 28212
rect 2685 28203 2743 28209
rect 2685 28200 2697 28203
rect 2556 28172 2697 28200
rect 2556 28160 2562 28172
rect 2685 28169 2697 28172
rect 2731 28169 2743 28203
rect 2685 28163 2743 28169
rect 4890 28160 4896 28212
rect 4948 28200 4954 28212
rect 5077 28203 5135 28209
rect 5077 28200 5089 28203
rect 4948 28172 5089 28200
rect 4948 28160 4954 28172
rect 5077 28169 5089 28172
rect 5123 28200 5135 28203
rect 5442 28200 5448 28212
rect 5123 28172 5448 28200
rect 5123 28169 5135 28172
rect 5077 28163 5135 28169
rect 5442 28160 5448 28172
rect 5500 28160 5506 28212
rect 6178 28200 6184 28212
rect 6139 28172 6184 28200
rect 6178 28160 6184 28172
rect 6236 28160 6242 28212
rect 6822 28200 6828 28212
rect 6748 28172 6828 28200
rect 1762 28132 1768 28144
rect 1723 28104 1768 28132
rect 1762 28092 1768 28104
rect 1820 28092 1826 28144
rect 6748 28132 6776 28172
rect 6822 28160 6828 28172
rect 6880 28160 6886 28212
rect 7374 28160 7380 28212
rect 7432 28160 7438 28212
rect 7926 28200 7932 28212
rect 7887 28172 7932 28200
rect 7926 28160 7932 28172
rect 7984 28160 7990 28212
rect 10137 28203 10195 28209
rect 10137 28169 10149 28203
rect 10183 28200 10195 28203
rect 11330 28200 11336 28212
rect 10183 28172 11336 28200
rect 10183 28169 10195 28172
rect 10137 28163 10195 28169
rect 11330 28160 11336 28172
rect 11388 28160 11394 28212
rect 12802 28160 12808 28212
rect 12860 28200 12866 28212
rect 17221 28203 17279 28209
rect 17221 28200 17233 28203
rect 12860 28172 17233 28200
rect 12860 28160 12866 28172
rect 7392 28132 7420 28160
rect 6104 28104 6776 28132
rect 6840 28104 7420 28132
rect 3142 28064 3148 28076
rect 3103 28036 3148 28064
rect 3142 28024 3148 28036
rect 3200 28024 3206 28076
rect 3786 28024 3792 28076
rect 3844 28064 3850 28076
rect 3844 28036 4936 28064
rect 3844 28024 3850 28036
rect 1946 27996 1952 28008
rect 1907 27968 1952 27996
rect 1946 27956 1952 27968
rect 2004 27956 2010 28008
rect 4246 27996 4252 28008
rect 4207 27968 4252 27996
rect 4246 27956 4252 27968
rect 4304 27956 4310 28008
rect 4908 28005 4936 28036
rect 6104 28005 6132 28104
rect 4893 27999 4951 28005
rect 4893 27965 4905 27999
rect 4939 27965 4951 27999
rect 4893 27959 4951 27965
rect 6089 27999 6147 28005
rect 6089 27965 6101 27999
rect 6135 27965 6147 27999
rect 6089 27959 6147 27965
rect 6273 27999 6331 28005
rect 6273 27965 6285 27999
rect 6319 27996 6331 27999
rect 6730 27996 6736 28008
rect 6319 27968 6736 27996
rect 6319 27965 6331 27968
rect 6273 27959 6331 27965
rect 6730 27956 6736 27968
rect 6788 27956 6794 28008
rect 3234 27928 3240 27940
rect 3195 27900 3240 27928
rect 3234 27888 3240 27900
rect 3292 27888 3298 27940
rect 3142 27860 3148 27872
rect 3103 27832 3148 27860
rect 3142 27820 3148 27832
rect 3200 27820 3206 27872
rect 4338 27860 4344 27872
rect 4299 27832 4344 27860
rect 4338 27820 4344 27832
rect 4396 27820 4402 27872
rect 6733 27863 6791 27869
rect 6733 27829 6745 27863
rect 6779 27860 6791 27863
rect 6840 27860 6868 28104
rect 11422 28092 11428 28144
rect 11480 28132 11486 28144
rect 12253 28135 12311 28141
rect 12253 28132 12265 28135
rect 11480 28104 12265 28132
rect 11480 28092 11486 28104
rect 12253 28101 12265 28104
rect 12299 28101 12311 28135
rect 12253 28095 12311 28101
rect 14642 28092 14648 28144
rect 14700 28132 14706 28144
rect 14918 28132 14924 28144
rect 14700 28104 14924 28132
rect 14700 28092 14706 28104
rect 14918 28092 14924 28104
rect 14976 28092 14982 28144
rect 7374 28024 7380 28076
rect 7432 28064 7438 28076
rect 10781 28067 10839 28073
rect 7432 28036 10548 28064
rect 7432 28024 7438 28036
rect 6917 27999 6975 28005
rect 6917 27965 6929 27999
rect 6963 27965 6975 27999
rect 7098 27996 7104 28008
rect 7059 27968 7104 27996
rect 6917 27959 6975 27965
rect 6932 27928 6960 27959
rect 7098 27956 7104 27968
rect 7156 27956 7162 28008
rect 7190 27956 7196 28008
rect 7248 27996 7254 28008
rect 7650 27996 7656 28008
rect 7248 27968 7293 27996
rect 7611 27968 7656 27996
rect 7248 27956 7254 27968
rect 7650 27956 7656 27968
rect 7708 27956 7714 28008
rect 8754 27956 8760 28008
rect 8812 27996 8818 28008
rect 9490 27996 9496 28008
rect 8812 27968 9496 27996
rect 8812 27956 8818 27968
rect 9490 27956 9496 27968
rect 9548 27956 9554 28008
rect 10520 28005 10548 28036
rect 10781 28033 10793 28067
rect 10827 28064 10839 28067
rect 11054 28064 11060 28076
rect 10827 28036 11060 28064
rect 10827 28033 10839 28036
rect 10781 28027 10839 28033
rect 11054 28024 11060 28036
rect 11112 28064 11118 28076
rect 11330 28064 11336 28076
rect 11112 28036 11336 28064
rect 11112 28024 11118 28036
rect 11330 28024 11336 28036
rect 11388 28024 11394 28076
rect 12069 28067 12127 28073
rect 12069 28033 12081 28067
rect 12115 28064 12127 28067
rect 12342 28064 12348 28076
rect 12115 28036 12348 28064
rect 12115 28033 12127 28036
rect 12069 28027 12127 28033
rect 12342 28024 12348 28036
rect 12400 28024 12406 28076
rect 12526 28024 12532 28076
rect 12584 28064 12590 28076
rect 14090 28064 14096 28076
rect 12584 28036 14096 28064
rect 12584 28024 12590 28036
rect 14090 28024 14096 28036
rect 14148 28024 14154 28076
rect 16206 28024 16212 28076
rect 16264 28064 16270 28076
rect 16669 28067 16727 28073
rect 16669 28064 16681 28067
rect 16264 28036 16681 28064
rect 16264 28024 16270 28036
rect 16669 28033 16681 28036
rect 16715 28033 16727 28067
rect 16669 28027 16727 28033
rect 10505 27999 10563 28005
rect 10505 27965 10517 27999
rect 10551 27965 10563 27999
rect 10505 27959 10563 27965
rect 11422 27956 11428 28008
rect 11480 27996 11486 28008
rect 11606 27996 11612 28008
rect 11480 27968 11612 27996
rect 11480 27956 11486 27968
rect 11606 27956 11612 27968
rect 11664 27956 11670 28008
rect 11974 27996 11980 28008
rect 11935 27968 11980 27996
rect 11974 27956 11980 27968
rect 12032 27956 12038 28008
rect 13081 27999 13139 28005
rect 13081 27965 13093 27999
rect 13127 27996 13139 27999
rect 13262 27996 13268 28008
rect 13127 27968 13268 27996
rect 13127 27965 13139 27968
rect 13081 27959 13139 27965
rect 13262 27956 13268 27968
rect 13320 27956 13326 28008
rect 15194 27956 15200 28008
rect 15252 27996 15258 28008
rect 15289 27999 15347 28005
rect 15289 27996 15301 27999
rect 15252 27968 15301 27996
rect 15252 27956 15258 27968
rect 15289 27965 15301 27968
rect 15335 27965 15347 27999
rect 15562 27996 15568 28008
rect 15523 27968 15568 27996
rect 15289 27959 15347 27965
rect 15562 27956 15568 27968
rect 15620 27956 15626 28008
rect 17144 27996 17172 28172
rect 17221 28169 17233 28172
rect 17267 28169 17279 28203
rect 17221 28163 17279 28169
rect 19429 28203 19487 28209
rect 19429 28169 19441 28203
rect 19475 28200 19487 28203
rect 20162 28200 20168 28212
rect 19475 28172 20168 28200
rect 19475 28169 19487 28172
rect 19429 28163 19487 28169
rect 20162 28160 20168 28172
rect 20220 28160 20226 28212
rect 24213 28203 24271 28209
rect 24213 28169 24225 28203
rect 24259 28200 24271 28203
rect 25130 28200 25136 28212
rect 24259 28172 25136 28200
rect 24259 28169 24271 28172
rect 24213 28163 24271 28169
rect 25130 28160 25136 28172
rect 25188 28160 25194 28212
rect 27982 28200 27988 28212
rect 27943 28172 27988 28200
rect 27982 28160 27988 28172
rect 28040 28160 28046 28212
rect 17494 28132 17500 28144
rect 17420 28104 17500 28132
rect 17218 28024 17224 28076
rect 17276 28064 17282 28076
rect 17420 28064 17448 28104
rect 17494 28092 17500 28104
rect 17552 28092 17558 28144
rect 17276 28050 17448 28064
rect 19984 28076 20036 28082
rect 17276 28036 17434 28050
rect 17276 28024 17282 28036
rect 25222 28064 25228 28076
rect 19984 28018 20036 28024
rect 23860 28036 25228 28064
rect 17862 27996 17868 28008
rect 17144 27968 17868 27996
rect 17862 27956 17868 27968
rect 17920 27956 17926 28008
rect 18064 27968 19932 27996
rect 6932 27900 8248 27928
rect 8220 27872 8248 27900
rect 9214 27888 9220 27940
rect 9272 27928 9278 27940
rect 10597 27931 10655 27937
rect 10597 27928 10609 27931
rect 9272 27900 10609 27928
rect 9272 27888 9278 27900
rect 10597 27897 10609 27900
rect 10643 27928 10655 27931
rect 10643 27900 15240 27928
rect 10643 27897 10655 27900
rect 10597 27891 10655 27897
rect 6779 27832 6868 27860
rect 6779 27829 6791 27832
rect 6733 27823 6791 27829
rect 6914 27820 6920 27872
rect 6972 27860 6978 27872
rect 7742 27860 7748 27872
rect 6972 27832 7748 27860
rect 6972 27820 6978 27832
rect 7742 27820 7748 27832
rect 7800 27860 7806 27872
rect 8113 27863 8171 27869
rect 8113 27860 8125 27863
rect 7800 27832 8125 27860
rect 7800 27820 7806 27832
rect 8113 27829 8125 27832
rect 8159 27829 8171 27863
rect 8113 27823 8171 27829
rect 8202 27820 8208 27872
rect 8260 27860 8266 27872
rect 9585 27863 9643 27869
rect 9585 27860 9597 27863
rect 8260 27832 9597 27860
rect 8260 27820 8266 27832
rect 9585 27829 9597 27832
rect 9631 27829 9643 27863
rect 11606 27860 11612 27872
rect 11567 27832 11612 27860
rect 9585 27823 9643 27829
rect 11606 27820 11612 27832
rect 11664 27820 11670 27872
rect 12526 27820 12532 27872
rect 12584 27860 12590 27872
rect 13173 27863 13231 27869
rect 13173 27860 13185 27863
rect 12584 27832 13185 27860
rect 12584 27820 12590 27832
rect 13173 27829 13185 27832
rect 13219 27860 13231 27863
rect 13446 27860 13452 27872
rect 13219 27832 13452 27860
rect 13219 27829 13231 27832
rect 13173 27823 13231 27829
rect 13446 27820 13452 27832
rect 13504 27860 13510 27872
rect 13814 27860 13820 27872
rect 13504 27832 13820 27860
rect 13504 27820 13510 27832
rect 13814 27820 13820 27832
rect 13872 27820 13878 27872
rect 15212 27860 15240 27900
rect 17678 27888 17684 27940
rect 17736 27928 17742 27940
rect 17957 27931 18015 27937
rect 17957 27928 17969 27931
rect 17736 27900 17969 27928
rect 17736 27888 17742 27900
rect 17957 27897 17969 27900
rect 18003 27897 18015 27931
rect 17957 27891 18015 27897
rect 17589 27863 17647 27869
rect 17589 27860 17601 27863
rect 15212 27832 17601 27860
rect 17589 27829 17601 27832
rect 17635 27860 17647 27863
rect 18064 27860 18092 27968
rect 18325 27931 18383 27937
rect 18325 27897 18337 27931
rect 18371 27928 18383 27931
rect 19429 27931 19487 27937
rect 19429 27928 19441 27931
rect 18371 27900 19441 27928
rect 18371 27897 18383 27900
rect 18325 27891 18383 27897
rect 19429 27897 19441 27900
rect 19475 27897 19487 27931
rect 19429 27891 19487 27897
rect 17635 27832 18092 27860
rect 17635 27829 17647 27832
rect 17589 27823 17647 27829
rect 18506 27820 18512 27872
rect 18564 27860 18570 27872
rect 18693 27863 18751 27869
rect 18693 27860 18705 27863
rect 18564 27832 18705 27860
rect 18564 27820 18570 27832
rect 18693 27829 18705 27832
rect 18739 27829 18751 27863
rect 18874 27860 18880 27872
rect 18835 27832 18880 27860
rect 18693 27823 18751 27829
rect 18874 27820 18880 27832
rect 18932 27820 18938 27872
rect 19904 27860 19932 27968
rect 20070 27956 20076 28008
rect 20128 27996 20134 28008
rect 20901 27999 20959 28005
rect 20901 27996 20913 27999
rect 20128 27968 20913 27996
rect 20128 27956 20134 27968
rect 20901 27965 20913 27968
rect 20947 27996 20959 27999
rect 21358 27996 21364 28008
rect 20947 27968 21364 27996
rect 20947 27965 20959 27968
rect 20901 27959 20959 27965
rect 21358 27956 21364 27968
rect 21416 27956 21422 28008
rect 23860 28005 23888 28036
rect 25222 28024 25228 28036
rect 25280 28024 25286 28076
rect 27982 28064 27988 28076
rect 25700 28008 25728 28050
rect 27172 28036 27988 28064
rect 24026 28005 24032 28008
rect 23845 27999 23903 28005
rect 23845 27965 23857 27999
rect 23891 27965 23903 27999
rect 23845 27959 23903 27965
rect 23983 27999 24032 28005
rect 23983 27965 23995 27999
rect 24029 27965 24032 27999
rect 23983 27959 24032 27965
rect 24026 27956 24032 27959
rect 24084 27956 24090 28008
rect 24118 27956 24124 28008
rect 24176 27996 24182 28008
rect 24305 27999 24363 28005
rect 24176 27968 24221 27996
rect 24176 27956 24182 27968
rect 24305 27965 24317 27999
rect 24351 27996 24363 27999
rect 24854 27996 24860 28008
rect 24351 27968 24860 27996
rect 24351 27965 24363 27968
rect 24305 27959 24363 27965
rect 24854 27956 24860 27968
rect 24912 27956 24918 28008
rect 25682 27956 25688 28008
rect 25740 27956 25746 28008
rect 26329 27999 26387 28005
rect 25792 27968 26280 27996
rect 20162 27928 20168 27940
rect 20123 27900 20168 27928
rect 20162 27888 20168 27900
rect 20220 27888 20226 27940
rect 20438 27928 20444 27940
rect 20399 27900 20444 27928
rect 20438 27888 20444 27900
rect 20496 27888 20502 27940
rect 20530 27888 20536 27940
rect 20588 27928 20594 27940
rect 21266 27928 21272 27940
rect 20588 27900 20633 27928
rect 21227 27900 21272 27928
rect 20588 27888 20594 27900
rect 21266 27888 21272 27900
rect 21324 27888 21330 27940
rect 25792 27928 25820 27968
rect 22066 27900 25820 27928
rect 25869 27931 25927 27937
rect 21082 27860 21088 27872
rect 19904 27832 21088 27860
rect 21082 27820 21088 27832
rect 21140 27820 21146 27872
rect 21453 27863 21511 27869
rect 21453 27829 21465 27863
rect 21499 27860 21511 27863
rect 21634 27860 21640 27872
rect 21499 27832 21640 27860
rect 21499 27829 21511 27832
rect 21453 27823 21511 27829
rect 21634 27820 21640 27832
rect 21692 27820 21698 27872
rect 21726 27820 21732 27872
rect 21784 27860 21790 27872
rect 22066 27860 22094 27900
rect 25869 27897 25881 27931
rect 25915 27897 25927 27931
rect 25869 27891 25927 27897
rect 21784 27832 22094 27860
rect 21784 27820 21790 27832
rect 23382 27820 23388 27872
rect 23440 27860 23446 27872
rect 23566 27860 23572 27872
rect 23440 27832 23572 27860
rect 23440 27820 23446 27832
rect 23566 27820 23572 27832
rect 23624 27860 23630 27872
rect 25590 27860 25596 27872
rect 23624 27832 25596 27860
rect 23624 27820 23630 27832
rect 25590 27820 25596 27832
rect 25648 27820 25654 27872
rect 25884 27860 25912 27891
rect 25958 27888 25964 27940
rect 26016 27928 26022 27940
rect 26252 27928 26280 27968
rect 26329 27965 26341 27999
rect 26375 27996 26387 27999
rect 26694 27996 26700 28008
rect 26375 27968 26700 27996
rect 26375 27965 26387 27968
rect 26329 27959 26387 27965
rect 26694 27956 26700 27968
rect 26752 27956 26758 28008
rect 27172 27928 27200 28036
rect 27982 28024 27988 28036
rect 28040 28024 28046 28076
rect 27522 27956 27528 28008
rect 27580 27996 27586 28008
rect 27709 27999 27767 28005
rect 27709 27996 27721 27999
rect 27580 27968 27721 27996
rect 27580 27956 27586 27968
rect 27709 27965 27721 27968
rect 27755 27965 27767 27999
rect 27709 27959 27767 27965
rect 26016 27900 26061 27928
rect 26252 27900 27200 27928
rect 26016 27888 26022 27900
rect 27246 27888 27252 27940
rect 27304 27928 27310 27940
rect 27433 27931 27491 27937
rect 27433 27928 27445 27931
rect 27304 27900 27445 27928
rect 27304 27888 27310 27900
rect 27433 27897 27445 27900
rect 27479 27897 27491 27931
rect 27798 27928 27804 27940
rect 27433 27891 27491 27897
rect 27540 27900 27804 27928
rect 26050 27860 26056 27872
rect 25884 27832 26056 27860
rect 26050 27820 26056 27832
rect 26108 27820 26114 27872
rect 26234 27820 26240 27872
rect 26292 27860 26298 27872
rect 26697 27863 26755 27869
rect 26697 27860 26709 27863
rect 26292 27832 26709 27860
rect 26292 27820 26298 27832
rect 26697 27829 26709 27832
rect 26743 27829 26755 27863
rect 26697 27823 26755 27829
rect 26881 27863 26939 27869
rect 26881 27829 26893 27863
rect 26927 27860 26939 27863
rect 27540 27860 27568 27900
rect 27798 27888 27804 27900
rect 27856 27888 27862 27940
rect 26927 27832 27568 27860
rect 26927 27829 26939 27832
rect 26881 27823 26939 27829
rect 27614 27820 27620 27872
rect 27672 27860 27678 27872
rect 27672 27832 27717 27860
rect 27672 27820 27678 27832
rect 1104 27770 28888 27792
rect 1104 27718 10246 27770
rect 10298 27718 10310 27770
rect 10362 27718 10374 27770
rect 10426 27718 10438 27770
rect 10490 27718 19510 27770
rect 19562 27718 19574 27770
rect 19626 27718 19638 27770
rect 19690 27718 19702 27770
rect 19754 27718 28888 27770
rect 1104 27696 28888 27718
rect 1581 27659 1639 27665
rect 1581 27625 1593 27659
rect 1627 27656 1639 27659
rect 2038 27656 2044 27668
rect 1627 27628 2044 27656
rect 1627 27625 1639 27628
rect 1581 27619 1639 27625
rect 2038 27616 2044 27628
rect 2096 27616 2102 27668
rect 3142 27616 3148 27668
rect 3200 27656 3206 27668
rect 3421 27659 3479 27665
rect 3421 27656 3433 27659
rect 3200 27628 3433 27656
rect 3200 27616 3206 27628
rect 3421 27625 3433 27628
rect 3467 27625 3479 27659
rect 7190 27656 7196 27668
rect 7151 27628 7196 27656
rect 3421 27619 3479 27625
rect 7190 27616 7196 27628
rect 7248 27616 7254 27668
rect 7650 27616 7656 27668
rect 7708 27616 7714 27668
rect 8294 27616 8300 27668
rect 8352 27656 8358 27668
rect 9125 27659 9183 27665
rect 9125 27656 9137 27659
rect 8352 27628 9137 27656
rect 8352 27616 8358 27628
rect 9125 27625 9137 27628
rect 9171 27625 9183 27659
rect 9125 27619 9183 27625
rect 11992 27628 12664 27656
rect 1762 27548 1768 27600
rect 1820 27588 1826 27600
rect 2685 27591 2743 27597
rect 2685 27588 2697 27591
rect 1820 27560 2697 27588
rect 1820 27548 1826 27560
rect 2685 27557 2697 27560
rect 2731 27557 2743 27591
rect 2685 27551 2743 27557
rect 3789 27591 3847 27597
rect 3789 27557 3801 27591
rect 3835 27588 3847 27591
rect 4338 27588 4344 27600
rect 3835 27560 4344 27588
rect 3835 27557 3847 27560
rect 3789 27551 3847 27557
rect 4338 27548 4344 27560
rect 4396 27548 4402 27600
rect 6914 27588 6920 27600
rect 6875 27560 6920 27588
rect 6914 27548 6920 27560
rect 6972 27548 6978 27600
rect 7006 27548 7012 27600
rect 7064 27588 7070 27600
rect 7101 27591 7159 27597
rect 7101 27588 7113 27591
rect 7064 27560 7113 27588
rect 7064 27548 7070 27560
rect 7101 27557 7113 27560
rect 7147 27557 7159 27591
rect 7668 27588 7696 27616
rect 8478 27588 8484 27600
rect 7668 27560 8340 27588
rect 8439 27560 8484 27588
rect 7101 27551 7159 27557
rect 1670 27480 1676 27532
rect 1728 27520 1734 27532
rect 1857 27523 1915 27529
rect 1857 27520 1869 27523
rect 1728 27492 1869 27520
rect 1728 27480 1734 27492
rect 1857 27489 1869 27492
rect 1903 27489 1915 27523
rect 1857 27483 1915 27489
rect 1949 27523 2007 27529
rect 1949 27489 1961 27523
rect 1995 27520 2007 27523
rect 2038 27520 2044 27532
rect 1995 27492 2044 27520
rect 1995 27489 2007 27492
rect 1949 27483 2007 27489
rect 2038 27480 2044 27492
rect 2096 27480 2102 27532
rect 2317 27523 2375 27529
rect 2317 27489 2329 27523
rect 2363 27520 2375 27523
rect 2406 27520 2412 27532
rect 2363 27492 2412 27520
rect 2363 27489 2375 27492
rect 2317 27483 2375 27489
rect 2406 27480 2412 27492
rect 2464 27480 2470 27532
rect 7190 27480 7196 27532
rect 7248 27520 7254 27532
rect 7653 27523 7711 27529
rect 7248 27492 7293 27520
rect 7248 27480 7254 27492
rect 7653 27489 7665 27523
rect 7699 27520 7711 27523
rect 8202 27520 8208 27532
rect 7699 27492 8208 27520
rect 7699 27489 7711 27492
rect 7653 27483 7711 27489
rect 8202 27480 8208 27492
rect 8260 27480 8266 27532
rect 8312 27520 8340 27560
rect 8478 27548 8484 27560
rect 8536 27588 8542 27600
rect 8536 27560 9260 27588
rect 8536 27548 8542 27560
rect 8389 27523 8447 27529
rect 8389 27520 8401 27523
rect 8312 27492 8401 27520
rect 8389 27489 8401 27492
rect 8435 27489 8447 27523
rect 8389 27483 8447 27489
rect 8662 27480 8668 27532
rect 8720 27520 8726 27532
rect 9232 27529 9260 27560
rect 10870 27548 10876 27600
rect 10928 27588 10934 27600
rect 11992 27588 12020 27628
rect 10928 27560 12020 27588
rect 12069 27591 12127 27597
rect 10928 27548 10934 27560
rect 12069 27557 12081 27591
rect 12115 27588 12127 27591
rect 12636 27588 12664 27628
rect 17862 27616 17868 27668
rect 17920 27656 17926 27668
rect 17920 27628 20024 27656
rect 17920 27616 17926 27628
rect 12713 27591 12771 27597
rect 12713 27588 12725 27591
rect 12115 27560 12572 27588
rect 12636 27560 12725 27588
rect 12115 27557 12127 27560
rect 12069 27551 12127 27557
rect 9033 27523 9091 27529
rect 9033 27520 9045 27523
rect 8720 27492 9045 27520
rect 8720 27480 8726 27492
rect 9033 27489 9045 27492
rect 9079 27489 9091 27523
rect 9033 27483 9091 27489
rect 9217 27523 9275 27529
rect 9217 27489 9229 27523
rect 9263 27489 9275 27523
rect 9217 27483 9275 27489
rect 11698 27480 11704 27532
rect 11756 27520 11762 27532
rect 12437 27523 12495 27529
rect 12437 27520 12449 27523
rect 11756 27492 12449 27520
rect 11756 27480 11762 27492
rect 12437 27489 12449 27492
rect 12483 27489 12495 27523
rect 12544 27520 12572 27560
rect 12713 27557 12725 27560
rect 12759 27557 12771 27591
rect 13814 27588 13820 27600
rect 12713 27551 12771 27557
rect 13372 27560 13820 27588
rect 12544 27492 12664 27520
rect 12437 27483 12495 27489
rect 2682 27452 2688 27464
rect 2622 27424 2688 27452
rect 2682 27412 2688 27424
rect 2740 27412 2746 27464
rect 3878 27452 3884 27464
rect 3839 27424 3884 27452
rect 3878 27412 3884 27424
rect 3936 27412 3942 27464
rect 3973 27455 4031 27461
rect 3973 27421 3985 27455
rect 4019 27421 4031 27455
rect 3973 27415 4031 27421
rect 3510 27344 3516 27396
rect 3568 27384 3574 27396
rect 3988 27384 4016 27415
rect 6822 27412 6828 27464
rect 6880 27452 6886 27464
rect 11517 27455 11575 27461
rect 11517 27452 11529 27455
rect 6880 27424 11529 27452
rect 6880 27412 6886 27424
rect 11517 27421 11529 27424
rect 11563 27421 11575 27455
rect 11517 27415 11575 27421
rect 12342 27412 12348 27464
rect 12400 27452 12406 27464
rect 12529 27455 12587 27461
rect 12529 27452 12541 27455
rect 12400 27424 12541 27452
rect 12400 27412 12406 27424
rect 12529 27421 12541 27424
rect 12575 27421 12587 27455
rect 12636 27452 12664 27492
rect 12802 27480 12808 27532
rect 12860 27520 12866 27532
rect 13170 27520 13176 27532
rect 12860 27492 13176 27520
rect 12860 27480 12866 27492
rect 13170 27480 13176 27492
rect 13228 27520 13234 27532
rect 13372 27529 13400 27560
rect 13814 27548 13820 27560
rect 13872 27548 13878 27600
rect 14918 27548 14924 27600
rect 14976 27588 14982 27600
rect 16209 27591 16267 27597
rect 16209 27588 16221 27591
rect 14976 27560 16221 27588
rect 14976 27548 14982 27560
rect 16209 27557 16221 27560
rect 16255 27588 16267 27591
rect 16390 27588 16396 27600
rect 16255 27560 16396 27588
rect 16255 27557 16267 27560
rect 16209 27551 16267 27557
rect 16390 27548 16396 27560
rect 16448 27548 16454 27600
rect 18874 27588 18880 27600
rect 18340 27560 18880 27588
rect 13265 27523 13323 27529
rect 13265 27520 13277 27523
rect 13228 27492 13277 27520
rect 13228 27480 13234 27492
rect 13265 27489 13277 27492
rect 13311 27489 13323 27523
rect 13265 27483 13323 27489
rect 13357 27523 13415 27529
rect 13357 27489 13369 27523
rect 13403 27489 13415 27523
rect 13357 27483 13415 27489
rect 13446 27480 13452 27532
rect 13504 27529 13510 27532
rect 13504 27523 13519 27529
rect 13507 27489 13519 27523
rect 13504 27483 13519 27489
rect 14645 27523 14703 27529
rect 14645 27489 14657 27523
rect 14691 27520 14703 27523
rect 17402 27520 17408 27532
rect 14691 27492 17408 27520
rect 14691 27489 14703 27492
rect 14645 27483 14703 27489
rect 13504 27480 13510 27483
rect 17402 27480 17408 27492
rect 17460 27480 17466 27532
rect 17494 27480 17500 27532
rect 17552 27520 17558 27532
rect 18340 27529 18368 27560
rect 18874 27548 18880 27560
rect 18932 27548 18938 27600
rect 19996 27588 20024 27628
rect 20070 27616 20076 27668
rect 20128 27656 20134 27668
rect 20165 27659 20223 27665
rect 20165 27656 20177 27659
rect 20128 27628 20177 27656
rect 20128 27616 20134 27628
rect 20165 27625 20177 27628
rect 20211 27625 20223 27659
rect 20165 27619 20223 27625
rect 20254 27616 20260 27668
rect 20312 27656 20318 27668
rect 20349 27659 20407 27665
rect 20349 27656 20361 27659
rect 20312 27628 20361 27656
rect 20312 27616 20318 27628
rect 20349 27625 20361 27628
rect 20395 27625 20407 27659
rect 21726 27656 21732 27668
rect 20349 27619 20407 27625
rect 20456 27628 21732 27656
rect 20456 27588 20484 27628
rect 21726 27616 21732 27628
rect 21784 27616 21790 27668
rect 23845 27659 23903 27665
rect 22664 27628 23060 27656
rect 19996 27560 20484 27588
rect 22554 27548 22560 27600
rect 22612 27588 22618 27600
rect 22664 27588 22692 27628
rect 22612 27560 22692 27588
rect 22741 27591 22799 27597
rect 22612 27548 22618 27560
rect 22741 27557 22753 27591
rect 22787 27588 22799 27591
rect 22922 27588 22928 27600
rect 22787 27560 22928 27588
rect 22787 27557 22799 27560
rect 22741 27551 22799 27557
rect 22922 27548 22928 27560
rect 22980 27548 22986 27600
rect 23032 27588 23060 27628
rect 23845 27625 23857 27659
rect 23891 27656 23903 27659
rect 23934 27656 23940 27668
rect 23891 27628 23940 27656
rect 23891 27625 23903 27628
rect 23845 27619 23903 27625
rect 23934 27616 23940 27628
rect 23992 27616 23998 27668
rect 24670 27616 24676 27668
rect 24728 27656 24734 27668
rect 24765 27659 24823 27665
rect 24765 27656 24777 27659
rect 24728 27628 24777 27656
rect 24728 27616 24734 27628
rect 24765 27625 24777 27628
rect 24811 27625 24823 27659
rect 24765 27619 24823 27625
rect 24857 27659 24915 27665
rect 24857 27625 24869 27659
rect 24903 27656 24915 27659
rect 24903 27628 25360 27656
rect 24903 27625 24915 27628
rect 24857 27619 24915 27625
rect 23566 27597 23572 27600
rect 23109 27591 23167 27597
rect 23109 27588 23121 27591
rect 23032 27560 23121 27588
rect 23109 27557 23121 27560
rect 23155 27557 23167 27591
rect 23109 27551 23167 27557
rect 23523 27591 23572 27597
rect 23523 27557 23535 27591
rect 23569 27557 23572 27591
rect 23523 27551 23572 27557
rect 23566 27548 23572 27551
rect 23624 27548 23630 27600
rect 24026 27548 24032 27600
rect 24084 27588 24090 27600
rect 24581 27591 24639 27597
rect 24581 27588 24593 27591
rect 24084 27560 24593 27588
rect 24084 27548 24090 27560
rect 24581 27557 24593 27560
rect 24627 27557 24639 27591
rect 25332 27588 25360 27628
rect 25958 27616 25964 27668
rect 26016 27656 26022 27668
rect 26142 27656 26148 27668
rect 26016 27628 26148 27656
rect 26016 27616 26022 27628
rect 26142 27616 26148 27628
rect 26200 27616 26206 27668
rect 27522 27616 27528 27668
rect 27580 27656 27586 27668
rect 28006 27659 28064 27665
rect 28006 27656 28018 27659
rect 27580 27628 28018 27656
rect 27580 27616 27586 27628
rect 28006 27625 28018 27628
rect 28052 27625 28064 27659
rect 28006 27619 28064 27625
rect 25685 27591 25743 27597
rect 25332 27560 25636 27588
rect 24581 27551 24639 27557
rect 17681 27523 17739 27529
rect 17681 27520 17693 27523
rect 17552 27492 17693 27520
rect 17552 27480 17558 27492
rect 17681 27489 17693 27492
rect 17727 27489 17739 27523
rect 17681 27483 17739 27489
rect 18325 27523 18383 27529
rect 18325 27489 18337 27523
rect 18371 27489 18383 27523
rect 18325 27483 18383 27489
rect 18509 27523 18567 27529
rect 18509 27489 18521 27523
rect 18555 27489 18567 27523
rect 18509 27483 18567 27489
rect 13633 27455 13691 27461
rect 13633 27452 13645 27455
rect 12636 27424 13645 27452
rect 12529 27415 12587 27421
rect 13633 27421 13645 27424
rect 13679 27421 13691 27455
rect 13633 27415 13691 27421
rect 14550 27412 14556 27464
rect 14608 27452 14614 27464
rect 15102 27452 15108 27464
rect 14608 27424 15108 27452
rect 14608 27412 14614 27424
rect 15102 27412 15108 27424
rect 15160 27412 15166 27464
rect 17773 27455 17831 27461
rect 17773 27421 17785 27455
rect 17819 27452 17831 27455
rect 18524 27452 18552 27483
rect 18782 27480 18788 27532
rect 18840 27520 18846 27532
rect 18969 27523 19027 27529
rect 18969 27520 18981 27523
rect 18840 27492 18981 27520
rect 18840 27480 18846 27492
rect 18969 27489 18981 27492
rect 19015 27489 19027 27523
rect 18969 27483 19027 27489
rect 19242 27480 19248 27532
rect 19300 27520 19306 27532
rect 20073 27523 20131 27529
rect 20073 27520 20085 27523
rect 19300 27492 20085 27520
rect 19300 27480 19306 27492
rect 20073 27489 20085 27492
rect 20119 27489 20131 27523
rect 20073 27483 20131 27489
rect 20625 27523 20683 27529
rect 20625 27489 20637 27523
rect 20671 27489 20683 27523
rect 20625 27483 20683 27489
rect 18598 27452 18604 27464
rect 17819 27424 18604 27452
rect 17819 27421 17831 27424
rect 17773 27415 17831 27421
rect 18598 27412 18604 27424
rect 18656 27412 18662 27464
rect 19613 27455 19671 27461
rect 19613 27421 19625 27455
rect 19659 27452 19671 27455
rect 20346 27452 20352 27464
rect 19659 27424 20352 27452
rect 19659 27421 19671 27424
rect 19613 27415 19671 27421
rect 20346 27412 20352 27424
rect 20404 27452 20410 27464
rect 20640 27452 20668 27483
rect 21082 27480 21088 27532
rect 21140 27520 21146 27532
rect 23017 27523 23075 27529
rect 23017 27520 23029 27523
rect 21140 27492 23029 27520
rect 21140 27480 21146 27492
rect 23017 27489 23029 27492
rect 23063 27520 23075 27523
rect 23290 27520 23296 27532
rect 23063 27492 23296 27520
rect 23063 27489 23075 27492
rect 23017 27483 23075 27489
rect 23290 27480 23296 27492
rect 23348 27480 23354 27532
rect 24949 27523 25007 27529
rect 24949 27489 24961 27523
rect 24995 27520 25007 27523
rect 24995 27492 25084 27520
rect 24995 27489 25007 27492
rect 24949 27483 25007 27489
rect 20404 27424 20668 27452
rect 20404 27412 20410 27424
rect 22462 27412 22468 27464
rect 22520 27452 22526 27464
rect 22520 27424 22586 27452
rect 22520 27412 22526 27424
rect 5074 27384 5080 27396
rect 3568 27356 4016 27384
rect 4080 27356 5080 27384
rect 3568 27344 3574 27356
rect 2869 27319 2927 27325
rect 2869 27285 2881 27319
rect 2915 27316 2927 27319
rect 4080 27316 4108 27356
rect 5074 27344 5080 27356
rect 5132 27344 5138 27396
rect 6362 27344 6368 27396
rect 6420 27384 6426 27396
rect 21450 27384 21456 27396
rect 6420 27356 21456 27384
rect 6420 27344 6426 27356
rect 21450 27344 21456 27356
rect 21508 27344 21514 27396
rect 24029 27387 24087 27393
rect 24029 27353 24041 27387
rect 24075 27384 24087 27387
rect 24854 27384 24860 27396
rect 24075 27356 24860 27384
rect 24075 27353 24087 27356
rect 24029 27347 24087 27353
rect 24854 27344 24860 27356
rect 24912 27384 24918 27396
rect 25056 27384 25084 27492
rect 24912 27356 25084 27384
rect 25133 27387 25191 27393
rect 24912 27344 24918 27356
rect 25133 27353 25145 27387
rect 25179 27384 25191 27387
rect 25179 27356 25360 27384
rect 25179 27353 25191 27356
rect 25133 27347 25191 27353
rect 25332 27328 25360 27356
rect 2915 27288 4108 27316
rect 2915 27285 2927 27288
rect 2869 27279 2927 27285
rect 4154 27276 4160 27328
rect 4212 27316 4218 27328
rect 5902 27316 5908 27328
rect 4212 27288 5908 27316
rect 4212 27276 4218 27288
rect 5902 27276 5908 27288
rect 5960 27276 5966 27328
rect 6730 27276 6736 27328
rect 6788 27316 6794 27328
rect 7374 27316 7380 27328
rect 6788 27288 7380 27316
rect 6788 27276 6794 27288
rect 7374 27276 7380 27288
rect 7432 27316 7438 27328
rect 7837 27319 7895 27325
rect 7837 27316 7849 27319
rect 7432 27288 7849 27316
rect 7432 27276 7438 27288
rect 7837 27285 7849 27288
rect 7883 27285 7895 27319
rect 7837 27279 7895 27285
rect 9674 27276 9680 27328
rect 9732 27316 9738 27328
rect 9950 27316 9956 27328
rect 9732 27288 9956 27316
rect 9732 27276 9738 27288
rect 9950 27276 9956 27288
rect 10008 27276 10014 27328
rect 11517 27319 11575 27325
rect 11517 27285 11529 27319
rect 11563 27316 11575 27319
rect 16114 27316 16120 27328
rect 11563 27288 16120 27316
rect 11563 27285 11575 27288
rect 11517 27279 11575 27285
rect 16114 27276 16120 27288
rect 16172 27276 16178 27328
rect 17862 27276 17868 27328
rect 17920 27316 17926 27328
rect 19518 27316 19524 27328
rect 17920 27288 19524 27316
rect 17920 27276 17926 27288
rect 19518 27276 19524 27288
rect 19576 27276 19582 27328
rect 20530 27316 20536 27328
rect 20491 27288 20536 27316
rect 20530 27276 20536 27288
rect 20588 27276 20594 27328
rect 25314 27276 25320 27328
rect 25372 27276 25378 27328
rect 25516 27316 25544 27560
rect 25608 27529 25636 27560
rect 25685 27557 25697 27591
rect 25731 27588 25743 27591
rect 26326 27588 26332 27600
rect 25731 27560 26332 27588
rect 25731 27557 25743 27560
rect 25685 27551 25743 27557
rect 26326 27548 26332 27560
rect 26384 27548 26390 27600
rect 26694 27588 26700 27600
rect 26655 27560 26700 27588
rect 26694 27548 26700 27560
rect 26752 27548 26758 27600
rect 27246 27548 27252 27600
rect 27304 27588 27310 27600
rect 27801 27591 27859 27597
rect 27801 27588 27813 27591
rect 27304 27560 27813 27588
rect 27304 27548 27310 27560
rect 27801 27557 27813 27560
rect 27847 27557 27859 27591
rect 27801 27551 27859 27557
rect 25593 27523 25651 27529
rect 25593 27489 25605 27523
rect 25639 27489 25651 27523
rect 25819 27523 25877 27529
rect 25819 27520 25831 27523
rect 25593 27483 25651 27489
rect 25792 27489 25831 27520
rect 25865 27489 25877 27523
rect 25792 27483 25877 27489
rect 25961 27523 26019 27529
rect 25961 27489 25973 27523
rect 26007 27520 26019 27523
rect 26234 27520 26240 27532
rect 26007 27492 26240 27520
rect 26007 27489 26019 27492
rect 25961 27483 26019 27489
rect 25792 27396 25820 27483
rect 26234 27480 26240 27492
rect 26292 27480 26298 27532
rect 25774 27344 25780 27396
rect 25832 27344 25838 27396
rect 25961 27387 26019 27393
rect 25961 27353 25973 27387
rect 26007 27384 26019 27387
rect 26418 27384 26424 27396
rect 26007 27356 26424 27384
rect 26007 27353 26019 27356
rect 25961 27347 26019 27353
rect 26418 27344 26424 27356
rect 26476 27344 26482 27396
rect 26234 27316 26240 27328
rect 25516 27288 26240 27316
rect 26234 27276 26240 27288
rect 26292 27276 26298 27328
rect 26786 27316 26792 27328
rect 26747 27288 26792 27316
rect 26786 27276 26792 27288
rect 26844 27276 26850 27328
rect 27614 27276 27620 27328
rect 27672 27316 27678 27328
rect 27985 27319 28043 27325
rect 27985 27316 27997 27319
rect 27672 27288 27997 27316
rect 27672 27276 27678 27288
rect 27985 27285 27997 27288
rect 28031 27285 28043 27319
rect 28166 27316 28172 27328
rect 28127 27288 28172 27316
rect 27985 27279 28043 27285
rect 28166 27276 28172 27288
rect 28224 27276 28230 27328
rect 1104 27226 28888 27248
rect 1104 27174 5614 27226
rect 5666 27174 5678 27226
rect 5730 27174 5742 27226
rect 5794 27174 5806 27226
rect 5858 27174 14878 27226
rect 14930 27174 14942 27226
rect 14994 27174 15006 27226
rect 15058 27174 15070 27226
rect 15122 27174 24142 27226
rect 24194 27174 24206 27226
rect 24258 27174 24270 27226
rect 24322 27174 24334 27226
rect 24386 27174 28888 27226
rect 1104 27152 28888 27174
rect 2409 27115 2467 27121
rect 2409 27081 2421 27115
rect 2455 27112 2467 27115
rect 4154 27112 4160 27124
rect 2455 27084 4160 27112
rect 2455 27081 2467 27084
rect 2409 27075 2467 27081
rect 4154 27072 4160 27084
rect 4212 27072 4218 27124
rect 5997 27115 6055 27121
rect 5997 27081 6009 27115
rect 6043 27112 6055 27115
rect 7282 27112 7288 27124
rect 6043 27084 7288 27112
rect 6043 27081 6055 27084
rect 5997 27075 6055 27081
rect 7282 27072 7288 27084
rect 7340 27072 7346 27124
rect 11054 27112 11060 27124
rect 9646 27084 11060 27112
rect 1670 27004 1676 27056
rect 1728 27044 1734 27056
rect 3237 27047 3295 27053
rect 3237 27044 3249 27047
rect 1728 27016 3249 27044
rect 1728 27004 1734 27016
rect 3237 27013 3249 27016
rect 3283 27044 3295 27047
rect 3283 27016 4476 27044
rect 3283 27013 3295 27016
rect 3237 27007 3295 27013
rect 1946 26908 1952 26920
rect 1907 26880 1952 26908
rect 1946 26868 1952 26880
rect 2004 26868 2010 26920
rect 2593 26911 2651 26917
rect 2593 26877 2605 26911
rect 2639 26908 2651 26911
rect 2774 26908 2780 26920
rect 2639 26880 2780 26908
rect 2639 26877 2651 26880
rect 2593 26871 2651 26877
rect 2774 26868 2780 26880
rect 2832 26868 2838 26920
rect 3050 26908 3056 26920
rect 3011 26880 3056 26908
rect 3050 26868 3056 26880
rect 3108 26868 3114 26920
rect 4448 26908 4476 27016
rect 6362 27004 6368 27056
rect 6420 27044 6426 27056
rect 9646 27044 9674 27084
rect 11054 27072 11060 27084
rect 11112 27072 11118 27124
rect 11606 27072 11612 27124
rect 11664 27112 11670 27124
rect 12345 27115 12403 27121
rect 12345 27112 12357 27115
rect 11664 27084 12357 27112
rect 11664 27072 11670 27084
rect 12345 27081 12357 27084
rect 12391 27081 12403 27115
rect 12345 27075 12403 27081
rect 12989 27115 13047 27121
rect 12989 27081 13001 27115
rect 13035 27112 13047 27115
rect 13538 27112 13544 27124
rect 13035 27084 13544 27112
rect 13035 27081 13047 27084
rect 12989 27075 13047 27081
rect 13538 27072 13544 27084
rect 13596 27072 13602 27124
rect 13633 27115 13691 27121
rect 13633 27081 13645 27115
rect 13679 27112 13691 27115
rect 13722 27112 13728 27124
rect 13679 27084 13728 27112
rect 13679 27081 13691 27084
rect 13633 27075 13691 27081
rect 13722 27072 13728 27084
rect 13780 27072 13786 27124
rect 17494 27112 17500 27124
rect 17455 27084 17500 27112
rect 17494 27072 17500 27084
rect 17552 27072 17558 27124
rect 18785 27115 18843 27121
rect 18785 27081 18797 27115
rect 18831 27112 18843 27115
rect 20530 27112 20536 27124
rect 18831 27084 20536 27112
rect 18831 27081 18843 27084
rect 18785 27075 18843 27081
rect 20530 27072 20536 27084
rect 20588 27072 20594 27124
rect 23934 27072 23940 27124
rect 23992 27112 23998 27124
rect 25774 27112 25780 27124
rect 23992 27084 25780 27112
rect 23992 27072 23998 27084
rect 25774 27072 25780 27084
rect 25832 27072 25838 27124
rect 27525 27115 27583 27121
rect 27525 27081 27537 27115
rect 27571 27112 27583 27115
rect 27706 27112 27712 27124
rect 27571 27084 27712 27112
rect 27571 27081 27583 27084
rect 27525 27075 27583 27081
rect 27706 27072 27712 27084
rect 27764 27072 27770 27124
rect 6420 27016 9674 27044
rect 6420 27004 6426 27016
rect 9950 27004 9956 27056
rect 10008 27044 10014 27056
rect 10594 27044 10600 27056
rect 10008 27016 10600 27044
rect 10008 27004 10014 27016
rect 10594 27004 10600 27016
rect 10652 27004 10658 27056
rect 12158 27004 12164 27056
rect 12216 27044 12222 27056
rect 14829 27047 14887 27053
rect 14829 27044 14841 27047
rect 12216 27016 12664 27044
rect 12216 27004 12222 27016
rect 6270 26976 6276 26988
rect 5750 26948 6276 26976
rect 6270 26936 6276 26948
rect 6328 26976 6334 26988
rect 11606 26976 11612 26988
rect 6328 26948 11612 26976
rect 6328 26936 6334 26948
rect 11606 26936 11612 26948
rect 11664 26936 11670 26988
rect 11882 26936 11888 26988
rect 11940 26976 11946 26988
rect 12526 26976 12532 26988
rect 11940 26948 12020 26976
rect 11940 26936 11946 26948
rect 4448 26880 6132 26908
rect 1780 26812 4844 26840
rect 1780 26781 1808 26812
rect 1765 26775 1823 26781
rect 1765 26741 1777 26775
rect 1811 26741 1823 26775
rect 1765 26735 1823 26741
rect 3970 26732 3976 26784
rect 4028 26772 4034 26784
rect 4709 26775 4767 26781
rect 4709 26772 4721 26775
rect 4028 26744 4721 26772
rect 4028 26732 4034 26744
rect 4709 26741 4721 26744
rect 4755 26741 4767 26775
rect 4816 26772 4844 26812
rect 4890 26800 4896 26852
rect 4948 26840 4954 26852
rect 4985 26843 5043 26849
rect 4985 26840 4997 26843
rect 4948 26812 4997 26840
rect 4948 26800 4954 26812
rect 4985 26809 4997 26812
rect 5031 26809 5043 26843
rect 4985 26803 5043 26809
rect 5074 26800 5080 26852
rect 5132 26840 5138 26852
rect 5445 26843 5503 26849
rect 5132 26812 5177 26840
rect 5132 26800 5138 26812
rect 5445 26809 5457 26843
rect 5491 26840 5503 26843
rect 6104 26840 6132 26880
rect 10778 26868 10784 26920
rect 10836 26908 10842 26920
rect 11992 26917 12020 26948
rect 12084 26948 12532 26976
rect 12084 26917 12112 26948
rect 12526 26936 12532 26948
rect 12584 26936 12590 26988
rect 10873 26911 10931 26917
rect 10873 26908 10885 26911
rect 10836 26880 10885 26908
rect 10836 26868 10842 26880
rect 10873 26877 10885 26880
rect 10919 26877 10931 26911
rect 10873 26871 10931 26877
rect 11977 26911 12035 26917
rect 11977 26877 11989 26911
rect 12023 26877 12035 26911
rect 11977 26871 12035 26877
rect 12069 26911 12127 26917
rect 12069 26877 12081 26911
rect 12115 26877 12127 26911
rect 12069 26871 12127 26877
rect 12161 26911 12219 26917
rect 12161 26877 12173 26911
rect 12207 26877 12219 26911
rect 12161 26871 12219 26877
rect 5491 26812 6040 26840
rect 6104 26812 11836 26840
rect 5491 26809 5503 26812
rect 5445 26803 5503 26809
rect 5813 26775 5871 26781
rect 5813 26772 5825 26775
rect 4816 26744 5825 26772
rect 4709 26735 4767 26741
rect 5813 26741 5825 26744
rect 5859 26741 5871 26775
rect 6012 26772 6040 26812
rect 6638 26772 6644 26784
rect 6012 26744 6644 26772
rect 5813 26735 5871 26741
rect 6638 26732 6644 26744
rect 6696 26732 6702 26784
rect 10870 26732 10876 26784
rect 10928 26772 10934 26784
rect 10965 26775 11023 26781
rect 10965 26772 10977 26775
rect 10928 26744 10977 26772
rect 10928 26732 10934 26744
rect 10965 26741 10977 26744
rect 11011 26741 11023 26775
rect 11808 26772 11836 26812
rect 11882 26800 11888 26852
rect 11940 26840 11946 26852
rect 12176 26840 12204 26871
rect 11940 26812 12204 26840
rect 11940 26800 11946 26812
rect 12526 26800 12532 26852
rect 12584 26840 12590 26852
rect 12636 26840 12664 27016
rect 13096 27016 14841 27044
rect 13096 26985 13124 27016
rect 14829 27013 14841 27016
rect 14875 27013 14887 27047
rect 14829 27007 14887 27013
rect 18509 27047 18567 27053
rect 18509 27013 18521 27047
rect 18555 27044 18567 27047
rect 18966 27044 18972 27056
rect 18555 27016 18972 27044
rect 18555 27013 18567 27016
rect 18509 27007 18567 27013
rect 18966 27004 18972 27016
rect 19024 27004 19030 27056
rect 23566 27044 23572 27056
rect 23527 27016 23572 27044
rect 23566 27004 23572 27016
rect 23624 27004 23630 27056
rect 26326 27044 26332 27056
rect 24780 27016 26332 27044
rect 13081 26979 13139 26985
rect 13081 26945 13093 26979
rect 13127 26945 13139 26979
rect 13814 26976 13820 26988
rect 13775 26948 13820 26976
rect 13081 26939 13139 26945
rect 13814 26936 13820 26948
rect 13872 26936 13878 26988
rect 17218 26936 17224 26988
rect 17276 26976 17282 26988
rect 17494 26976 17500 26988
rect 17276 26948 17500 26976
rect 17276 26936 17282 26948
rect 17494 26936 17500 26948
rect 17552 26936 17558 26988
rect 22462 26936 22468 26988
rect 22520 26936 22526 26988
rect 12802 26908 12808 26920
rect 12763 26880 12808 26908
rect 12802 26868 12808 26880
rect 12860 26868 12866 26920
rect 12897 26911 12955 26917
rect 12897 26877 12909 26911
rect 12943 26877 12955 26911
rect 13538 26908 13544 26920
rect 13499 26880 13544 26908
rect 12897 26871 12955 26877
rect 12584 26812 12664 26840
rect 12584 26800 12590 26812
rect 12710 26772 12716 26784
rect 11808 26744 12716 26772
rect 10965 26735 11023 26741
rect 12710 26732 12716 26744
rect 12768 26732 12774 26784
rect 12912 26772 12940 26871
rect 13538 26868 13544 26880
rect 13596 26868 13602 26920
rect 15013 26911 15071 26917
rect 15013 26877 15025 26911
rect 15059 26908 15071 26911
rect 15838 26908 15844 26920
rect 15059 26880 15844 26908
rect 15059 26877 15071 26880
rect 15013 26871 15071 26877
rect 15838 26868 15844 26880
rect 15896 26868 15902 26920
rect 16114 26868 16120 26920
rect 16172 26908 16178 26920
rect 16485 26911 16543 26917
rect 16485 26908 16497 26911
rect 16172 26880 16497 26908
rect 16172 26868 16178 26880
rect 16485 26877 16497 26880
rect 16531 26877 16543 26911
rect 16485 26871 16543 26877
rect 16577 26911 16635 26917
rect 16577 26877 16589 26911
rect 16623 26908 16635 26911
rect 17678 26908 17684 26920
rect 16623 26880 17684 26908
rect 16623 26877 16635 26880
rect 16577 26871 16635 26877
rect 17678 26868 17684 26880
rect 17736 26868 17742 26920
rect 17862 26868 17868 26920
rect 17920 26908 17926 26920
rect 18782 26908 18788 26920
rect 17920 26880 18276 26908
rect 18743 26880 18788 26908
rect 17920 26868 17926 26880
rect 13078 26800 13084 26852
rect 13136 26840 13142 26852
rect 13817 26843 13875 26849
rect 13817 26840 13829 26843
rect 13136 26812 13829 26840
rect 13136 26800 13142 26812
rect 13817 26809 13829 26812
rect 13863 26809 13875 26843
rect 14734 26840 14740 26852
rect 14695 26812 14740 26840
rect 13817 26803 13875 26809
rect 14734 26800 14740 26812
rect 14792 26800 14798 26852
rect 14826 26800 14832 26852
rect 14884 26840 14890 26852
rect 14921 26843 14979 26849
rect 14921 26840 14933 26843
rect 14884 26812 14933 26840
rect 14884 26800 14890 26812
rect 14921 26809 14933 26812
rect 14967 26809 14979 26843
rect 14921 26803 14979 26809
rect 15930 26800 15936 26852
rect 15988 26840 15994 26852
rect 16209 26843 16267 26849
rect 16209 26840 16221 26843
rect 15988 26812 16221 26840
rect 15988 26800 15994 26812
rect 16209 26809 16221 26812
rect 16255 26809 16267 26843
rect 16209 26803 16267 26809
rect 16945 26843 17003 26849
rect 16945 26809 16957 26843
rect 16991 26840 17003 26843
rect 18248 26840 18276 26880
rect 18782 26868 18788 26880
rect 18840 26868 18846 26920
rect 18874 26868 18880 26920
rect 18932 26908 18938 26920
rect 18969 26911 19027 26917
rect 18969 26908 18981 26911
rect 18932 26880 18981 26908
rect 18932 26868 18938 26880
rect 18969 26877 18981 26880
rect 19015 26877 19027 26911
rect 18969 26871 19027 26877
rect 19518 26868 19524 26920
rect 19576 26908 19582 26920
rect 24780 26908 24808 27016
rect 26326 27004 26332 27016
rect 26384 27004 26390 27056
rect 27249 27047 27307 27053
rect 27249 27013 27261 27047
rect 27295 27044 27307 27047
rect 28350 27044 28356 27056
rect 27295 27016 28356 27044
rect 27295 27013 27307 27016
rect 27249 27007 27307 27013
rect 28350 27004 28356 27016
rect 28408 27004 28414 27056
rect 24854 26936 24860 26988
rect 24912 26976 24918 26988
rect 25406 26976 25412 26988
rect 24912 26948 25412 26976
rect 24912 26936 24918 26948
rect 25406 26936 25412 26948
rect 25464 26936 25470 26988
rect 28166 26976 28172 26988
rect 27540 26948 28172 26976
rect 25314 26908 25320 26920
rect 19576 26880 23428 26908
rect 19576 26868 19582 26880
rect 22557 26843 22615 26849
rect 22557 26840 22569 26843
rect 16991 26812 18184 26840
rect 18248 26812 22569 26840
rect 16991 26809 17003 26812
rect 16945 26803 17003 26809
rect 13722 26772 13728 26784
rect 12912 26744 13728 26772
rect 13722 26732 13728 26744
rect 13780 26732 13786 26784
rect 14274 26732 14280 26784
rect 14332 26772 14338 26784
rect 14844 26772 14872 26800
rect 14332 26744 14872 26772
rect 14332 26732 14338 26744
rect 17034 26732 17040 26784
rect 17092 26772 17098 26784
rect 17313 26775 17371 26781
rect 17313 26772 17325 26775
rect 17092 26744 17325 26772
rect 17092 26732 17098 26744
rect 17313 26741 17325 26744
rect 17359 26741 17371 26775
rect 18156 26772 18184 26812
rect 22557 26809 22569 26812
rect 22603 26809 22615 26843
rect 22557 26803 22615 26809
rect 20162 26772 20168 26784
rect 18156 26744 20168 26772
rect 17313 26735 17371 26741
rect 20162 26732 20168 26744
rect 20220 26732 20226 26784
rect 21910 26732 21916 26784
rect 21968 26772 21974 26784
rect 22281 26775 22339 26781
rect 22281 26772 22293 26775
rect 21968 26744 22293 26772
rect 21968 26732 21974 26744
rect 22281 26741 22293 26744
rect 22327 26741 22339 26775
rect 22572 26772 22600 26803
rect 22646 26800 22652 26852
rect 22704 26840 22710 26852
rect 23014 26840 23020 26852
rect 22704 26812 22749 26840
rect 22975 26812 23020 26840
rect 22704 26800 22710 26812
rect 23014 26800 23020 26812
rect 23072 26800 23078 26852
rect 23400 26849 23428 26880
rect 23768 26880 24808 26908
rect 25275 26880 25320 26908
rect 23385 26843 23443 26849
rect 23385 26809 23397 26843
rect 23431 26809 23443 26843
rect 23385 26803 23443 26809
rect 23768 26772 23796 26880
rect 25314 26868 25320 26880
rect 25372 26868 25378 26920
rect 27540 26917 27568 26948
rect 28166 26936 28172 26948
rect 28224 26936 28230 26988
rect 27525 26911 27583 26917
rect 27525 26877 27537 26911
rect 27571 26877 27583 26911
rect 27525 26871 27583 26877
rect 27709 26911 27767 26917
rect 27709 26877 27721 26911
rect 27755 26908 27767 26911
rect 27798 26908 27804 26920
rect 27755 26880 27804 26908
rect 27755 26877 27767 26880
rect 27709 26871 27767 26877
rect 27798 26868 27804 26880
rect 27856 26868 27862 26920
rect 24026 26800 24032 26852
rect 24084 26840 24090 26852
rect 25501 26843 25559 26849
rect 25501 26840 25513 26843
rect 24084 26812 25513 26840
rect 24084 26800 24090 26812
rect 25501 26809 25513 26812
rect 25547 26840 25559 26843
rect 26418 26840 26424 26852
rect 25547 26812 26424 26840
rect 25547 26809 25559 26812
rect 25501 26803 25559 26809
rect 26418 26800 26424 26812
rect 26476 26800 26482 26852
rect 26602 26840 26608 26852
rect 26563 26812 26608 26840
rect 26602 26800 26608 26812
rect 26660 26800 26666 26852
rect 22572 26744 23796 26772
rect 22281 26735 22339 26741
rect 24946 26732 24952 26784
rect 25004 26772 25010 26784
rect 25314 26772 25320 26784
rect 25004 26744 25320 26772
rect 25004 26732 25010 26744
rect 25314 26732 25320 26744
rect 25372 26732 25378 26784
rect 26694 26772 26700 26784
rect 26655 26744 26700 26772
rect 26694 26732 26700 26744
rect 26752 26732 26758 26784
rect 1104 26682 28888 26704
rect 1104 26630 10246 26682
rect 10298 26630 10310 26682
rect 10362 26630 10374 26682
rect 10426 26630 10438 26682
rect 10490 26630 19510 26682
rect 19562 26630 19574 26682
rect 19626 26630 19638 26682
rect 19690 26630 19702 26682
rect 19754 26630 28888 26682
rect 1104 26608 28888 26630
rect 1762 26568 1768 26580
rect 1723 26540 1768 26568
rect 1762 26528 1768 26540
rect 1820 26528 1826 26580
rect 2406 26528 2412 26580
rect 2464 26568 2470 26580
rect 2501 26571 2559 26577
rect 2501 26568 2513 26571
rect 2464 26540 2513 26568
rect 2464 26528 2470 26540
rect 2501 26537 2513 26540
rect 2547 26568 2559 26571
rect 2958 26568 2964 26580
rect 2547 26540 2964 26568
rect 2547 26537 2559 26540
rect 2501 26531 2559 26537
rect 2958 26528 2964 26540
rect 3016 26528 3022 26580
rect 3237 26571 3295 26577
rect 3237 26537 3249 26571
rect 3283 26537 3295 26571
rect 3237 26531 3295 26537
rect 4525 26571 4583 26577
rect 4525 26537 4537 26571
rect 4571 26568 4583 26571
rect 4614 26568 4620 26580
rect 4571 26540 4620 26568
rect 4571 26537 4583 26540
rect 4525 26531 4583 26537
rect 3252 26500 3280 26531
rect 4614 26528 4620 26540
rect 4672 26528 4678 26580
rect 5902 26528 5908 26580
rect 5960 26568 5966 26580
rect 6822 26568 6828 26580
rect 5960 26540 6828 26568
rect 5960 26528 5966 26540
rect 6822 26528 6828 26540
rect 6880 26528 6886 26580
rect 9858 26568 9864 26580
rect 9819 26540 9864 26568
rect 9858 26528 9864 26540
rect 9916 26568 9922 26580
rect 11698 26568 11704 26580
rect 9916 26540 11704 26568
rect 9916 26528 9922 26540
rect 11698 26528 11704 26540
rect 11756 26528 11762 26580
rect 12342 26528 12348 26580
rect 12400 26568 12406 26580
rect 12710 26568 12716 26580
rect 12400 26540 12716 26568
rect 12400 26528 12406 26540
rect 12710 26528 12716 26540
rect 12768 26528 12774 26580
rect 12989 26571 13047 26577
rect 12989 26537 13001 26571
rect 13035 26568 13047 26571
rect 13262 26568 13268 26580
rect 13035 26540 13268 26568
rect 13035 26537 13047 26540
rect 12989 26531 13047 26537
rect 13262 26528 13268 26540
rect 13320 26528 13326 26580
rect 13814 26528 13820 26580
rect 13872 26568 13878 26580
rect 15197 26571 15255 26577
rect 15197 26568 15209 26571
rect 13872 26540 15209 26568
rect 13872 26528 13878 26540
rect 15197 26537 15209 26540
rect 15243 26537 15255 26571
rect 15197 26531 15255 26537
rect 15470 26528 15476 26580
rect 15528 26568 15534 26580
rect 15933 26571 15991 26577
rect 15933 26568 15945 26571
rect 15528 26540 15945 26568
rect 15528 26528 15534 26540
rect 15933 26537 15945 26540
rect 15979 26537 15991 26571
rect 15933 26531 15991 26537
rect 18509 26571 18567 26577
rect 18509 26537 18521 26571
rect 18555 26568 18567 26571
rect 18782 26568 18788 26580
rect 18555 26540 18788 26568
rect 18555 26537 18567 26540
rect 18509 26531 18567 26537
rect 18782 26528 18788 26540
rect 18840 26528 18846 26580
rect 20254 26528 20260 26580
rect 20312 26568 20318 26580
rect 26602 26568 26608 26580
rect 20312 26540 26608 26568
rect 20312 26528 20318 26540
rect 26602 26528 26608 26540
rect 26660 26528 26666 26580
rect 10962 26500 10968 26512
rect 2746 26472 9444 26500
rect 10923 26472 10968 26500
rect 1946 26432 1952 26444
rect 1907 26404 1952 26432
rect 1946 26392 1952 26404
rect 2004 26392 2010 26444
rect 2409 26435 2467 26441
rect 2409 26401 2421 26435
rect 2455 26432 2467 26435
rect 2498 26432 2504 26444
rect 2455 26404 2504 26432
rect 2455 26401 2467 26404
rect 2409 26395 2467 26401
rect 2498 26392 2504 26404
rect 2556 26392 2562 26444
rect 2222 26256 2228 26308
rect 2280 26296 2286 26308
rect 2746 26296 2774 26472
rect 3050 26432 3056 26444
rect 3011 26404 3056 26432
rect 3050 26392 3056 26404
rect 3108 26392 3114 26444
rect 4154 26392 4160 26444
rect 4212 26432 4218 26444
rect 5353 26435 5411 26441
rect 5353 26432 5365 26435
rect 4212 26404 5365 26432
rect 4212 26392 4218 26404
rect 5353 26401 5365 26404
rect 5399 26401 5411 26435
rect 8018 26432 8024 26444
rect 7979 26404 8024 26432
rect 5353 26395 5411 26401
rect 8018 26392 8024 26404
rect 8076 26392 8082 26444
rect 9030 26432 9036 26444
rect 8991 26404 9036 26432
rect 9030 26392 9036 26404
rect 9088 26392 9094 26444
rect 9217 26435 9275 26441
rect 9217 26401 9229 26435
rect 9263 26401 9275 26435
rect 9217 26395 9275 26401
rect 9309 26435 9367 26441
rect 9309 26401 9321 26435
rect 9355 26401 9367 26435
rect 9309 26395 9367 26401
rect 4614 26364 4620 26376
rect 4575 26336 4620 26364
rect 4614 26324 4620 26336
rect 4672 26324 4678 26376
rect 4801 26367 4859 26373
rect 4801 26333 4813 26367
rect 4847 26364 4859 26367
rect 4890 26364 4896 26376
rect 4847 26336 4896 26364
rect 4847 26333 4859 26336
rect 4801 26327 4859 26333
rect 4890 26324 4896 26336
rect 4948 26324 4954 26376
rect 8110 26364 8116 26376
rect 8071 26336 8116 26364
rect 8110 26324 8116 26336
rect 8168 26324 8174 26376
rect 8389 26367 8447 26373
rect 8389 26333 8401 26367
rect 8435 26364 8447 26367
rect 9232 26364 9260 26395
rect 8435 26336 9260 26364
rect 8435 26333 8447 26336
rect 8389 26327 8447 26333
rect 2280 26268 2774 26296
rect 4157 26299 4215 26305
rect 2280 26256 2286 26268
rect 4157 26265 4169 26299
rect 4203 26296 4215 26299
rect 5166 26296 5172 26308
rect 4203 26268 5172 26296
rect 4203 26265 4215 26268
rect 4157 26259 4215 26265
rect 5166 26256 5172 26268
rect 5224 26256 5230 26308
rect 5537 26299 5595 26305
rect 5537 26265 5549 26299
rect 5583 26296 5595 26299
rect 6086 26296 6092 26308
rect 5583 26268 6092 26296
rect 5583 26265 5595 26268
rect 5537 26259 5595 26265
rect 6086 26256 6092 26268
rect 6144 26256 6150 26308
rect 9324 26296 9352 26395
rect 9416 26364 9444 26472
rect 10962 26460 10968 26472
rect 11020 26460 11026 26512
rect 11057 26503 11115 26509
rect 11057 26469 11069 26503
rect 11103 26500 11115 26503
rect 12250 26500 12256 26512
rect 11103 26472 12256 26500
rect 11103 26469 11115 26472
rect 11057 26463 11115 26469
rect 9769 26435 9827 26441
rect 9769 26401 9781 26435
rect 9815 26432 9827 26435
rect 10134 26432 10140 26444
rect 9815 26404 10140 26432
rect 9815 26401 9827 26404
rect 9769 26395 9827 26401
rect 10134 26392 10140 26404
rect 10192 26392 10198 26444
rect 10778 26432 10784 26444
rect 10739 26404 10784 26432
rect 10778 26392 10784 26404
rect 10836 26392 10842 26444
rect 11164 26376 11192 26472
rect 12250 26460 12256 26472
rect 12308 26460 12314 26512
rect 13998 26460 14004 26512
rect 14056 26500 14062 26512
rect 14826 26500 14832 26512
rect 14056 26472 14832 26500
rect 14056 26460 14062 26472
rect 14826 26460 14832 26472
rect 14884 26500 14890 26512
rect 15289 26503 15347 26509
rect 15289 26500 15301 26503
rect 14884 26472 15301 26500
rect 14884 26460 14890 26472
rect 15289 26469 15301 26472
rect 15335 26500 15347 26503
rect 16025 26503 16083 26509
rect 16025 26500 16037 26503
rect 15335 26472 16037 26500
rect 15335 26469 15347 26472
rect 15289 26463 15347 26469
rect 16025 26469 16037 26472
rect 16071 26469 16083 26503
rect 16025 26463 16083 26469
rect 17402 26460 17408 26512
rect 17460 26500 17466 26512
rect 17460 26472 22968 26500
rect 17460 26460 17466 26472
rect 12526 26392 12532 26444
rect 12584 26432 12590 26444
rect 12805 26435 12863 26441
rect 12805 26432 12817 26435
rect 12584 26404 12817 26432
rect 12584 26392 12590 26404
rect 12805 26401 12817 26404
rect 12851 26401 12863 26435
rect 12805 26395 12863 26401
rect 13262 26392 13268 26444
rect 13320 26432 13326 26444
rect 13538 26432 13544 26444
rect 13320 26404 13544 26432
rect 13320 26392 13326 26404
rect 13538 26392 13544 26404
rect 13596 26392 13602 26444
rect 14461 26435 14519 26441
rect 14461 26401 14473 26435
rect 14507 26432 14519 26435
rect 14550 26432 14556 26444
rect 14507 26404 14556 26432
rect 14507 26401 14519 26404
rect 14461 26395 14519 26401
rect 14550 26392 14556 26404
rect 14608 26392 14614 26444
rect 14642 26392 14648 26444
rect 14700 26432 14706 26444
rect 15105 26435 15163 26441
rect 15105 26432 15117 26435
rect 14700 26404 15117 26432
rect 14700 26392 14706 26404
rect 15105 26401 15117 26404
rect 15151 26401 15163 26435
rect 15105 26395 15163 26401
rect 15381 26435 15439 26441
rect 15381 26401 15393 26435
rect 15427 26401 15439 26435
rect 15381 26395 15439 26401
rect 10410 26364 10416 26376
rect 9416 26336 10416 26364
rect 10410 26324 10416 26336
rect 10468 26324 10474 26376
rect 11146 26324 11152 26376
rect 11204 26324 11210 26376
rect 15396 26364 15424 26395
rect 15470 26392 15476 26444
rect 15528 26432 15534 26444
rect 15841 26435 15899 26441
rect 15841 26432 15853 26435
rect 15528 26404 15853 26432
rect 15528 26392 15534 26404
rect 15841 26401 15853 26404
rect 15887 26401 15899 26435
rect 15841 26395 15899 26401
rect 16117 26435 16175 26441
rect 16117 26401 16129 26435
rect 16163 26401 16175 26435
rect 16117 26395 16175 26401
rect 15930 26364 15936 26376
rect 15396 26336 15936 26364
rect 15930 26324 15936 26336
rect 15988 26364 15994 26376
rect 16132 26364 16160 26395
rect 18322 26392 18328 26444
rect 18380 26432 18386 26444
rect 18417 26435 18475 26441
rect 18417 26432 18429 26435
rect 18380 26404 18429 26432
rect 18380 26392 18386 26404
rect 18417 26401 18429 26404
rect 18463 26401 18475 26435
rect 18598 26432 18604 26444
rect 18559 26404 18604 26432
rect 18417 26395 18475 26401
rect 15988 26336 16160 26364
rect 18432 26364 18460 26395
rect 18598 26392 18604 26404
rect 18656 26392 18662 26444
rect 22940 26432 22968 26472
rect 23014 26460 23020 26512
rect 23072 26500 23078 26512
rect 25961 26503 26019 26509
rect 25961 26500 25973 26503
rect 23072 26472 25973 26500
rect 23072 26460 23078 26472
rect 25961 26469 25973 26472
rect 26007 26469 26019 26503
rect 25961 26463 26019 26469
rect 26142 26460 26148 26512
rect 26200 26500 26206 26512
rect 26881 26503 26939 26509
rect 26881 26500 26893 26503
rect 26200 26472 26893 26500
rect 26200 26460 26206 26472
rect 26881 26469 26893 26472
rect 26927 26469 26939 26503
rect 27982 26500 27988 26512
rect 27943 26472 27988 26500
rect 26881 26463 26939 26469
rect 27982 26460 27988 26472
rect 28040 26460 28046 26512
rect 25225 26435 25283 26441
rect 22940 26404 24808 26432
rect 18782 26364 18788 26376
rect 18432 26336 18788 26364
rect 15988 26324 15994 26336
rect 18782 26324 18788 26336
rect 18840 26324 18846 26376
rect 9674 26296 9680 26308
rect 9324 26268 9680 26296
rect 9674 26256 9680 26268
rect 9732 26256 9738 26308
rect 10505 26299 10563 26305
rect 10505 26265 10517 26299
rect 10551 26296 10563 26299
rect 22278 26296 22284 26308
rect 10551 26268 22284 26296
rect 10551 26265 10563 26268
rect 10505 26259 10563 26265
rect 22278 26256 22284 26268
rect 22336 26256 22342 26308
rect 22646 26256 22652 26308
rect 22704 26296 22710 26308
rect 23290 26296 23296 26308
rect 22704 26268 23296 26296
rect 22704 26256 22710 26268
rect 23290 26256 23296 26268
rect 23348 26256 23354 26308
rect 24780 26296 24808 26404
rect 25225 26401 25237 26435
rect 25271 26401 25283 26435
rect 25225 26395 25283 26401
rect 25240 26364 25268 26395
rect 26050 26392 26056 26444
rect 26108 26432 26114 26444
rect 26697 26435 26755 26441
rect 26697 26432 26709 26435
rect 26108 26404 26709 26432
rect 26108 26392 26114 26404
rect 26697 26401 26709 26404
rect 26743 26401 26755 26435
rect 26697 26395 26755 26401
rect 26234 26364 26240 26376
rect 25240 26336 26240 26364
rect 26234 26324 26240 26336
rect 26292 26324 26298 26376
rect 25406 26296 25412 26308
rect 24780 26268 25268 26296
rect 25367 26268 25412 26296
rect 9033 26231 9091 26237
rect 9033 26197 9045 26231
rect 9079 26228 9091 26231
rect 9582 26228 9588 26240
rect 9079 26200 9588 26228
rect 9079 26197 9091 26200
rect 9033 26191 9091 26197
rect 9582 26188 9588 26200
rect 9640 26188 9646 26240
rect 13354 26188 13360 26240
rect 13412 26228 13418 26240
rect 13538 26228 13544 26240
rect 13412 26200 13544 26228
rect 13412 26188 13418 26200
rect 13538 26188 13544 26200
rect 13596 26188 13602 26240
rect 13722 26188 13728 26240
rect 13780 26228 13786 26240
rect 14090 26228 14096 26240
rect 13780 26200 14096 26228
rect 13780 26188 13786 26200
rect 14090 26188 14096 26200
rect 14148 26188 14154 26240
rect 14274 26188 14280 26240
rect 14332 26228 14338 26240
rect 14553 26231 14611 26237
rect 14553 26228 14565 26231
rect 14332 26200 14565 26228
rect 14332 26188 14338 26200
rect 14553 26197 14565 26200
rect 14599 26197 14611 26231
rect 25240 26228 25268 26268
rect 25406 26256 25412 26268
rect 25464 26256 25470 26308
rect 25682 26296 25688 26308
rect 25516 26268 25688 26296
rect 25516 26228 25544 26268
rect 25682 26256 25688 26268
rect 25740 26256 25746 26308
rect 26142 26296 26148 26308
rect 26103 26268 26148 26296
rect 26142 26256 26148 26268
rect 26200 26256 26206 26308
rect 28166 26296 28172 26308
rect 28127 26268 28172 26296
rect 28166 26256 28172 26268
rect 28224 26256 28230 26308
rect 25240 26200 25544 26228
rect 14553 26191 14611 26197
rect 1104 26138 28888 26160
rect 1104 26086 5614 26138
rect 5666 26086 5678 26138
rect 5730 26086 5742 26138
rect 5794 26086 5806 26138
rect 5858 26086 14878 26138
rect 14930 26086 14942 26138
rect 14994 26086 15006 26138
rect 15058 26086 15070 26138
rect 15122 26086 24142 26138
rect 24194 26086 24206 26138
rect 24258 26086 24270 26138
rect 24322 26086 24334 26138
rect 24386 26086 28888 26138
rect 1104 26064 28888 26086
rect 6454 26024 6460 26036
rect 4448 25996 6460 26024
rect 1762 25848 1768 25900
rect 1820 25888 1826 25900
rect 2038 25888 2044 25900
rect 1820 25860 2044 25888
rect 1820 25848 1826 25860
rect 2038 25848 2044 25860
rect 2096 25848 2102 25900
rect 4448 25897 4476 25996
rect 6454 25984 6460 25996
rect 6512 25984 6518 26036
rect 6733 26027 6791 26033
rect 6733 25993 6745 26027
rect 6779 26024 6791 26027
rect 7190 26024 7196 26036
rect 6779 25996 7196 26024
rect 6779 25993 6791 25996
rect 6733 25987 6791 25993
rect 7190 25984 7196 25996
rect 7248 25984 7254 26036
rect 7466 26024 7472 26036
rect 7427 25996 7472 26024
rect 7466 25984 7472 25996
rect 7524 25984 7530 26036
rect 10962 25984 10968 26036
rect 11020 26024 11026 26036
rect 11425 26027 11483 26033
rect 11425 26024 11437 26027
rect 11020 25996 11437 26024
rect 11020 25984 11026 25996
rect 11425 25993 11437 25996
rect 11471 25993 11483 26027
rect 11425 25987 11483 25993
rect 12342 25984 12348 26036
rect 12400 26024 12406 26036
rect 12618 26024 12624 26036
rect 12400 25996 12624 26024
rect 12400 25984 12406 25996
rect 12618 25984 12624 25996
rect 12676 25984 12682 26036
rect 12710 25984 12716 26036
rect 12768 26024 12774 26036
rect 13265 26027 13323 26033
rect 13265 26024 13277 26027
rect 12768 25996 13277 26024
rect 12768 25984 12774 25996
rect 13265 25993 13277 25996
rect 13311 26024 13323 26027
rect 13354 26024 13360 26036
rect 13311 25996 13360 26024
rect 13311 25993 13323 25996
rect 13265 25987 13323 25993
rect 13354 25984 13360 25996
rect 13412 25984 13418 26036
rect 16114 25984 16120 26036
rect 16172 26024 16178 26036
rect 17402 26024 17408 26036
rect 16172 25996 17408 26024
rect 16172 25984 16178 25996
rect 17402 25984 17408 25996
rect 17460 25984 17466 26036
rect 20162 25984 20168 26036
rect 20220 26024 20226 26036
rect 23842 26024 23848 26036
rect 20220 25996 23848 26024
rect 20220 25984 20226 25996
rect 23842 25984 23848 25996
rect 23900 26024 23906 26036
rect 25682 26024 25688 26036
rect 23900 25996 25688 26024
rect 23900 25984 23906 25996
rect 25682 25984 25688 25996
rect 25740 25984 25746 26036
rect 26329 26027 26387 26033
rect 26329 25993 26341 26027
rect 26375 26024 26387 26027
rect 27798 26024 27804 26036
rect 26375 25996 27804 26024
rect 26375 25993 26387 25996
rect 26329 25987 26387 25993
rect 27798 25984 27804 25996
rect 27856 25984 27862 26036
rect 11330 25916 11336 25968
rect 11388 25956 11394 25968
rect 11388 25928 12020 25956
rect 11388 25916 11394 25928
rect 6184 25900 6236 25906
rect 4433 25891 4491 25897
rect 4433 25857 4445 25891
rect 4479 25857 4491 25891
rect 4433 25851 4491 25857
rect 10870 25848 10876 25900
rect 10928 25888 10934 25900
rect 11992 25897 12020 25928
rect 12250 25916 12256 25968
rect 12308 25956 12314 25968
rect 14918 25956 14924 25968
rect 12308 25928 14924 25956
rect 12308 25916 12314 25928
rect 14918 25916 14924 25928
rect 14976 25956 14982 25968
rect 16206 25956 16212 25968
rect 14976 25928 16212 25956
rect 14976 25916 14982 25928
rect 16206 25916 16212 25928
rect 16264 25916 16270 25968
rect 17494 25916 17500 25968
rect 17552 25956 17558 25968
rect 17681 25959 17739 25965
rect 17681 25956 17693 25959
rect 17552 25928 17693 25956
rect 17552 25916 17558 25928
rect 17681 25925 17693 25928
rect 17727 25925 17739 25959
rect 19334 25956 19340 25968
rect 17681 25919 17739 25925
rect 17788 25928 19340 25956
rect 11885 25891 11943 25897
rect 11885 25888 11897 25891
rect 10928 25860 11897 25888
rect 10928 25848 10934 25860
rect 11885 25857 11897 25860
rect 11931 25857 11943 25891
rect 11885 25851 11943 25857
rect 11977 25891 12035 25897
rect 11977 25857 11989 25891
rect 12023 25888 12035 25891
rect 15470 25888 15476 25900
rect 12023 25860 15476 25888
rect 12023 25857 12035 25860
rect 11977 25851 12035 25857
rect 15470 25848 15476 25860
rect 15528 25848 15534 25900
rect 16301 25891 16359 25897
rect 16301 25857 16313 25891
rect 16347 25888 16359 25891
rect 17788 25888 17816 25928
rect 19334 25916 19340 25928
rect 19392 25916 19398 25968
rect 24670 25956 24676 25968
rect 23860 25928 24676 25956
rect 23860 25900 23888 25928
rect 24670 25916 24676 25928
rect 24728 25916 24734 25968
rect 16347 25860 17816 25888
rect 18693 25891 18751 25897
rect 16347 25857 16359 25860
rect 16301 25851 16359 25857
rect 18693 25857 18705 25891
rect 18739 25888 18751 25891
rect 18782 25888 18788 25900
rect 18739 25860 18788 25888
rect 18739 25857 18751 25860
rect 18693 25851 18751 25857
rect 18782 25848 18788 25860
rect 18840 25848 18846 25900
rect 18966 25888 18972 25900
rect 18927 25860 18972 25888
rect 18966 25848 18972 25860
rect 19024 25848 19030 25900
rect 23842 25848 23848 25900
rect 23900 25848 23906 25900
rect 24305 25891 24363 25897
rect 24305 25857 24317 25891
rect 24351 25888 24363 25891
rect 24946 25888 24952 25900
rect 24351 25860 24952 25888
rect 24351 25857 24363 25860
rect 24305 25851 24363 25857
rect 24946 25848 24952 25860
rect 25004 25848 25010 25900
rect 26053 25891 26111 25897
rect 26053 25857 26065 25891
rect 26099 25888 26111 25891
rect 26099 25860 26924 25888
rect 26099 25857 26111 25860
rect 26053 25851 26111 25857
rect 6184 25842 6236 25848
rect 1854 25820 1860 25832
rect 1815 25792 1860 25820
rect 1854 25780 1860 25792
rect 1912 25780 1918 25832
rect 2961 25823 3019 25829
rect 2961 25789 2973 25823
rect 3007 25820 3019 25823
rect 4246 25820 4252 25832
rect 3007 25792 4252 25820
rect 3007 25789 3019 25792
rect 2961 25783 3019 25789
rect 4246 25780 4252 25792
rect 4304 25780 4310 25832
rect 5166 25780 5172 25832
rect 5224 25780 5230 25832
rect 6914 25820 6920 25832
rect 6875 25792 6920 25820
rect 6914 25780 6920 25792
rect 6972 25780 6978 25832
rect 7374 25820 7380 25832
rect 7335 25792 7380 25820
rect 7374 25780 7380 25792
rect 7432 25780 7438 25832
rect 7742 25820 7748 25832
rect 7703 25792 7748 25820
rect 7742 25780 7748 25792
rect 7800 25780 7806 25832
rect 8294 25820 8300 25832
rect 8255 25792 8300 25820
rect 8294 25780 8300 25792
rect 8352 25780 8358 25832
rect 9490 25820 9496 25832
rect 9451 25792 9496 25820
rect 9490 25780 9496 25792
rect 9548 25780 9554 25832
rect 9582 25780 9588 25832
rect 9640 25820 9646 25832
rect 9749 25823 9807 25829
rect 9749 25820 9761 25823
rect 9640 25792 9761 25820
rect 9640 25780 9646 25792
rect 9749 25789 9761 25792
rect 9795 25789 9807 25823
rect 9749 25783 9807 25789
rect 11698 25780 11704 25832
rect 11756 25820 11762 25832
rect 11793 25823 11851 25829
rect 11793 25820 11805 25823
rect 11756 25792 11805 25820
rect 11756 25780 11762 25792
rect 11793 25789 11805 25792
rect 11839 25789 11851 25823
rect 11793 25783 11851 25789
rect 14550 25780 14556 25832
rect 14608 25820 14614 25832
rect 14737 25823 14795 25829
rect 14737 25820 14749 25823
rect 14608 25792 14749 25820
rect 14608 25780 14614 25792
rect 14737 25789 14749 25792
rect 14783 25789 14795 25823
rect 16574 25820 16580 25832
rect 16535 25792 16580 25820
rect 14737 25783 14795 25789
rect 16574 25780 16580 25792
rect 16632 25780 16638 25832
rect 18598 25820 18604 25832
rect 18559 25792 18604 25820
rect 18598 25780 18604 25792
rect 18656 25780 18662 25832
rect 19334 25780 19340 25832
rect 19392 25820 19398 25832
rect 21177 25823 21235 25829
rect 21177 25820 21189 25823
rect 19392 25792 21189 25820
rect 19392 25780 19398 25792
rect 21177 25789 21189 25792
rect 21223 25789 21235 25823
rect 21177 25783 21235 25789
rect 24026 25780 24032 25832
rect 24084 25820 24090 25832
rect 24486 25820 24492 25832
rect 24084 25792 24492 25820
rect 24084 25780 24090 25792
rect 24486 25780 24492 25792
rect 24544 25780 24550 25832
rect 25961 25823 26019 25829
rect 25961 25789 25973 25823
rect 26007 25820 26019 25823
rect 26694 25820 26700 25832
rect 26007 25792 26700 25820
rect 26007 25789 26019 25792
rect 25961 25783 26019 25789
rect 26694 25780 26700 25792
rect 26752 25780 26758 25832
rect 26789 25823 26847 25829
rect 26789 25789 26801 25823
rect 26835 25789 26847 25823
rect 26896 25820 26924 25860
rect 27982 25820 27988 25832
rect 26896 25792 27988 25820
rect 26789 25783 26847 25789
rect 2038 25752 2044 25764
rect 1999 25724 2044 25752
rect 2038 25712 2044 25724
rect 2096 25712 2102 25764
rect 6638 25752 6644 25764
rect 6599 25724 6644 25752
rect 6638 25712 6644 25724
rect 6696 25712 6702 25764
rect 6825 25755 6883 25761
rect 6825 25721 6837 25755
rect 6871 25752 6883 25755
rect 7558 25752 7564 25764
rect 6871 25724 7564 25752
rect 6871 25721 6883 25724
rect 6825 25715 6883 25721
rect 7558 25712 7564 25724
rect 7616 25712 7622 25764
rect 13078 25712 13084 25764
rect 13136 25712 13142 25764
rect 13173 25755 13231 25761
rect 13173 25721 13185 25755
rect 13219 25752 13231 25755
rect 13262 25752 13268 25764
rect 13219 25724 13268 25752
rect 13219 25721 13231 25724
rect 13173 25715 13231 25721
rect 13262 25712 13268 25724
rect 13320 25712 13326 25764
rect 13814 25712 13820 25764
rect 13872 25752 13878 25764
rect 15657 25755 15715 25761
rect 15657 25752 15669 25755
rect 13872 25724 15669 25752
rect 13872 25712 13878 25724
rect 15657 25721 15669 25724
rect 15703 25721 15715 25755
rect 15657 25715 15715 25721
rect 15841 25755 15899 25761
rect 15841 25721 15853 25755
rect 15887 25752 15899 25755
rect 16114 25752 16120 25764
rect 15887 25724 16120 25752
rect 15887 25721 15899 25724
rect 15841 25715 15899 25721
rect 2314 25644 2320 25696
rect 2372 25684 2378 25696
rect 3145 25687 3203 25693
rect 3145 25684 3157 25687
rect 2372 25656 3157 25684
rect 2372 25644 2378 25656
rect 3145 25653 3157 25656
rect 3191 25653 3203 25687
rect 3145 25647 3203 25653
rect 4798 25644 4804 25696
rect 4856 25684 4862 25696
rect 5445 25687 5503 25693
rect 5445 25684 5457 25687
rect 4856 25656 5457 25684
rect 4856 25644 4862 25656
rect 5445 25653 5457 25656
rect 5491 25653 5503 25687
rect 10870 25684 10876 25696
rect 10831 25656 10876 25684
rect 5445 25647 5503 25653
rect 10870 25644 10876 25656
rect 10928 25644 10934 25696
rect 11698 25644 11704 25696
rect 11756 25684 11762 25696
rect 11974 25684 11980 25696
rect 11756 25656 11980 25684
rect 11756 25644 11762 25656
rect 11974 25644 11980 25656
rect 12032 25644 12038 25696
rect 12710 25644 12716 25696
rect 12768 25684 12774 25696
rect 13096 25684 13124 25712
rect 14921 25687 14979 25693
rect 14921 25684 14933 25687
rect 12768 25656 14933 25684
rect 12768 25644 12774 25656
rect 14921 25653 14933 25656
rect 14967 25653 14979 25687
rect 15672 25684 15700 25715
rect 16114 25712 16120 25724
rect 16172 25712 16178 25764
rect 21266 25712 21272 25764
rect 21324 25752 21330 25764
rect 21422 25755 21480 25761
rect 21422 25752 21434 25755
rect 21324 25724 21434 25752
rect 21324 25712 21330 25724
rect 21422 25721 21434 25724
rect 21468 25721 21480 25755
rect 21422 25715 21480 25721
rect 24121 25755 24179 25761
rect 24121 25721 24133 25755
rect 24167 25721 24179 25755
rect 24121 25715 24179 25721
rect 18046 25684 18052 25696
rect 15672 25656 18052 25684
rect 14921 25647 14979 25653
rect 18046 25644 18052 25656
rect 18104 25644 18110 25696
rect 22554 25684 22560 25696
rect 22515 25656 22560 25684
rect 22554 25644 22560 25656
rect 22612 25684 22618 25696
rect 23014 25684 23020 25696
rect 22612 25656 23020 25684
rect 22612 25644 22618 25656
rect 23014 25644 23020 25656
rect 23072 25644 23078 25696
rect 24136 25684 24164 25715
rect 26050 25712 26056 25764
rect 26108 25752 26114 25764
rect 26804 25752 26832 25783
rect 27982 25780 27988 25792
rect 28040 25780 28046 25832
rect 26108 25724 26832 25752
rect 27056 25755 27114 25761
rect 26108 25712 26114 25724
rect 27056 25721 27068 25755
rect 27102 25752 27114 25755
rect 27430 25752 27436 25764
rect 27102 25724 27436 25752
rect 27102 25721 27114 25724
rect 27056 25715 27114 25721
rect 27430 25712 27436 25724
rect 27488 25712 27494 25764
rect 28074 25684 28080 25696
rect 24136 25656 28080 25684
rect 28074 25644 28080 25656
rect 28132 25684 28138 25696
rect 28169 25687 28227 25693
rect 28169 25684 28181 25687
rect 28132 25656 28181 25684
rect 28132 25644 28138 25656
rect 28169 25653 28181 25656
rect 28215 25653 28227 25687
rect 28169 25647 28227 25653
rect 1104 25594 28888 25616
rect 1104 25542 10246 25594
rect 10298 25542 10310 25594
rect 10362 25542 10374 25594
rect 10426 25542 10438 25594
rect 10490 25542 19510 25594
rect 19562 25542 19574 25594
rect 19626 25542 19638 25594
rect 19690 25542 19702 25594
rect 19754 25542 28888 25594
rect 1104 25520 28888 25542
rect 4798 25480 4804 25492
rect 4759 25452 4804 25480
rect 4798 25440 4804 25452
rect 4856 25440 4862 25492
rect 5350 25440 5356 25492
rect 5408 25480 5414 25492
rect 5442 25480 5448 25492
rect 5408 25452 5448 25480
rect 5408 25440 5414 25452
rect 5442 25440 5448 25452
rect 5500 25440 5506 25492
rect 7929 25483 7987 25489
rect 7929 25449 7941 25483
rect 7975 25480 7987 25483
rect 8018 25480 8024 25492
rect 7975 25452 8024 25480
rect 7975 25449 7987 25452
rect 7929 25443 7987 25449
rect 8018 25440 8024 25452
rect 8076 25440 8082 25492
rect 8110 25440 8116 25492
rect 8168 25480 8174 25492
rect 8481 25483 8539 25489
rect 8481 25480 8493 25483
rect 8168 25452 8493 25480
rect 8168 25440 8174 25452
rect 8481 25449 8493 25452
rect 8527 25449 8539 25483
rect 8481 25443 8539 25449
rect 9030 25440 9036 25492
rect 9088 25480 9094 25492
rect 9309 25483 9367 25489
rect 9309 25480 9321 25483
rect 9088 25452 9321 25480
rect 9088 25440 9094 25452
rect 9309 25449 9321 25452
rect 9355 25449 9367 25483
rect 9309 25443 9367 25449
rect 10689 25483 10747 25489
rect 10689 25449 10701 25483
rect 10735 25480 10747 25483
rect 10778 25480 10784 25492
rect 10735 25452 10784 25480
rect 10735 25449 10747 25452
rect 10689 25443 10747 25449
rect 10778 25440 10784 25452
rect 10836 25440 10842 25492
rect 12526 25440 12532 25492
rect 12584 25480 12590 25492
rect 13173 25483 13231 25489
rect 13173 25480 13185 25483
rect 12584 25452 13185 25480
rect 12584 25440 12590 25452
rect 13173 25449 13185 25452
rect 13219 25480 13231 25483
rect 13814 25480 13820 25492
rect 13219 25452 13820 25480
rect 13219 25449 13231 25452
rect 13173 25443 13231 25449
rect 13814 25440 13820 25452
rect 13872 25440 13878 25492
rect 14182 25480 14188 25492
rect 13924 25452 14188 25480
rect 1762 25412 1768 25424
rect 1723 25384 1768 25412
rect 1762 25372 1768 25384
rect 1820 25372 1826 25424
rect 2130 25372 2136 25424
rect 2188 25412 2194 25424
rect 2188 25384 2636 25412
rect 2188 25372 2194 25384
rect 2608 25356 2636 25384
rect 7374 25372 7380 25424
rect 7432 25412 7438 25424
rect 10134 25412 10140 25424
rect 7432 25384 8432 25412
rect 7432 25372 7438 25384
rect 2498 25344 2504 25356
rect 2459 25316 2504 25344
rect 2498 25304 2504 25316
rect 2556 25304 2562 25356
rect 2590 25304 2596 25356
rect 2648 25344 2654 25356
rect 2777 25347 2835 25353
rect 2777 25344 2789 25347
rect 2648 25316 2789 25344
rect 2648 25304 2654 25316
rect 2777 25313 2789 25316
rect 2823 25313 2835 25347
rect 2777 25307 2835 25313
rect 3973 25347 4031 25353
rect 3973 25313 3985 25347
rect 4019 25344 4031 25347
rect 4246 25344 4252 25356
rect 4019 25316 4252 25344
rect 4019 25313 4031 25316
rect 3973 25307 4031 25313
rect 4246 25304 4252 25316
rect 4304 25304 4310 25356
rect 4709 25347 4767 25353
rect 4709 25313 4721 25347
rect 4755 25344 4767 25347
rect 5442 25344 5448 25356
rect 4755 25316 5448 25344
rect 4755 25313 4767 25316
rect 4709 25307 4767 25313
rect 5442 25304 5448 25316
rect 5500 25304 5506 25356
rect 7558 25304 7564 25356
rect 7616 25344 7622 25356
rect 7745 25347 7803 25353
rect 7745 25344 7757 25347
rect 7616 25316 7757 25344
rect 7616 25304 7622 25316
rect 7745 25313 7757 25316
rect 7791 25313 7803 25347
rect 7745 25307 7803 25313
rect 7834 25304 7840 25356
rect 7892 25344 7898 25356
rect 8404 25353 8432 25384
rect 9232 25384 10140 25412
rect 9232 25356 9260 25384
rect 10134 25372 10140 25384
rect 10192 25412 10198 25424
rect 10870 25412 10876 25424
rect 10192 25384 10876 25412
rect 10192 25372 10198 25384
rect 10870 25372 10876 25384
rect 10928 25372 10934 25424
rect 13924 25412 13952 25452
rect 14182 25440 14188 25452
rect 14240 25440 14246 25492
rect 15381 25483 15439 25489
rect 15381 25449 15393 25483
rect 15427 25480 15439 25483
rect 15562 25480 15568 25492
rect 15427 25452 15568 25480
rect 15427 25449 15439 25452
rect 15381 25443 15439 25449
rect 15562 25440 15568 25452
rect 15620 25440 15626 25492
rect 18325 25483 18383 25489
rect 18325 25449 18337 25483
rect 18371 25449 18383 25483
rect 18325 25443 18383 25449
rect 18693 25483 18751 25489
rect 18693 25449 18705 25483
rect 18739 25480 18751 25483
rect 18966 25480 18972 25492
rect 18739 25452 18972 25480
rect 18739 25449 18751 25452
rect 18693 25443 18751 25449
rect 14274 25412 14280 25424
rect 13832 25384 13952 25412
rect 14108 25384 14280 25412
rect 7929 25347 7987 25353
rect 7929 25344 7941 25347
rect 7892 25316 7941 25344
rect 7892 25304 7898 25316
rect 7929 25313 7941 25316
rect 7975 25313 7987 25347
rect 7929 25307 7987 25313
rect 8389 25347 8447 25353
rect 8389 25313 8401 25347
rect 8435 25313 8447 25347
rect 8389 25307 8447 25313
rect 8573 25347 8631 25353
rect 8573 25313 8585 25347
rect 8619 25313 8631 25347
rect 9214 25344 9220 25356
rect 9175 25316 9220 25344
rect 8573 25307 8631 25313
rect 3418 25276 3424 25288
rect 3379 25248 3424 25276
rect 3418 25236 3424 25248
rect 3476 25236 3482 25288
rect 8294 25236 8300 25288
rect 8352 25276 8358 25288
rect 8588 25276 8616 25307
rect 9214 25304 9220 25316
rect 9272 25304 9278 25356
rect 9398 25344 9404 25356
rect 9359 25316 9404 25344
rect 9398 25304 9404 25316
rect 9456 25304 9462 25356
rect 10594 25344 10600 25356
rect 10555 25316 10600 25344
rect 10594 25304 10600 25316
rect 10652 25304 10658 25356
rect 13081 25347 13139 25353
rect 13081 25313 13093 25347
rect 13127 25344 13139 25347
rect 13262 25344 13268 25356
rect 13127 25316 13268 25344
rect 13127 25313 13139 25316
rect 13081 25307 13139 25313
rect 13262 25304 13268 25316
rect 13320 25304 13326 25356
rect 8352 25248 8616 25276
rect 8352 25236 8358 25248
rect 11054 25236 11060 25288
rect 11112 25276 11118 25288
rect 13832 25276 13860 25384
rect 14108 25353 14136 25384
rect 14274 25372 14280 25384
rect 14332 25372 14338 25424
rect 18340 25412 18368 25443
rect 18966 25440 18972 25452
rect 19024 25440 19030 25492
rect 26605 25483 26663 25489
rect 26605 25480 26617 25483
rect 22066 25452 26617 25480
rect 19766 25415 19824 25421
rect 19766 25412 19778 25415
rect 18340 25384 19778 25412
rect 19766 25381 19778 25384
rect 19812 25381 19824 25415
rect 19766 25375 19824 25381
rect 21453 25415 21511 25421
rect 21453 25381 21465 25415
rect 21499 25412 21511 25415
rect 21818 25412 21824 25424
rect 21499 25384 21824 25412
rect 21499 25381 21511 25384
rect 21453 25375 21511 25381
rect 21818 25372 21824 25384
rect 21876 25372 21882 25424
rect 13981 25347 14039 25353
rect 13981 25313 13993 25347
rect 14027 25344 14039 25347
rect 14074 25347 14136 25353
rect 14027 25313 14044 25344
rect 13981 25307 14044 25313
rect 14074 25313 14086 25347
rect 14120 25316 14136 25347
rect 14190 25347 14248 25353
rect 14120 25313 14132 25316
rect 14074 25307 14132 25313
rect 14190 25313 14202 25347
rect 14236 25344 14248 25347
rect 14369 25347 14427 25353
rect 14236 25313 14249 25344
rect 14190 25307 14249 25313
rect 14369 25313 14381 25347
rect 14415 25313 14427 25347
rect 14369 25307 14427 25313
rect 14016 25276 14044 25307
rect 14221 25276 14249 25307
rect 11112 25248 14044 25276
rect 14108 25248 14249 25276
rect 11112 25236 11118 25248
rect 1578 25168 1584 25220
rect 1636 25208 1642 25220
rect 1949 25211 2007 25217
rect 1949 25208 1961 25211
rect 1636 25180 1961 25208
rect 1636 25168 1642 25180
rect 1949 25177 1961 25180
rect 1995 25208 2007 25211
rect 6362 25208 6368 25220
rect 1995 25180 6368 25208
rect 1995 25177 2007 25180
rect 1949 25171 2007 25177
rect 6362 25168 6368 25180
rect 6420 25168 6426 25220
rect 12618 25168 12624 25220
rect 12676 25208 12682 25220
rect 13170 25208 13176 25220
rect 12676 25180 13176 25208
rect 12676 25168 12682 25180
rect 13170 25168 13176 25180
rect 13228 25168 13234 25220
rect 14108 25152 14136 25248
rect 14274 25168 14280 25220
rect 14332 25208 14338 25220
rect 14384 25208 14412 25307
rect 14918 25304 14924 25356
rect 14976 25344 14982 25356
rect 15657 25347 15715 25353
rect 15657 25344 15669 25347
rect 14976 25316 15669 25344
rect 14976 25304 14982 25316
rect 15657 25313 15669 25316
rect 15703 25313 15715 25347
rect 15657 25307 15715 25313
rect 15749 25347 15807 25353
rect 15749 25313 15761 25347
rect 15795 25313 15807 25347
rect 15749 25307 15807 25313
rect 15194 25236 15200 25288
rect 15252 25276 15258 25288
rect 15470 25276 15476 25288
rect 15252 25248 15476 25276
rect 15252 25236 15258 25248
rect 15470 25236 15476 25248
rect 15528 25236 15534 25288
rect 15764 25276 15792 25307
rect 15838 25304 15844 25356
rect 15896 25344 15902 25356
rect 16022 25344 16028 25356
rect 15896 25316 15941 25344
rect 15983 25316 16028 25344
rect 15896 25304 15902 25316
rect 16022 25304 16028 25316
rect 16080 25304 16086 25356
rect 17310 25304 17316 25356
rect 17368 25344 17374 25356
rect 22066 25344 22094 25452
rect 26605 25449 26617 25452
rect 26651 25449 26663 25483
rect 26605 25443 26663 25449
rect 26694 25440 26700 25492
rect 26752 25480 26758 25492
rect 26789 25483 26847 25489
rect 26789 25480 26801 25483
rect 26752 25452 26801 25480
rect 26752 25440 26758 25452
rect 26789 25449 26801 25452
rect 26835 25480 26847 25483
rect 27522 25480 27528 25492
rect 26835 25452 27528 25480
rect 26835 25449 26847 25452
rect 26789 25443 26847 25449
rect 27522 25440 27528 25452
rect 27580 25440 27586 25492
rect 23014 25372 23020 25424
rect 23072 25412 23078 25424
rect 25501 25415 25559 25421
rect 25501 25412 25513 25415
rect 23072 25384 25513 25412
rect 23072 25372 23078 25384
rect 25501 25381 25513 25384
rect 25547 25381 25559 25415
rect 25501 25375 25559 25381
rect 25866 25372 25872 25424
rect 25924 25412 25930 25424
rect 26234 25412 26240 25424
rect 25924 25384 25969 25412
rect 26195 25384 26240 25412
rect 25924 25372 25930 25384
rect 26234 25372 26240 25384
rect 26292 25372 26298 25424
rect 17368 25316 22094 25344
rect 17368 25304 17374 25316
rect 22278 25304 22284 25356
rect 22336 25344 22342 25356
rect 22557 25347 22615 25353
rect 22557 25344 22569 25347
rect 22336 25316 22569 25344
rect 22336 25304 22342 25316
rect 22557 25313 22569 25316
rect 22603 25313 22615 25347
rect 22557 25307 22615 25313
rect 22649 25347 22707 25353
rect 22649 25313 22661 25347
rect 22695 25313 22707 25347
rect 22649 25307 22707 25313
rect 17034 25276 17040 25288
rect 15764 25248 17040 25276
rect 17034 25236 17040 25248
rect 17092 25236 17098 25288
rect 18785 25279 18843 25285
rect 18785 25245 18797 25279
rect 18831 25245 18843 25279
rect 18785 25239 18843 25245
rect 18969 25279 19027 25285
rect 18969 25245 18981 25279
rect 19015 25276 19027 25279
rect 19242 25276 19248 25288
rect 19015 25248 19248 25276
rect 19015 25245 19027 25248
rect 18969 25239 19027 25245
rect 14332 25180 14412 25208
rect 14332 25168 14338 25180
rect 15286 25168 15292 25220
rect 15344 25208 15350 25220
rect 15562 25208 15568 25220
rect 15344 25180 15568 25208
rect 15344 25168 15350 25180
rect 15562 25168 15568 25180
rect 15620 25168 15626 25220
rect 4157 25143 4215 25149
rect 4157 25109 4169 25143
rect 4203 25140 4215 25143
rect 4522 25140 4528 25152
rect 4203 25112 4528 25140
rect 4203 25109 4215 25112
rect 4157 25103 4215 25109
rect 4522 25100 4528 25112
rect 4580 25100 4586 25152
rect 5258 25100 5264 25152
rect 5316 25140 5322 25152
rect 6270 25140 6276 25152
rect 5316 25112 6276 25140
rect 5316 25100 5322 25112
rect 6270 25100 6276 25112
rect 6328 25100 6334 25152
rect 13722 25140 13728 25152
rect 13683 25112 13728 25140
rect 13722 25100 13728 25112
rect 13780 25100 13786 25152
rect 14090 25100 14096 25152
rect 14148 25100 14154 25152
rect 15194 25100 15200 25152
rect 15252 25140 15258 25152
rect 15378 25140 15384 25152
rect 15252 25112 15384 25140
rect 15252 25100 15258 25112
rect 15378 25100 15384 25112
rect 15436 25100 15442 25152
rect 18800 25140 18828 25239
rect 19242 25236 19248 25248
rect 19300 25236 19306 25288
rect 19334 25236 19340 25288
rect 19392 25276 19398 25288
rect 19521 25279 19579 25285
rect 19521 25276 19533 25279
rect 19392 25248 19533 25276
rect 19392 25236 19398 25248
rect 19521 25245 19533 25248
rect 19567 25245 19579 25279
rect 22664 25276 22692 25307
rect 22738 25304 22744 25356
rect 22796 25344 22802 25356
rect 23109 25347 23167 25353
rect 23109 25344 23121 25347
rect 22796 25316 23121 25344
rect 22796 25304 22802 25316
rect 23109 25313 23121 25316
rect 23155 25313 23167 25347
rect 24486 25344 24492 25356
rect 24447 25316 24492 25344
rect 23109 25307 23167 25313
rect 24486 25304 24492 25316
rect 24544 25304 24550 25356
rect 25682 25304 25688 25356
rect 25740 25344 25746 25356
rect 25777 25347 25835 25353
rect 25777 25344 25789 25347
rect 25740 25316 25789 25344
rect 25740 25304 25746 25316
rect 25777 25313 25789 25316
rect 25823 25344 25835 25347
rect 27985 25347 28043 25353
rect 27985 25344 27997 25347
rect 25823 25316 27997 25344
rect 25823 25313 25835 25316
rect 25777 25307 25835 25313
rect 27985 25313 27997 25316
rect 28031 25313 28043 25347
rect 27985 25307 28043 25313
rect 23382 25276 23388 25288
rect 22664 25248 23388 25276
rect 19521 25239 19579 25245
rect 23382 25236 23388 25248
rect 23440 25236 23446 25288
rect 24581 25279 24639 25285
rect 24581 25245 24593 25279
rect 24627 25245 24639 25279
rect 24581 25239 24639 25245
rect 24765 25279 24823 25285
rect 24765 25245 24777 25279
rect 24811 25276 24823 25279
rect 24946 25276 24952 25288
rect 24811 25248 24952 25276
rect 24811 25245 24823 25248
rect 24765 25239 24823 25245
rect 19058 25168 19064 25220
rect 19116 25208 19122 25220
rect 19352 25208 19380 25236
rect 19116 25180 19380 25208
rect 21637 25211 21695 25217
rect 19116 25168 19122 25180
rect 21637 25177 21649 25211
rect 21683 25208 21695 25211
rect 22094 25208 22100 25220
rect 21683 25180 22100 25208
rect 21683 25177 21695 25180
rect 21637 25171 21695 25177
rect 22094 25168 22100 25180
rect 22152 25168 22158 25220
rect 24596 25208 24624 25239
rect 24946 25236 24952 25248
rect 25004 25276 25010 25288
rect 25130 25276 25136 25288
rect 25004 25248 25136 25276
rect 25004 25236 25010 25248
rect 25130 25236 25136 25248
rect 25188 25236 25194 25288
rect 25498 25236 25504 25288
rect 25556 25236 25562 25288
rect 24596 25180 25176 25208
rect 25148 25152 25176 25180
rect 20898 25140 20904 25152
rect 18800 25112 20904 25140
rect 20898 25100 20904 25112
rect 20956 25100 20962 25152
rect 22922 25140 22928 25152
rect 22883 25112 22928 25140
rect 22922 25100 22928 25112
rect 22980 25100 22986 25152
rect 23014 25100 23020 25152
rect 23072 25140 23078 25152
rect 24121 25143 24179 25149
rect 23072 25112 23117 25140
rect 23072 25100 23078 25112
rect 24121 25109 24133 25143
rect 24167 25140 24179 25143
rect 24762 25140 24768 25152
rect 24167 25112 24768 25140
rect 24167 25109 24179 25112
rect 24121 25103 24179 25109
rect 24762 25100 24768 25112
rect 24820 25100 24826 25152
rect 25130 25100 25136 25152
rect 25188 25100 25194 25152
rect 27522 25100 27528 25152
rect 27580 25140 27586 25152
rect 28077 25143 28135 25149
rect 28077 25140 28089 25143
rect 27580 25112 28089 25140
rect 27580 25100 27586 25112
rect 28077 25109 28089 25112
rect 28123 25109 28135 25143
rect 28077 25103 28135 25109
rect 1104 25050 28888 25072
rect 1104 24998 5614 25050
rect 5666 24998 5678 25050
rect 5730 24998 5742 25050
rect 5794 24998 5806 25050
rect 5858 24998 14878 25050
rect 14930 24998 14942 25050
rect 14994 24998 15006 25050
rect 15058 24998 15070 25050
rect 15122 24998 24142 25050
rect 24194 24998 24206 25050
rect 24258 24998 24270 25050
rect 24322 24998 24334 25050
rect 24386 24998 28888 25050
rect 1104 24976 28888 24998
rect 10229 24939 10287 24945
rect 10229 24905 10241 24939
rect 10275 24936 10287 24939
rect 10594 24936 10600 24948
rect 10275 24908 10600 24936
rect 10275 24905 10287 24908
rect 10229 24899 10287 24905
rect 10594 24896 10600 24908
rect 10652 24896 10658 24948
rect 10870 24896 10876 24948
rect 10928 24936 10934 24948
rect 13173 24939 13231 24945
rect 13173 24936 13185 24939
rect 10928 24908 13185 24936
rect 10928 24896 10934 24908
rect 13173 24905 13185 24908
rect 13219 24905 13231 24939
rect 13173 24899 13231 24905
rect 13725 24939 13783 24945
rect 13725 24905 13737 24939
rect 13771 24936 13783 24939
rect 14274 24936 14280 24948
rect 13771 24908 14280 24936
rect 13771 24905 13783 24908
rect 13725 24899 13783 24905
rect 14274 24896 14280 24908
rect 14332 24896 14338 24948
rect 15565 24939 15623 24945
rect 15565 24905 15577 24939
rect 15611 24936 15623 24939
rect 16022 24936 16028 24948
rect 15611 24908 16028 24936
rect 15611 24905 15623 24908
rect 15565 24899 15623 24905
rect 16022 24896 16028 24908
rect 16080 24896 16086 24948
rect 16117 24939 16175 24945
rect 16117 24905 16129 24939
rect 16163 24936 16175 24939
rect 16574 24936 16580 24948
rect 16163 24908 16580 24936
rect 16163 24905 16175 24908
rect 16117 24899 16175 24905
rect 16574 24896 16580 24908
rect 16632 24896 16638 24948
rect 23382 24896 23388 24948
rect 23440 24936 23446 24948
rect 24121 24939 24179 24945
rect 24121 24936 24133 24939
rect 23440 24908 24133 24936
rect 23440 24896 23446 24908
rect 24121 24905 24133 24908
rect 24167 24905 24179 24939
rect 24121 24899 24179 24905
rect 25130 24896 25136 24948
rect 25188 24936 25194 24948
rect 26234 24936 26240 24948
rect 25188 24908 26240 24936
rect 25188 24896 25194 24908
rect 26234 24896 26240 24908
rect 26292 24936 26298 24948
rect 26605 24939 26663 24945
rect 26605 24936 26617 24939
rect 26292 24908 26617 24936
rect 26292 24896 26298 24908
rect 26605 24905 26617 24908
rect 26651 24905 26663 24939
rect 27430 24936 27436 24948
rect 27391 24908 27436 24936
rect 26605 24899 26663 24905
rect 27430 24896 27436 24908
rect 27488 24896 27494 24948
rect 6086 24868 6092 24880
rect 5828 24840 6092 24868
rect 1857 24735 1915 24741
rect 1857 24701 1869 24735
rect 1903 24732 1915 24735
rect 2222 24732 2228 24744
rect 1903 24704 2228 24732
rect 1903 24701 1915 24704
rect 1857 24695 1915 24701
rect 2222 24692 2228 24704
rect 2280 24692 2286 24744
rect 2498 24692 2504 24744
rect 2556 24732 2562 24744
rect 2608 24732 2636 24786
rect 5258 24760 5264 24812
rect 5316 24760 5322 24812
rect 5828 24744 5856 24840
rect 6086 24828 6092 24840
rect 6144 24828 6150 24880
rect 11330 24868 11336 24880
rect 10796 24840 11336 24868
rect 10796 24812 10824 24840
rect 11330 24828 11336 24840
rect 11388 24828 11394 24880
rect 12710 24868 12716 24880
rect 11992 24840 12716 24868
rect 5920 24772 6408 24800
rect 2682 24732 2688 24744
rect 2556 24704 2688 24732
rect 2556 24692 2562 24704
rect 2682 24692 2688 24704
rect 2740 24732 2746 24744
rect 4890 24732 4896 24744
rect 2740 24704 4896 24732
rect 2740 24692 2746 24704
rect 4890 24692 4896 24704
rect 4948 24692 4954 24744
rect 5074 24732 5080 24744
rect 5035 24704 5080 24732
rect 5074 24692 5080 24704
rect 5132 24692 5138 24744
rect 5810 24732 5816 24744
rect 5368 24704 5816 24732
rect 1578 24664 1584 24676
rect 1539 24636 1584 24664
rect 1578 24624 1584 24636
rect 1636 24624 1642 24676
rect 1762 24624 1768 24676
rect 1820 24664 1826 24676
rect 1949 24667 2007 24673
rect 1949 24664 1961 24667
rect 1820 24636 1961 24664
rect 1820 24624 1826 24636
rect 1949 24633 1961 24636
rect 1995 24633 2007 24667
rect 1949 24627 2007 24633
rect 2038 24624 2044 24676
rect 2096 24664 2102 24676
rect 2317 24667 2375 24673
rect 2317 24664 2329 24667
rect 2096 24636 2329 24664
rect 2096 24624 2102 24636
rect 2317 24633 2329 24636
rect 2363 24664 2375 24667
rect 4709 24667 4767 24673
rect 4709 24664 4721 24667
rect 2363 24636 4721 24664
rect 2363 24633 2375 24636
rect 2317 24627 2375 24633
rect 4709 24633 4721 24636
rect 4755 24633 4767 24667
rect 4709 24627 4767 24633
rect 4985 24667 5043 24673
rect 4985 24633 4997 24667
rect 5031 24664 5043 24667
rect 5368 24664 5396 24704
rect 5810 24692 5816 24704
rect 5868 24692 5874 24744
rect 5031 24636 5396 24664
rect 5445 24667 5503 24673
rect 5031 24633 5043 24636
rect 4985 24627 5043 24633
rect 5445 24633 5457 24667
rect 5491 24664 5503 24667
rect 5534 24664 5540 24676
rect 5491 24636 5540 24664
rect 5491 24633 5503 24636
rect 5445 24627 5503 24633
rect 1486 24556 1492 24608
rect 1544 24596 1550 24608
rect 2498 24596 2504 24608
rect 1544 24568 2504 24596
rect 1544 24556 1550 24568
rect 2498 24556 2504 24568
rect 2556 24556 2562 24608
rect 2682 24596 2688 24608
rect 2643 24568 2688 24596
rect 2682 24556 2688 24568
rect 2740 24556 2746 24608
rect 2869 24599 2927 24605
rect 2869 24565 2881 24599
rect 2915 24596 2927 24599
rect 3694 24596 3700 24608
rect 2915 24568 3700 24596
rect 2915 24565 2927 24568
rect 2869 24559 2927 24565
rect 3694 24556 3700 24568
rect 3752 24556 3758 24608
rect 4724 24596 4752 24627
rect 5534 24624 5540 24636
rect 5592 24624 5598 24676
rect 5920 24664 5948 24772
rect 6380 24732 6408 24772
rect 6454 24760 6460 24812
rect 6512 24800 6518 24812
rect 9214 24800 9220 24812
rect 6512 24772 9220 24800
rect 6512 24760 6518 24772
rect 9214 24760 9220 24772
rect 9272 24760 9278 24812
rect 9950 24760 9956 24812
rect 10008 24800 10014 24812
rect 10689 24803 10747 24809
rect 10689 24800 10701 24803
rect 10008 24772 10701 24800
rect 10008 24760 10014 24772
rect 10689 24769 10701 24772
rect 10735 24769 10747 24803
rect 10689 24763 10747 24769
rect 10778 24760 10784 24812
rect 10836 24800 10842 24812
rect 10836 24772 10881 24800
rect 10836 24760 10842 24772
rect 10502 24732 10508 24744
rect 6380 24704 10508 24732
rect 10502 24692 10508 24704
rect 10560 24692 10566 24744
rect 11992 24741 12020 24840
rect 12710 24828 12716 24840
rect 12768 24868 12774 24880
rect 12768 24840 13308 24868
rect 12768 24828 12774 24840
rect 12250 24760 12256 24812
rect 12308 24760 12314 24812
rect 11977 24735 12035 24741
rect 11977 24701 11989 24735
rect 12023 24701 12035 24735
rect 11977 24695 12035 24701
rect 12069 24735 12127 24741
rect 12069 24701 12081 24735
rect 12115 24701 12127 24735
rect 12069 24695 12127 24701
rect 12161 24735 12219 24741
rect 12161 24701 12173 24735
rect 12207 24732 12219 24735
rect 12268 24732 12296 24760
rect 12207 24704 12296 24732
rect 12345 24735 12403 24741
rect 12207 24701 12219 24704
rect 12161 24695 12219 24701
rect 12345 24701 12357 24735
rect 12391 24732 12403 24735
rect 12710 24732 12716 24744
rect 12391 24704 12716 24732
rect 12391 24701 12403 24704
rect 12345 24695 12403 24701
rect 7650 24664 7656 24676
rect 5644 24636 5948 24664
rect 6012 24636 7656 24664
rect 5644 24596 5672 24636
rect 5810 24596 5816 24608
rect 4724 24568 5672 24596
rect 5771 24568 5816 24596
rect 5810 24556 5816 24568
rect 5868 24556 5874 24608
rect 6012 24605 6040 24636
rect 7650 24624 7656 24636
rect 7708 24624 7714 24676
rect 12084 24664 12112 24695
rect 12710 24692 12716 24704
rect 12768 24692 12774 24744
rect 13280 24732 13308 24840
rect 13354 24828 13360 24880
rect 13412 24868 13418 24880
rect 17494 24868 17500 24880
rect 13412 24840 13492 24868
rect 13412 24828 13418 24840
rect 13464 24741 13492 24840
rect 16408 24840 17500 24868
rect 16114 24800 16120 24812
rect 15304 24772 16120 24800
rect 13357 24735 13415 24741
rect 13357 24732 13369 24735
rect 13280 24704 13369 24732
rect 13357 24701 13369 24704
rect 13403 24701 13415 24735
rect 13357 24695 13415 24701
rect 13449 24735 13507 24741
rect 13449 24701 13461 24735
rect 13495 24701 13507 24735
rect 13449 24695 13507 24701
rect 13541 24735 13599 24741
rect 13541 24701 13553 24735
rect 13587 24701 13599 24735
rect 13541 24695 13599 24701
rect 12250 24664 12256 24676
rect 12084 24636 12256 24664
rect 12250 24624 12256 24636
rect 12308 24624 12314 24676
rect 13556 24664 13584 24695
rect 15102 24692 15108 24744
rect 15160 24741 15166 24744
rect 15304 24741 15332 24772
rect 16114 24760 16120 24772
rect 16172 24760 16178 24812
rect 15160 24735 15219 24741
rect 15160 24701 15173 24735
rect 15207 24701 15219 24735
rect 15160 24695 15219 24701
rect 15289 24735 15347 24741
rect 15289 24701 15301 24735
rect 15335 24701 15347 24735
rect 15289 24695 15347 24701
rect 15160 24692 15166 24695
rect 15378 24692 15384 24744
rect 15436 24732 15442 24744
rect 15654 24732 15660 24744
rect 15436 24704 15660 24732
rect 15436 24692 15442 24704
rect 15654 24692 15660 24704
rect 15712 24692 15718 24744
rect 16206 24692 16212 24744
rect 16264 24732 16270 24744
rect 16408 24741 16436 24840
rect 17494 24828 17500 24840
rect 17552 24828 17558 24880
rect 22278 24868 22284 24880
rect 22239 24840 22284 24868
rect 22278 24828 22284 24840
rect 22336 24828 22342 24880
rect 27890 24828 27896 24880
rect 27948 24868 27954 24880
rect 27948 24840 28028 24868
rect 27948 24828 27954 24840
rect 19984 24812 20036 24818
rect 17034 24800 17040 24812
rect 16500 24772 17040 24800
rect 16500 24741 16528 24772
rect 17034 24760 17040 24772
rect 17092 24800 17098 24812
rect 17773 24803 17831 24809
rect 17773 24800 17785 24803
rect 17092 24772 17785 24800
rect 17092 24760 17098 24772
rect 17773 24769 17785 24772
rect 17819 24769 17831 24803
rect 17773 24763 17831 24769
rect 21818 24760 21824 24812
rect 21876 24800 21882 24812
rect 28000 24809 28028 24840
rect 27985 24803 28043 24809
rect 21876 24772 22140 24800
rect 21876 24760 21882 24772
rect 19984 24754 20036 24760
rect 16393 24735 16451 24741
rect 16393 24732 16405 24735
rect 16264 24704 16405 24732
rect 16264 24692 16270 24704
rect 16393 24701 16405 24704
rect 16439 24701 16451 24735
rect 16393 24695 16451 24701
rect 16485 24735 16543 24741
rect 16485 24701 16497 24735
rect 16531 24701 16543 24735
rect 16485 24695 16543 24701
rect 16577 24735 16635 24741
rect 16577 24701 16589 24735
rect 16623 24701 16635 24735
rect 16577 24695 16635 24701
rect 16761 24735 16819 24741
rect 16761 24701 16773 24735
rect 16807 24701 16819 24735
rect 16761 24695 16819 24701
rect 12452 24636 13584 24664
rect 5997 24599 6055 24605
rect 5997 24565 6009 24599
rect 6043 24565 6055 24599
rect 5997 24559 6055 24565
rect 6086 24556 6092 24608
rect 6144 24596 6150 24608
rect 10597 24599 10655 24605
rect 10597 24596 10609 24599
rect 6144 24568 10609 24596
rect 6144 24556 6150 24568
rect 10597 24565 10609 24568
rect 10643 24565 10655 24599
rect 10597 24559 10655 24565
rect 11330 24556 11336 24608
rect 11388 24596 11394 24608
rect 11514 24596 11520 24608
rect 11388 24568 11520 24596
rect 11388 24556 11394 24568
rect 11514 24556 11520 24568
rect 11572 24596 11578 24608
rect 12452 24596 12480 24636
rect 15838 24624 15844 24676
rect 15896 24664 15902 24676
rect 16592 24664 16620 24695
rect 15896 24636 16620 24664
rect 15896 24624 15902 24636
rect 16666 24624 16672 24676
rect 16724 24664 16730 24676
rect 16776 24664 16804 24695
rect 17310 24692 17316 24744
rect 17368 24732 17374 24744
rect 17589 24735 17647 24741
rect 17589 24732 17601 24735
rect 17368 24704 17601 24732
rect 17368 24692 17374 24704
rect 17589 24701 17601 24704
rect 17635 24701 17647 24735
rect 20438 24732 20444 24744
rect 17589 24695 17647 24701
rect 20272 24704 20444 24732
rect 20162 24664 20168 24676
rect 16724 24636 16804 24664
rect 20123 24636 20168 24664
rect 16724 24624 16730 24636
rect 20162 24624 20168 24636
rect 20220 24624 20226 24676
rect 11572 24568 12480 24596
rect 13173 24599 13231 24605
rect 11572 24556 11578 24568
rect 13173 24565 13185 24599
rect 13219 24596 13231 24599
rect 20272 24596 20300 24704
rect 20438 24692 20444 24704
rect 20496 24692 20502 24744
rect 20898 24732 20904 24744
rect 20811 24704 20904 24732
rect 20898 24692 20904 24704
rect 20956 24732 20962 24744
rect 21910 24732 21916 24744
rect 20956 24704 21916 24732
rect 20956 24692 20962 24704
rect 21910 24692 21916 24704
rect 21968 24692 21974 24744
rect 22112 24741 22140 24772
rect 27985 24769 27997 24803
rect 28031 24769 28043 24803
rect 27985 24763 28043 24769
rect 22097 24735 22155 24741
rect 22097 24701 22109 24735
rect 22143 24701 22155 24735
rect 22097 24695 22155 24701
rect 22741 24735 22799 24741
rect 22741 24701 22753 24735
rect 22787 24732 22799 24735
rect 25225 24735 25283 24741
rect 25225 24732 25237 24735
rect 22787 24704 25237 24732
rect 22787 24701 22799 24704
rect 22741 24695 22799 24701
rect 25225 24701 25237 24704
rect 25271 24732 25283 24735
rect 25958 24732 25964 24744
rect 25271 24704 25964 24732
rect 25271 24701 25283 24704
rect 25225 24695 25283 24701
rect 25958 24692 25964 24704
rect 26016 24692 26022 24744
rect 27798 24732 27804 24744
rect 27759 24704 27804 24732
rect 27798 24692 27804 24704
rect 27856 24692 27862 24744
rect 27893 24735 27951 24741
rect 27893 24701 27905 24735
rect 27939 24732 27951 24735
rect 28074 24732 28080 24744
rect 27939 24704 28080 24732
rect 27939 24701 27951 24704
rect 27893 24695 27951 24701
rect 28074 24692 28080 24704
rect 28132 24692 28138 24744
rect 20530 24664 20536 24676
rect 20491 24636 20536 24664
rect 20530 24624 20536 24636
rect 20588 24624 20594 24676
rect 21726 24624 21732 24676
rect 21784 24664 21790 24676
rect 22278 24664 22284 24676
rect 21784 24636 22284 24664
rect 21784 24624 21790 24636
rect 22278 24624 22284 24636
rect 22336 24664 22342 24676
rect 22646 24664 22652 24676
rect 22336 24636 22652 24664
rect 22336 24624 22342 24636
rect 22646 24624 22652 24636
rect 22704 24624 22710 24676
rect 22922 24624 22928 24676
rect 22980 24673 22986 24676
rect 22980 24667 23044 24673
rect 22980 24633 22998 24667
rect 23032 24633 23044 24667
rect 22980 24627 23044 24633
rect 22980 24624 22986 24627
rect 24762 24624 24768 24676
rect 24820 24664 24826 24676
rect 25470 24667 25528 24673
rect 25470 24664 25482 24667
rect 24820 24636 25482 24664
rect 24820 24624 24826 24636
rect 25470 24633 25482 24636
rect 25516 24633 25528 24667
rect 25470 24627 25528 24633
rect 13219 24568 20300 24596
rect 13219 24565 13231 24568
rect 13173 24559 13231 24565
rect 20714 24556 20720 24608
rect 20772 24596 20778 24608
rect 21269 24599 21327 24605
rect 21269 24596 21281 24599
rect 20772 24568 21281 24596
rect 20772 24556 20778 24568
rect 21269 24565 21281 24568
rect 21315 24565 21327 24599
rect 21450 24596 21456 24608
rect 21411 24568 21456 24596
rect 21269 24559 21327 24565
rect 21450 24556 21456 24568
rect 21508 24556 21514 24608
rect 1104 24506 28888 24528
rect 1104 24454 10246 24506
rect 10298 24454 10310 24506
rect 10362 24454 10374 24506
rect 10426 24454 10438 24506
rect 10490 24454 19510 24506
rect 19562 24454 19574 24506
rect 19626 24454 19638 24506
rect 19690 24454 19702 24506
rect 19754 24454 28888 24506
rect 1104 24432 28888 24454
rect 1765 24395 1823 24401
rect 1765 24361 1777 24395
rect 1811 24392 1823 24395
rect 5810 24392 5816 24404
rect 1811 24364 5816 24392
rect 1811 24361 1823 24364
rect 1765 24355 1823 24361
rect 5810 24352 5816 24364
rect 5868 24352 5874 24404
rect 6917 24395 6975 24401
rect 6917 24361 6929 24395
rect 6963 24392 6975 24395
rect 7374 24392 7380 24404
rect 6963 24364 7380 24392
rect 6963 24361 6975 24364
rect 6917 24355 6975 24361
rect 7374 24352 7380 24364
rect 7432 24352 7438 24404
rect 13262 24392 13268 24404
rect 13223 24364 13268 24392
rect 13262 24352 13268 24364
rect 13320 24352 13326 24404
rect 14090 24392 14096 24404
rect 13372 24364 14096 24392
rect 2498 24284 2504 24336
rect 2556 24324 2562 24336
rect 5169 24327 5227 24333
rect 5169 24324 5181 24327
rect 2556 24296 5181 24324
rect 2556 24284 2562 24296
rect 5169 24293 5181 24296
rect 5215 24293 5227 24327
rect 5169 24287 5227 24293
rect 5261 24327 5319 24333
rect 5261 24293 5273 24327
rect 5307 24324 5319 24327
rect 6454 24324 6460 24336
rect 5307 24296 6460 24324
rect 5307 24293 5319 24296
rect 5261 24287 5319 24293
rect 6454 24284 6460 24296
rect 6512 24284 6518 24336
rect 6638 24284 6644 24336
rect 6696 24324 6702 24336
rect 13372 24324 13400 24364
rect 14090 24352 14096 24364
rect 14148 24352 14154 24404
rect 14182 24352 14188 24404
rect 14240 24392 14246 24404
rect 15197 24395 15255 24401
rect 15197 24392 15209 24395
rect 14240 24364 15209 24392
rect 14240 24352 14246 24364
rect 15197 24361 15209 24364
rect 15243 24361 15255 24395
rect 15197 24355 15255 24361
rect 15470 24352 15476 24404
rect 15528 24392 15534 24404
rect 15838 24392 15844 24404
rect 15528 24364 15844 24392
rect 15528 24352 15534 24364
rect 15838 24352 15844 24364
rect 15896 24352 15902 24404
rect 16393 24395 16451 24401
rect 16393 24361 16405 24395
rect 16439 24392 16451 24395
rect 16666 24392 16672 24404
rect 16439 24364 16672 24392
rect 16439 24361 16451 24364
rect 16393 24355 16451 24361
rect 16666 24352 16672 24364
rect 16724 24352 16730 24404
rect 21361 24395 21419 24401
rect 21361 24361 21373 24395
rect 21407 24392 21419 24395
rect 23014 24392 23020 24404
rect 21407 24364 23020 24392
rect 21407 24361 21419 24364
rect 21361 24355 21419 24361
rect 23014 24352 23020 24364
rect 23072 24352 23078 24404
rect 23952 24364 28028 24392
rect 6696 24296 7420 24324
rect 6696 24284 6702 24296
rect 1946 24256 1952 24268
rect 1907 24228 1952 24256
rect 1946 24216 1952 24228
rect 2004 24216 2010 24268
rect 3142 24265 3148 24268
rect 3136 24219 3148 24265
rect 3200 24256 3206 24268
rect 6822 24256 6828 24268
rect 3200 24228 3236 24256
rect 6783 24228 6828 24256
rect 3142 24216 3148 24219
rect 3200 24216 3206 24228
rect 6822 24216 6828 24228
rect 6880 24216 6886 24268
rect 7392 24265 7420 24296
rect 12544 24296 13400 24324
rect 7377 24259 7435 24265
rect 7377 24225 7389 24259
rect 7423 24225 7435 24259
rect 7377 24219 7435 24225
rect 11698 24216 11704 24268
rect 11756 24256 11762 24268
rect 12066 24256 12072 24268
rect 11756 24228 12072 24256
rect 11756 24216 11762 24228
rect 12066 24216 12072 24228
rect 12124 24256 12130 24268
rect 12544 24265 12572 24296
rect 13538 24284 13544 24336
rect 13596 24284 13602 24336
rect 16574 24324 16580 24336
rect 16004 24296 16580 24324
rect 12345 24259 12403 24265
rect 12345 24256 12357 24259
rect 12124 24228 12357 24256
rect 12124 24216 12130 24228
rect 12345 24225 12357 24228
rect 12391 24225 12403 24259
rect 12345 24219 12403 24225
rect 12437 24259 12495 24265
rect 12437 24225 12449 24259
rect 12483 24225 12495 24259
rect 12437 24219 12495 24225
rect 12529 24259 12587 24265
rect 12529 24225 12541 24259
rect 12575 24225 12587 24259
rect 12710 24256 12716 24268
rect 12671 24228 12716 24256
rect 12529 24219 12587 24225
rect 2866 24188 2872 24200
rect 2827 24160 2872 24188
rect 2866 24148 2872 24160
rect 2924 24148 2930 24200
rect 4798 24148 4804 24200
rect 4856 24188 4862 24200
rect 5258 24188 5264 24200
rect 4856 24160 5264 24188
rect 4856 24148 4862 24160
rect 5258 24148 5264 24160
rect 5316 24188 5322 24200
rect 5353 24191 5411 24197
rect 5353 24188 5365 24191
rect 5316 24160 5365 24188
rect 5316 24148 5322 24160
rect 5353 24157 5365 24160
rect 5399 24157 5411 24191
rect 5353 24151 5411 24157
rect 7006 24148 7012 24200
rect 7064 24188 7070 24200
rect 7653 24191 7711 24197
rect 7653 24188 7665 24191
rect 7064 24160 7665 24188
rect 7064 24148 7070 24160
rect 7653 24157 7665 24160
rect 7699 24157 7711 24191
rect 12452 24188 12480 24219
rect 12710 24216 12716 24228
rect 12768 24216 12774 24268
rect 13170 24256 13176 24268
rect 13131 24228 13176 24256
rect 13170 24216 13176 24228
rect 13228 24216 13234 24268
rect 13354 24256 13360 24268
rect 13315 24228 13360 24256
rect 13354 24216 13360 24228
rect 13412 24256 13418 24268
rect 13556 24256 13584 24284
rect 13412 24228 13584 24256
rect 13412 24216 13418 24228
rect 13722 24216 13728 24268
rect 13780 24256 13786 24268
rect 14093 24259 14151 24265
rect 14093 24256 14105 24259
rect 13780 24228 14105 24256
rect 13780 24216 13786 24228
rect 14093 24225 14105 24228
rect 14139 24225 14151 24259
rect 14093 24219 14151 24225
rect 15102 24216 15108 24268
rect 15160 24256 15166 24268
rect 16004 24265 16032 24296
rect 16574 24284 16580 24296
rect 16632 24284 16638 24336
rect 19705 24327 19763 24333
rect 19705 24293 19717 24327
rect 19751 24324 19763 24327
rect 19978 24324 19984 24336
rect 19751 24296 19984 24324
rect 19751 24293 19763 24296
rect 19705 24287 19763 24293
rect 19978 24284 19984 24296
rect 20036 24284 20042 24336
rect 20438 24284 20444 24336
rect 20496 24324 20502 24336
rect 23952 24324 23980 24364
rect 25961 24327 26019 24333
rect 25961 24324 25973 24327
rect 20496 24296 23980 24324
rect 24044 24296 25973 24324
rect 20496 24284 20502 24296
rect 15989 24259 16047 24265
rect 15989 24256 16001 24259
rect 15160 24228 16001 24256
rect 15160 24216 15166 24228
rect 15989 24225 16001 24228
rect 16035 24225 16047 24259
rect 16114 24256 16120 24268
rect 16075 24228 16120 24256
rect 15989 24219 16047 24225
rect 16114 24216 16120 24228
rect 16172 24216 16178 24268
rect 16209 24259 16267 24265
rect 16209 24225 16221 24259
rect 16255 24256 16267 24259
rect 18049 24259 18107 24265
rect 16255 24228 17632 24256
rect 16255 24225 16267 24228
rect 16209 24219 16267 24225
rect 13538 24188 13544 24200
rect 12452 24160 13544 24188
rect 7653 24151 7711 24157
rect 13538 24148 13544 24160
rect 13596 24148 13602 24200
rect 13817 24191 13875 24197
rect 13817 24157 13829 24191
rect 13863 24188 13875 24191
rect 14182 24188 14188 24200
rect 13863 24160 14188 24188
rect 13863 24157 13875 24160
rect 13817 24151 13875 24157
rect 14182 24148 14188 24160
rect 14240 24188 14246 24200
rect 15286 24188 15292 24200
rect 14240 24160 15292 24188
rect 14240 24148 14246 24160
rect 15286 24148 15292 24160
rect 15344 24148 15350 24200
rect 15838 24148 15844 24200
rect 15896 24188 15902 24200
rect 16390 24188 16396 24200
rect 15896 24160 16396 24188
rect 15896 24148 15902 24160
rect 16390 24148 16396 24160
rect 16448 24148 16454 24200
rect 16666 24148 16672 24200
rect 16724 24188 16730 24200
rect 17034 24188 17040 24200
rect 16724 24160 17040 24188
rect 16724 24148 16730 24160
rect 17034 24148 17040 24160
rect 17092 24148 17098 24200
rect 4890 24080 4896 24132
rect 4948 24120 4954 24132
rect 11054 24120 11060 24132
rect 4948 24092 11060 24120
rect 4948 24080 4954 24092
rect 11054 24080 11060 24092
rect 11112 24080 11118 24132
rect 12710 24080 12716 24132
rect 12768 24120 12774 24132
rect 13354 24120 13360 24132
rect 12768 24092 13360 24120
rect 12768 24080 12774 24092
rect 13354 24080 13360 24092
rect 13412 24080 13418 24132
rect 4246 24052 4252 24064
rect 4207 24024 4252 24052
rect 4246 24012 4252 24024
rect 4304 24012 4310 24064
rect 4801 24055 4859 24061
rect 4801 24021 4813 24055
rect 4847 24052 4859 24055
rect 5994 24052 6000 24064
rect 4847 24024 6000 24052
rect 4847 24021 4859 24024
rect 4801 24015 4859 24021
rect 5994 24012 6000 24024
rect 6052 24012 6058 24064
rect 11698 24012 11704 24064
rect 11756 24052 11762 24064
rect 12069 24055 12127 24061
rect 12069 24052 12081 24055
rect 11756 24024 12081 24052
rect 11756 24012 11762 24024
rect 12069 24021 12081 24024
rect 12115 24021 12127 24055
rect 12069 24015 12127 24021
rect 12342 24012 12348 24064
rect 12400 24052 12406 24064
rect 13262 24052 13268 24064
rect 12400 24024 13268 24052
rect 12400 24012 12406 24024
rect 13262 24012 13268 24024
rect 13320 24012 13326 24064
rect 17604 24052 17632 24228
rect 18049 24225 18061 24259
rect 18095 24256 18107 24259
rect 19058 24256 19064 24268
rect 18095 24228 19064 24256
rect 18095 24225 18107 24228
rect 18049 24219 18107 24225
rect 19058 24216 19064 24228
rect 19116 24216 19122 24268
rect 21174 24216 21180 24268
rect 21232 24256 21238 24268
rect 21453 24259 21511 24265
rect 21453 24256 21465 24259
rect 21232 24228 21465 24256
rect 21232 24216 21238 24228
rect 21453 24225 21465 24228
rect 21499 24225 21511 24259
rect 21634 24256 21640 24268
rect 21595 24228 21640 24256
rect 21453 24219 21511 24225
rect 21634 24216 21640 24228
rect 21692 24216 21698 24268
rect 22554 24256 22560 24268
rect 22515 24228 22560 24256
rect 22554 24216 22560 24228
rect 22612 24216 22618 24268
rect 22646 24216 22652 24268
rect 22704 24256 22710 24268
rect 22741 24259 22799 24265
rect 22741 24256 22753 24259
rect 22704 24228 22753 24256
rect 22704 24216 22710 24228
rect 22741 24225 22753 24228
rect 22787 24225 22799 24259
rect 22741 24219 22799 24225
rect 18322 24188 18328 24200
rect 18283 24160 18328 24188
rect 18322 24148 18328 24160
rect 18380 24148 18386 24200
rect 21358 24148 21364 24200
rect 21416 24188 21422 24200
rect 21818 24188 21824 24200
rect 21416 24160 21824 24188
rect 21416 24148 21422 24160
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 21910 24148 21916 24200
rect 21968 24188 21974 24200
rect 24044 24188 24072 24296
rect 25961 24293 25973 24296
rect 26007 24293 26019 24327
rect 26142 24324 26148 24336
rect 26103 24296 26148 24324
rect 25961 24287 26019 24293
rect 26142 24284 26148 24296
rect 26200 24284 26206 24336
rect 26326 24284 26332 24336
rect 26384 24324 26390 24336
rect 28000 24333 28028 24364
rect 26697 24327 26755 24333
rect 26697 24324 26709 24327
rect 26384 24296 26709 24324
rect 26384 24284 26390 24296
rect 26697 24293 26709 24296
rect 26743 24293 26755 24327
rect 26697 24287 26755 24293
rect 27985 24327 28043 24333
rect 27985 24293 27997 24327
rect 28031 24293 28043 24327
rect 27985 24287 28043 24293
rect 24121 24259 24179 24265
rect 24121 24225 24133 24259
rect 24167 24225 24179 24259
rect 24121 24219 24179 24225
rect 21968 24160 24072 24188
rect 21968 24148 21974 24160
rect 21177 24123 21235 24129
rect 21177 24089 21189 24123
rect 21223 24120 21235 24123
rect 22094 24120 22100 24132
rect 21223 24092 22100 24120
rect 21223 24089 21235 24092
rect 21177 24083 21235 24089
rect 22094 24080 22100 24092
rect 22152 24080 22158 24132
rect 23566 24080 23572 24132
rect 23624 24120 23630 24132
rect 24136 24120 24164 24219
rect 24213 24191 24271 24197
rect 24213 24157 24225 24191
rect 24259 24157 24271 24191
rect 24486 24188 24492 24200
rect 24447 24160 24492 24188
rect 24213 24151 24271 24157
rect 23624 24092 24164 24120
rect 24228 24120 24256 24151
rect 24486 24148 24492 24160
rect 24544 24148 24550 24200
rect 24762 24120 24768 24132
rect 24228 24092 24768 24120
rect 23624 24080 23630 24092
rect 24762 24080 24768 24092
rect 24820 24080 24826 24132
rect 28166 24120 28172 24132
rect 28127 24092 28172 24120
rect 28166 24080 28172 24092
rect 28224 24080 28230 24132
rect 18230 24052 18236 24064
rect 17604 24024 18236 24052
rect 18230 24012 18236 24024
rect 18288 24012 18294 24064
rect 22646 24052 22652 24064
rect 22607 24024 22652 24052
rect 22646 24012 22652 24024
rect 22704 24012 22710 24064
rect 26786 24052 26792 24064
rect 26747 24024 26792 24052
rect 26786 24012 26792 24024
rect 26844 24012 26850 24064
rect 1104 23962 28888 23984
rect 1104 23910 5614 23962
rect 5666 23910 5678 23962
rect 5730 23910 5742 23962
rect 5794 23910 5806 23962
rect 5858 23910 14878 23962
rect 14930 23910 14942 23962
rect 14994 23910 15006 23962
rect 15058 23910 15070 23962
rect 15122 23910 24142 23962
rect 24194 23910 24206 23962
rect 24258 23910 24270 23962
rect 24322 23910 24334 23962
rect 24386 23910 28888 23962
rect 1104 23888 28888 23910
rect 2498 23848 2504 23860
rect 2459 23820 2504 23848
rect 2498 23808 2504 23820
rect 2556 23808 2562 23860
rect 3145 23851 3203 23857
rect 3145 23817 3157 23851
rect 3191 23848 3203 23851
rect 6086 23848 6092 23860
rect 3191 23820 6092 23848
rect 3191 23817 3203 23820
rect 3145 23811 3203 23817
rect 6086 23808 6092 23820
rect 6144 23808 6150 23860
rect 6638 23808 6644 23860
rect 6696 23848 6702 23860
rect 7101 23851 7159 23857
rect 7101 23848 7113 23851
rect 6696 23820 7113 23848
rect 6696 23808 6702 23820
rect 7101 23817 7113 23820
rect 7147 23817 7159 23851
rect 17773 23851 17831 23857
rect 7101 23811 7159 23817
rect 8036 23820 12434 23848
rect 4522 23740 4528 23792
rect 4580 23780 4586 23792
rect 4890 23780 4896 23792
rect 4580 23752 4896 23780
rect 4580 23740 4586 23752
rect 4890 23740 4896 23752
rect 4948 23740 4954 23792
rect 5902 23740 5908 23792
rect 5960 23780 5966 23792
rect 6457 23783 6515 23789
rect 5960 23752 6316 23780
rect 5960 23740 5966 23752
rect 1854 23672 1860 23724
rect 1912 23712 1918 23724
rect 1912 23684 6224 23712
rect 1912 23672 1918 23684
rect 2685 23647 2743 23653
rect 2685 23613 2697 23647
rect 2731 23644 2743 23647
rect 2774 23644 2780 23656
rect 2731 23616 2780 23644
rect 2731 23613 2743 23616
rect 2685 23607 2743 23613
rect 2774 23604 2780 23616
rect 2832 23604 2838 23656
rect 3326 23644 3332 23656
rect 3287 23616 3332 23644
rect 3326 23604 3332 23616
rect 3384 23604 3390 23656
rect 4249 23647 4307 23653
rect 4249 23613 4261 23647
rect 4295 23644 4307 23647
rect 4522 23644 4528 23656
rect 4295 23616 4528 23644
rect 4295 23613 4307 23616
rect 4249 23607 4307 23613
rect 4522 23604 4528 23616
rect 4580 23604 4586 23656
rect 1578 23536 1584 23588
rect 1636 23576 1642 23588
rect 1857 23579 1915 23585
rect 1857 23576 1869 23579
rect 1636 23548 1869 23576
rect 1636 23536 1642 23548
rect 1857 23545 1869 23548
rect 1903 23545 1915 23579
rect 1857 23539 1915 23545
rect 2041 23579 2099 23585
rect 2041 23545 2053 23579
rect 2087 23576 2099 23579
rect 2130 23576 2136 23588
rect 2087 23548 2136 23576
rect 2087 23545 2099 23548
rect 2041 23539 2099 23545
rect 2130 23536 2136 23548
rect 2188 23536 2194 23588
rect 6086 23576 6092 23588
rect 6047 23548 6092 23576
rect 6086 23536 6092 23548
rect 6144 23536 6150 23588
rect 4433 23511 4491 23517
rect 4433 23477 4445 23511
rect 4479 23508 4491 23511
rect 4798 23508 4804 23520
rect 4479 23480 4804 23508
rect 4479 23477 4491 23480
rect 4433 23471 4491 23477
rect 4798 23468 4804 23480
rect 4856 23468 4862 23520
rect 6196 23508 6224 23684
rect 6288 23576 6316 23752
rect 6457 23749 6469 23783
rect 6503 23780 6515 23783
rect 6730 23780 6736 23792
rect 6503 23752 6736 23780
rect 6503 23749 6515 23752
rect 6457 23743 6515 23749
rect 6730 23740 6736 23752
rect 6788 23780 6794 23792
rect 7929 23783 7987 23789
rect 7929 23780 7941 23783
rect 6788 23752 7941 23780
rect 6788 23740 6794 23752
rect 7929 23749 7941 23752
rect 7975 23749 7987 23783
rect 7929 23743 7987 23749
rect 6549 23715 6607 23721
rect 6549 23681 6561 23715
rect 6595 23712 6607 23715
rect 6595 23684 7052 23712
rect 6595 23681 6607 23684
rect 6549 23675 6607 23681
rect 7024 23653 7052 23684
rect 7009 23647 7067 23653
rect 7009 23613 7021 23647
rect 7055 23613 7067 23647
rect 7009 23607 7067 23613
rect 8036 23576 8064 23820
rect 12406 23780 12434 23820
rect 17773 23817 17785 23851
rect 17819 23848 17831 23851
rect 18322 23848 18328 23860
rect 17819 23820 18328 23848
rect 17819 23817 17831 23820
rect 17773 23811 17831 23817
rect 18322 23808 18328 23820
rect 18380 23808 18386 23860
rect 21266 23848 21272 23860
rect 21227 23820 21272 23848
rect 21266 23808 21272 23820
rect 21324 23808 21330 23860
rect 27982 23848 27988 23860
rect 27943 23820 27988 23848
rect 27982 23808 27988 23820
rect 28040 23808 28046 23860
rect 20714 23780 20720 23792
rect 12406 23752 20720 23780
rect 20714 23740 20720 23752
rect 20772 23740 20778 23792
rect 8389 23715 8447 23721
rect 8389 23681 8401 23715
rect 8435 23712 8447 23715
rect 8478 23712 8484 23724
rect 8435 23684 8484 23712
rect 8435 23681 8447 23684
rect 8389 23675 8447 23681
rect 8478 23672 8484 23684
rect 8536 23672 8542 23724
rect 11698 23712 11704 23724
rect 11659 23684 11704 23712
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 12066 23672 12072 23724
rect 12124 23712 12130 23724
rect 12805 23715 12863 23721
rect 12805 23712 12817 23715
rect 12124 23684 12817 23712
rect 12124 23672 12130 23684
rect 12805 23681 12817 23684
rect 12851 23681 12863 23715
rect 14182 23712 14188 23724
rect 12805 23675 12863 23681
rect 13280 23684 14188 23712
rect 11425 23647 11483 23653
rect 6288 23548 8064 23576
rect 8220 23616 11376 23644
rect 8220 23508 8248 23616
rect 8481 23579 8539 23585
rect 8481 23545 8493 23579
rect 8527 23576 8539 23579
rect 8570 23576 8576 23588
rect 8527 23548 8576 23576
rect 8527 23545 8539 23548
rect 8481 23539 8539 23545
rect 8570 23536 8576 23548
rect 8628 23576 8634 23588
rect 9122 23576 9128 23588
rect 8628 23548 9128 23576
rect 8628 23536 8634 23548
rect 9122 23536 9128 23548
rect 9180 23536 9186 23588
rect 8386 23508 8392 23520
rect 6196 23480 8248 23508
rect 8347 23480 8392 23508
rect 8386 23468 8392 23480
rect 8444 23468 8450 23520
rect 11348 23508 11376 23616
rect 11425 23613 11437 23647
rect 11471 23644 11483 23647
rect 13280 23644 13308 23684
rect 14182 23672 14188 23684
rect 14240 23672 14246 23724
rect 16022 23672 16028 23724
rect 16080 23712 16086 23724
rect 17313 23715 17371 23721
rect 16080 23684 17080 23712
rect 16080 23672 16086 23684
rect 11471 23616 13308 23644
rect 13633 23647 13691 23653
rect 11471 23613 11483 23616
rect 11425 23607 11483 23613
rect 13633 23613 13645 23647
rect 13679 23644 13691 23647
rect 14274 23644 14280 23656
rect 13679 23616 14280 23644
rect 13679 23613 13691 23616
rect 13633 23607 13691 23613
rect 14274 23604 14280 23616
rect 14332 23604 14338 23656
rect 14734 23604 14740 23656
rect 14792 23644 14798 23656
rect 15473 23647 15531 23653
rect 15473 23644 15485 23647
rect 14792 23616 15485 23644
rect 14792 23604 14798 23616
rect 15473 23613 15485 23616
rect 15519 23613 15531 23647
rect 15473 23607 15531 23613
rect 16574 23604 16580 23656
rect 16632 23644 16638 23656
rect 17052 23653 17080 23684
rect 17313 23681 17325 23715
rect 17359 23712 17371 23715
rect 21266 23712 21272 23724
rect 17359 23684 18460 23712
rect 17359 23681 17371 23684
rect 17313 23675 17371 23681
rect 16945 23647 17003 23653
rect 16945 23644 16957 23647
rect 16632 23616 16957 23644
rect 16632 23604 16638 23616
rect 16945 23613 16957 23616
rect 16991 23613 17003 23647
rect 16945 23607 17003 23613
rect 17037 23647 17095 23653
rect 17037 23613 17049 23647
rect 17083 23613 17095 23647
rect 17037 23607 17095 23613
rect 17129 23647 17187 23653
rect 17129 23613 17141 23647
rect 17175 23644 17187 23647
rect 17218 23644 17224 23656
rect 17175 23616 17224 23644
rect 17175 23613 17187 23616
rect 17129 23607 17187 23613
rect 17218 23604 17224 23616
rect 17276 23604 17282 23656
rect 18046 23644 18052 23656
rect 18007 23616 18052 23644
rect 18046 23604 18052 23616
rect 18104 23604 18110 23656
rect 18141 23647 18199 23653
rect 18141 23613 18153 23647
rect 18187 23613 18199 23647
rect 18141 23607 18199 23613
rect 18233 23647 18291 23653
rect 18233 23613 18245 23647
rect 18279 23644 18291 23647
rect 18322 23644 18328 23656
rect 18279 23616 18328 23644
rect 18279 23613 18291 23616
rect 18233 23607 18291 23613
rect 15657 23579 15715 23585
rect 15657 23545 15669 23579
rect 15703 23576 15715 23579
rect 16390 23576 16396 23588
rect 15703 23548 16396 23576
rect 15703 23545 15715 23548
rect 15657 23539 15715 23545
rect 16390 23536 16396 23548
rect 16448 23536 16454 23588
rect 16666 23536 16672 23588
rect 16724 23576 16730 23588
rect 18156 23576 18184 23607
rect 18322 23604 18328 23616
rect 18380 23604 18386 23656
rect 18432 23653 18460 23684
rect 20916 23684 21272 23712
rect 20916 23653 20944 23684
rect 21266 23672 21272 23684
rect 21324 23712 21330 23724
rect 21726 23712 21732 23724
rect 21324 23684 21732 23712
rect 21324 23672 21330 23684
rect 21726 23672 21732 23684
rect 21784 23672 21790 23724
rect 26237 23715 26295 23721
rect 26237 23681 26249 23715
rect 26283 23712 26295 23715
rect 26326 23712 26332 23724
rect 26283 23684 26332 23712
rect 26283 23681 26295 23684
rect 26237 23675 26295 23681
rect 26326 23672 26332 23684
rect 26384 23672 26390 23724
rect 27614 23712 27620 23724
rect 26712 23684 27620 23712
rect 18417 23647 18475 23653
rect 18417 23613 18429 23647
rect 18463 23613 18475 23647
rect 18417 23607 18475 23613
rect 20901 23647 20959 23653
rect 20901 23613 20913 23647
rect 20947 23613 20959 23647
rect 20901 23607 20959 23613
rect 20990 23604 20996 23656
rect 21048 23653 21054 23656
rect 21048 23647 21097 23653
rect 21048 23613 21051 23647
rect 21085 23613 21097 23647
rect 21174 23644 21180 23656
rect 21135 23616 21180 23644
rect 21048 23607 21097 23613
rect 21048 23604 21054 23607
rect 21174 23604 21180 23616
rect 21232 23604 21238 23656
rect 21361 23647 21419 23653
rect 21361 23613 21373 23647
rect 21407 23644 21419 23647
rect 22646 23644 22652 23656
rect 21407 23616 22652 23644
rect 21407 23613 21419 23616
rect 21361 23607 21419 23613
rect 22646 23604 22652 23616
rect 22704 23604 22710 23656
rect 26510 23604 26516 23656
rect 26568 23644 26574 23656
rect 26712 23653 26740 23684
rect 27614 23672 27620 23684
rect 27672 23672 27678 23724
rect 26697 23647 26755 23653
rect 26697 23644 26709 23647
rect 26568 23616 26709 23644
rect 26568 23604 26574 23616
rect 26697 23613 26709 23616
rect 26743 23613 26755 23647
rect 26878 23644 26884 23656
rect 26839 23616 26884 23644
rect 26697 23607 26755 23613
rect 26878 23604 26884 23616
rect 26936 23604 26942 23656
rect 27154 23604 27160 23656
rect 27212 23644 27218 23656
rect 27341 23647 27399 23653
rect 27341 23644 27353 23647
rect 27212 23616 27353 23644
rect 27212 23604 27218 23616
rect 27341 23613 27353 23616
rect 27387 23613 27399 23647
rect 27341 23607 27399 23613
rect 16724 23548 18184 23576
rect 18340 23576 18368 23604
rect 20070 23576 20076 23588
rect 18340 23548 20076 23576
rect 16724 23536 16730 23548
rect 20070 23536 20076 23548
rect 20128 23536 20134 23588
rect 26053 23579 26111 23585
rect 26053 23545 26065 23579
rect 26099 23576 26111 23579
rect 26234 23576 26240 23588
rect 26099 23548 26240 23576
rect 26099 23545 26111 23548
rect 26053 23539 26111 23545
rect 26234 23536 26240 23548
rect 26292 23536 26298 23588
rect 12066 23508 12072 23520
rect 11348 23480 12072 23508
rect 12066 23468 12072 23480
rect 12124 23468 12130 23520
rect 13354 23468 13360 23520
rect 13412 23508 13418 23520
rect 13538 23508 13544 23520
rect 13412 23480 13544 23508
rect 13412 23468 13418 23480
rect 13538 23468 13544 23480
rect 13596 23508 13602 23520
rect 13725 23511 13783 23517
rect 13725 23508 13737 23511
rect 13596 23480 13737 23508
rect 13596 23468 13602 23480
rect 13725 23477 13737 23480
rect 13771 23477 13783 23511
rect 13725 23471 13783 23477
rect 16942 23468 16948 23520
rect 17000 23508 17006 23520
rect 17218 23508 17224 23520
rect 17000 23480 17224 23508
rect 17000 23468 17006 23480
rect 17218 23468 17224 23480
rect 17276 23468 17282 23520
rect 18046 23468 18052 23520
rect 18104 23508 18110 23520
rect 19978 23508 19984 23520
rect 18104 23480 19984 23508
rect 18104 23468 18110 23480
rect 19978 23468 19984 23480
rect 20036 23468 20042 23520
rect 1104 23418 28888 23440
rect 1104 23366 10246 23418
rect 10298 23366 10310 23418
rect 10362 23366 10374 23418
rect 10426 23366 10438 23418
rect 10490 23366 19510 23418
rect 19562 23366 19574 23418
rect 19626 23366 19638 23418
rect 19690 23366 19702 23418
rect 19754 23366 28888 23418
rect 1104 23344 28888 23366
rect 2501 23307 2559 23313
rect 2501 23273 2513 23307
rect 2547 23304 2559 23307
rect 2682 23304 2688 23316
rect 2547 23276 2688 23304
rect 2547 23273 2559 23276
rect 2501 23267 2559 23273
rect 2682 23264 2688 23276
rect 2740 23264 2746 23316
rect 3142 23264 3148 23316
rect 3200 23304 3206 23316
rect 3237 23307 3295 23313
rect 3237 23304 3249 23307
rect 3200 23276 3249 23304
rect 3200 23264 3206 23276
rect 3237 23273 3249 23276
rect 3283 23273 3295 23307
rect 3237 23267 3295 23273
rect 3605 23307 3663 23313
rect 3605 23273 3617 23307
rect 3651 23304 3663 23307
rect 4246 23304 4252 23316
rect 3651 23276 4252 23304
rect 3651 23273 3663 23276
rect 3605 23267 3663 23273
rect 4246 23264 4252 23276
rect 4304 23264 4310 23316
rect 4706 23264 4712 23316
rect 4764 23304 4770 23316
rect 4801 23307 4859 23313
rect 4801 23304 4813 23307
rect 4764 23276 4813 23304
rect 4764 23264 4770 23276
rect 4801 23273 4813 23276
rect 4847 23273 4859 23307
rect 4801 23267 4859 23273
rect 6822 23264 6828 23316
rect 6880 23304 6886 23316
rect 7285 23307 7343 23313
rect 7285 23304 7297 23307
rect 6880 23276 7297 23304
rect 6880 23264 6886 23276
rect 7285 23273 7297 23276
rect 7331 23273 7343 23307
rect 7285 23267 7343 23273
rect 8386 23264 8392 23316
rect 8444 23304 8450 23316
rect 9677 23307 9735 23313
rect 9677 23304 9689 23307
rect 8444 23276 9689 23304
rect 8444 23264 8450 23276
rect 9677 23273 9689 23276
rect 9723 23273 9735 23307
rect 9677 23267 9735 23273
rect 12250 23264 12256 23316
rect 12308 23304 12314 23316
rect 13633 23307 13691 23313
rect 13633 23304 13645 23307
rect 12308 23276 13645 23304
rect 12308 23264 12314 23276
rect 13633 23273 13645 23276
rect 13679 23273 13691 23307
rect 13633 23267 13691 23273
rect 14090 23264 14096 23316
rect 14148 23304 14154 23316
rect 14369 23307 14427 23313
rect 14369 23304 14381 23307
rect 14148 23276 14381 23304
rect 14148 23264 14154 23276
rect 14369 23273 14381 23276
rect 14415 23273 14427 23307
rect 17218 23304 17224 23316
rect 14369 23267 14427 23273
rect 14476 23276 17224 23304
rect 1762 23196 1768 23248
rect 1820 23236 1826 23248
rect 2041 23239 2099 23245
rect 2041 23236 2053 23239
rect 1820 23208 2053 23236
rect 1820 23196 1826 23208
rect 2041 23205 2053 23208
rect 2087 23236 2099 23239
rect 14476 23236 14504 23276
rect 17218 23264 17224 23276
rect 17276 23264 17282 23316
rect 28074 23304 28080 23316
rect 24964 23276 28080 23304
rect 2087 23208 14504 23236
rect 2087 23205 2099 23208
rect 2041 23199 2099 23205
rect 1394 23128 1400 23180
rect 1452 23168 1458 23180
rect 1857 23171 1915 23177
rect 1857 23168 1869 23171
rect 1452 23140 1869 23168
rect 1452 23128 1458 23140
rect 1857 23137 1869 23140
rect 1903 23137 1915 23171
rect 1857 23131 1915 23137
rect 2685 23171 2743 23177
rect 2685 23137 2697 23171
rect 2731 23168 2743 23171
rect 2774 23168 2780 23180
rect 2731 23140 2780 23168
rect 2731 23137 2743 23140
rect 2685 23131 2743 23137
rect 2774 23128 2780 23140
rect 2832 23128 2838 23180
rect 3697 23171 3755 23177
rect 3697 23137 3709 23171
rect 3743 23168 3755 23171
rect 4154 23168 4160 23180
rect 3743 23140 4160 23168
rect 3743 23137 3755 23140
rect 3697 23131 3755 23137
rect 4154 23128 4160 23140
rect 4212 23128 4218 23180
rect 4724 23177 4752 23208
rect 14550 23196 14556 23248
rect 14608 23236 14614 23248
rect 14608 23208 15700 23236
rect 14608 23196 14614 23208
rect 4709 23171 4767 23177
rect 4709 23137 4721 23171
rect 4755 23137 4767 23171
rect 4709 23131 4767 23137
rect 6730 23128 6736 23180
rect 6788 23168 6794 23180
rect 8110 23177 8116 23180
rect 6825 23171 6883 23177
rect 6825 23168 6837 23171
rect 6788 23140 6837 23168
rect 6788 23128 6794 23140
rect 6825 23137 6837 23140
rect 6871 23137 6883 23171
rect 6825 23131 6883 23137
rect 8104 23131 8116 23177
rect 8168 23168 8174 23180
rect 8168 23140 8204 23168
rect 8110 23128 8116 23131
rect 8168 23128 8174 23140
rect 9582 23128 9588 23180
rect 9640 23168 9646 23180
rect 10045 23171 10103 23177
rect 10045 23168 10057 23171
rect 9640 23140 10057 23168
rect 9640 23128 9646 23140
rect 10045 23137 10057 23140
rect 10091 23137 10103 23171
rect 10045 23131 10103 23137
rect 10137 23171 10195 23177
rect 10137 23137 10149 23171
rect 10183 23168 10195 23171
rect 10594 23168 10600 23180
rect 10183 23140 10600 23168
rect 10183 23137 10195 23140
rect 10137 23131 10195 23137
rect 10594 23128 10600 23140
rect 10652 23128 10658 23180
rect 10870 23168 10876 23180
rect 10831 23140 10876 23168
rect 10870 23128 10876 23140
rect 10928 23168 10934 23180
rect 10928 23140 12434 23168
rect 10928 23128 10934 23140
rect 3881 23103 3939 23109
rect 3881 23069 3893 23103
rect 3927 23100 3939 23103
rect 4338 23100 4344 23112
rect 3927 23072 4344 23100
rect 3927 23069 3939 23072
rect 3881 23063 3939 23069
rect 4338 23060 4344 23072
rect 4396 23060 4402 23112
rect 7837 23103 7895 23109
rect 7837 23069 7849 23103
rect 7883 23069 7895 23103
rect 7837 23063 7895 23069
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23069 10287 23103
rect 12406 23100 12434 23140
rect 12618 23128 12624 23180
rect 12676 23168 12682 23180
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 12676 23140 13553 23168
rect 12676 23128 12682 23140
rect 13541 23137 13553 23140
rect 13587 23137 13599 23171
rect 13541 23131 13599 23137
rect 14277 23171 14335 23177
rect 14277 23137 14289 23171
rect 14323 23168 14335 23171
rect 14734 23168 14740 23180
rect 14323 23140 14740 23168
rect 14323 23137 14335 23140
rect 14277 23131 14335 23137
rect 14734 23128 14740 23140
rect 14792 23168 14798 23180
rect 15672 23177 15700 23208
rect 16390 23196 16396 23248
rect 16448 23236 16454 23248
rect 17681 23239 17739 23245
rect 17681 23236 17693 23239
rect 16448 23208 17693 23236
rect 16448 23196 16454 23208
rect 17681 23205 17693 23208
rect 17727 23205 17739 23239
rect 17681 23199 17739 23205
rect 17865 23239 17923 23245
rect 17865 23205 17877 23239
rect 17911 23236 17923 23239
rect 18322 23236 18328 23248
rect 17911 23208 18328 23236
rect 17911 23205 17923 23208
rect 17865 23199 17923 23205
rect 18322 23196 18328 23208
rect 18380 23196 18386 23248
rect 24964 23245 24992 23276
rect 28074 23264 28080 23276
rect 28132 23264 28138 23316
rect 24949 23239 25007 23245
rect 24949 23205 24961 23239
rect 24995 23205 25007 23239
rect 27985 23239 28043 23245
rect 27985 23236 27997 23239
rect 24949 23199 25007 23205
rect 25148 23208 27997 23236
rect 15013 23171 15071 23177
rect 15013 23168 15025 23171
rect 14792 23140 15025 23168
rect 14792 23128 14798 23140
rect 15013 23137 15025 23140
rect 15059 23137 15071 23171
rect 15013 23131 15071 23137
rect 15657 23171 15715 23177
rect 15657 23137 15669 23171
rect 15703 23137 15715 23171
rect 15657 23131 15715 23137
rect 17034 23128 17040 23180
rect 17092 23168 17098 23180
rect 17310 23168 17316 23180
rect 17092 23140 17316 23168
rect 17092 23128 17098 23140
rect 17310 23128 17316 23140
rect 17368 23128 17374 23180
rect 17402 23128 17408 23180
rect 17460 23168 17466 23180
rect 25148 23168 25176 23208
rect 27985 23205 27997 23208
rect 28031 23205 28043 23239
rect 27985 23199 28043 23205
rect 17460 23140 25176 23168
rect 17460 23128 17466 23140
rect 25590 23128 25596 23180
rect 25648 23168 25654 23180
rect 25685 23171 25743 23177
rect 25685 23168 25697 23171
rect 25648 23140 25697 23168
rect 25648 23128 25654 23140
rect 25685 23137 25697 23140
rect 25731 23137 25743 23171
rect 26510 23168 26516 23180
rect 26471 23140 26516 23168
rect 25685 23131 25743 23137
rect 26510 23128 26516 23140
rect 26568 23128 26574 23180
rect 26418 23100 26424 23112
rect 12406 23072 26424 23100
rect 10229 23063 10287 23069
rect 6086 22992 6092 23044
rect 6144 23032 6150 23044
rect 6638 23032 6644 23044
rect 6144 23004 6644 23032
rect 6144 22992 6150 23004
rect 6638 22992 6644 23004
rect 6696 23032 6702 23044
rect 7101 23035 7159 23041
rect 7101 23032 7113 23035
rect 6696 23004 7113 23032
rect 6696 22992 6702 23004
rect 7101 23001 7113 23004
rect 7147 23001 7159 23035
rect 7101 22995 7159 23001
rect 2866 22924 2872 22976
rect 2924 22964 2930 22976
rect 7852 22964 7880 23063
rect 8938 23032 8944 23044
rect 8772 23004 8944 23032
rect 8772 22964 8800 23004
rect 8938 22992 8944 23004
rect 8996 23032 9002 23044
rect 9490 23032 9496 23044
rect 8996 23004 9496 23032
rect 8996 22992 9002 23004
rect 9490 22992 9496 23004
rect 9548 22992 9554 23044
rect 9766 22992 9772 23044
rect 9824 23032 9830 23044
rect 10244 23032 10272 23063
rect 26418 23060 26424 23072
rect 26476 23060 26482 23112
rect 26605 23103 26663 23109
rect 26605 23069 26617 23103
rect 26651 23100 26663 23103
rect 26694 23100 26700 23112
rect 26651 23072 26700 23100
rect 26651 23069 26663 23072
rect 26605 23063 26663 23069
rect 26694 23060 26700 23072
rect 26752 23100 26758 23112
rect 27246 23100 27252 23112
rect 26752 23072 27252 23100
rect 26752 23060 26758 23072
rect 27246 23060 27252 23072
rect 27304 23060 27310 23112
rect 9824 23004 10272 23032
rect 15197 23035 15255 23041
rect 9824 22992 9830 23004
rect 10152 22976 10180 23004
rect 15197 23001 15209 23035
rect 15243 23032 15255 23035
rect 15470 23032 15476 23044
rect 15243 23004 15476 23032
rect 15243 23001 15255 23004
rect 15197 22995 15255 23001
rect 15470 22992 15476 23004
rect 15528 22992 15534 23044
rect 15562 22992 15568 23044
rect 15620 23032 15626 23044
rect 15841 23035 15899 23041
rect 15841 23032 15853 23035
rect 15620 23004 15853 23032
rect 15620 22992 15626 23004
rect 15841 23001 15853 23004
rect 15887 23032 15899 23035
rect 16574 23032 16580 23044
rect 15887 23004 16580 23032
rect 15887 23001 15899 23004
rect 15841 22995 15899 23001
rect 16574 22992 16580 23004
rect 16632 22992 16638 23044
rect 25130 23032 25136 23044
rect 25091 23004 25136 23032
rect 25130 22992 25136 23004
rect 25188 22992 25194 23044
rect 25866 23032 25872 23044
rect 25827 23004 25872 23032
rect 25866 22992 25872 23004
rect 25924 22992 25930 23044
rect 28166 23032 28172 23044
rect 28127 23004 28172 23032
rect 28166 22992 28172 23004
rect 28224 22992 28230 23044
rect 9214 22964 9220 22976
rect 2924 22936 8800 22964
rect 9175 22936 9220 22964
rect 2924 22924 2930 22936
rect 9214 22924 9220 22936
rect 9272 22924 9278 22976
rect 10134 22924 10140 22976
rect 10192 22924 10198 22976
rect 10965 22967 11023 22973
rect 10965 22933 10977 22967
rect 11011 22964 11023 22967
rect 12526 22964 12532 22976
rect 11011 22936 12532 22964
rect 11011 22933 11023 22936
rect 10965 22927 11023 22933
rect 12526 22924 12532 22936
rect 12584 22924 12590 22976
rect 26881 22967 26939 22973
rect 26881 22933 26893 22967
rect 26927 22964 26939 22967
rect 27798 22964 27804 22976
rect 26927 22936 27804 22964
rect 26927 22933 26939 22936
rect 26881 22927 26939 22933
rect 27798 22924 27804 22936
rect 27856 22924 27862 22976
rect 1104 22874 28888 22896
rect 1104 22822 5614 22874
rect 5666 22822 5678 22874
rect 5730 22822 5742 22874
rect 5794 22822 5806 22874
rect 5858 22822 14878 22874
rect 14930 22822 14942 22874
rect 14994 22822 15006 22874
rect 15058 22822 15070 22874
rect 15122 22822 24142 22874
rect 24194 22822 24206 22874
rect 24258 22822 24270 22874
rect 24322 22822 24334 22874
rect 24386 22822 28888 22874
rect 1104 22800 28888 22822
rect 2038 22720 2044 22772
rect 2096 22760 2102 22772
rect 2590 22760 2596 22772
rect 2096 22732 2596 22760
rect 2096 22720 2102 22732
rect 2590 22720 2596 22732
rect 2648 22720 2654 22772
rect 8478 22760 8484 22772
rect 8439 22732 8484 22760
rect 8478 22720 8484 22732
rect 8536 22720 8542 22772
rect 9582 22760 9588 22772
rect 9543 22732 9588 22760
rect 9582 22720 9588 22732
rect 9640 22720 9646 22772
rect 23106 22760 23112 22772
rect 11624 22732 23112 22760
rect 4062 22652 4068 22704
rect 4120 22692 4126 22704
rect 10870 22692 10876 22704
rect 4120 22664 10876 22692
rect 4120 22652 4126 22664
rect 10870 22652 10876 22664
rect 10928 22652 10934 22704
rect 5534 22584 5540 22636
rect 5592 22624 5598 22636
rect 6270 22624 6276 22636
rect 5592 22596 6276 22624
rect 5592 22584 5598 22596
rect 6270 22584 6276 22596
rect 6328 22584 6334 22636
rect 6454 22584 6460 22636
rect 6512 22624 6518 22636
rect 6730 22624 6736 22636
rect 6512 22596 6736 22624
rect 6512 22584 6518 22596
rect 6730 22584 6736 22596
rect 6788 22584 6794 22636
rect 8662 22624 8668 22636
rect 8404 22596 8668 22624
rect 8404 22568 8432 22596
rect 8662 22584 8668 22596
rect 8720 22584 8726 22636
rect 10594 22584 10600 22636
rect 10652 22624 10658 22636
rect 11624 22633 11652 22732
rect 23106 22720 23112 22732
rect 23164 22720 23170 22772
rect 24486 22720 24492 22772
rect 24544 22760 24550 22772
rect 24762 22760 24768 22772
rect 24544 22732 24768 22760
rect 24544 22720 24550 22732
rect 24762 22720 24768 22732
rect 24820 22760 24826 22772
rect 25501 22763 25559 22769
rect 25501 22760 25513 22763
rect 24820 22732 25513 22760
rect 24820 22720 24826 22732
rect 25501 22729 25513 22732
rect 25547 22729 25559 22763
rect 25501 22723 25559 22729
rect 25958 22720 25964 22772
rect 26016 22760 26022 22772
rect 26016 22732 26464 22760
rect 26016 22720 26022 22732
rect 16022 22692 16028 22704
rect 15672 22664 16028 22692
rect 11609 22627 11667 22633
rect 10652 22596 11284 22624
rect 10652 22584 10658 22596
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 2866 22556 2872 22568
rect 1443 22528 2872 22556
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 4246 22556 4252 22568
rect 4207 22528 4252 22556
rect 4246 22516 4252 22528
rect 4304 22516 4310 22568
rect 6638 22556 6644 22568
rect 6599 22528 6644 22556
rect 6638 22516 6644 22528
rect 6696 22516 6702 22568
rect 8386 22556 8392 22568
rect 8299 22528 8392 22556
rect 8386 22516 8392 22528
rect 8444 22516 8450 22568
rect 8570 22556 8576 22568
rect 8531 22528 8576 22556
rect 8570 22516 8576 22528
rect 8628 22516 8634 22568
rect 9493 22559 9551 22565
rect 9493 22525 9505 22559
rect 9539 22525 9551 22559
rect 10870 22556 10876 22568
rect 10831 22528 10876 22556
rect 9493 22519 9551 22525
rect 1664 22491 1722 22497
rect 1664 22457 1676 22491
rect 1710 22488 1722 22491
rect 2038 22488 2044 22500
rect 1710 22460 2044 22488
rect 1710 22457 1722 22460
rect 1664 22451 1722 22457
rect 2038 22448 2044 22460
rect 2096 22448 2102 22500
rect 8478 22448 8484 22500
rect 8536 22488 8542 22500
rect 9214 22488 9220 22500
rect 8536 22460 9220 22488
rect 8536 22448 8542 22460
rect 9214 22448 9220 22460
rect 9272 22488 9278 22500
rect 9508 22488 9536 22519
rect 10870 22516 10876 22528
rect 10928 22516 10934 22568
rect 10965 22559 11023 22565
rect 10965 22525 10977 22559
rect 11011 22525 11023 22559
rect 11146 22556 11152 22568
rect 11107 22528 11152 22556
rect 10965 22519 11023 22525
rect 9272 22460 9536 22488
rect 9272 22448 9278 22460
rect 2774 22380 2780 22432
rect 2832 22420 2838 22432
rect 4338 22420 4344 22432
rect 2832 22392 2877 22420
rect 4299 22392 4344 22420
rect 2832 22380 2838 22392
rect 4338 22380 4344 22392
rect 4396 22380 4402 22432
rect 7466 22420 7472 22432
rect 7427 22392 7472 22420
rect 7466 22380 7472 22392
rect 7524 22380 7530 22432
rect 10980 22420 11008 22519
rect 11146 22516 11152 22528
rect 11204 22516 11210 22568
rect 11256 22556 11284 22596
rect 11609 22593 11621 22627
rect 11655 22593 11667 22627
rect 12526 22624 12532 22636
rect 12487 22596 12532 22624
rect 11609 22587 11667 22593
rect 12526 22584 12532 22596
rect 12584 22584 12590 22636
rect 12713 22627 12771 22633
rect 12713 22593 12725 22627
rect 12759 22624 12771 22627
rect 13814 22624 13820 22636
rect 12759 22596 13820 22624
rect 12759 22593 12771 22596
rect 12713 22587 12771 22593
rect 12437 22559 12495 22565
rect 12437 22556 12449 22559
rect 11256 22528 12449 22556
rect 12437 22525 12449 22528
rect 12483 22525 12495 22559
rect 12437 22519 12495 22525
rect 11514 22448 11520 22500
rect 11572 22488 11578 22500
rect 12728 22488 12756 22587
rect 13814 22584 13820 22596
rect 13872 22584 13878 22636
rect 15562 22556 15568 22568
rect 15523 22528 15568 22556
rect 15562 22516 15568 22528
rect 15620 22516 15626 22568
rect 15672 22565 15700 22664
rect 16022 22652 16028 22664
rect 16080 22652 16086 22704
rect 17678 22652 17684 22704
rect 17736 22692 17742 22704
rect 17773 22695 17831 22701
rect 17773 22692 17785 22695
rect 17736 22664 17785 22692
rect 17736 22652 17742 22664
rect 17773 22661 17785 22664
rect 17819 22661 17831 22695
rect 17773 22655 17831 22661
rect 18046 22652 18052 22704
rect 18104 22692 18110 22704
rect 19058 22692 19064 22704
rect 18104 22664 19064 22692
rect 18104 22652 18110 22664
rect 19058 22652 19064 22664
rect 19116 22692 19122 22704
rect 20165 22695 20223 22701
rect 20165 22692 20177 22695
rect 19116 22664 20177 22692
rect 19116 22652 19122 22664
rect 20165 22661 20177 22664
rect 20211 22661 20223 22695
rect 20165 22655 20223 22661
rect 22186 22652 22192 22704
rect 22244 22692 22250 22704
rect 22738 22692 22744 22704
rect 22244 22664 22744 22692
rect 22244 22652 22250 22664
rect 22738 22652 22744 22664
rect 22796 22652 22802 22704
rect 23842 22652 23848 22704
rect 23900 22692 23906 22704
rect 24213 22695 24271 22701
rect 23900 22664 24164 22692
rect 23900 22652 23906 22664
rect 17310 22624 17316 22636
rect 15764 22596 17316 22624
rect 15764 22565 15792 22596
rect 17310 22584 17316 22596
rect 17368 22584 17374 22636
rect 22922 22584 22928 22636
rect 22980 22624 22986 22636
rect 24029 22627 24087 22633
rect 24029 22624 24041 22627
rect 22980 22596 24041 22624
rect 22980 22584 22986 22596
rect 24029 22593 24041 22596
rect 24075 22593 24087 22627
rect 24029 22587 24087 22593
rect 15657 22559 15715 22565
rect 15657 22525 15669 22559
rect 15703 22525 15715 22559
rect 15657 22519 15715 22525
rect 15749 22559 15807 22565
rect 15749 22525 15761 22559
rect 15795 22525 15807 22559
rect 15749 22519 15807 22525
rect 16393 22559 16451 22565
rect 16393 22525 16405 22559
rect 16439 22556 16451 22559
rect 16666 22556 16672 22568
rect 16439 22528 16528 22556
rect 16627 22528 16672 22556
rect 16439 22525 16451 22528
rect 16393 22519 16451 22525
rect 11572 22460 12756 22488
rect 11572 22448 11578 22460
rect 14734 22448 14740 22500
rect 14792 22488 14798 22500
rect 15672 22488 15700 22519
rect 14792 22460 15700 22488
rect 14792 22448 14798 22460
rect 12069 22423 12127 22429
rect 12069 22420 12081 22423
rect 10980 22392 12081 22420
rect 12069 22389 12081 22392
rect 12115 22389 12127 22423
rect 12069 22383 12127 22389
rect 15933 22423 15991 22429
rect 15933 22389 15945 22423
rect 15979 22420 15991 22423
rect 16298 22420 16304 22432
rect 15979 22392 16304 22420
rect 15979 22389 15991 22392
rect 15933 22383 15991 22389
rect 16298 22380 16304 22392
rect 16356 22380 16362 22432
rect 16500 22420 16528 22528
rect 16666 22516 16672 22528
rect 16724 22516 16730 22568
rect 20349 22559 20407 22565
rect 20349 22525 20361 22559
rect 20395 22556 20407 22559
rect 20438 22556 20444 22568
rect 20395 22528 20444 22556
rect 20395 22525 20407 22528
rect 20349 22519 20407 22525
rect 20438 22516 20444 22528
rect 20496 22516 20502 22568
rect 21634 22556 21640 22568
rect 21595 22528 21640 22556
rect 21634 22516 21640 22528
rect 21692 22516 21698 22568
rect 23842 22556 23848 22568
rect 23803 22528 23848 22556
rect 23842 22516 23848 22528
rect 23900 22516 23906 22568
rect 23934 22516 23940 22568
rect 23992 22516 23998 22568
rect 24136 22556 24164 22664
rect 24213 22661 24225 22695
rect 24259 22692 24271 22695
rect 25363 22695 25421 22701
rect 25363 22692 25375 22695
rect 24259 22664 25375 22692
rect 24259 22661 24271 22664
rect 24213 22655 24271 22661
rect 25363 22661 25375 22664
rect 25409 22661 25421 22695
rect 25363 22655 25421 22661
rect 26068 22664 26372 22692
rect 25958 22624 25964 22636
rect 25240 22596 25964 22624
rect 24210 22556 24216 22568
rect 24123 22528 24216 22556
rect 24210 22516 24216 22528
rect 24268 22516 24274 22568
rect 24946 22516 24952 22568
rect 25004 22556 25010 22568
rect 25240 22565 25268 22596
rect 25958 22584 25964 22596
rect 26016 22624 26022 22636
rect 26068 22624 26096 22664
rect 26234 22624 26240 22636
rect 26016 22596 26096 22624
rect 26160 22596 26240 22624
rect 26016 22584 26022 22596
rect 25225 22559 25283 22565
rect 25225 22556 25237 22559
rect 25004 22528 25237 22556
rect 25004 22516 25010 22528
rect 25225 22525 25237 22528
rect 25271 22525 25283 22559
rect 25498 22556 25504 22568
rect 25225 22519 25283 22525
rect 25424 22528 25504 22556
rect 21358 22488 21364 22500
rect 21319 22460 21364 22488
rect 21358 22448 21364 22460
rect 21416 22448 21422 22500
rect 21450 22448 21456 22500
rect 21508 22488 21514 22500
rect 21545 22491 21603 22497
rect 21545 22488 21557 22491
rect 21508 22460 21557 22488
rect 21508 22448 21514 22460
rect 21545 22457 21557 22460
rect 21591 22457 21603 22491
rect 21545 22451 21603 22457
rect 21913 22491 21971 22497
rect 21913 22457 21925 22491
rect 21959 22488 21971 22491
rect 22557 22491 22615 22497
rect 22557 22488 22569 22491
rect 21959 22460 22569 22488
rect 21959 22457 21971 22460
rect 21913 22451 21971 22457
rect 22557 22457 22569 22460
rect 22603 22457 22615 22491
rect 23952 22488 23980 22516
rect 24670 22488 24676 22500
rect 23952 22460 24676 22488
rect 22557 22451 22615 22457
rect 24670 22448 24676 22460
rect 24728 22448 24734 22500
rect 25424 22488 25452 22528
rect 25498 22516 25504 22528
rect 25556 22516 25562 22568
rect 26160 22565 26188 22596
rect 26234 22584 26240 22596
rect 26292 22584 26298 22636
rect 26344 22565 26372 22664
rect 26436 22624 26464 22732
rect 28074 22720 28080 22772
rect 28132 22760 28138 22772
rect 28169 22763 28227 22769
rect 28169 22760 28181 22763
rect 28132 22732 28181 22760
rect 28132 22720 28138 22732
rect 28169 22729 28181 22732
rect 28215 22729 28227 22763
rect 28169 22723 28227 22729
rect 26789 22627 26847 22633
rect 26789 22624 26801 22627
rect 26436 22596 26801 22624
rect 26789 22593 26801 22596
rect 26835 22593 26847 22627
rect 26789 22587 26847 22593
rect 25685 22559 25743 22565
rect 25685 22525 25697 22559
rect 25731 22525 25743 22559
rect 25685 22519 25743 22525
rect 26145 22559 26203 22565
rect 26145 22525 26157 22559
rect 26191 22525 26203 22559
rect 26145 22519 26203 22525
rect 26329 22559 26387 22565
rect 26329 22525 26341 22559
rect 26375 22525 26387 22559
rect 26329 22519 26387 22525
rect 24964 22460 25452 22488
rect 25700 22488 25728 22519
rect 26237 22491 26295 22497
rect 26237 22488 26249 22491
rect 25700 22460 26249 22488
rect 18046 22420 18052 22432
rect 16500 22392 18052 22420
rect 18046 22380 18052 22392
rect 18104 22380 18110 22432
rect 20714 22380 20720 22432
rect 20772 22420 20778 22432
rect 21468 22420 21496 22448
rect 24964 22432 24992 22460
rect 26237 22457 26249 22460
rect 26283 22457 26295 22491
rect 26237 22451 26295 22457
rect 27056 22491 27114 22497
rect 27056 22457 27068 22491
rect 27102 22488 27114 22491
rect 27430 22488 27436 22500
rect 27102 22460 27436 22488
rect 27102 22457 27114 22460
rect 27056 22451 27114 22457
rect 27430 22448 27436 22460
rect 27488 22448 27494 22500
rect 21726 22420 21732 22432
rect 20772 22392 21496 22420
rect 21687 22392 21732 22420
rect 20772 22380 20778 22392
rect 21726 22380 21732 22392
rect 21784 22380 21790 22432
rect 23934 22420 23940 22432
rect 23895 22392 23940 22420
rect 23934 22380 23940 22392
rect 23992 22380 23998 22432
rect 24946 22380 24952 22432
rect 25004 22380 25010 22432
rect 25498 22380 25504 22432
rect 25556 22420 25562 22432
rect 25593 22423 25651 22429
rect 25593 22420 25605 22423
rect 25556 22392 25605 22420
rect 25556 22380 25562 22392
rect 25593 22389 25605 22392
rect 25639 22389 25651 22423
rect 25593 22383 25651 22389
rect 1104 22330 28888 22352
rect 1104 22278 10246 22330
rect 10298 22278 10310 22330
rect 10362 22278 10374 22330
rect 10426 22278 10438 22330
rect 10490 22278 19510 22330
rect 19562 22278 19574 22330
rect 19626 22278 19638 22330
rect 19690 22278 19702 22330
rect 19754 22278 28888 22330
rect 1104 22256 28888 22278
rect 2038 22216 2044 22228
rect 1999 22188 2044 22216
rect 2038 22176 2044 22188
rect 2096 22176 2102 22228
rect 2409 22219 2467 22225
rect 2409 22185 2421 22219
rect 2455 22216 2467 22219
rect 2774 22216 2780 22228
rect 2455 22188 2780 22216
rect 2455 22185 2467 22188
rect 2409 22179 2467 22185
rect 2774 22176 2780 22188
rect 2832 22176 2838 22228
rect 5074 22216 5080 22228
rect 4816 22188 5080 22216
rect 2130 22108 2136 22160
rect 2188 22148 2194 22160
rect 4062 22148 4068 22160
rect 2188 22120 4068 22148
rect 2188 22108 2194 22120
rect 4062 22108 4068 22120
rect 4120 22148 4126 22160
rect 4433 22151 4491 22157
rect 4433 22148 4445 22151
rect 4120 22120 4445 22148
rect 4120 22108 4126 22120
rect 4433 22117 4445 22120
rect 4479 22117 4491 22151
rect 4706 22148 4712 22160
rect 4667 22120 4712 22148
rect 4433 22111 4491 22117
rect 4706 22108 4712 22120
rect 4764 22108 4770 22160
rect 4816 22157 4844 22188
rect 5074 22176 5080 22188
rect 5132 22216 5138 22228
rect 5626 22216 5632 22228
rect 5132 22188 5632 22216
rect 5132 22176 5138 22188
rect 5626 22176 5632 22188
rect 5684 22176 5690 22228
rect 5721 22219 5779 22225
rect 5721 22185 5733 22219
rect 5767 22216 5779 22219
rect 8110 22216 8116 22228
rect 5767 22188 6684 22216
rect 8071 22188 8116 22216
rect 5767 22185 5779 22188
rect 5721 22179 5779 22185
rect 6656 22160 6684 22188
rect 8110 22176 8116 22188
rect 8168 22176 8174 22228
rect 8570 22216 8576 22228
rect 8531 22188 8576 22216
rect 8570 22176 8576 22188
rect 8628 22176 8634 22228
rect 9766 22176 9772 22228
rect 9824 22216 9830 22228
rect 10229 22219 10287 22225
rect 10229 22216 10241 22219
rect 9824 22188 10241 22216
rect 9824 22176 9830 22188
rect 10229 22185 10241 22188
rect 10275 22216 10287 22219
rect 10594 22216 10600 22228
rect 10275 22188 10600 22216
rect 10275 22185 10287 22188
rect 10229 22179 10287 22185
rect 10594 22176 10600 22188
rect 10652 22176 10658 22228
rect 10870 22216 10876 22228
rect 10831 22188 10876 22216
rect 10870 22176 10876 22188
rect 10928 22176 10934 22228
rect 11422 22176 11428 22228
rect 11480 22216 11486 22228
rect 14642 22216 14648 22228
rect 11480 22188 12388 22216
rect 14603 22188 14648 22216
rect 11480 22176 11486 22188
rect 4801 22151 4859 22157
rect 4801 22117 4813 22151
rect 4847 22117 4859 22151
rect 5537 22151 5595 22157
rect 4801 22111 4859 22117
rect 5000 22120 5304 22148
rect 1578 22080 1584 22092
rect 1539 22052 1584 22080
rect 1578 22040 1584 22052
rect 1636 22040 1642 22092
rect 2314 22040 2320 22092
rect 2372 22080 2378 22092
rect 2372 22052 2636 22080
rect 2372 22040 2378 22052
rect 2222 21972 2228 22024
rect 2280 22012 2286 22024
rect 2608 22021 2636 22052
rect 2774 22040 2780 22092
rect 2832 22080 2838 22092
rect 3237 22083 3295 22089
rect 3237 22080 3249 22083
rect 2832 22052 3249 22080
rect 2832 22040 2838 22052
rect 3237 22049 3249 22052
rect 3283 22049 3295 22083
rect 5000 22080 5028 22120
rect 5166 22080 5172 22092
rect 3237 22043 3295 22049
rect 3896 22052 5028 22080
rect 5127 22052 5172 22080
rect 2501 22015 2559 22021
rect 2501 22012 2513 22015
rect 2280 21984 2513 22012
rect 2280 21972 2286 21984
rect 2501 21981 2513 21984
rect 2547 21981 2559 22015
rect 2501 21975 2559 21981
rect 2593 22015 2651 22021
rect 2593 21981 2605 22015
rect 2639 21981 2651 22015
rect 2593 21975 2651 21981
rect 1397 21947 1455 21953
rect 1397 21913 1409 21947
rect 1443 21944 1455 21947
rect 3896 21944 3924 22052
rect 5166 22040 5172 22052
rect 5224 22040 5230 22092
rect 5276 22080 5304 22120
rect 5537 22117 5549 22151
rect 5583 22148 5595 22151
rect 5902 22148 5908 22160
rect 5583 22120 5908 22148
rect 5583 22117 5595 22120
rect 5537 22111 5595 22117
rect 5902 22108 5908 22120
rect 5960 22108 5966 22160
rect 6638 22108 6644 22160
rect 6696 22148 6702 22160
rect 8478 22148 8484 22160
rect 6696 22120 6914 22148
rect 8439 22120 8484 22148
rect 6696 22108 6702 22120
rect 6886 22080 6914 22120
rect 8478 22108 8484 22120
rect 8536 22108 8542 22160
rect 7009 22083 7067 22089
rect 7009 22080 7021 22083
rect 5276 22052 6776 22080
rect 6886 22052 7021 22080
rect 5534 22012 5540 22024
rect 5474 21984 5540 22012
rect 5534 21972 5540 21984
rect 5592 21972 5598 22024
rect 6748 22012 6776 22052
rect 7009 22049 7021 22052
rect 7055 22049 7067 22083
rect 7009 22043 7067 22049
rect 7098 22040 7104 22092
rect 7156 22080 7162 22092
rect 8588 22080 8616 22176
rect 9674 22108 9680 22160
rect 9732 22148 9738 22160
rect 10962 22148 10968 22160
rect 9732 22120 10968 22148
rect 9732 22108 9738 22120
rect 10962 22108 10968 22120
rect 11020 22108 11026 22160
rect 7156 22052 8616 22080
rect 10137 22083 10195 22089
rect 7156 22040 7162 22052
rect 10137 22049 10149 22083
rect 10183 22049 10195 22083
rect 10137 22043 10195 22049
rect 8662 22012 8668 22024
rect 6748 21984 8668 22012
rect 8662 21972 8668 21984
rect 8720 21972 8726 22024
rect 8757 22015 8815 22021
rect 8757 21981 8769 22015
rect 8803 22012 8815 22015
rect 9398 22012 9404 22024
rect 8803 21984 9404 22012
rect 8803 21981 8815 21984
rect 8757 21975 8815 21981
rect 9398 21972 9404 21984
rect 9456 21972 9462 22024
rect 1443 21916 3924 21944
rect 1443 21913 1455 21916
rect 1397 21907 1455 21913
rect 5626 21904 5632 21956
rect 5684 21944 5690 21956
rect 5994 21944 6000 21956
rect 5684 21916 6000 21944
rect 5684 21904 5690 21916
rect 5994 21904 6000 21916
rect 6052 21904 6058 21956
rect 6270 21904 6276 21956
rect 6328 21944 6334 21956
rect 10152 21944 10180 22043
rect 10226 22040 10232 22092
rect 10284 22080 10290 22092
rect 10781 22083 10839 22089
rect 10781 22080 10793 22083
rect 10284 22052 10793 22080
rect 10284 22040 10290 22052
rect 10781 22049 10793 22052
rect 10827 22049 10839 22083
rect 11606 22080 11612 22092
rect 10781 22043 10839 22049
rect 11348 22052 11612 22080
rect 11054 21972 11060 22024
rect 11112 22012 11118 22024
rect 11348 22012 11376 22052
rect 11606 22040 11612 22052
rect 11664 22040 11670 22092
rect 12066 22040 12072 22092
rect 12124 22089 12130 22092
rect 12124 22083 12183 22089
rect 12124 22049 12137 22083
rect 12171 22049 12183 22083
rect 12250 22080 12256 22092
rect 12211 22052 12256 22080
rect 12124 22043 12183 22049
rect 12124 22040 12130 22043
rect 12250 22040 12256 22052
rect 12308 22040 12314 22092
rect 12360 22089 12388 22188
rect 14642 22176 14648 22188
rect 14700 22176 14706 22228
rect 15749 22219 15807 22225
rect 15749 22185 15761 22219
rect 15795 22216 15807 22219
rect 16666 22216 16672 22228
rect 15795 22188 16672 22216
rect 15795 22185 15807 22188
rect 15749 22179 15807 22185
rect 16666 22176 16672 22188
rect 16724 22176 16730 22228
rect 17218 22176 17224 22228
rect 17276 22216 17282 22228
rect 23845 22219 23903 22225
rect 23845 22216 23857 22219
rect 17276 22188 23857 22216
rect 17276 22176 17282 22188
rect 23845 22185 23857 22188
rect 23891 22185 23903 22219
rect 24026 22216 24032 22228
rect 23939 22188 24032 22216
rect 23845 22179 23903 22185
rect 24026 22176 24032 22188
rect 24084 22216 24090 22228
rect 24210 22216 24216 22228
rect 24084 22188 24216 22216
rect 24084 22176 24090 22188
rect 24210 22176 24216 22188
rect 24268 22176 24274 22228
rect 25317 22219 25375 22225
rect 25317 22185 25329 22219
rect 25363 22216 25375 22219
rect 25590 22216 25596 22228
rect 25363 22188 25596 22216
rect 25363 22185 25375 22188
rect 25317 22179 25375 22185
rect 15470 22108 15476 22160
rect 15528 22148 15534 22160
rect 21726 22148 21732 22160
rect 15528 22120 16252 22148
rect 15528 22108 15534 22120
rect 12345 22083 12403 22089
rect 12345 22049 12357 22083
rect 12391 22049 12403 22083
rect 12345 22043 12403 22049
rect 13265 22083 13323 22089
rect 13265 22049 13277 22083
rect 13311 22080 13323 22083
rect 14182 22080 14188 22092
rect 13311 22052 14188 22080
rect 13311 22049 13323 22052
rect 13265 22043 13323 22049
rect 14182 22040 14188 22052
rect 14240 22040 14246 22092
rect 16111 22089 16117 22092
rect 16005 22083 16063 22089
rect 16005 22049 16017 22083
rect 16051 22049 16063 22083
rect 16005 22043 16063 22049
rect 16098 22083 16117 22089
rect 16098 22049 16110 22083
rect 16098 22043 16117 22049
rect 13538 22012 13544 22024
rect 11112 21984 11376 22012
rect 13499 21984 13544 22012
rect 11112 21972 11118 21984
rect 13538 21972 13544 21984
rect 13596 21972 13602 22024
rect 6328 21916 11192 21944
rect 6328 21904 6334 21916
rect 1486 21836 1492 21888
rect 1544 21876 1550 21888
rect 2406 21876 2412 21888
rect 1544 21848 2412 21876
rect 1544 21836 1550 21848
rect 2406 21836 2412 21848
rect 2464 21836 2470 21888
rect 3329 21879 3387 21885
rect 3329 21845 3341 21879
rect 3375 21876 3387 21879
rect 3694 21876 3700 21888
rect 3375 21848 3700 21876
rect 3375 21845 3387 21848
rect 3329 21839 3387 21845
rect 3694 21836 3700 21848
rect 3752 21836 3758 21888
rect 6012 21876 6040 21904
rect 11054 21876 11060 21888
rect 6012 21848 11060 21876
rect 11054 21836 11060 21848
rect 11112 21836 11118 21888
rect 11164 21876 11192 21916
rect 11606 21876 11612 21888
rect 11164 21848 11612 21876
rect 11606 21836 11612 21848
rect 11664 21836 11670 21888
rect 12158 21836 12164 21888
rect 12216 21876 12222 21888
rect 12342 21876 12348 21888
rect 12216 21848 12348 21876
rect 12216 21836 12222 21848
rect 12342 21836 12348 21848
rect 12400 21836 12406 21888
rect 12529 21879 12587 21885
rect 12529 21845 12541 21879
rect 12575 21876 12587 21879
rect 12710 21876 12716 21888
rect 12575 21848 12716 21876
rect 12575 21845 12587 21848
rect 12529 21839 12587 21845
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 15194 21836 15200 21888
rect 15252 21876 15258 21888
rect 15562 21876 15568 21888
rect 15252 21848 15568 21876
rect 15252 21836 15258 21848
rect 15562 21836 15568 21848
rect 15620 21836 15626 21888
rect 16020 21876 16048 22043
rect 16111 22040 16117 22043
rect 16169 22040 16175 22092
rect 16224 22089 16252 22120
rect 21376 22120 21732 22148
rect 16209 22083 16267 22089
rect 16209 22049 16221 22083
rect 16255 22049 16267 22083
rect 16209 22043 16267 22049
rect 16393 22083 16451 22089
rect 16393 22049 16405 22083
rect 16439 22049 16451 22083
rect 16393 22043 16451 22049
rect 16298 21904 16304 21956
rect 16356 21944 16362 21956
rect 16408 21944 16436 22043
rect 17862 22040 17868 22092
rect 17920 22080 17926 22092
rect 18046 22080 18052 22092
rect 17920 22052 18052 22080
rect 17920 22040 17926 22052
rect 18046 22040 18052 22052
rect 18104 22080 18110 22092
rect 18325 22083 18383 22089
rect 18325 22080 18337 22083
rect 18104 22052 18337 22080
rect 18104 22040 18110 22052
rect 18325 22049 18337 22052
rect 18371 22049 18383 22083
rect 18325 22043 18383 22049
rect 18592 22083 18650 22089
rect 18592 22049 18604 22083
rect 18638 22080 18650 22083
rect 19058 22080 19064 22092
rect 18638 22052 19064 22080
rect 18638 22049 18650 22052
rect 18592 22043 18650 22049
rect 19058 22040 19064 22052
rect 19116 22040 19122 22092
rect 20714 22080 20720 22092
rect 20675 22052 20720 22080
rect 20714 22040 20720 22052
rect 20772 22040 20778 22092
rect 20806 22040 20812 22092
rect 20864 22080 20870 22092
rect 21376 22089 21404 22120
rect 21726 22108 21732 22120
rect 21784 22108 21790 22160
rect 22462 22108 22468 22160
rect 22520 22148 22526 22160
rect 22520 22120 22692 22148
rect 22520 22108 22526 22120
rect 20901 22083 20959 22089
rect 20901 22080 20913 22083
rect 20864 22052 20913 22080
rect 20864 22040 20870 22052
rect 20901 22049 20913 22052
rect 20947 22049 20959 22083
rect 20901 22043 20959 22049
rect 21085 22083 21143 22089
rect 21085 22049 21097 22083
rect 21131 22049 21143 22083
rect 21085 22043 21143 22049
rect 21361 22083 21419 22089
rect 21361 22049 21373 22083
rect 21407 22080 21419 22083
rect 21634 22080 21640 22092
rect 21407 22052 21441 22080
rect 21595 22052 21640 22080
rect 21407 22049 21419 22052
rect 21361 22043 21419 22049
rect 20533 22015 20591 22021
rect 20533 21981 20545 22015
rect 20579 22012 20591 22015
rect 20990 22012 20996 22024
rect 20579 21984 20996 22012
rect 20579 21981 20591 21984
rect 20533 21975 20591 21981
rect 20990 21972 20996 21984
rect 21048 21972 21054 22024
rect 21100 22012 21128 22043
rect 21634 22040 21640 22052
rect 21692 22040 21698 22092
rect 22664 22080 22692 22120
rect 22738 22108 22744 22160
rect 22796 22148 22802 22160
rect 23106 22148 23112 22160
rect 22796 22120 22841 22148
rect 23019 22120 23112 22148
rect 22796 22108 22802 22120
rect 23106 22108 23112 22120
rect 23164 22148 23170 22160
rect 23290 22148 23296 22160
rect 23164 22120 23296 22148
rect 23164 22108 23170 22120
rect 23290 22108 23296 22120
rect 23348 22108 23354 22160
rect 23477 22151 23535 22157
rect 23477 22117 23489 22151
rect 23523 22148 23535 22151
rect 23566 22148 23572 22160
rect 23523 22120 23572 22148
rect 23523 22117 23535 22120
rect 23477 22111 23535 22117
rect 23566 22108 23572 22120
rect 23624 22148 23630 22160
rect 25332 22148 25360 22179
rect 25590 22176 25596 22188
rect 25648 22176 25654 22228
rect 26602 22216 26608 22228
rect 26252 22188 26608 22216
rect 26252 22160 26280 22188
rect 26602 22176 26608 22188
rect 26660 22176 26666 22228
rect 26694 22176 26700 22228
rect 26752 22216 26758 22228
rect 27893 22219 27951 22225
rect 27893 22216 27905 22219
rect 26752 22188 27905 22216
rect 26752 22176 26758 22188
rect 27893 22185 27905 22188
rect 27939 22185 27951 22219
rect 27893 22179 27951 22185
rect 23624 22120 25360 22148
rect 26053 22151 26111 22157
rect 23624 22108 23630 22120
rect 26053 22117 26065 22151
rect 26099 22148 26111 22151
rect 26234 22148 26240 22160
rect 26099 22120 26240 22148
rect 26099 22117 26111 22120
rect 26053 22111 26111 22117
rect 26234 22108 26240 22120
rect 26292 22108 26298 22160
rect 26418 22148 26424 22160
rect 26379 22120 26424 22148
rect 26418 22108 26424 22120
rect 26476 22108 26482 22160
rect 23017 22083 23075 22089
rect 23017 22080 23029 22083
rect 22664 22052 23029 22080
rect 23017 22049 23029 22052
rect 23063 22049 23075 22083
rect 23017 22043 23075 22049
rect 24854 22040 24860 22092
rect 24912 22080 24918 22092
rect 25593 22083 25651 22089
rect 25593 22080 25605 22083
rect 24912 22052 25605 22080
rect 24912 22040 24918 22052
rect 25593 22049 25605 22052
rect 25639 22049 25651 22083
rect 25593 22043 25651 22049
rect 25682 22040 25688 22092
rect 25740 22080 25746 22092
rect 25740 22052 25785 22080
rect 25740 22040 25746 22052
rect 26878 22040 26884 22092
rect 26936 22080 26942 22092
rect 27801 22083 27859 22089
rect 27801 22080 27813 22083
rect 26936 22052 27813 22080
rect 26936 22040 26942 22052
rect 27801 22049 27813 22052
rect 27847 22049 27859 22083
rect 27801 22043 27859 22049
rect 27985 22083 28043 22089
rect 27985 22049 27997 22083
rect 28031 22049 28043 22083
rect 27985 22043 28043 22049
rect 22560 22024 22612 22030
rect 21910 22012 21916 22024
rect 21100 21984 21916 22012
rect 21910 21972 21916 21984
rect 21968 21972 21974 22024
rect 24946 21972 24952 22024
rect 25004 22012 25010 22024
rect 25004 21984 25162 22012
rect 25004 21972 25010 21984
rect 27154 21972 27160 22024
rect 27212 22012 27218 22024
rect 28000 22012 28028 22043
rect 27212 21984 28028 22012
rect 27212 21972 27218 21984
rect 22560 21966 22612 21972
rect 16666 21944 16672 21956
rect 16356 21916 16436 21944
rect 16500 21916 16672 21944
rect 16356 21904 16362 21916
rect 16500 21876 16528 21916
rect 16666 21904 16672 21916
rect 16724 21944 16730 21956
rect 17678 21944 17684 21956
rect 16724 21916 17684 21944
rect 16724 21904 16730 21916
rect 17678 21904 17684 21916
rect 17736 21904 17742 21956
rect 26510 21904 26516 21956
rect 26568 21944 26574 21956
rect 26605 21947 26663 21953
rect 26605 21944 26617 21947
rect 26568 21916 26617 21944
rect 26568 21904 26574 21916
rect 26605 21913 26617 21916
rect 26651 21913 26663 21947
rect 26605 21907 26663 21913
rect 16020 21848 16528 21876
rect 19705 21879 19763 21885
rect 19705 21845 19717 21879
rect 19751 21876 19763 21879
rect 20898 21876 20904 21888
rect 19751 21848 20904 21876
rect 19751 21845 19763 21848
rect 19705 21839 19763 21845
rect 20898 21836 20904 21848
rect 20956 21836 20962 21888
rect 1104 21786 28888 21808
rect 1104 21734 5614 21786
rect 5666 21734 5678 21786
rect 5730 21734 5742 21786
rect 5794 21734 5806 21786
rect 5858 21734 14878 21786
rect 14930 21734 14942 21786
rect 14994 21734 15006 21786
rect 15058 21734 15070 21786
rect 15122 21734 24142 21786
rect 24194 21734 24206 21786
rect 24258 21734 24270 21786
rect 24322 21734 24334 21786
rect 24386 21734 28888 21786
rect 1104 21712 28888 21734
rect 4709 21675 4767 21681
rect 4709 21641 4721 21675
rect 4755 21672 4767 21675
rect 4982 21672 4988 21684
rect 4755 21644 4988 21672
rect 4755 21641 4767 21644
rect 4709 21635 4767 21641
rect 4982 21632 4988 21644
rect 5040 21632 5046 21684
rect 6822 21632 6828 21684
rect 6880 21672 6886 21684
rect 6917 21675 6975 21681
rect 6917 21672 6929 21675
rect 6880 21644 6929 21672
rect 6880 21632 6886 21644
rect 6917 21641 6929 21644
rect 6963 21641 6975 21675
rect 6917 21635 6975 21641
rect 7009 21675 7067 21681
rect 7009 21641 7021 21675
rect 7055 21672 7067 21675
rect 7098 21672 7104 21684
rect 7055 21644 7104 21672
rect 7055 21641 7067 21644
rect 7009 21635 7067 21641
rect 7098 21632 7104 21644
rect 7156 21632 7162 21684
rect 10226 21672 10232 21684
rect 10187 21644 10232 21672
rect 10226 21632 10232 21644
rect 10284 21632 10290 21684
rect 11054 21632 11060 21684
rect 11112 21672 11118 21684
rect 12158 21672 12164 21684
rect 11112 21644 12164 21672
rect 11112 21632 11118 21644
rect 12158 21632 12164 21644
rect 12216 21632 12222 21684
rect 12526 21672 12532 21684
rect 12487 21644 12532 21672
rect 12526 21632 12532 21644
rect 12584 21632 12590 21684
rect 12989 21675 13047 21681
rect 12989 21641 13001 21675
rect 13035 21672 13047 21675
rect 13538 21672 13544 21684
rect 13035 21644 13544 21672
rect 13035 21641 13047 21644
rect 12989 21635 13047 21641
rect 13538 21632 13544 21644
rect 13596 21632 13602 21684
rect 13630 21632 13636 21684
rect 13688 21672 13694 21684
rect 14274 21672 14280 21684
rect 13688 21644 14280 21672
rect 13688 21632 13694 21644
rect 14274 21632 14280 21644
rect 14332 21632 14338 21684
rect 15286 21632 15292 21684
rect 15344 21672 15350 21684
rect 15930 21672 15936 21684
rect 15344 21644 15936 21672
rect 15344 21632 15350 21644
rect 15930 21632 15936 21644
rect 15988 21632 15994 21684
rect 19058 21672 19064 21684
rect 19019 21644 19064 21672
rect 19058 21632 19064 21644
rect 19116 21632 19122 21684
rect 19794 21632 19800 21684
rect 19852 21672 19858 21684
rect 20162 21672 20168 21684
rect 19852 21644 20168 21672
rect 19852 21632 19858 21644
rect 20162 21632 20168 21644
rect 20220 21632 20226 21684
rect 21453 21675 21511 21681
rect 21453 21641 21465 21675
rect 21499 21672 21511 21675
rect 21726 21672 21732 21684
rect 21499 21644 21732 21672
rect 21499 21641 21511 21644
rect 21453 21635 21511 21641
rect 21726 21632 21732 21644
rect 21784 21632 21790 21684
rect 23566 21632 23572 21684
rect 23624 21672 23630 21684
rect 23753 21675 23811 21681
rect 23753 21672 23765 21675
rect 23624 21644 23765 21672
rect 23624 21632 23630 21644
rect 23753 21641 23765 21644
rect 23799 21641 23811 21675
rect 26602 21672 26608 21684
rect 26563 21644 26608 21672
rect 23753 21635 23811 21641
rect 26602 21632 26608 21644
rect 26660 21632 26666 21684
rect 27430 21672 27436 21684
rect 27391 21644 27436 21672
rect 27430 21632 27436 21644
rect 27488 21632 27494 21684
rect 2869 21607 2927 21613
rect 2869 21604 2881 21607
rect 2700 21576 2881 21604
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1670 21428 1676 21480
rect 1728 21468 1734 21480
rect 2700 21468 2728 21576
rect 2869 21573 2881 21576
rect 2915 21573 2927 21607
rect 2869 21567 2927 21573
rect 6362 21564 6368 21616
rect 6420 21604 6426 21616
rect 6420 21576 6960 21604
rect 6420 21564 6426 21576
rect 4246 21496 4252 21548
rect 4304 21536 4310 21548
rect 5353 21539 5411 21545
rect 5353 21536 5365 21539
rect 4304 21508 5365 21536
rect 4304 21496 4310 21508
rect 5353 21505 5365 21508
rect 5399 21536 5411 21539
rect 5810 21536 5816 21548
rect 5399 21508 5816 21536
rect 5399 21505 5411 21508
rect 5353 21499 5411 21505
rect 5810 21496 5816 21508
rect 5868 21536 5874 21548
rect 5868 21508 6408 21536
rect 5868 21496 5874 21508
rect 1728 21440 2728 21468
rect 5169 21471 5227 21477
rect 1728 21428 1734 21440
rect 5169 21437 5181 21471
rect 5215 21468 5227 21471
rect 6270 21468 6276 21480
rect 5215 21440 6276 21468
rect 5215 21437 5227 21440
rect 5169 21431 5227 21437
rect 6270 21428 6276 21440
rect 6328 21428 6334 21480
rect 1581 21403 1639 21409
rect 1581 21369 1593 21403
rect 1627 21400 1639 21403
rect 1762 21400 1768 21412
rect 1627 21372 1768 21400
rect 1627 21369 1639 21372
rect 1581 21363 1639 21369
rect 1762 21360 1768 21372
rect 1820 21360 1826 21412
rect 1857 21403 1915 21409
rect 1857 21369 1869 21403
rect 1903 21369 1915 21403
rect 1857 21363 1915 21369
rect 1949 21403 2007 21409
rect 1949 21369 1961 21403
rect 1995 21400 2007 21403
rect 2038 21400 2044 21412
rect 1995 21372 2044 21400
rect 1995 21369 2007 21372
rect 1949 21363 2007 21369
rect 1872 21332 1900 21363
rect 2038 21360 2044 21372
rect 2096 21360 2102 21412
rect 2130 21360 2136 21412
rect 2188 21400 2194 21412
rect 2317 21403 2375 21409
rect 2317 21400 2329 21403
rect 2188 21372 2329 21400
rect 2188 21360 2194 21372
rect 2317 21369 2329 21372
rect 2363 21369 2375 21403
rect 3326 21400 3332 21412
rect 2317 21363 2375 21369
rect 2424 21372 3332 21400
rect 2424 21332 2452 21372
rect 3326 21360 3332 21372
rect 3384 21360 3390 21412
rect 4798 21360 4804 21412
rect 4856 21400 4862 21412
rect 6380 21400 6408 21508
rect 6638 21496 6644 21548
rect 6696 21536 6702 21548
rect 6932 21545 6960 21576
rect 9858 21564 9864 21616
rect 9916 21604 9922 21616
rect 10594 21604 10600 21616
rect 9916 21576 10600 21604
rect 9916 21564 9922 21576
rect 10594 21564 10600 21576
rect 10652 21564 10658 21616
rect 13722 21604 13728 21616
rect 12820 21576 13728 21604
rect 6733 21539 6791 21545
rect 6733 21536 6745 21539
rect 6696 21508 6745 21536
rect 6696 21496 6702 21508
rect 6733 21505 6745 21508
rect 6779 21505 6791 21539
rect 6733 21499 6791 21505
rect 6917 21539 6975 21545
rect 6917 21505 6929 21539
rect 6963 21505 6975 21539
rect 6917 21499 6975 21505
rect 10778 21496 10784 21548
rect 10836 21536 10842 21548
rect 10873 21539 10931 21545
rect 10873 21536 10885 21539
rect 10836 21508 10885 21536
rect 10836 21496 10842 21508
rect 10873 21505 10885 21508
rect 10919 21536 10931 21539
rect 11054 21536 11060 21548
rect 10919 21508 11060 21536
rect 10919 21505 10931 21508
rect 10873 21499 10931 21505
rect 11054 21496 11060 21508
rect 11112 21536 11118 21548
rect 11514 21536 11520 21548
rect 11112 21508 11520 21536
rect 11112 21496 11118 21508
rect 11514 21496 11520 21508
rect 11572 21496 11578 21548
rect 6454 21428 6460 21480
rect 6512 21468 6518 21480
rect 7101 21471 7159 21477
rect 7101 21468 7113 21471
rect 6512 21440 7113 21468
rect 6512 21428 6518 21440
rect 7101 21437 7113 21440
rect 7147 21437 7159 21471
rect 7101 21431 7159 21437
rect 8662 21428 8668 21480
rect 8720 21468 8726 21480
rect 10597 21471 10655 21477
rect 10597 21468 10609 21471
rect 8720 21440 10609 21468
rect 8720 21428 8726 21440
rect 10597 21437 10609 21440
rect 10643 21437 10655 21471
rect 10597 21431 10655 21437
rect 10689 21471 10747 21477
rect 10689 21437 10701 21471
rect 10735 21468 10747 21471
rect 11238 21468 11244 21480
rect 10735 21440 11244 21468
rect 10735 21437 10747 21440
rect 10689 21431 10747 21437
rect 11238 21428 11244 21440
rect 11296 21428 11302 21480
rect 12066 21428 12072 21480
rect 12124 21477 12130 21480
rect 12124 21471 12183 21477
rect 12124 21437 12137 21471
rect 12171 21437 12183 21471
rect 12250 21468 12256 21480
rect 12211 21440 12256 21468
rect 12124 21431 12183 21437
rect 12124 21428 12130 21431
rect 12250 21428 12256 21440
rect 12308 21428 12314 21480
rect 12345 21471 12403 21477
rect 12345 21437 12357 21471
rect 12391 21468 12403 21471
rect 12820 21468 12848 21576
rect 13722 21564 13728 21576
rect 13780 21564 13786 21616
rect 13814 21564 13820 21616
rect 13872 21604 13878 21616
rect 17034 21604 17040 21616
rect 13872 21576 17040 21604
rect 13872 21564 13878 21576
rect 14642 21536 14648 21548
rect 13234 21508 14648 21536
rect 13234 21477 13262 21508
rect 14642 21496 14648 21508
rect 14700 21496 14706 21548
rect 12391 21440 12848 21468
rect 13219 21471 13277 21477
rect 12391 21437 12403 21440
rect 12345 21431 12403 21437
rect 13219 21437 13231 21471
rect 13265 21437 13277 21471
rect 13354 21468 13360 21480
rect 13315 21440 13360 21468
rect 13219 21431 13277 21437
rect 13234 21400 13262 21431
rect 13354 21428 13360 21440
rect 13412 21428 13418 21480
rect 15580 21477 15608 21576
rect 17034 21564 17040 21576
rect 17092 21564 17098 21616
rect 20070 21604 20076 21616
rect 19996 21576 20076 21604
rect 16114 21536 16120 21548
rect 15672 21508 16120 21536
rect 15672 21477 15700 21508
rect 16114 21496 16120 21508
rect 16172 21536 16178 21548
rect 16574 21536 16580 21548
rect 16172 21508 16580 21536
rect 16172 21496 16178 21508
rect 16574 21496 16580 21508
rect 16632 21496 16638 21548
rect 18785 21539 18843 21545
rect 18785 21505 18797 21539
rect 18831 21536 18843 21539
rect 19242 21536 19248 21548
rect 18831 21508 19248 21536
rect 18831 21505 18843 21508
rect 18785 21499 18843 21505
rect 19242 21496 19248 21508
rect 19300 21496 19306 21548
rect 19334 21496 19340 21548
rect 19392 21536 19398 21548
rect 19996 21536 20024 21576
rect 20070 21564 20076 21576
rect 20128 21564 20134 21616
rect 27982 21536 27988 21548
rect 19392 21522 20024 21536
rect 19392 21508 20010 21522
rect 22066 21508 22508 21536
rect 27943 21508 27988 21536
rect 19392 21496 19398 21508
rect 13449 21471 13507 21477
rect 13449 21437 13461 21471
rect 13495 21437 13507 21471
rect 13449 21431 13507 21437
rect 13627 21471 13685 21477
rect 13627 21437 13639 21471
rect 13673 21437 13685 21471
rect 13627 21431 13685 21437
rect 15565 21471 15623 21477
rect 15565 21437 15577 21471
rect 15611 21437 15623 21471
rect 15565 21431 15623 21437
rect 15657 21471 15715 21477
rect 15657 21437 15669 21471
rect 15703 21437 15715 21471
rect 15657 21431 15715 21437
rect 15749 21471 15807 21477
rect 15749 21437 15761 21471
rect 15795 21437 15807 21471
rect 15930 21468 15936 21480
rect 15891 21440 15936 21468
rect 15749 21431 15807 21437
rect 4856 21372 5212 21400
rect 6380 21372 13262 21400
rect 4856 21360 4862 21372
rect 2682 21332 2688 21344
rect 1872 21304 2452 21332
rect 2643 21304 2688 21332
rect 2682 21292 2688 21304
rect 2740 21292 2746 21344
rect 4154 21292 4160 21344
rect 4212 21332 4218 21344
rect 5077 21335 5135 21341
rect 5077 21332 5089 21335
rect 4212 21304 5089 21332
rect 4212 21292 4218 21304
rect 5077 21301 5089 21304
rect 5123 21301 5135 21335
rect 5184 21332 5212 21372
rect 11790 21332 11796 21344
rect 5184 21304 11796 21332
rect 5077 21295 5135 21301
rect 11790 21292 11796 21304
rect 11848 21292 11854 21344
rect 12894 21292 12900 21344
rect 12952 21332 12958 21344
rect 13464 21332 13492 21431
rect 13648 21400 13676 21431
rect 13722 21400 13728 21412
rect 13648 21372 13728 21400
rect 13722 21360 13728 21372
rect 13780 21360 13786 21412
rect 15194 21360 15200 21412
rect 15252 21400 15258 21412
rect 15470 21400 15476 21412
rect 15252 21372 15476 21400
rect 15252 21360 15258 21372
rect 15470 21360 15476 21372
rect 15528 21400 15534 21412
rect 15764 21400 15792 21431
rect 15930 21428 15936 21440
rect 15988 21428 15994 21480
rect 18877 21471 18935 21477
rect 18877 21437 18889 21471
rect 18923 21468 18935 21471
rect 18923 21440 20944 21468
rect 18923 21437 18935 21440
rect 18877 21431 18935 21437
rect 20916 21412 20944 21440
rect 20990 21428 20996 21480
rect 21048 21468 21054 21480
rect 22066 21468 22094 21508
rect 22370 21468 22376 21480
rect 21048 21440 22094 21468
rect 22331 21440 22376 21468
rect 21048 21428 21054 21440
rect 22370 21428 22376 21440
rect 22428 21428 22434 21480
rect 22480 21468 22508 21508
rect 27982 21496 27988 21508
rect 28040 21496 28046 21548
rect 24854 21468 24860 21480
rect 22480 21440 24860 21468
rect 24854 21428 24860 21440
rect 24912 21428 24918 21480
rect 25498 21477 25504 21480
rect 25225 21471 25283 21477
rect 25225 21437 25237 21471
rect 25271 21437 25283 21471
rect 25225 21431 25283 21437
rect 25492 21431 25504 21477
rect 25556 21468 25562 21480
rect 27798 21468 27804 21480
rect 25556 21440 25592 21468
rect 27759 21440 27804 21468
rect 15528 21372 15792 21400
rect 15528 21360 15534 21372
rect 20070 21360 20076 21412
rect 20128 21400 20134 21412
rect 20441 21403 20499 21409
rect 20441 21400 20453 21403
rect 20128 21372 20453 21400
rect 20128 21360 20134 21372
rect 20441 21369 20453 21372
rect 20487 21369 20499 21403
rect 20441 21363 20499 21369
rect 20530 21360 20536 21412
rect 20588 21400 20594 21412
rect 20898 21400 20904 21412
rect 20588 21372 20633 21400
rect 20811 21372 20904 21400
rect 20588 21360 20594 21372
rect 20898 21360 20904 21372
rect 20956 21400 20962 21412
rect 22278 21400 22284 21412
rect 20956 21372 22284 21400
rect 20956 21360 20962 21372
rect 22278 21360 22284 21372
rect 22336 21360 22342 21412
rect 22554 21360 22560 21412
rect 22612 21409 22618 21412
rect 22612 21403 22676 21409
rect 22612 21369 22630 21403
rect 22664 21369 22676 21403
rect 22612 21363 22676 21369
rect 22612 21360 22618 21363
rect 23290 21360 23296 21412
rect 23348 21400 23354 21412
rect 25240 21400 25268 21431
rect 25498 21428 25504 21431
rect 25556 21428 25562 21440
rect 27798 21428 27804 21440
rect 27856 21428 27862 21480
rect 27893 21471 27951 21477
rect 27893 21437 27905 21471
rect 27939 21468 27951 21471
rect 28074 21468 28080 21480
rect 27939 21440 28080 21468
rect 27939 21437 27951 21440
rect 27893 21431 27951 21437
rect 28074 21428 28080 21440
rect 28132 21428 28138 21480
rect 26050 21400 26056 21412
rect 23348 21372 26056 21400
rect 23348 21360 23354 21372
rect 26050 21360 26056 21372
rect 26108 21360 26114 21412
rect 14090 21332 14096 21344
rect 12952 21304 14096 21332
rect 12952 21292 12958 21304
rect 14090 21292 14096 21304
rect 14148 21292 14154 21344
rect 15289 21335 15347 21341
rect 15289 21301 15301 21335
rect 15335 21332 15347 21335
rect 16390 21332 16396 21344
rect 15335 21304 16396 21332
rect 15335 21301 15347 21304
rect 15289 21295 15347 21301
rect 16390 21292 16396 21304
rect 16448 21292 16454 21344
rect 18230 21292 18236 21344
rect 18288 21332 18294 21344
rect 18417 21335 18475 21341
rect 18417 21332 18429 21335
rect 18288 21304 18429 21332
rect 18288 21292 18294 21304
rect 18417 21301 18429 21304
rect 18463 21301 18475 21335
rect 18417 21295 18475 21301
rect 19058 21292 19064 21344
rect 19116 21332 19122 21344
rect 20165 21335 20223 21341
rect 20165 21332 20177 21335
rect 19116 21304 20177 21332
rect 19116 21292 19122 21304
rect 20165 21301 20177 21304
rect 20211 21301 20223 21335
rect 20165 21295 20223 21301
rect 20254 21292 20260 21344
rect 20312 21332 20318 21344
rect 21269 21335 21327 21341
rect 21269 21332 21281 21335
rect 20312 21304 21281 21332
rect 20312 21292 20318 21304
rect 21269 21301 21281 21304
rect 21315 21301 21327 21335
rect 22296 21332 22324 21360
rect 22738 21332 22744 21344
rect 22296 21304 22744 21332
rect 21269 21295 21327 21301
rect 22738 21292 22744 21304
rect 22796 21292 22802 21344
rect 1104 21242 28888 21264
rect 1104 21190 10246 21242
rect 10298 21190 10310 21242
rect 10362 21190 10374 21242
rect 10426 21190 10438 21242
rect 10490 21190 19510 21242
rect 19562 21190 19574 21242
rect 19626 21190 19638 21242
rect 19690 21190 19702 21242
rect 19754 21190 28888 21242
rect 1104 21168 28888 21190
rect 1489 21131 1547 21137
rect 1489 21097 1501 21131
rect 1535 21097 1547 21131
rect 1489 21091 1547 21097
rect 2685 21131 2743 21137
rect 2685 21097 2697 21131
rect 2731 21128 2743 21131
rect 3329 21131 3387 21137
rect 3329 21128 3341 21131
rect 2731 21100 3341 21128
rect 2731 21097 2743 21100
rect 2685 21091 2743 21097
rect 3329 21097 3341 21100
rect 3375 21097 3387 21131
rect 3694 21128 3700 21140
rect 3655 21100 3700 21128
rect 3329 21091 3387 21097
rect 1504 21060 1532 21091
rect 3694 21088 3700 21100
rect 3752 21088 3758 21140
rect 3789 21131 3847 21137
rect 3789 21097 3801 21131
rect 3835 21128 3847 21131
rect 5350 21128 5356 21140
rect 3835 21100 5356 21128
rect 3835 21097 3847 21100
rect 3789 21091 3847 21097
rect 5350 21088 5356 21100
rect 5408 21088 5414 21140
rect 6914 21088 6920 21140
rect 6972 21128 6978 21140
rect 7009 21131 7067 21137
rect 7009 21128 7021 21131
rect 6972 21100 7021 21128
rect 6972 21088 6978 21100
rect 7009 21097 7021 21100
rect 7055 21097 7067 21131
rect 7009 21091 7067 21097
rect 9674 21088 9680 21140
rect 9732 21128 9738 21140
rect 10778 21128 10784 21140
rect 9732 21100 10784 21128
rect 9732 21088 9738 21100
rect 10778 21088 10784 21100
rect 10836 21088 10842 21140
rect 12250 21128 12256 21140
rect 10980 21100 12256 21128
rect 5902 21060 5908 21072
rect 1504 21032 5908 21060
rect 5902 21020 5908 21032
rect 5960 21020 5966 21072
rect 10980 21060 11008 21100
rect 12250 21088 12256 21100
rect 12308 21128 12314 21140
rect 15381 21131 15439 21137
rect 12308 21100 13676 21128
rect 12308 21088 12314 21100
rect 10888 21032 11008 21060
rect 1670 20992 1676 21004
rect 1631 20964 1676 20992
rect 1670 20952 1676 20964
rect 1728 20952 1734 21004
rect 2777 20995 2835 21001
rect 2777 20961 2789 20995
rect 2823 20992 2835 20995
rect 3234 20992 3240 21004
rect 2823 20964 3240 20992
rect 2823 20961 2835 20964
rect 2777 20955 2835 20961
rect 3234 20952 3240 20964
rect 3292 20952 3298 21004
rect 3510 20952 3516 21004
rect 3568 20992 3574 21004
rect 6822 20992 6828 21004
rect 3568 20964 3924 20992
rect 6783 20964 6828 20992
rect 3568 20952 3574 20964
rect 2685 20927 2743 20933
rect 2685 20893 2697 20927
rect 2731 20893 2743 20927
rect 2685 20887 2743 20893
rect 2700 20856 2728 20887
rect 2958 20856 2964 20868
rect 2700 20828 2964 20856
rect 2958 20816 2964 20828
rect 3016 20816 3022 20868
rect 3252 20856 3280 20952
rect 3896 20936 3924 20964
rect 6822 20952 6828 20964
rect 6880 20952 6886 21004
rect 7098 20992 7104 21004
rect 7059 20964 7104 20992
rect 7098 20952 7104 20964
rect 7156 20952 7162 21004
rect 7282 20992 7288 21004
rect 7243 20964 7288 20992
rect 7282 20952 7288 20964
rect 7340 20952 7346 21004
rect 9217 20995 9275 21001
rect 9217 20961 9229 20995
rect 9263 20961 9275 20995
rect 9674 20992 9680 21004
rect 9635 20964 9680 20992
rect 9217 20955 9275 20961
rect 3878 20884 3884 20936
rect 3936 20924 3942 20936
rect 3936 20896 4029 20924
rect 3936 20884 3942 20896
rect 4798 20856 4804 20868
rect 3252 20828 4804 20856
rect 4798 20816 4804 20828
rect 4856 20816 4862 20868
rect 9232 20856 9260 20955
rect 9674 20952 9680 20964
rect 9732 20952 9738 21004
rect 10888 21001 10916 21032
rect 11146 21020 11152 21072
rect 11204 21060 11210 21072
rect 11514 21060 11520 21072
rect 11204 21032 11520 21060
rect 11204 21020 11210 21032
rect 11514 21020 11520 21032
rect 11572 21020 11578 21072
rect 12066 21020 12072 21072
rect 12124 21060 12130 21072
rect 12124 21032 13584 21060
rect 12124 21020 12130 21032
rect 10781 20995 10839 21001
rect 10781 20961 10793 20995
rect 10827 20961 10839 20995
rect 10781 20955 10839 20961
rect 10873 20995 10931 21001
rect 10873 20961 10885 20995
rect 10919 20961 10931 20995
rect 10873 20955 10931 20961
rect 9950 20924 9956 20936
rect 9911 20896 9956 20924
rect 9950 20884 9956 20896
rect 10008 20884 10014 20936
rect 10796 20924 10824 20955
rect 10962 20952 10968 21004
rect 11020 20992 11026 21004
rect 11020 20964 11065 20992
rect 11020 20952 11026 20964
rect 12084 20924 12112 21020
rect 12158 20952 12164 21004
rect 12216 20992 12222 21004
rect 12345 20995 12403 21001
rect 12345 20992 12357 20995
rect 12216 20964 12357 20992
rect 12216 20952 12222 20964
rect 12345 20961 12357 20964
rect 12391 20961 12403 20995
rect 12345 20955 12403 20961
rect 12437 20995 12495 21001
rect 12437 20961 12449 20995
rect 12483 20961 12495 20995
rect 12437 20955 12495 20961
rect 12534 20995 12592 21001
rect 12534 20961 12546 20995
rect 12580 20961 12592 20995
rect 12710 20992 12716 21004
rect 12671 20964 12716 20992
rect 12534 20955 12592 20961
rect 10796 20896 12112 20924
rect 10962 20856 10968 20868
rect 9232 20828 10968 20856
rect 10962 20816 10968 20828
rect 11020 20816 11026 20868
rect 12452 20856 12480 20955
rect 12549 20924 12577 20955
rect 12710 20952 12716 20964
rect 12768 20952 12774 21004
rect 13556 21001 13584 21032
rect 13648 21001 13676 21100
rect 15381 21097 15393 21131
rect 15427 21128 15439 21131
rect 15930 21128 15936 21140
rect 15427 21100 15936 21128
rect 15427 21097 15439 21100
rect 15381 21091 15439 21097
rect 15930 21088 15936 21100
rect 15988 21088 15994 21140
rect 18230 21128 18236 21140
rect 18191 21100 18236 21128
rect 18230 21088 18236 21100
rect 18288 21088 18294 21140
rect 19794 21088 19800 21140
rect 19852 21128 19858 21140
rect 20530 21128 20536 21140
rect 19852 21100 20536 21128
rect 19852 21088 19858 21100
rect 20530 21088 20536 21100
rect 20588 21088 20594 21140
rect 20714 21088 20720 21140
rect 20772 21128 20778 21140
rect 21085 21131 21143 21137
rect 21085 21128 21097 21131
rect 20772 21100 21097 21128
rect 20772 21088 20778 21100
rect 21085 21097 21097 21100
rect 21131 21097 21143 21131
rect 21085 21091 21143 21097
rect 21174 21088 21180 21140
rect 21232 21128 21238 21140
rect 21453 21131 21511 21137
rect 21453 21128 21465 21131
rect 21232 21100 21465 21128
rect 21232 21088 21238 21100
rect 21453 21097 21465 21100
rect 21499 21097 21511 21131
rect 22554 21128 22560 21140
rect 22515 21100 22560 21128
rect 21453 21091 21511 21097
rect 22554 21088 22560 21100
rect 22612 21088 22618 21140
rect 22922 21088 22928 21140
rect 22980 21088 22986 21140
rect 23017 21131 23075 21137
rect 23017 21097 23029 21131
rect 23063 21128 23075 21131
rect 23566 21128 23572 21140
rect 23063 21100 23572 21128
rect 23063 21097 23075 21100
rect 23017 21091 23075 21097
rect 23566 21088 23572 21100
rect 23624 21088 23630 21140
rect 24026 21088 24032 21140
rect 24084 21128 24090 21140
rect 24305 21131 24363 21137
rect 24305 21128 24317 21131
rect 24084 21100 24317 21128
rect 24084 21088 24090 21100
rect 24305 21097 24317 21100
rect 24351 21097 24363 21131
rect 24486 21128 24492 21140
rect 24447 21100 24492 21128
rect 24305 21091 24363 21097
rect 24486 21088 24492 21100
rect 24544 21088 24550 21140
rect 24854 21088 24860 21140
rect 24912 21128 24918 21140
rect 24912 21100 26740 21128
rect 24912 21088 24918 21100
rect 14734 21020 14740 21072
rect 14792 21060 14798 21072
rect 17954 21060 17960 21072
rect 14792 21032 15148 21060
rect 14792 21020 14798 21032
rect 13541 20995 13599 21001
rect 13541 20961 13553 20995
rect 13587 20961 13599 20995
rect 13541 20955 13599 20961
rect 13633 20995 13691 21001
rect 13633 20961 13645 20995
rect 13679 20961 13691 20995
rect 13633 20955 13691 20961
rect 12894 20924 12900 20936
rect 12549 20896 12900 20924
rect 12728 20868 12756 20896
rect 12894 20884 12900 20896
rect 12952 20884 12958 20936
rect 13556 20924 13584 20955
rect 13722 20952 13728 21004
rect 13780 20992 13786 21004
rect 14274 20992 14280 21004
rect 13780 20964 14280 20992
rect 13780 20952 13786 20964
rect 14274 20952 14280 20964
rect 14332 20952 14338 21004
rect 15120 21001 15148 21032
rect 15212 21032 15332 21060
rect 17915 21032 17960 21060
rect 15212 21001 15240 21032
rect 15013 20995 15071 21001
rect 15013 20992 15025 20995
rect 14384 20964 15025 20992
rect 14384 20924 14412 20964
rect 15013 20961 15025 20964
rect 15059 20961 15071 20995
rect 15013 20955 15071 20961
rect 15105 20995 15163 21001
rect 15105 20961 15117 20995
rect 15151 20961 15163 20995
rect 15105 20955 15163 20961
rect 15197 20995 15255 21001
rect 15197 20961 15209 20995
rect 15243 20961 15255 20995
rect 15304 20992 15332 21032
rect 17954 21020 17960 21032
rect 18012 21020 18018 21072
rect 18046 21020 18052 21072
rect 18104 21060 18110 21072
rect 18141 21063 18199 21069
rect 18141 21060 18153 21063
rect 18104 21032 18153 21060
rect 18104 21020 18110 21032
rect 18141 21029 18153 21032
rect 18187 21060 18199 21063
rect 18782 21060 18788 21072
rect 18187 21032 18788 21060
rect 18187 21029 18199 21032
rect 18141 21023 18199 21029
rect 18782 21020 18788 21032
rect 18840 21020 18846 21072
rect 19058 21020 19064 21072
rect 19116 21060 19122 21072
rect 20990 21060 20996 21072
rect 19116 21032 20996 21060
rect 19116 21020 19122 21032
rect 20990 21020 20996 21032
rect 21048 21020 21054 21072
rect 21294 21063 21352 21069
rect 21294 21029 21306 21063
rect 21340 21060 21352 21063
rect 21726 21060 21732 21072
rect 21340 21032 21732 21060
rect 21340 21029 21352 21032
rect 21294 21023 21352 21029
rect 21726 21020 21732 21032
rect 21784 21020 21790 21072
rect 22940 21060 22968 21088
rect 22940 21032 23244 21060
rect 15470 20992 15476 21004
rect 15304 20964 15476 20992
rect 15197 20955 15255 20961
rect 13556 20896 14412 20924
rect 15028 20924 15056 20955
rect 15470 20952 15476 20964
rect 15528 20952 15534 21004
rect 15562 20952 15568 21004
rect 15620 20992 15626 21004
rect 15841 20995 15899 21001
rect 15841 20992 15853 20995
rect 15620 20964 15853 20992
rect 15620 20952 15626 20964
rect 15841 20961 15853 20964
rect 15887 20961 15899 20995
rect 15841 20955 15899 20961
rect 17972 20924 18000 21020
rect 18230 20992 18236 21004
rect 18191 20964 18236 20992
rect 18230 20952 18236 20964
rect 18288 20952 18294 21004
rect 20898 20952 20904 21004
rect 20956 20992 20962 21004
rect 21177 20995 21235 21001
rect 21177 20992 21189 20995
rect 20956 20964 21189 20992
rect 20956 20952 20962 20964
rect 21177 20961 21189 20964
rect 21223 20961 21235 20995
rect 22922 20992 22928 21004
rect 22883 20964 22928 20992
rect 21177 20955 21235 20961
rect 22922 20952 22928 20964
rect 22980 20952 22986 21004
rect 18782 20924 18788 20936
rect 15028 20896 16068 20924
rect 17972 20896 18788 20924
rect 12526 20856 12532 20868
rect 11992 20828 12388 20856
rect 12452 20828 12532 20856
rect 2130 20748 2136 20800
rect 2188 20788 2194 20800
rect 2225 20791 2283 20797
rect 2225 20788 2237 20791
rect 2188 20760 2237 20788
rect 2188 20748 2194 20760
rect 2225 20757 2237 20760
rect 2271 20757 2283 20791
rect 2225 20751 2283 20757
rect 8478 20748 8484 20800
rect 8536 20788 8542 20800
rect 8938 20788 8944 20800
rect 8536 20760 8944 20788
rect 8536 20748 8542 20760
rect 8938 20748 8944 20760
rect 8996 20788 9002 20800
rect 9033 20791 9091 20797
rect 9033 20788 9045 20791
rect 8996 20760 9045 20788
rect 8996 20748 9002 20760
rect 9033 20757 9045 20760
rect 9079 20757 9091 20791
rect 9766 20788 9772 20800
rect 9727 20760 9772 20788
rect 9033 20751 9091 20757
rect 9766 20748 9772 20760
rect 9824 20748 9830 20800
rect 9861 20791 9919 20797
rect 9861 20757 9873 20791
rect 9907 20788 9919 20791
rect 10042 20788 10048 20800
rect 9907 20760 10048 20788
rect 9907 20757 9919 20760
rect 9861 20751 9919 20757
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 11149 20791 11207 20797
rect 11149 20757 11161 20791
rect 11195 20788 11207 20791
rect 11992 20788 12020 20828
rect 11195 20760 12020 20788
rect 12069 20791 12127 20797
rect 11195 20757 11207 20760
rect 11149 20751 11207 20757
rect 12069 20757 12081 20791
rect 12115 20788 12127 20791
rect 12250 20788 12256 20800
rect 12115 20760 12256 20788
rect 12115 20757 12127 20760
rect 12069 20751 12127 20757
rect 12250 20748 12256 20760
rect 12308 20748 12314 20800
rect 12360 20788 12388 20828
rect 12526 20816 12532 20828
rect 12584 20816 12590 20868
rect 12710 20816 12716 20868
rect 12768 20816 12774 20868
rect 14550 20816 14556 20868
rect 14608 20856 14614 20868
rect 15562 20856 15568 20868
rect 14608 20828 15568 20856
rect 14608 20816 14614 20828
rect 15562 20816 15568 20828
rect 15620 20816 15626 20868
rect 16040 20865 16068 20896
rect 18782 20884 18788 20896
rect 18840 20884 18846 20936
rect 20806 20924 20812 20936
rect 20767 20896 20812 20924
rect 20806 20884 20812 20896
rect 20864 20884 20870 20936
rect 22094 20884 22100 20936
rect 22152 20924 22158 20936
rect 23014 20924 23020 20936
rect 22152 20896 23020 20924
rect 22152 20884 22158 20896
rect 23014 20884 23020 20896
rect 23072 20924 23078 20936
rect 23109 20927 23167 20933
rect 23109 20924 23121 20927
rect 23072 20896 23121 20924
rect 23072 20884 23078 20896
rect 23109 20893 23121 20896
rect 23155 20893 23167 20927
rect 23109 20887 23167 20893
rect 16025 20859 16083 20865
rect 16025 20825 16037 20859
rect 16071 20825 16083 20859
rect 16025 20819 16083 20825
rect 16114 20816 16120 20868
rect 16172 20856 16178 20868
rect 23216 20856 23244 21032
rect 23842 21020 23848 21072
rect 23900 21060 23906 21072
rect 24213 21063 24271 21069
rect 24213 21060 24225 21063
rect 23900 21032 24225 21060
rect 23900 21020 23906 21032
rect 24213 21029 24225 21032
rect 24259 21029 24271 21063
rect 24213 21023 24271 21029
rect 25593 21063 25651 21069
rect 25593 21029 25605 21063
rect 25639 21060 25651 21063
rect 25958 21060 25964 21072
rect 25639 21032 25964 21060
rect 25639 21029 25651 21032
rect 25593 21023 25651 21029
rect 25958 21020 25964 21032
rect 26016 21020 26022 21072
rect 26712 21069 26740 21100
rect 26697 21063 26755 21069
rect 26697 21029 26709 21063
rect 26743 21029 26755 21063
rect 26697 21023 26755 21029
rect 23934 20952 23940 21004
rect 23992 20952 23998 21004
rect 24121 20995 24179 21001
rect 24121 20961 24133 20995
rect 24167 20961 24179 20995
rect 25406 20992 25412 21004
rect 25367 20964 25412 20992
rect 24121 20955 24179 20961
rect 23566 20884 23572 20936
rect 23624 20924 23630 20936
rect 23952 20924 23980 20952
rect 24136 20924 24164 20955
rect 25406 20952 25412 20964
rect 25464 20952 25470 21004
rect 26878 20992 26884 21004
rect 26839 20964 26884 20992
rect 26878 20952 26884 20964
rect 26936 20952 26942 21004
rect 27985 20995 28043 21001
rect 27985 20961 27997 20995
rect 28031 20961 28043 20995
rect 27985 20955 28043 20961
rect 28000 20924 28028 20955
rect 23624 20896 24164 20924
rect 24872 20896 28028 20924
rect 23624 20884 23630 20896
rect 23937 20859 23995 20865
rect 23937 20856 23949 20859
rect 16172 20828 22094 20856
rect 23216 20828 23949 20856
rect 16172 20816 16178 20828
rect 12894 20788 12900 20800
rect 12360 20760 12900 20788
rect 12894 20748 12900 20760
rect 12952 20748 12958 20800
rect 13906 20788 13912 20800
rect 13867 20760 13912 20788
rect 13906 20748 13912 20760
rect 13964 20748 13970 20800
rect 14090 20748 14096 20800
rect 14148 20788 14154 20800
rect 20254 20788 20260 20800
rect 14148 20760 20260 20788
rect 14148 20748 14154 20760
rect 20254 20748 20260 20760
rect 20312 20748 20318 20800
rect 22066 20788 22094 20828
rect 23937 20825 23949 20828
rect 23983 20856 23995 20859
rect 24762 20856 24768 20868
rect 23983 20828 24768 20856
rect 23983 20825 23995 20828
rect 23937 20819 23995 20825
rect 24762 20816 24768 20828
rect 24820 20816 24826 20868
rect 22462 20788 22468 20800
rect 22066 20760 22468 20788
rect 22462 20748 22468 20760
rect 22520 20788 22526 20800
rect 24872 20788 24900 20896
rect 28074 20788 28080 20800
rect 22520 20760 24900 20788
rect 28035 20760 28080 20788
rect 22520 20748 22526 20760
rect 28074 20748 28080 20760
rect 28132 20748 28138 20800
rect 1104 20698 28888 20720
rect 1104 20646 5614 20698
rect 5666 20646 5678 20698
rect 5730 20646 5742 20698
rect 5794 20646 5806 20698
rect 5858 20646 14878 20698
rect 14930 20646 14942 20698
rect 14994 20646 15006 20698
rect 15058 20646 15070 20698
rect 15122 20646 24142 20698
rect 24194 20646 24206 20698
rect 24258 20646 24270 20698
rect 24322 20646 24334 20698
rect 24386 20646 28888 20698
rect 1104 20624 28888 20646
rect 1765 20587 1823 20593
rect 1765 20553 1777 20587
rect 1811 20584 1823 20587
rect 2682 20584 2688 20596
rect 1811 20556 2688 20584
rect 1811 20553 1823 20556
rect 1765 20547 1823 20553
rect 2682 20544 2688 20556
rect 2740 20544 2746 20596
rect 2958 20584 2964 20596
rect 2919 20556 2964 20584
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 4525 20587 4583 20593
rect 4525 20553 4537 20587
rect 4571 20584 4583 20587
rect 4614 20584 4620 20596
rect 4571 20556 4620 20584
rect 4571 20553 4583 20556
rect 4525 20547 4583 20553
rect 4614 20544 4620 20556
rect 4672 20544 4678 20596
rect 11333 20587 11391 20593
rect 11333 20553 11345 20587
rect 11379 20584 11391 20587
rect 11606 20584 11612 20596
rect 11379 20556 11612 20584
rect 11379 20553 11391 20556
rect 11333 20547 11391 20553
rect 11606 20544 11612 20556
rect 11664 20544 11670 20596
rect 13265 20587 13323 20593
rect 13265 20553 13277 20587
rect 13311 20584 13323 20587
rect 14182 20584 14188 20596
rect 13311 20556 14188 20584
rect 13311 20553 13323 20556
rect 13265 20547 13323 20553
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 20438 20544 20444 20596
rect 20496 20584 20502 20596
rect 20809 20587 20867 20593
rect 20809 20584 20821 20587
rect 20496 20556 20821 20584
rect 20496 20544 20502 20556
rect 20809 20553 20821 20556
rect 20855 20553 20867 20587
rect 20809 20547 20867 20553
rect 22005 20587 22063 20593
rect 22005 20553 22017 20587
rect 22051 20584 22063 20587
rect 22922 20584 22928 20596
rect 22051 20556 22928 20584
rect 22051 20553 22063 20556
rect 22005 20547 22063 20553
rect 12526 20476 12532 20528
rect 12584 20476 12590 20528
rect 13354 20476 13360 20528
rect 13412 20476 13418 20528
rect 13906 20476 13912 20528
rect 13964 20516 13970 20528
rect 13964 20488 15332 20516
rect 13964 20476 13970 20488
rect 2958 20448 2964 20460
rect 2871 20420 2964 20448
rect 1946 20380 1952 20392
rect 1907 20352 1952 20380
rect 1946 20340 1952 20352
rect 2004 20340 2010 20392
rect 2884 20389 2912 20420
rect 2958 20408 2964 20420
rect 3016 20448 3022 20460
rect 3786 20448 3792 20460
rect 3016 20420 3792 20448
rect 3016 20408 3022 20420
rect 3786 20408 3792 20420
rect 3844 20408 3850 20460
rect 7650 20448 7656 20460
rect 7611 20420 7656 20448
rect 7650 20408 7656 20420
rect 7708 20408 7714 20460
rect 8113 20451 8171 20457
rect 8113 20417 8125 20451
rect 8159 20448 8171 20451
rect 9858 20448 9864 20460
rect 8159 20420 9864 20448
rect 8159 20417 8171 20420
rect 8113 20411 8171 20417
rect 9858 20408 9864 20420
rect 9916 20408 9922 20460
rect 12549 20448 12577 20476
rect 13372 20448 13400 20476
rect 15304 20448 15332 20488
rect 16022 20476 16028 20528
rect 16080 20476 16086 20528
rect 20824 20516 20852 20547
rect 22922 20544 22928 20556
rect 22980 20544 22986 20596
rect 24486 20544 24492 20596
rect 24544 20584 24550 20596
rect 26142 20584 26148 20596
rect 24544 20556 26148 20584
rect 24544 20544 24550 20556
rect 26142 20544 26148 20556
rect 26200 20544 26206 20596
rect 27341 20587 27399 20593
rect 27341 20553 27353 20587
rect 27387 20584 27399 20587
rect 27522 20584 27528 20596
rect 27387 20556 27528 20584
rect 27387 20553 27399 20556
rect 27341 20547 27399 20553
rect 27522 20544 27528 20556
rect 27580 20544 27586 20596
rect 20824 20488 22094 20516
rect 12549 20420 15148 20448
rect 15304 20420 15424 20448
rect 2869 20383 2927 20389
rect 2869 20349 2881 20383
rect 2915 20349 2927 20383
rect 2869 20343 2927 20349
rect 3053 20383 3111 20389
rect 3053 20349 3065 20383
rect 3099 20349 3111 20383
rect 3053 20343 3111 20349
rect 4433 20383 4491 20389
rect 4433 20349 4445 20383
rect 4479 20380 4491 20383
rect 5074 20380 5080 20392
rect 4479 20352 5080 20380
rect 4479 20349 4491 20352
rect 4433 20343 4491 20349
rect 2222 20272 2228 20324
rect 2280 20312 2286 20324
rect 3068 20312 3096 20343
rect 5074 20340 5080 20352
rect 5132 20340 5138 20392
rect 6086 20380 6092 20392
rect 6047 20352 6092 20380
rect 6086 20340 6092 20352
rect 6144 20340 6150 20392
rect 6362 20380 6368 20392
rect 6323 20352 6368 20380
rect 6362 20340 6368 20352
rect 6420 20340 6426 20392
rect 7466 20340 7472 20392
rect 7524 20380 7530 20392
rect 7745 20383 7803 20389
rect 7745 20380 7757 20383
rect 7524 20352 7757 20380
rect 7524 20340 7530 20352
rect 7745 20349 7757 20352
rect 7791 20349 7803 20383
rect 7745 20343 7803 20349
rect 8478 20340 8484 20392
rect 8536 20380 8542 20392
rect 9953 20383 10011 20389
rect 9953 20380 9965 20383
rect 8536 20352 9965 20380
rect 8536 20340 8542 20352
rect 9953 20349 9965 20352
rect 9999 20349 10011 20383
rect 9953 20343 10011 20349
rect 10042 20340 10048 20392
rect 10100 20380 10106 20392
rect 10209 20383 10267 20389
rect 10209 20380 10221 20383
rect 10100 20352 10221 20380
rect 10100 20340 10106 20352
rect 10209 20349 10221 20352
rect 10255 20349 10267 20383
rect 10209 20343 10267 20349
rect 12342 20340 12348 20392
rect 12400 20389 12406 20392
rect 12549 20389 12577 20420
rect 12400 20383 12449 20389
rect 12400 20349 12403 20383
rect 12437 20349 12449 20383
rect 12400 20343 12449 20349
rect 12510 20383 12577 20389
rect 12510 20349 12522 20383
rect 12556 20352 12577 20383
rect 12621 20383 12679 20389
rect 12556 20349 12568 20352
rect 12510 20343 12568 20349
rect 12621 20349 12633 20383
rect 12667 20380 12679 20383
rect 12710 20380 12716 20392
rect 12667 20352 12716 20380
rect 12667 20349 12679 20352
rect 12621 20343 12679 20349
rect 12400 20340 12406 20343
rect 12710 20340 12716 20352
rect 12768 20340 12774 20392
rect 12805 20383 12863 20389
rect 12805 20349 12817 20383
rect 12851 20380 12863 20383
rect 12894 20380 12900 20392
rect 12851 20352 12900 20380
rect 12851 20349 12863 20352
rect 12805 20343 12863 20349
rect 12894 20340 12900 20352
rect 12952 20340 12958 20392
rect 13354 20340 13360 20392
rect 13412 20380 13418 20392
rect 13449 20383 13507 20389
rect 13449 20380 13461 20383
rect 13412 20352 13461 20380
rect 13412 20340 13418 20352
rect 13449 20349 13461 20352
rect 13495 20349 13507 20383
rect 15010 20380 15016 20392
rect 14971 20352 15016 20380
rect 13449 20343 13507 20349
rect 15010 20340 15016 20352
rect 15068 20340 15074 20392
rect 15120 20389 15148 20420
rect 15105 20383 15163 20389
rect 15105 20349 15117 20383
rect 15151 20349 15163 20383
rect 15105 20343 15163 20349
rect 15194 20340 15200 20392
rect 15252 20380 15258 20392
rect 15396 20389 15424 20420
rect 15746 20408 15752 20460
rect 15804 20448 15810 20460
rect 16040 20448 16068 20476
rect 15804 20420 16146 20448
rect 15804 20408 15810 20420
rect 21358 20408 21364 20460
rect 21416 20448 21422 20460
rect 21545 20451 21603 20457
rect 21545 20448 21557 20451
rect 21416 20420 21557 20448
rect 21416 20408 21422 20420
rect 21545 20417 21557 20420
rect 21591 20417 21603 20451
rect 21545 20411 21603 20417
rect 15381 20383 15439 20389
rect 15252 20352 15297 20380
rect 15252 20340 15258 20352
rect 15381 20349 15393 20383
rect 15427 20349 15439 20383
rect 15381 20343 15439 20349
rect 16022 20340 16028 20392
rect 16080 20380 16086 20392
rect 16666 20380 16672 20392
rect 16080 20352 16672 20380
rect 16080 20340 16086 20352
rect 16666 20340 16672 20352
rect 16724 20340 16730 20392
rect 17037 20383 17095 20389
rect 17037 20349 17049 20383
rect 17083 20380 17095 20383
rect 19058 20380 19064 20392
rect 17083 20352 19064 20380
rect 17083 20349 17095 20352
rect 17037 20343 17095 20349
rect 19058 20340 19064 20352
rect 19116 20340 19122 20392
rect 20990 20380 20996 20392
rect 20951 20352 20996 20380
rect 20990 20340 20996 20352
rect 21048 20340 21054 20392
rect 21634 20380 21640 20392
rect 21595 20352 21640 20380
rect 21634 20340 21640 20352
rect 21692 20340 21698 20392
rect 22066 20380 22094 20488
rect 22370 20476 22376 20528
rect 22428 20516 22434 20528
rect 22465 20519 22523 20525
rect 22465 20516 22477 20519
rect 22428 20488 22477 20516
rect 22428 20476 22434 20488
rect 22465 20485 22477 20488
rect 22511 20516 22523 20519
rect 23290 20516 23296 20528
rect 22511 20488 23296 20516
rect 22511 20485 22523 20488
rect 22465 20479 22523 20485
rect 23290 20476 23296 20488
rect 23348 20476 23354 20528
rect 22278 20408 22284 20460
rect 22336 20448 22342 20460
rect 22336 20420 27292 20448
rect 22336 20408 22342 20420
rect 27264 20389 27292 20420
rect 22649 20383 22707 20389
rect 22649 20380 22661 20383
rect 22066 20352 22661 20380
rect 22649 20349 22661 20352
rect 22695 20349 22707 20383
rect 27249 20383 27307 20389
rect 22649 20343 22707 20349
rect 25056 20352 26832 20380
rect 2280 20284 3096 20312
rect 2280 20272 2286 20284
rect 5166 20272 5172 20324
rect 5224 20312 5230 20324
rect 16574 20312 16580 20324
rect 5224 20284 16580 20312
rect 5224 20272 5230 20284
rect 16574 20272 16580 20284
rect 16632 20272 16638 20324
rect 20070 20272 20076 20324
rect 20128 20312 20134 20324
rect 25056 20312 25084 20352
rect 20128 20284 25084 20312
rect 25777 20315 25835 20321
rect 20128 20272 20134 20284
rect 25777 20281 25789 20315
rect 25823 20281 25835 20315
rect 25958 20312 25964 20324
rect 25919 20284 25964 20312
rect 25777 20275 25835 20281
rect 6733 20247 6791 20253
rect 6733 20213 6745 20247
rect 6779 20244 6791 20247
rect 7466 20244 7472 20256
rect 6779 20216 7472 20244
rect 6779 20213 6791 20216
rect 6733 20207 6791 20213
rect 7466 20204 7472 20216
rect 7524 20204 7530 20256
rect 12158 20244 12164 20256
rect 12119 20216 12164 20244
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 14734 20244 14740 20256
rect 14695 20216 14740 20244
rect 14734 20204 14740 20216
rect 14792 20204 14798 20256
rect 16114 20204 16120 20256
rect 16172 20244 16178 20256
rect 16301 20247 16359 20253
rect 16301 20244 16313 20247
rect 16172 20216 16313 20244
rect 16172 20204 16178 20216
rect 16301 20213 16313 20216
rect 16347 20213 16359 20247
rect 17402 20244 17408 20256
rect 17363 20216 17408 20244
rect 16301 20207 16359 20213
rect 17402 20204 17408 20216
rect 17460 20204 17466 20256
rect 17589 20247 17647 20253
rect 17589 20213 17601 20247
rect 17635 20244 17647 20247
rect 17954 20244 17960 20256
rect 17635 20216 17960 20244
rect 17635 20213 17647 20216
rect 17589 20207 17647 20213
rect 17954 20204 17960 20216
rect 18012 20204 18018 20256
rect 25792 20244 25820 20275
rect 25958 20272 25964 20284
rect 26016 20272 26022 20324
rect 26234 20272 26240 20324
rect 26292 20312 26298 20324
rect 26513 20315 26571 20321
rect 26513 20312 26525 20315
rect 26292 20284 26525 20312
rect 26292 20272 26298 20284
rect 26513 20281 26525 20284
rect 26559 20281 26571 20315
rect 26694 20312 26700 20324
rect 26655 20284 26700 20312
rect 26513 20275 26571 20281
rect 26694 20272 26700 20284
rect 26752 20272 26758 20324
rect 26804 20312 26832 20352
rect 27249 20349 27261 20383
rect 27295 20349 27307 20383
rect 27249 20343 27307 20349
rect 27985 20315 28043 20321
rect 27985 20312 27997 20315
rect 26804 20284 27997 20312
rect 27985 20281 27997 20284
rect 28031 20281 28043 20315
rect 28166 20312 28172 20324
rect 28127 20284 28172 20312
rect 27985 20275 28043 20281
rect 28166 20272 28172 20284
rect 28224 20272 28230 20324
rect 28074 20244 28080 20256
rect 25792 20216 28080 20244
rect 28074 20204 28080 20216
rect 28132 20204 28138 20256
rect 1104 20154 28888 20176
rect 1104 20102 10246 20154
rect 10298 20102 10310 20154
rect 10362 20102 10374 20154
rect 10426 20102 10438 20154
rect 10490 20102 19510 20154
rect 19562 20102 19574 20154
rect 19626 20102 19638 20154
rect 19690 20102 19702 20154
rect 19754 20102 28888 20154
rect 1104 20080 28888 20102
rect 2501 20043 2559 20049
rect 2501 20009 2513 20043
rect 2547 20040 2559 20043
rect 4154 20040 4160 20052
rect 2547 20012 4160 20040
rect 2547 20009 2559 20012
rect 2501 20003 2559 20009
rect 4154 20000 4160 20012
rect 4212 20000 4218 20052
rect 4338 20000 4344 20052
rect 4396 20040 4402 20052
rect 4525 20043 4583 20049
rect 4525 20040 4537 20043
rect 4396 20012 4537 20040
rect 4396 20000 4402 20012
rect 4525 20009 4537 20012
rect 4571 20009 4583 20043
rect 4525 20003 4583 20009
rect 9950 20000 9956 20052
rect 10008 20040 10014 20052
rect 10045 20043 10103 20049
rect 10045 20040 10057 20043
rect 10008 20012 10057 20040
rect 10008 20000 10014 20012
rect 10045 20009 10057 20012
rect 10091 20009 10103 20043
rect 10045 20003 10103 20009
rect 17313 20043 17371 20049
rect 17313 20009 17325 20043
rect 17359 20040 17371 20043
rect 20070 20040 20076 20052
rect 17359 20012 20076 20040
rect 17359 20009 17371 20012
rect 17313 20003 17371 20009
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 4617 19975 4675 19981
rect 4617 19941 4629 19975
rect 4663 19972 4675 19975
rect 4706 19972 4712 19984
rect 4663 19944 4712 19972
rect 4663 19941 4675 19944
rect 4617 19935 4675 19941
rect 4706 19932 4712 19944
rect 4764 19932 4770 19984
rect 7374 19972 7380 19984
rect 7300 19944 7380 19972
rect 1854 19904 1860 19916
rect 1815 19876 1860 19904
rect 1854 19864 1860 19876
rect 1912 19864 1918 19916
rect 2685 19907 2743 19913
rect 2685 19873 2697 19907
rect 2731 19904 2743 19907
rect 2774 19904 2780 19916
rect 2731 19876 2780 19904
rect 2731 19873 2743 19876
rect 2685 19867 2743 19873
rect 2774 19864 2780 19876
rect 2832 19864 2838 19916
rect 3142 19904 3148 19916
rect 3103 19876 3148 19904
rect 3142 19864 3148 19876
rect 3200 19864 3206 19916
rect 7300 19913 7328 19944
rect 7374 19932 7380 19944
rect 7432 19932 7438 19984
rect 8205 19975 8263 19981
rect 8205 19941 8217 19975
rect 8251 19972 8263 19975
rect 8294 19972 8300 19984
rect 8251 19944 8300 19972
rect 8251 19941 8263 19944
rect 8205 19935 8263 19941
rect 8294 19932 8300 19944
rect 8352 19932 8358 19984
rect 8662 19932 8668 19984
rect 8720 19972 8726 19984
rect 9030 19972 9036 19984
rect 8720 19944 9036 19972
rect 8720 19932 8726 19944
rect 9030 19932 9036 19944
rect 9088 19932 9094 19984
rect 9309 19975 9367 19981
rect 9309 19941 9321 19975
rect 9355 19972 9367 19975
rect 9490 19972 9496 19984
rect 9355 19944 9496 19972
rect 9355 19941 9367 19944
rect 9309 19935 9367 19941
rect 9490 19932 9496 19944
rect 9548 19932 9554 19984
rect 9858 19932 9864 19984
rect 9916 19972 9922 19984
rect 9916 19944 10180 19972
rect 9916 19932 9922 19944
rect 7285 19907 7343 19913
rect 7285 19873 7297 19907
rect 7331 19873 7343 19907
rect 7466 19904 7472 19916
rect 7427 19876 7472 19904
rect 7285 19867 7343 19873
rect 7466 19864 7472 19876
rect 7524 19864 7530 19916
rect 8110 19904 8116 19916
rect 8071 19876 8116 19904
rect 8110 19864 8116 19876
rect 8168 19864 8174 19916
rect 9122 19904 9128 19916
rect 9083 19876 9128 19904
rect 9122 19864 9128 19876
rect 9180 19864 9186 19916
rect 9214 19864 9220 19916
rect 9272 19904 9278 19916
rect 9401 19907 9459 19913
rect 9401 19904 9413 19907
rect 9272 19876 9413 19904
rect 9272 19864 9278 19876
rect 9401 19873 9413 19876
rect 9447 19873 9459 19907
rect 9401 19867 9459 19873
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 10152 19913 10180 19944
rect 11238 19932 11244 19984
rect 11296 19972 11302 19984
rect 15010 19972 15016 19984
rect 11296 19944 15016 19972
rect 11296 19932 11302 19944
rect 15010 19932 15016 19944
rect 15068 19972 15074 19984
rect 16114 19972 16120 19984
rect 15068 19944 16120 19972
rect 15068 19932 15074 19944
rect 16114 19932 16120 19944
rect 16172 19932 16178 19984
rect 16574 19932 16580 19984
rect 16632 19972 16638 19984
rect 27985 19975 28043 19981
rect 27985 19972 27997 19975
rect 16632 19944 27997 19972
rect 16632 19932 16638 19944
rect 27985 19941 27997 19944
rect 28031 19941 28043 19975
rect 27985 19935 28043 19941
rect 9953 19907 10011 19913
rect 9953 19904 9965 19907
rect 9732 19876 9965 19904
rect 9732 19864 9738 19876
rect 9953 19873 9965 19876
rect 9999 19873 10011 19907
rect 9953 19867 10011 19873
rect 10137 19907 10195 19913
rect 10137 19873 10149 19907
rect 10183 19873 10195 19907
rect 17586 19904 17592 19916
rect 17547 19876 17592 19904
rect 10137 19867 10195 19873
rect 3878 19796 3884 19848
rect 3936 19836 3942 19848
rect 4709 19839 4767 19845
rect 4709 19836 4721 19839
rect 3936 19808 4721 19836
rect 3936 19796 3942 19808
rect 4709 19805 4721 19808
rect 4755 19805 4767 19839
rect 9968 19836 9996 19867
rect 17586 19864 17592 19876
rect 17644 19864 17650 19916
rect 18322 19864 18328 19916
rect 18380 19904 18386 19916
rect 18857 19907 18915 19913
rect 18857 19904 18869 19907
rect 18380 19876 18869 19904
rect 18380 19864 18386 19876
rect 18857 19873 18869 19876
rect 18903 19873 18915 19907
rect 18857 19867 18915 19873
rect 24949 19907 25007 19913
rect 24949 19873 24961 19907
rect 24995 19904 25007 19907
rect 25222 19904 25228 19916
rect 24995 19876 25228 19904
rect 24995 19873 25007 19876
rect 24949 19867 25007 19873
rect 25222 19864 25228 19876
rect 25280 19864 25286 19916
rect 25682 19904 25688 19916
rect 25643 19876 25688 19904
rect 25682 19864 25688 19876
rect 25740 19864 25746 19916
rect 26510 19904 26516 19916
rect 26471 19876 26516 19904
rect 26510 19864 26516 19876
rect 26568 19904 26574 19916
rect 26786 19904 26792 19916
rect 26568 19876 26792 19904
rect 26568 19864 26574 19876
rect 26786 19864 26792 19876
rect 26844 19864 26850 19916
rect 11146 19836 11152 19848
rect 4709 19799 4767 19805
rect 6196 19808 8984 19836
rect 9968 19808 11152 19836
rect 2041 19771 2099 19777
rect 2041 19737 2053 19771
rect 2087 19768 2099 19771
rect 2406 19768 2412 19780
rect 2087 19740 2412 19768
rect 2087 19737 2099 19740
rect 2041 19731 2099 19737
rect 2406 19728 2412 19740
rect 2464 19728 2470 19780
rect 3326 19768 3332 19780
rect 3239 19740 3332 19768
rect 3326 19728 3332 19740
rect 3384 19768 3390 19780
rect 6196 19768 6224 19808
rect 3384 19740 6224 19768
rect 3384 19728 3390 19740
rect 6362 19728 6368 19780
rect 6420 19768 6426 19780
rect 8849 19771 8907 19777
rect 8849 19768 8861 19771
rect 6420 19740 8861 19768
rect 6420 19728 6426 19740
rect 8849 19737 8861 19740
rect 8895 19737 8907 19771
rect 8956 19768 8984 19808
rect 11146 19796 11152 19808
rect 11204 19796 11210 19848
rect 12342 19796 12348 19848
rect 12400 19836 12406 19848
rect 12526 19836 12532 19848
rect 12400 19808 12532 19836
rect 12400 19796 12406 19808
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 16574 19796 16580 19848
rect 16632 19836 16638 19848
rect 17678 19836 17684 19848
rect 16632 19808 17540 19836
rect 17639 19808 17684 19836
rect 16632 19796 16638 19808
rect 17402 19768 17408 19780
rect 8956 19740 17408 19768
rect 8849 19731 8907 19737
rect 17402 19728 17408 19740
rect 17460 19728 17466 19780
rect 17512 19768 17540 19808
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 17862 19796 17868 19848
rect 17920 19836 17926 19848
rect 18601 19839 18659 19845
rect 18601 19836 18613 19839
rect 17920 19808 18613 19836
rect 17920 19796 17926 19808
rect 18601 19805 18613 19808
rect 18647 19805 18659 19839
rect 18601 19799 18659 19805
rect 20530 19796 20536 19848
rect 20588 19836 20594 19848
rect 23382 19836 23388 19848
rect 20588 19808 23388 19836
rect 20588 19796 20594 19808
rect 23382 19796 23388 19808
rect 23440 19796 23446 19848
rect 26605 19839 26663 19845
rect 26605 19805 26617 19839
rect 26651 19805 26663 19839
rect 26605 19799 26663 19805
rect 17880 19768 17908 19796
rect 25866 19768 25872 19780
rect 17512 19740 17908 19768
rect 25827 19740 25872 19768
rect 25866 19728 25872 19740
rect 25924 19728 25930 19780
rect 26620 19768 26648 19799
rect 26786 19768 26792 19780
rect 26620 19740 26792 19768
rect 26786 19728 26792 19740
rect 26844 19768 26850 19780
rect 27154 19768 27160 19780
rect 26844 19740 27160 19768
rect 26844 19728 26850 19740
rect 27154 19728 27160 19740
rect 27212 19728 27218 19780
rect 28166 19768 28172 19780
rect 28127 19740 28172 19768
rect 28166 19728 28172 19740
rect 28224 19728 28230 19780
rect 4154 19700 4160 19712
rect 4115 19672 4160 19700
rect 4154 19660 4160 19672
rect 4212 19660 4218 19712
rect 6178 19660 6184 19712
rect 6236 19700 6242 19712
rect 11238 19700 11244 19712
rect 6236 19672 11244 19700
rect 6236 19660 6242 19672
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 11606 19660 11612 19712
rect 11664 19700 11670 19712
rect 17313 19703 17371 19709
rect 17313 19700 17325 19703
rect 11664 19672 17325 19700
rect 11664 19660 11670 19672
rect 17313 19669 17325 19672
rect 17359 19669 17371 19703
rect 17313 19663 17371 19669
rect 17862 19660 17868 19712
rect 17920 19700 17926 19712
rect 17957 19703 18015 19709
rect 17957 19700 17969 19703
rect 17920 19672 17969 19700
rect 17920 19660 17926 19672
rect 17957 19669 17969 19672
rect 18003 19669 18015 19703
rect 19978 19700 19984 19712
rect 19939 19672 19984 19700
rect 17957 19663 18015 19669
rect 19978 19660 19984 19672
rect 20036 19660 20042 19712
rect 25041 19703 25099 19709
rect 25041 19669 25053 19703
rect 25087 19700 25099 19703
rect 25406 19700 25412 19712
rect 25087 19672 25412 19700
rect 25087 19669 25099 19672
rect 25041 19663 25099 19669
rect 25406 19660 25412 19672
rect 25464 19700 25470 19712
rect 25774 19700 25780 19712
rect 25464 19672 25780 19700
rect 25464 19660 25470 19672
rect 25774 19660 25780 19672
rect 25832 19660 25838 19712
rect 26881 19703 26939 19709
rect 26881 19669 26893 19703
rect 26927 19700 26939 19703
rect 27798 19700 27804 19712
rect 26927 19672 27804 19700
rect 26927 19669 26939 19672
rect 26881 19663 26939 19669
rect 27798 19660 27804 19672
rect 27856 19660 27862 19712
rect 1104 19610 28888 19632
rect 1104 19558 5614 19610
rect 5666 19558 5678 19610
rect 5730 19558 5742 19610
rect 5794 19558 5806 19610
rect 5858 19558 14878 19610
rect 14930 19558 14942 19610
rect 14994 19558 15006 19610
rect 15058 19558 15070 19610
rect 15122 19558 24142 19610
rect 24194 19558 24206 19610
rect 24258 19558 24270 19610
rect 24322 19558 24334 19610
rect 24386 19558 28888 19610
rect 1104 19536 28888 19558
rect 7193 19499 7251 19505
rect 7193 19465 7205 19499
rect 7239 19496 7251 19499
rect 7650 19496 7656 19508
rect 7239 19468 7656 19496
rect 7239 19465 7251 19468
rect 7193 19459 7251 19465
rect 7650 19456 7656 19468
rect 7708 19456 7714 19508
rect 9490 19496 9496 19508
rect 9451 19468 9496 19496
rect 9490 19456 9496 19468
rect 9548 19456 9554 19508
rect 10962 19456 10968 19508
rect 11020 19496 11026 19508
rect 11885 19499 11943 19505
rect 11885 19496 11897 19499
rect 11020 19468 11897 19496
rect 11020 19456 11026 19468
rect 11885 19465 11897 19468
rect 11931 19496 11943 19499
rect 13354 19496 13360 19508
rect 11931 19468 13360 19496
rect 11931 19465 11943 19468
rect 11885 19459 11943 19465
rect 13354 19456 13360 19468
rect 13412 19456 13418 19508
rect 16114 19496 16120 19508
rect 16075 19468 16120 19496
rect 16114 19456 16120 19468
rect 16172 19456 16178 19508
rect 17034 19456 17040 19508
rect 17092 19496 17098 19508
rect 18233 19499 18291 19505
rect 18233 19496 18245 19499
rect 17092 19468 18245 19496
rect 17092 19456 17098 19468
rect 18233 19465 18245 19468
rect 18279 19465 18291 19499
rect 18233 19459 18291 19465
rect 21358 19456 21364 19508
rect 21416 19496 21422 19508
rect 21453 19499 21511 19505
rect 21453 19496 21465 19499
rect 21416 19468 21465 19496
rect 21416 19456 21422 19468
rect 21453 19465 21465 19468
rect 21499 19465 21511 19499
rect 21453 19459 21511 19465
rect 28074 19456 28080 19508
rect 28132 19496 28138 19508
rect 28169 19499 28227 19505
rect 28169 19496 28181 19499
rect 28132 19468 28181 19496
rect 28132 19456 28138 19468
rect 28169 19465 28181 19468
rect 28215 19465 28227 19499
rect 28169 19459 28227 19465
rect 6086 19388 6092 19440
rect 6144 19428 6150 19440
rect 6273 19431 6331 19437
rect 6273 19428 6285 19431
rect 6144 19400 6285 19428
rect 6144 19388 6150 19400
rect 6273 19397 6285 19400
rect 6319 19397 6331 19431
rect 6273 19391 6331 19397
rect 14734 19388 14740 19440
rect 14792 19388 14798 19440
rect 21726 19428 21732 19440
rect 21560 19400 21732 19428
rect 4154 19320 4160 19372
rect 4212 19360 4218 19372
rect 4709 19363 4767 19369
rect 4709 19360 4721 19363
rect 4212 19332 4721 19360
rect 4212 19320 4218 19332
rect 4709 19329 4721 19332
rect 4755 19329 4767 19363
rect 4709 19323 4767 19329
rect 4798 19320 4804 19372
rect 4856 19360 4862 19372
rect 5997 19363 6055 19369
rect 4856 19332 4901 19360
rect 4856 19320 4862 19332
rect 5997 19329 6009 19363
rect 6043 19360 6055 19363
rect 6362 19360 6368 19372
rect 6043 19332 6368 19360
rect 6043 19329 6055 19332
rect 5997 19323 6055 19329
rect 6362 19320 6368 19332
rect 6420 19320 6426 19372
rect 10134 19360 10140 19372
rect 6840 19332 7972 19360
rect 10095 19332 10140 19360
rect 2501 19295 2559 19301
rect 2501 19261 2513 19295
rect 2547 19292 2559 19295
rect 2866 19292 2872 19304
rect 2547 19264 2872 19292
rect 2547 19261 2559 19264
rect 2501 19255 2559 19261
rect 2866 19252 2872 19264
rect 2924 19252 2930 19304
rect 2958 19252 2964 19304
rect 3016 19292 3022 19304
rect 3145 19295 3203 19301
rect 3145 19292 3157 19295
rect 3016 19264 3157 19292
rect 3016 19252 3022 19264
rect 3145 19261 3157 19264
rect 3191 19261 3203 19295
rect 3145 19255 3203 19261
rect 3329 19295 3387 19301
rect 3329 19261 3341 19295
rect 3375 19292 3387 19295
rect 4246 19292 4252 19304
rect 3375 19264 4252 19292
rect 3375 19261 3387 19264
rect 3329 19255 3387 19261
rect 4246 19252 4252 19264
rect 4304 19252 4310 19304
rect 5166 19252 5172 19304
rect 5224 19292 5230 19304
rect 6840 19292 6868 19332
rect 5224 19264 6868 19292
rect 6917 19295 6975 19301
rect 5224 19252 5230 19264
rect 6917 19261 6929 19295
rect 6963 19292 6975 19295
rect 7006 19292 7012 19304
rect 6963 19264 7012 19292
rect 6963 19261 6975 19264
rect 6917 19255 6975 19261
rect 7006 19252 7012 19264
rect 7064 19252 7070 19304
rect 7098 19252 7104 19304
rect 7156 19292 7162 19304
rect 7193 19295 7251 19301
rect 7193 19292 7205 19295
rect 7156 19264 7205 19292
rect 7156 19252 7162 19264
rect 7193 19261 7205 19264
rect 7239 19261 7251 19295
rect 7374 19292 7380 19304
rect 7335 19264 7380 19292
rect 7193 19255 7251 19261
rect 7374 19252 7380 19264
rect 7432 19252 7438 19304
rect 7466 19252 7472 19304
rect 7524 19292 7530 19304
rect 7837 19295 7895 19301
rect 7837 19292 7849 19295
rect 7524 19264 7849 19292
rect 7524 19252 7530 19264
rect 7837 19261 7849 19264
rect 7883 19261 7895 19295
rect 7944 19292 7972 19332
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 14752 19360 14780 19388
rect 21560 19372 21588 19400
rect 21726 19388 21732 19400
rect 21784 19428 21790 19440
rect 25406 19428 25412 19440
rect 21784 19400 22232 19428
rect 21784 19388 21790 19400
rect 15013 19363 15071 19369
rect 15013 19360 15025 19363
rect 14752 19332 15025 19360
rect 15013 19329 15025 19332
rect 15059 19329 15071 19363
rect 15013 19323 15071 19329
rect 16574 19320 16580 19372
rect 16632 19360 16638 19372
rect 21294 19363 21352 19369
rect 16632 19332 16896 19360
rect 16632 19320 16638 19332
rect 8941 19295 8999 19301
rect 7944 19264 8064 19292
rect 7837 19255 7895 19261
rect 1854 19224 1860 19236
rect 1815 19196 1860 19224
rect 1854 19184 1860 19196
rect 1912 19184 1918 19236
rect 2041 19227 2099 19233
rect 2041 19193 2053 19227
rect 2087 19224 2099 19227
rect 3237 19227 3295 19233
rect 2087 19196 3188 19224
rect 2087 19193 2099 19196
rect 2041 19187 2099 19193
rect 1578 19116 1584 19168
rect 1636 19156 1642 19168
rect 2056 19156 2084 19187
rect 2682 19156 2688 19168
rect 1636 19128 2084 19156
rect 2643 19128 2688 19156
rect 1636 19116 1642 19128
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 3160 19156 3188 19196
rect 3237 19193 3249 19227
rect 3283 19224 3295 19227
rect 4617 19227 4675 19233
rect 4617 19224 4629 19227
rect 3283 19196 4629 19224
rect 3283 19193 3295 19196
rect 3237 19187 3295 19193
rect 4617 19193 4629 19196
rect 4663 19193 4675 19227
rect 4617 19187 4675 19193
rect 4982 19184 4988 19236
rect 5040 19224 5046 19236
rect 5258 19224 5264 19236
rect 5040 19196 5264 19224
rect 5040 19184 5046 19196
rect 5258 19184 5264 19196
rect 5316 19184 5322 19236
rect 7392 19224 7420 19252
rect 7929 19227 7987 19233
rect 7929 19224 7941 19227
rect 6380 19196 7328 19224
rect 7392 19196 7941 19224
rect 4062 19156 4068 19168
rect 3160 19128 4068 19156
rect 4062 19116 4068 19128
rect 4120 19116 4126 19168
rect 4246 19156 4252 19168
rect 4207 19128 4252 19156
rect 4246 19116 4252 19128
rect 4304 19116 4310 19168
rect 4522 19116 4528 19168
rect 4580 19156 4586 19168
rect 6380 19156 6408 19196
rect 4580 19128 6408 19156
rect 6457 19159 6515 19165
rect 4580 19116 4586 19128
rect 6457 19125 6469 19159
rect 6503 19156 6515 19159
rect 6914 19156 6920 19168
rect 6503 19128 6920 19156
rect 6503 19125 6515 19128
rect 6457 19119 6515 19125
rect 6914 19116 6920 19128
rect 6972 19116 6978 19168
rect 7300 19156 7328 19196
rect 7929 19193 7941 19196
rect 7975 19193 7987 19227
rect 8036 19224 8064 19264
rect 8941 19261 8953 19295
rect 8987 19292 8999 19295
rect 11241 19295 11299 19301
rect 11241 19292 11253 19295
rect 8987 19264 11253 19292
rect 8987 19261 8999 19264
rect 8941 19255 8999 19261
rect 11241 19261 11253 19264
rect 11287 19261 11299 19295
rect 11241 19255 11299 19261
rect 12069 19295 12127 19301
rect 12069 19261 12081 19295
rect 12115 19292 12127 19295
rect 13354 19292 13360 19304
rect 12115 19264 13360 19292
rect 12115 19261 12127 19264
rect 12069 19255 12127 19261
rect 10962 19224 10968 19236
rect 8036 19196 10968 19224
rect 7929 19187 7987 19193
rect 10962 19184 10968 19196
rect 11020 19184 11026 19236
rect 11256 19224 11284 19255
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 14737 19295 14795 19301
rect 14737 19261 14749 19295
rect 14783 19292 14795 19295
rect 16592 19292 16620 19320
rect 16868 19301 16896 19332
rect 18616 19332 19472 19360
rect 14783 19264 16620 19292
rect 16853 19295 16911 19301
rect 14783 19261 14795 19264
rect 14737 19255 14795 19261
rect 16853 19261 16865 19295
rect 16899 19261 16911 19295
rect 17129 19295 17187 19301
rect 17129 19292 17141 19295
rect 16853 19255 16911 19261
rect 16960 19264 17141 19292
rect 14826 19224 14832 19236
rect 11256 19196 14832 19224
rect 14826 19184 14832 19196
rect 14884 19184 14890 19236
rect 16040 19196 16252 19224
rect 8941 19159 8999 19165
rect 8941 19156 8953 19159
rect 7300 19128 8953 19156
rect 8941 19125 8953 19128
rect 8987 19125 8999 19159
rect 9858 19156 9864 19168
rect 9819 19128 9864 19156
rect 8941 19119 8999 19125
rect 9858 19116 9864 19128
rect 9916 19116 9922 19168
rect 9950 19116 9956 19168
rect 10008 19156 10014 19168
rect 10008 19128 10053 19156
rect 10008 19116 10014 19128
rect 10870 19116 10876 19168
rect 10928 19156 10934 19168
rect 11333 19159 11391 19165
rect 11333 19156 11345 19159
rect 10928 19128 11345 19156
rect 10928 19116 10934 19128
rect 11333 19125 11345 19128
rect 11379 19125 11391 19159
rect 11333 19119 11391 19125
rect 11606 19116 11612 19168
rect 11664 19156 11670 19168
rect 16040 19156 16068 19196
rect 11664 19128 16068 19156
rect 16224 19156 16252 19196
rect 16390 19184 16396 19236
rect 16448 19224 16454 19236
rect 16960 19224 16988 19264
rect 17129 19261 17141 19264
rect 17175 19261 17187 19295
rect 17129 19255 17187 19261
rect 17218 19252 17224 19304
rect 17276 19292 17282 19304
rect 18616 19292 18644 19332
rect 17276 19264 18644 19292
rect 17276 19252 17282 19264
rect 18690 19252 18696 19304
rect 18748 19292 18754 19304
rect 19334 19292 19340 19304
rect 18748 19264 19340 19292
rect 18748 19252 18754 19264
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 19444 19292 19472 19332
rect 21294 19329 21306 19363
rect 21340 19360 21352 19363
rect 21542 19360 21548 19372
rect 21340 19332 21548 19360
rect 21340 19329 21352 19332
rect 21294 19323 21352 19329
rect 21542 19320 21548 19332
rect 21600 19320 21606 19372
rect 21910 19320 21916 19372
rect 21968 19360 21974 19372
rect 21968 19332 22140 19360
rect 21968 19320 21974 19332
rect 20530 19292 20536 19304
rect 19444 19264 20536 19292
rect 20530 19252 20536 19264
rect 20588 19252 20594 19304
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 22112 19301 22140 19332
rect 22204 19301 22232 19400
rect 23768 19400 25412 19428
rect 20809 19295 20867 19301
rect 20809 19292 20821 19295
rect 20772 19264 20821 19292
rect 20772 19252 20778 19264
rect 20809 19261 20821 19264
rect 20855 19261 20867 19295
rect 22097 19295 22155 19301
rect 20809 19255 20867 19261
rect 20916 19264 22048 19292
rect 20916 19224 20944 19264
rect 21913 19227 21971 19233
rect 21913 19224 21925 19227
rect 16448 19196 16988 19224
rect 17788 19196 20944 19224
rect 21100 19196 21925 19224
rect 16448 19184 16454 19196
rect 17788 19156 17816 19196
rect 16224 19128 17816 19156
rect 11664 19116 11670 19128
rect 19058 19116 19064 19168
rect 19116 19156 19122 19168
rect 20622 19156 20628 19168
rect 19116 19128 20628 19156
rect 19116 19116 19122 19128
rect 20622 19116 20628 19128
rect 20680 19116 20686 19168
rect 20898 19116 20904 19168
rect 20956 19156 20962 19168
rect 21100 19165 21128 19196
rect 21913 19193 21925 19196
rect 21959 19193 21971 19227
rect 22020 19224 22048 19264
rect 22097 19261 22109 19295
rect 22143 19261 22155 19295
rect 22097 19255 22155 19261
rect 22189 19295 22247 19301
rect 22189 19261 22201 19295
rect 22235 19261 22247 19295
rect 22189 19255 22247 19261
rect 23474 19252 23480 19304
rect 23532 19292 23538 19304
rect 23768 19292 23796 19400
rect 25406 19388 25412 19400
rect 25464 19428 25470 19440
rect 26234 19428 26240 19440
rect 25464 19400 26240 19428
rect 25464 19388 25470 19400
rect 26234 19388 26240 19400
rect 26292 19388 26298 19440
rect 23845 19363 23903 19369
rect 23845 19329 23857 19363
rect 23891 19360 23903 19363
rect 24305 19363 24363 19369
rect 23891 19332 24072 19360
rect 23891 19329 23903 19332
rect 23845 19323 23903 19329
rect 24044 19304 24072 19332
rect 24305 19329 24317 19363
rect 24351 19329 24363 19363
rect 25774 19360 25780 19372
rect 25735 19332 25780 19360
rect 24305 19323 24363 19329
rect 23934 19292 23940 19304
rect 23532 19264 23796 19292
rect 23895 19264 23940 19292
rect 23532 19252 23538 19264
rect 23934 19252 23940 19264
rect 23992 19252 23998 19304
rect 24026 19252 24032 19304
rect 24084 19252 24090 19304
rect 24320 19292 24348 19323
rect 25774 19320 25780 19332
rect 25832 19320 25838 19372
rect 25593 19295 25651 19301
rect 25593 19292 25605 19295
rect 24320 19264 25605 19292
rect 25593 19261 25605 19264
rect 25639 19261 25651 19295
rect 25593 19255 25651 19261
rect 26050 19252 26056 19304
rect 26108 19292 26114 19304
rect 26789 19295 26847 19301
rect 26789 19292 26801 19295
rect 26108 19264 26801 19292
rect 26108 19252 26114 19264
rect 26789 19261 26801 19264
rect 26835 19261 26847 19295
rect 26789 19255 26847 19261
rect 23842 19224 23848 19236
rect 22020 19196 23848 19224
rect 21913 19187 21971 19193
rect 23842 19184 23848 19196
rect 23900 19184 23906 19236
rect 26326 19224 26332 19236
rect 23952 19196 26332 19224
rect 21085 19159 21143 19165
rect 21085 19156 21097 19159
rect 20956 19128 21097 19156
rect 20956 19116 20962 19128
rect 21085 19125 21097 19128
rect 21131 19125 21143 19159
rect 21085 19119 21143 19125
rect 21174 19116 21180 19168
rect 21232 19156 21238 19168
rect 21232 19128 21277 19156
rect 21232 19116 21238 19128
rect 21542 19116 21548 19168
rect 21600 19156 21606 19168
rect 22011 19159 22069 19165
rect 22011 19156 22023 19159
rect 21600 19128 22023 19156
rect 21600 19116 21606 19128
rect 22011 19125 22023 19128
rect 22057 19125 22069 19159
rect 22011 19119 22069 19125
rect 23014 19116 23020 19168
rect 23072 19156 23078 19168
rect 23952 19156 23980 19196
rect 26326 19184 26332 19196
rect 26384 19184 26390 19236
rect 27056 19227 27114 19233
rect 27056 19193 27068 19227
rect 27102 19224 27114 19227
rect 27430 19224 27436 19236
rect 27102 19196 27436 19224
rect 27102 19193 27114 19196
rect 27056 19187 27114 19193
rect 27430 19184 27436 19196
rect 27488 19184 27494 19236
rect 23072 19128 23980 19156
rect 25225 19159 25283 19165
rect 23072 19116 23078 19128
rect 25225 19125 25237 19159
rect 25271 19156 25283 19159
rect 25314 19156 25320 19168
rect 25271 19128 25320 19156
rect 25271 19125 25283 19128
rect 25225 19119 25283 19125
rect 25314 19116 25320 19128
rect 25372 19116 25378 19168
rect 25682 19156 25688 19168
rect 25595 19128 25688 19156
rect 25682 19116 25688 19128
rect 25740 19156 25746 19168
rect 26142 19156 26148 19168
rect 25740 19128 26148 19156
rect 25740 19116 25746 19128
rect 26142 19116 26148 19128
rect 26200 19116 26206 19168
rect 1104 19066 28888 19088
rect 1104 19014 10246 19066
rect 10298 19014 10310 19066
rect 10362 19014 10374 19066
rect 10426 19014 10438 19066
rect 10490 19014 19510 19066
rect 19562 19014 19574 19066
rect 19626 19014 19638 19066
rect 19690 19014 19702 19066
rect 19754 19014 28888 19066
rect 1104 18992 28888 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 2590 18952 2596 18964
rect 1688 18924 2596 18952
rect 1688 18816 1716 18924
rect 2590 18912 2596 18924
rect 2648 18912 2654 18964
rect 2774 18912 2780 18964
rect 2832 18952 2838 18964
rect 2869 18955 2927 18961
rect 2869 18952 2881 18955
rect 2832 18924 2881 18952
rect 2832 18912 2838 18924
rect 2869 18921 2881 18924
rect 2915 18921 2927 18955
rect 2869 18915 2927 18921
rect 3605 18955 3663 18961
rect 3605 18921 3617 18955
rect 3651 18952 3663 18955
rect 5445 18955 5503 18961
rect 3651 18924 4660 18952
rect 3651 18921 3663 18924
rect 3605 18915 3663 18921
rect 1762 18844 1768 18896
rect 1820 18884 1826 18896
rect 2685 18887 2743 18893
rect 2685 18884 2697 18887
rect 1820 18856 2697 18884
rect 1820 18844 1826 18856
rect 2685 18853 2697 18856
rect 2731 18853 2743 18887
rect 4341 18887 4399 18893
rect 4341 18884 4353 18887
rect 2685 18847 2743 18853
rect 3252 18856 4353 18884
rect 1857 18819 1915 18825
rect 1857 18816 1869 18819
rect 1688 18788 1869 18816
rect 1857 18785 1869 18788
rect 1903 18785 1915 18819
rect 1857 18779 1915 18785
rect 1949 18819 2007 18825
rect 1949 18785 1961 18819
rect 1995 18816 2007 18819
rect 2038 18816 2044 18828
rect 1995 18788 2044 18816
rect 1995 18785 2007 18788
rect 1949 18779 2007 18785
rect 2038 18776 2044 18788
rect 2096 18776 2102 18828
rect 2317 18819 2375 18825
rect 2317 18785 2329 18819
rect 2363 18816 2375 18819
rect 2406 18816 2412 18828
rect 2363 18788 2412 18816
rect 2363 18785 2375 18788
rect 2317 18779 2375 18785
rect 2406 18776 2412 18788
rect 2464 18816 2470 18828
rect 3252 18816 3280 18856
rect 4341 18853 4353 18856
rect 4387 18884 4399 18887
rect 4522 18884 4528 18896
rect 4387 18856 4528 18884
rect 4387 18853 4399 18856
rect 4341 18847 4399 18853
rect 4522 18844 4528 18856
rect 4580 18844 4586 18896
rect 4632 18893 4660 18924
rect 5000 18924 5304 18952
rect 4617 18887 4675 18893
rect 4617 18853 4629 18887
rect 4663 18884 4675 18887
rect 5000 18884 5028 18924
rect 4663 18856 5028 18884
rect 5077 18887 5135 18893
rect 4663 18853 4675 18856
rect 4617 18847 4675 18853
rect 5077 18853 5089 18887
rect 5123 18884 5135 18887
rect 5166 18884 5172 18896
rect 5123 18856 5172 18884
rect 5123 18853 5135 18856
rect 5077 18847 5135 18853
rect 5166 18844 5172 18856
rect 5224 18844 5230 18896
rect 5276 18884 5304 18924
rect 5445 18921 5457 18955
rect 5491 18952 5503 18955
rect 5534 18952 5540 18964
rect 5491 18924 5540 18952
rect 5491 18921 5503 18924
rect 5445 18915 5503 18921
rect 5534 18912 5540 18924
rect 5592 18912 5598 18964
rect 5629 18955 5687 18961
rect 5629 18921 5641 18955
rect 5675 18952 5687 18955
rect 6086 18952 6092 18964
rect 5675 18924 6092 18952
rect 5675 18921 5687 18924
rect 5629 18915 5687 18921
rect 6086 18912 6092 18924
rect 6144 18912 6150 18964
rect 6638 18912 6644 18964
rect 6696 18952 6702 18964
rect 6917 18955 6975 18961
rect 6917 18952 6929 18955
rect 6696 18924 6929 18952
rect 6696 18912 6702 18924
rect 6917 18921 6929 18924
rect 6963 18921 6975 18955
rect 6917 18915 6975 18921
rect 8113 18955 8171 18961
rect 8113 18921 8125 18955
rect 8159 18952 8171 18955
rect 9122 18952 9128 18964
rect 8159 18924 9128 18952
rect 8159 18921 8171 18924
rect 8113 18915 8171 18921
rect 5276 18856 6040 18884
rect 3418 18816 3424 18828
rect 2464 18788 3280 18816
rect 3379 18788 3424 18816
rect 2464 18776 2470 18788
rect 3418 18776 3424 18788
rect 3476 18776 3482 18828
rect 4709 18819 4767 18825
rect 4709 18785 4721 18819
rect 4755 18816 4767 18819
rect 4755 18788 5948 18816
rect 4755 18785 4767 18788
rect 4709 18779 4767 18785
rect 1400 18760 1452 18766
rect 5166 18708 5172 18760
rect 5224 18708 5230 18760
rect 1400 18702 1452 18708
rect 5920 18612 5948 18788
rect 6012 18680 6040 18856
rect 6104 18816 6132 18912
rect 6932 18884 6960 18915
rect 9122 18912 9128 18924
rect 9180 18912 9186 18964
rect 9766 18912 9772 18964
rect 9824 18912 9830 18964
rect 9861 18955 9919 18961
rect 9861 18921 9873 18955
rect 9907 18952 9919 18955
rect 9950 18952 9956 18964
rect 9907 18924 9956 18952
rect 9907 18921 9919 18924
rect 9861 18915 9919 18921
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 10870 18952 10876 18964
rect 10831 18924 10876 18952
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 12526 18912 12532 18964
rect 12584 18952 12590 18964
rect 13633 18955 13691 18961
rect 13633 18952 13645 18955
rect 12584 18924 13645 18952
rect 12584 18912 12590 18924
rect 13633 18921 13645 18924
rect 13679 18921 13691 18955
rect 13633 18915 13691 18921
rect 13906 18912 13912 18964
rect 13964 18952 13970 18964
rect 14090 18952 14096 18964
rect 13964 18924 14096 18952
rect 13964 18912 13970 18924
rect 14090 18912 14096 18924
rect 14148 18952 14154 18964
rect 14642 18952 14648 18964
rect 14148 18924 14648 18952
rect 14148 18912 14154 18924
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 14826 18912 14832 18964
rect 14884 18952 14890 18964
rect 26513 18955 26571 18961
rect 26513 18952 26525 18955
rect 14884 18924 26525 18952
rect 14884 18912 14890 18924
rect 26513 18921 26525 18924
rect 26559 18921 26571 18955
rect 26513 18915 26571 18921
rect 9033 18887 9091 18893
rect 9033 18884 9045 18887
rect 6932 18856 9045 18884
rect 8128 18825 8156 18856
rect 9033 18853 9045 18856
rect 9079 18853 9091 18887
rect 9784 18884 9812 18912
rect 9033 18847 9091 18853
rect 9140 18856 9812 18884
rect 9968 18884 9996 18912
rect 10781 18887 10839 18893
rect 10781 18884 10793 18887
rect 9968 18856 10793 18884
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 6104 18788 6837 18816
rect 6825 18785 6837 18788
rect 6871 18785 6883 18819
rect 6825 18779 6883 18785
rect 7929 18819 7987 18825
rect 7929 18785 7941 18819
rect 7975 18785 7987 18819
rect 7929 18779 7987 18785
rect 8113 18819 8171 18825
rect 8113 18785 8125 18819
rect 8159 18785 8171 18819
rect 8938 18816 8944 18828
rect 8899 18788 8944 18816
rect 8113 18779 8171 18785
rect 7944 18748 7972 18779
rect 8938 18776 8944 18788
rect 8996 18776 9002 18828
rect 9140 18816 9168 18856
rect 10781 18853 10793 18856
rect 10827 18853 10839 18887
rect 10781 18847 10839 18853
rect 11790 18844 11796 18896
rect 11848 18884 11854 18896
rect 12342 18884 12348 18896
rect 11848 18856 12348 18884
rect 11848 18844 11854 18856
rect 12342 18844 12348 18856
rect 12400 18844 12406 18896
rect 14182 18844 14188 18896
rect 14240 18884 14246 18896
rect 14921 18887 14979 18893
rect 14921 18884 14933 18887
rect 14240 18856 14933 18884
rect 14240 18844 14246 18856
rect 14921 18853 14933 18856
rect 14967 18853 14979 18887
rect 17954 18884 17960 18896
rect 14921 18847 14979 18853
rect 17512 18856 17960 18884
rect 9048 18788 9168 18816
rect 9048 18760 9076 18788
rect 9490 18776 9496 18828
rect 9548 18816 9554 18828
rect 9769 18819 9827 18825
rect 9769 18816 9781 18819
rect 9548 18788 9781 18816
rect 9548 18776 9554 18788
rect 9769 18785 9781 18788
rect 9815 18816 9827 18819
rect 12066 18816 12072 18828
rect 9815 18788 12072 18816
rect 9815 18785 9827 18788
rect 9769 18779 9827 18785
rect 12066 18776 12072 18788
rect 12124 18776 12130 18828
rect 12158 18776 12164 18828
rect 12216 18816 12222 18828
rect 12529 18819 12587 18825
rect 12529 18816 12541 18819
rect 12216 18788 12541 18816
rect 12216 18776 12222 18788
rect 12529 18785 12541 18788
rect 12575 18785 12587 18819
rect 12529 18779 12587 18785
rect 13906 18776 13912 18828
rect 13964 18816 13970 18828
rect 14737 18819 14795 18825
rect 14737 18816 14749 18819
rect 13964 18788 14749 18816
rect 13964 18776 13970 18788
rect 14737 18785 14749 18788
rect 14783 18785 14795 18819
rect 14737 18779 14795 18785
rect 15838 18776 15844 18828
rect 15896 18816 15902 18828
rect 17512 18825 17540 18856
rect 17954 18844 17960 18856
rect 18012 18844 18018 18896
rect 18046 18844 18052 18896
rect 18104 18884 18110 18896
rect 18509 18887 18567 18893
rect 18509 18884 18521 18887
rect 18104 18856 18521 18884
rect 18104 18844 18110 18856
rect 18509 18853 18521 18856
rect 18555 18853 18567 18887
rect 18509 18847 18567 18853
rect 19058 18844 19064 18896
rect 19116 18884 19122 18896
rect 19245 18887 19303 18893
rect 19245 18884 19257 18887
rect 19116 18856 19257 18884
rect 19116 18844 19122 18856
rect 19245 18853 19257 18856
rect 19291 18853 19303 18887
rect 20349 18887 20407 18893
rect 20349 18884 20361 18887
rect 19245 18847 19303 18853
rect 19352 18856 20361 18884
rect 16301 18819 16359 18825
rect 16301 18816 16313 18819
rect 15896 18788 16313 18816
rect 15896 18776 15902 18788
rect 16301 18785 16313 18788
rect 16347 18785 16359 18819
rect 16301 18779 16359 18785
rect 17497 18819 17555 18825
rect 17497 18785 17509 18819
rect 17543 18785 17555 18819
rect 17497 18779 17555 18785
rect 17586 18776 17592 18828
rect 17644 18816 17650 18828
rect 17773 18819 17831 18825
rect 17773 18816 17785 18819
rect 17644 18788 17785 18816
rect 17644 18776 17650 18788
rect 17773 18785 17785 18788
rect 17819 18785 17831 18819
rect 17773 18779 17831 18785
rect 18141 18819 18199 18825
rect 18141 18785 18153 18819
rect 18187 18785 18199 18819
rect 19352 18816 19380 18856
rect 20349 18853 20361 18856
rect 20395 18853 20407 18887
rect 21542 18884 21548 18896
rect 20349 18847 20407 18853
rect 21468 18856 21548 18884
rect 19518 18816 19524 18828
rect 18141 18779 18199 18785
rect 18248 18788 19380 18816
rect 19479 18788 19524 18816
rect 9030 18748 9036 18760
rect 7944 18720 9036 18748
rect 9030 18708 9036 18720
rect 9088 18708 9094 18760
rect 9214 18748 9220 18760
rect 9175 18720 9220 18748
rect 9214 18708 9220 18720
rect 9272 18748 9278 18760
rect 9398 18748 9404 18760
rect 9272 18720 9404 18748
rect 9272 18708 9278 18720
rect 9398 18708 9404 18720
rect 9456 18708 9462 18760
rect 10965 18751 11023 18757
rect 10965 18717 10977 18751
rect 11011 18748 11023 18751
rect 11054 18748 11060 18760
rect 11011 18720 11060 18748
rect 11011 18717 11023 18720
rect 10965 18711 11023 18717
rect 11054 18708 11060 18720
rect 11112 18748 11118 18760
rect 11238 18748 11244 18760
rect 11112 18720 11244 18748
rect 11112 18708 11118 18720
rect 11238 18708 11244 18720
rect 11296 18708 11302 18760
rect 11698 18708 11704 18760
rect 11756 18748 11762 18760
rect 12253 18751 12311 18757
rect 11756 18720 12204 18748
rect 11756 18708 11762 18720
rect 12176 18692 12204 18720
rect 12253 18717 12265 18751
rect 12299 18748 12311 18751
rect 12710 18748 12716 18760
rect 12299 18720 12716 18748
rect 12299 18717 12311 18720
rect 12253 18711 12311 18717
rect 12710 18708 12716 18720
rect 12768 18748 12774 18760
rect 14274 18748 14280 18760
rect 12768 18720 14280 18748
rect 12768 18708 12774 18720
rect 14274 18708 14280 18720
rect 14332 18708 14338 18760
rect 15013 18751 15071 18757
rect 15013 18717 15025 18751
rect 15059 18717 15071 18751
rect 15013 18711 15071 18717
rect 11882 18680 11888 18692
rect 6012 18652 11888 18680
rect 11882 18640 11888 18652
rect 11940 18640 11946 18692
rect 12158 18640 12164 18692
rect 12216 18640 12222 18692
rect 13262 18640 13268 18692
rect 13320 18680 13326 18692
rect 14461 18683 14519 18689
rect 14461 18680 14473 18683
rect 13320 18652 14473 18680
rect 13320 18640 13326 18652
rect 14461 18649 14473 18652
rect 14507 18649 14519 18683
rect 14461 18643 14519 18649
rect 14642 18640 14648 18692
rect 14700 18680 14706 18692
rect 15028 18680 15056 18711
rect 15562 18708 15568 18760
rect 15620 18748 15626 18760
rect 17402 18748 17408 18760
rect 15620 18720 17408 18748
rect 15620 18708 15626 18720
rect 17402 18708 17408 18720
rect 17460 18708 17466 18760
rect 17678 18708 17684 18760
rect 17736 18748 17742 18760
rect 18156 18748 18184 18779
rect 17736 18720 18184 18748
rect 17736 18708 17742 18720
rect 14700 18652 15056 18680
rect 14700 18640 14706 18652
rect 15838 18640 15844 18692
rect 15896 18680 15902 18692
rect 18248 18680 18276 18788
rect 19518 18776 19524 18788
rect 19576 18776 19582 18828
rect 19610 18776 19616 18828
rect 19668 18816 19674 18828
rect 19978 18816 19984 18828
rect 19668 18788 19713 18816
rect 19891 18788 19984 18816
rect 19668 18776 19674 18788
rect 19978 18776 19984 18788
rect 20036 18816 20042 18828
rect 21177 18819 21235 18825
rect 20036 18788 21128 18816
rect 20036 18776 20042 18788
rect 18690 18708 18696 18760
rect 18748 18748 18754 18760
rect 18748 18720 19090 18748
rect 18748 18708 18754 18720
rect 15896 18652 18276 18680
rect 20533 18683 20591 18689
rect 15896 18640 15902 18652
rect 20533 18649 20545 18683
rect 20579 18680 20591 18683
rect 20898 18680 20904 18692
rect 20579 18652 20904 18680
rect 20579 18649 20591 18652
rect 20533 18643 20591 18649
rect 20898 18640 20904 18652
rect 20956 18640 20962 18692
rect 5994 18612 6000 18624
rect 5907 18584 6000 18612
rect 5994 18572 6000 18584
rect 6052 18612 6058 18624
rect 6270 18612 6276 18624
rect 6052 18584 6276 18612
rect 6052 18572 6058 18584
rect 6270 18572 6276 18584
rect 6328 18572 6334 18624
rect 8570 18612 8576 18624
rect 8531 18584 8576 18612
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 10413 18615 10471 18621
rect 10413 18581 10425 18615
rect 10459 18612 10471 18615
rect 11698 18612 11704 18624
rect 10459 18584 11704 18612
rect 10459 18581 10471 18584
rect 10413 18575 10471 18581
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 15194 18572 15200 18624
rect 15252 18612 15258 18624
rect 16117 18615 16175 18621
rect 16117 18612 16129 18615
rect 15252 18584 16129 18612
rect 15252 18572 15258 18584
rect 16117 18581 16129 18584
rect 16163 18581 16175 18615
rect 16117 18575 16175 18581
rect 16574 18572 16580 18624
rect 16632 18612 16638 18624
rect 19058 18612 19064 18624
rect 16632 18584 19064 18612
rect 16632 18572 16638 18584
rect 19058 18572 19064 18584
rect 19116 18572 19122 18624
rect 21100 18612 21128 18788
rect 21177 18785 21189 18819
rect 21223 18785 21235 18819
rect 21177 18779 21235 18785
rect 21315 18819 21373 18825
rect 21315 18785 21327 18819
rect 21361 18816 21373 18819
rect 21468 18816 21496 18856
rect 21542 18844 21548 18856
rect 21600 18844 21606 18896
rect 22738 18884 22744 18896
rect 21928 18856 22744 18884
rect 21634 18816 21640 18828
rect 21361 18788 21496 18816
rect 21595 18788 21640 18816
rect 21361 18785 21373 18788
rect 21315 18779 21373 18785
rect 21192 18748 21220 18779
rect 21634 18776 21640 18788
rect 21692 18776 21698 18828
rect 21453 18751 21511 18757
rect 21453 18748 21465 18751
rect 21192 18720 21312 18748
rect 21284 18692 21312 18720
rect 21376 18720 21465 18748
rect 21376 18692 21404 18720
rect 21453 18717 21465 18720
rect 21499 18717 21511 18751
rect 21928 18748 21956 18856
rect 22738 18844 22744 18856
rect 22796 18844 22802 18896
rect 23842 18884 23848 18896
rect 23803 18856 23848 18884
rect 23842 18844 23848 18856
rect 23900 18844 23906 18896
rect 23934 18844 23940 18896
rect 23992 18884 23998 18896
rect 24673 18887 24731 18893
rect 24673 18884 24685 18887
rect 23992 18856 24685 18884
rect 23992 18844 23998 18856
rect 24673 18853 24685 18856
rect 24719 18853 24731 18887
rect 25406 18884 25412 18896
rect 25367 18856 25412 18884
rect 24673 18847 24731 18853
rect 25406 18844 25412 18856
rect 25464 18844 25470 18896
rect 25682 18884 25688 18896
rect 25516 18856 25688 18884
rect 23014 18816 23020 18828
rect 21453 18711 21511 18717
rect 21560 18720 21956 18748
rect 22066 18788 23020 18816
rect 21266 18640 21272 18692
rect 21324 18640 21330 18692
rect 21358 18640 21364 18692
rect 21416 18640 21422 18692
rect 21560 18680 21588 18720
rect 21468 18652 21588 18680
rect 21468 18612 21496 18652
rect 21726 18640 21732 18692
rect 21784 18680 21790 18692
rect 22066 18680 22094 18788
rect 23014 18776 23020 18788
rect 23072 18776 23078 18828
rect 23106 18776 23112 18828
rect 23164 18816 23170 18828
rect 23474 18816 23480 18828
rect 23164 18788 23209 18816
rect 23435 18788 23480 18816
rect 23164 18776 23170 18788
rect 23474 18776 23480 18788
rect 23532 18776 23538 18828
rect 24118 18776 24124 18828
rect 24176 18816 24182 18828
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 24176 18788 24593 18816
rect 24176 18776 24182 18788
rect 24581 18785 24593 18788
rect 24627 18785 24639 18819
rect 25516 18816 25544 18856
rect 25682 18844 25688 18856
rect 25740 18844 25746 18896
rect 25777 18887 25835 18893
rect 25777 18853 25789 18887
rect 25823 18853 25835 18887
rect 25777 18847 25835 18853
rect 24581 18779 24639 18785
rect 24780 18788 25544 18816
rect 25792 18816 25820 18847
rect 25958 18816 25964 18828
rect 25792 18788 25964 18816
rect 22646 18708 22652 18760
rect 22704 18708 22710 18760
rect 24210 18708 24216 18760
rect 24268 18748 24274 18760
rect 24780 18748 24808 18788
rect 25958 18776 25964 18788
rect 26016 18776 26022 18828
rect 26142 18816 26148 18828
rect 26103 18788 26148 18816
rect 26142 18776 26148 18788
rect 26200 18776 26206 18828
rect 26234 18776 26240 18828
rect 26292 18816 26298 18828
rect 27985 18819 28043 18825
rect 27985 18816 27997 18819
rect 26292 18788 27997 18816
rect 26292 18776 26298 18788
rect 27985 18785 27997 18788
rect 28031 18785 28043 18819
rect 27985 18779 28043 18785
rect 24268 18720 24808 18748
rect 24268 18708 24274 18720
rect 25866 18708 25872 18760
rect 25924 18708 25930 18760
rect 21784 18652 22094 18680
rect 24029 18683 24087 18689
rect 21784 18640 21790 18652
rect 24029 18649 24041 18683
rect 24075 18680 24087 18683
rect 24118 18680 24124 18692
rect 24075 18652 24124 18680
rect 24075 18649 24087 18652
rect 24029 18643 24087 18649
rect 24118 18640 24124 18652
rect 24176 18640 24182 18692
rect 28166 18680 28172 18692
rect 28127 18652 28172 18680
rect 28166 18640 28172 18652
rect 28224 18640 28230 18692
rect 21100 18584 21496 18612
rect 21545 18615 21603 18621
rect 21545 18581 21557 18615
rect 21591 18612 21603 18615
rect 22370 18612 22376 18624
rect 21591 18584 22376 18612
rect 21591 18581 21603 18584
rect 21545 18575 21603 18581
rect 22370 18572 22376 18584
rect 22428 18572 22434 18624
rect 25038 18572 25044 18624
rect 25096 18612 25102 18624
rect 25406 18612 25412 18624
rect 25096 18584 25412 18612
rect 25096 18572 25102 18584
rect 25406 18572 25412 18584
rect 25464 18572 25470 18624
rect 26602 18572 26608 18624
rect 26660 18612 26666 18624
rect 26697 18615 26755 18621
rect 26697 18612 26709 18615
rect 26660 18584 26709 18612
rect 26660 18572 26666 18584
rect 26697 18581 26709 18584
rect 26743 18581 26755 18615
rect 26697 18575 26755 18581
rect 1104 18522 28888 18544
rect 1104 18470 5614 18522
rect 5666 18470 5678 18522
rect 5730 18470 5742 18522
rect 5794 18470 5806 18522
rect 5858 18470 14878 18522
rect 14930 18470 14942 18522
rect 14994 18470 15006 18522
rect 15058 18470 15070 18522
rect 15122 18470 24142 18522
rect 24194 18470 24206 18522
rect 24258 18470 24270 18522
rect 24322 18470 24334 18522
rect 24386 18470 28888 18522
rect 1104 18448 28888 18470
rect 2406 18368 2412 18420
rect 2464 18408 2470 18420
rect 4341 18411 4399 18417
rect 4341 18408 4353 18411
rect 2464 18380 4353 18408
rect 2464 18368 2470 18380
rect 4341 18377 4353 18380
rect 4387 18377 4399 18411
rect 5442 18408 5448 18420
rect 5403 18380 5448 18408
rect 4341 18371 4399 18377
rect 5442 18368 5448 18380
rect 5500 18368 5506 18420
rect 11790 18408 11796 18420
rect 7576 18380 11796 18408
rect 2682 18300 2688 18352
rect 2740 18340 2746 18352
rect 7576 18340 7604 18380
rect 11790 18368 11796 18380
rect 11848 18368 11854 18420
rect 11882 18368 11888 18420
rect 11940 18408 11946 18420
rect 15838 18408 15844 18420
rect 11940 18380 15844 18408
rect 11940 18368 11946 18380
rect 15838 18368 15844 18380
rect 15896 18368 15902 18420
rect 17129 18411 17187 18417
rect 17129 18377 17141 18411
rect 17175 18408 17187 18411
rect 17586 18408 17592 18420
rect 17175 18380 17592 18408
rect 17175 18377 17187 18380
rect 17129 18371 17187 18377
rect 17586 18368 17592 18380
rect 17644 18368 17650 18420
rect 18322 18408 18328 18420
rect 18283 18380 18328 18408
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 19518 18408 19524 18420
rect 18708 18380 19524 18408
rect 2740 18312 7604 18340
rect 2740 18300 2746 18312
rect 9214 18300 9220 18352
rect 9272 18340 9278 18352
rect 9677 18343 9735 18349
rect 9677 18340 9689 18343
rect 9272 18312 9689 18340
rect 9272 18300 9278 18312
rect 9677 18309 9689 18312
rect 9723 18309 9735 18343
rect 11606 18340 11612 18352
rect 9677 18303 9735 18309
rect 9784 18312 11612 18340
rect 2314 18232 2320 18284
rect 2372 18272 2378 18284
rect 2409 18275 2467 18281
rect 2409 18272 2421 18275
rect 2372 18244 2421 18272
rect 2372 18232 2378 18244
rect 2409 18241 2421 18244
rect 2455 18241 2467 18275
rect 2409 18235 2467 18241
rect 2976 18244 3280 18272
rect 2225 18139 2283 18145
rect 2225 18105 2237 18139
rect 2271 18136 2283 18139
rect 2774 18136 2780 18148
rect 2271 18108 2780 18136
rect 2271 18105 2283 18108
rect 2225 18099 2283 18105
rect 2774 18096 2780 18108
rect 2832 18096 2838 18148
rect 1854 18068 1860 18080
rect 1815 18040 1860 18068
rect 1854 18028 1860 18040
rect 1912 18028 1918 18080
rect 2314 18068 2320 18080
rect 2275 18040 2320 18068
rect 2314 18028 2320 18040
rect 2372 18068 2378 18080
rect 2976 18068 3004 18244
rect 3050 18164 3056 18216
rect 3108 18204 3114 18216
rect 3252 18213 3280 18244
rect 4798 18232 4804 18284
rect 4856 18272 4862 18284
rect 4893 18275 4951 18281
rect 4893 18272 4905 18275
rect 4856 18244 4905 18272
rect 4856 18232 4862 18244
rect 4893 18241 4905 18244
rect 4939 18241 4951 18275
rect 4893 18235 4951 18241
rect 5902 18232 5908 18284
rect 5960 18272 5966 18284
rect 5997 18275 6055 18281
rect 5997 18272 6009 18275
rect 5960 18244 6009 18272
rect 5960 18232 5966 18244
rect 5997 18241 6009 18244
rect 6043 18241 6055 18275
rect 9784 18272 9812 18312
rect 11606 18300 11612 18312
rect 11664 18300 11670 18352
rect 13814 18340 13820 18352
rect 11716 18312 13820 18340
rect 5997 18235 6055 18241
rect 6104 18244 9812 18272
rect 10965 18275 11023 18281
rect 3237 18207 3295 18213
rect 3108 18176 3153 18204
rect 3108 18164 3114 18176
rect 3237 18173 3249 18207
rect 3283 18173 3295 18207
rect 3237 18167 3295 18173
rect 4154 18164 4160 18216
rect 4212 18204 4218 18216
rect 5074 18204 5080 18216
rect 4212 18176 5080 18204
rect 4212 18164 4218 18176
rect 5074 18164 5080 18176
rect 5132 18204 5138 18216
rect 6104 18204 6132 18244
rect 10965 18241 10977 18275
rect 11011 18272 11023 18275
rect 11716 18272 11744 18312
rect 13814 18300 13820 18312
rect 13872 18300 13878 18352
rect 14829 18343 14887 18349
rect 14829 18340 14841 18343
rect 14200 18312 14841 18340
rect 11011 18244 11744 18272
rect 11011 18241 11023 18244
rect 10965 18235 11023 18241
rect 13078 18232 13084 18284
rect 13136 18272 13142 18284
rect 13906 18272 13912 18284
rect 13136 18244 13912 18272
rect 13136 18232 13142 18244
rect 13906 18232 13912 18244
rect 13964 18272 13970 18284
rect 14200 18272 14228 18312
rect 14829 18309 14841 18312
rect 14875 18309 14887 18343
rect 14829 18303 14887 18309
rect 17402 18300 17408 18352
rect 17460 18340 17466 18352
rect 18708 18340 18736 18380
rect 19518 18368 19524 18380
rect 19576 18408 19582 18420
rect 20806 18408 20812 18420
rect 19576 18380 20668 18408
rect 20767 18380 20812 18408
rect 19576 18368 19582 18380
rect 19978 18340 19984 18352
rect 17460 18312 18736 18340
rect 18800 18312 19984 18340
rect 17460 18300 17466 18312
rect 13964 18244 14228 18272
rect 13964 18232 13970 18244
rect 15838 18232 15844 18284
rect 15896 18232 15902 18284
rect 18800 18281 18828 18312
rect 19978 18300 19984 18312
rect 20036 18300 20042 18352
rect 20640 18340 20668 18380
rect 20806 18368 20812 18380
rect 20864 18368 20870 18420
rect 21266 18368 21272 18420
rect 21324 18408 21330 18420
rect 21542 18408 21548 18420
rect 21324 18380 21548 18408
rect 21324 18368 21330 18380
rect 21542 18368 21548 18380
rect 21600 18368 21606 18420
rect 24121 18411 24179 18417
rect 22066 18380 24072 18408
rect 22066 18340 22094 18380
rect 20640 18312 22094 18340
rect 23474 18300 23480 18352
rect 23532 18340 23538 18352
rect 23661 18343 23719 18349
rect 23661 18340 23673 18343
rect 23532 18312 23673 18340
rect 23532 18300 23538 18312
rect 23661 18309 23673 18312
rect 23707 18309 23719 18343
rect 24044 18340 24072 18380
rect 24121 18377 24133 18411
rect 24167 18408 24179 18411
rect 24670 18408 24676 18420
rect 24167 18380 24676 18408
rect 24167 18377 24179 18380
rect 24121 18371 24179 18377
rect 24670 18368 24676 18380
rect 24728 18368 24734 18420
rect 25958 18408 25964 18420
rect 25240 18380 25964 18408
rect 25038 18340 25044 18352
rect 24044 18312 25044 18340
rect 23661 18303 23719 18309
rect 25038 18300 25044 18312
rect 25096 18300 25102 18352
rect 18785 18275 18843 18281
rect 18785 18241 18797 18275
rect 18831 18241 18843 18275
rect 18785 18235 18843 18241
rect 18969 18275 19027 18281
rect 18969 18241 18981 18275
rect 19015 18272 19027 18275
rect 19242 18272 19248 18284
rect 19015 18244 19248 18272
rect 19015 18241 19027 18244
rect 18969 18235 19027 18241
rect 19242 18232 19248 18244
rect 19300 18232 19306 18284
rect 21726 18272 21732 18284
rect 19352 18244 21732 18272
rect 5132 18176 6132 18204
rect 5132 18164 5138 18176
rect 8754 18164 8760 18216
rect 8812 18204 8818 18216
rect 9398 18204 9404 18216
rect 8812 18176 9404 18204
rect 8812 18164 8818 18176
rect 9398 18164 9404 18176
rect 9456 18204 9462 18216
rect 9493 18207 9551 18213
rect 9493 18204 9505 18207
rect 9456 18176 9505 18204
rect 9456 18164 9462 18176
rect 9493 18173 9505 18176
rect 9539 18173 9551 18207
rect 9493 18167 9551 18173
rect 10134 18164 10140 18216
rect 10192 18204 10198 18216
rect 10229 18207 10287 18213
rect 10229 18204 10241 18207
rect 10192 18176 10241 18204
rect 10192 18164 10198 18176
rect 10229 18173 10241 18176
rect 10275 18173 10287 18207
rect 10229 18167 10287 18173
rect 11054 18164 11060 18216
rect 11112 18204 11118 18216
rect 11514 18204 11520 18216
rect 11112 18176 11520 18204
rect 11112 18164 11118 18176
rect 11514 18164 11520 18176
rect 11572 18204 11578 18216
rect 11609 18207 11667 18213
rect 11609 18204 11621 18207
rect 11572 18176 11621 18204
rect 11572 18164 11578 18176
rect 11609 18173 11621 18176
rect 11655 18173 11667 18207
rect 11609 18167 11667 18173
rect 11698 18164 11704 18216
rect 11756 18164 11762 18216
rect 14642 18164 14648 18216
rect 14700 18204 14706 18216
rect 14737 18207 14795 18213
rect 14737 18204 14749 18207
rect 14700 18176 14749 18204
rect 14700 18164 14706 18176
rect 14737 18173 14749 18176
rect 14783 18173 14795 18207
rect 14737 18167 14795 18173
rect 16022 18164 16028 18216
rect 16080 18204 16086 18216
rect 16209 18207 16267 18213
rect 16209 18204 16221 18207
rect 16080 18176 16221 18204
rect 16080 18164 16086 18176
rect 16209 18173 16221 18176
rect 16255 18173 16267 18207
rect 16209 18167 16267 18173
rect 16574 18164 16580 18216
rect 16632 18204 16638 18216
rect 16959 18207 17017 18213
rect 16959 18204 16971 18207
rect 16632 18176 16677 18204
rect 16776 18176 16971 18204
rect 16632 18164 16638 18176
rect 3145 18139 3203 18145
rect 3145 18105 3157 18139
rect 3191 18136 3203 18139
rect 4617 18139 4675 18145
rect 4617 18136 4629 18139
rect 3191 18108 4629 18136
rect 3191 18105 3203 18108
rect 3145 18099 3203 18105
rect 4617 18105 4629 18108
rect 4663 18105 4675 18139
rect 4617 18099 4675 18105
rect 5813 18139 5871 18145
rect 5813 18105 5825 18139
rect 5859 18136 5871 18139
rect 5994 18136 6000 18148
rect 5859 18108 6000 18136
rect 5859 18105 5871 18108
rect 5813 18099 5871 18105
rect 5994 18096 6000 18108
rect 6052 18096 6058 18148
rect 16117 18139 16175 18145
rect 16117 18105 16129 18139
rect 16163 18136 16175 18139
rect 16390 18136 16396 18148
rect 16163 18108 16396 18136
rect 16163 18105 16175 18108
rect 16117 18099 16175 18105
rect 16390 18096 16396 18108
rect 16448 18096 16454 18148
rect 16666 18096 16672 18148
rect 16724 18136 16730 18148
rect 16776 18136 16804 18176
rect 16959 18173 16971 18176
rect 17005 18173 17017 18207
rect 16959 18167 17017 18173
rect 17862 18164 17868 18216
rect 17920 18204 17926 18216
rect 18693 18207 18751 18213
rect 18693 18204 18705 18207
rect 17920 18176 18705 18204
rect 17920 18164 17926 18176
rect 18693 18173 18705 18176
rect 18739 18173 18751 18207
rect 18693 18167 18751 18173
rect 19352 18136 19380 18244
rect 21726 18232 21732 18244
rect 21784 18232 21790 18284
rect 22278 18272 22284 18284
rect 22239 18244 22284 18272
rect 22278 18232 22284 18244
rect 22336 18232 22342 18284
rect 23934 18232 23940 18284
rect 23992 18272 23998 18284
rect 25240 18281 25268 18380
rect 25958 18368 25964 18380
rect 26016 18368 26022 18420
rect 26142 18368 26148 18420
rect 26200 18408 26206 18420
rect 26605 18411 26663 18417
rect 26605 18408 26617 18411
rect 26200 18380 26617 18408
rect 26200 18368 26206 18380
rect 26605 18377 26617 18380
rect 26651 18377 26663 18411
rect 27430 18408 27436 18420
rect 27391 18380 27436 18408
rect 26605 18371 26663 18377
rect 27430 18368 27436 18380
rect 27488 18368 27494 18420
rect 28074 18408 28080 18420
rect 27908 18380 28080 18408
rect 27908 18281 27936 18380
rect 28074 18368 28080 18380
rect 28132 18368 28138 18420
rect 25225 18275 25283 18281
rect 23992 18244 24348 18272
rect 23992 18232 23998 18244
rect 20714 18204 20720 18216
rect 20627 18176 20720 18204
rect 20714 18164 20720 18176
rect 20772 18164 20778 18216
rect 20898 18204 20904 18216
rect 20859 18176 20904 18204
rect 20898 18164 20904 18176
rect 20956 18164 20962 18216
rect 21174 18204 21180 18216
rect 21135 18176 21180 18204
rect 21174 18164 21180 18176
rect 21232 18164 21238 18216
rect 22370 18164 22376 18216
rect 22428 18204 22434 18216
rect 24320 18213 24348 18244
rect 25225 18241 25237 18275
rect 25271 18241 25283 18275
rect 25225 18235 25283 18241
rect 27893 18275 27951 18281
rect 27893 18241 27905 18275
rect 27939 18241 27951 18275
rect 28074 18272 28080 18284
rect 28035 18244 28080 18272
rect 27893 18235 27951 18241
rect 28074 18232 28080 18244
rect 28132 18232 28138 18284
rect 22537 18207 22595 18213
rect 22537 18204 22549 18207
rect 22428 18176 22549 18204
rect 22428 18164 22434 18176
rect 22537 18173 22549 18176
rect 22583 18173 22595 18207
rect 24121 18207 24179 18213
rect 24121 18204 24133 18207
rect 22537 18167 22595 18173
rect 23952 18176 24133 18204
rect 16724 18108 16804 18136
rect 16868 18108 19380 18136
rect 20732 18136 20760 18164
rect 23952 18148 23980 18176
rect 24121 18173 24133 18176
rect 24167 18173 24179 18207
rect 24121 18167 24179 18173
rect 24305 18207 24363 18213
rect 24305 18173 24317 18207
rect 24351 18173 24363 18207
rect 24305 18167 24363 18173
rect 25314 18164 25320 18216
rect 25372 18204 25378 18216
rect 25481 18207 25539 18213
rect 25481 18204 25493 18207
rect 25372 18176 25493 18204
rect 25372 18164 25378 18176
rect 25481 18173 25493 18176
rect 25527 18173 25539 18207
rect 27798 18204 27804 18216
rect 27759 18176 27804 18204
rect 25481 18167 25539 18173
rect 27798 18164 27804 18176
rect 27856 18164 27862 18216
rect 21266 18136 21272 18148
rect 20732 18108 21272 18136
rect 16724 18096 16730 18108
rect 4798 18068 4804 18080
rect 2372 18040 3004 18068
rect 4759 18040 4804 18068
rect 2372 18028 2378 18040
rect 4798 18028 4804 18040
rect 4856 18028 4862 18080
rect 5905 18071 5963 18077
rect 5905 18037 5917 18071
rect 5951 18068 5963 18071
rect 8294 18068 8300 18080
rect 5951 18040 8300 18068
rect 5951 18037 5963 18040
rect 5905 18031 5963 18037
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 10321 18071 10379 18077
rect 10321 18037 10333 18071
rect 10367 18068 10379 18071
rect 11977 18071 12035 18077
rect 11977 18068 11989 18071
rect 10367 18040 11989 18068
rect 10367 18037 10379 18040
rect 10321 18031 10379 18037
rect 11977 18037 11989 18040
rect 12023 18037 12035 18071
rect 11977 18031 12035 18037
rect 12066 18028 12072 18080
rect 12124 18068 12130 18080
rect 15562 18068 15568 18080
rect 12124 18040 15568 18068
rect 12124 18028 12130 18040
rect 15562 18028 15568 18040
rect 15620 18028 15626 18080
rect 15746 18028 15752 18080
rect 15804 18068 15810 18080
rect 15841 18071 15899 18077
rect 15841 18068 15853 18071
rect 15804 18040 15853 18068
rect 15804 18028 15810 18040
rect 15841 18037 15853 18040
rect 15887 18068 15899 18071
rect 16868 18068 16896 18108
rect 21266 18096 21272 18108
rect 21324 18096 21330 18148
rect 22066 18108 23888 18136
rect 15887 18040 16896 18068
rect 15887 18037 15899 18040
rect 15841 18031 15899 18037
rect 17034 18028 17040 18080
rect 17092 18068 17098 18080
rect 22066 18068 22094 18108
rect 17092 18040 22094 18068
rect 23860 18068 23888 18108
rect 23934 18096 23940 18148
rect 23992 18096 23998 18148
rect 27706 18068 27712 18080
rect 23860 18040 27712 18068
rect 17092 18028 17098 18040
rect 27706 18028 27712 18040
rect 27764 18028 27770 18080
rect 1104 17978 28888 18000
rect 1104 17926 10246 17978
rect 10298 17926 10310 17978
rect 10362 17926 10374 17978
rect 10426 17926 10438 17978
rect 10490 17926 19510 17978
rect 19562 17926 19574 17978
rect 19626 17926 19638 17978
rect 19690 17926 19702 17978
rect 19754 17926 28888 17978
rect 1104 17904 28888 17926
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 3237 17867 3295 17873
rect 2832 17836 2877 17864
rect 2832 17824 2838 17836
rect 3237 17833 3249 17867
rect 3283 17864 3295 17867
rect 4798 17864 4804 17876
rect 3283 17836 4804 17864
rect 3283 17833 3295 17836
rect 3237 17827 3295 17833
rect 4798 17824 4804 17836
rect 4856 17824 4862 17876
rect 5251 17867 5309 17873
rect 5251 17833 5263 17867
rect 5297 17864 5309 17867
rect 8846 17864 8852 17876
rect 5297 17836 8852 17864
rect 5297 17833 5309 17836
rect 5251 17827 5309 17833
rect 8846 17824 8852 17836
rect 8904 17824 8910 17876
rect 8938 17824 8944 17876
rect 8996 17864 9002 17876
rect 9582 17864 9588 17876
rect 8996 17836 9588 17864
rect 8996 17824 9002 17836
rect 9582 17824 9588 17836
rect 9640 17864 9646 17876
rect 9677 17867 9735 17873
rect 9677 17864 9689 17867
rect 9640 17836 9689 17864
rect 9640 17824 9646 17836
rect 9677 17833 9689 17836
rect 9723 17833 9735 17867
rect 9677 17827 9735 17833
rect 10134 17824 10140 17876
rect 10192 17864 10198 17876
rect 10229 17867 10287 17873
rect 10229 17864 10241 17867
rect 10192 17836 10241 17864
rect 10192 17824 10198 17836
rect 10229 17833 10241 17836
rect 10275 17833 10287 17867
rect 10686 17864 10692 17876
rect 10647 17836 10692 17864
rect 10229 17827 10287 17833
rect 10686 17824 10692 17836
rect 10744 17824 10750 17876
rect 14182 17864 14188 17876
rect 10796 17836 13952 17864
rect 14143 17836 14188 17864
rect 1664 17799 1722 17805
rect 1664 17765 1676 17799
rect 1710 17796 1722 17799
rect 1854 17796 1860 17808
rect 1710 17768 1860 17796
rect 1710 17765 1722 17768
rect 1664 17759 1722 17765
rect 1854 17756 1860 17768
rect 1912 17756 1918 17808
rect 4338 17756 4344 17808
rect 4396 17796 4402 17808
rect 4525 17799 4583 17805
rect 4525 17796 4537 17799
rect 4396 17768 4537 17796
rect 4396 17756 4402 17768
rect 4525 17765 4537 17768
rect 4571 17765 4583 17799
rect 4525 17759 4583 17765
rect 5166 17756 5172 17808
rect 5224 17796 5230 17808
rect 5721 17799 5779 17805
rect 5721 17796 5733 17799
rect 5224 17768 5733 17796
rect 5224 17756 5230 17768
rect 5721 17765 5733 17768
rect 5767 17765 5779 17799
rect 5721 17759 5779 17765
rect 5813 17799 5871 17805
rect 5813 17765 5825 17799
rect 5859 17796 5871 17799
rect 6178 17796 6184 17808
rect 5859 17768 6184 17796
rect 5859 17765 5871 17768
rect 5813 17759 5871 17765
rect 6178 17756 6184 17768
rect 6236 17756 6242 17808
rect 8570 17805 8576 17808
rect 8564 17796 8576 17805
rect 8531 17768 8576 17796
rect 8564 17759 8576 17768
rect 8570 17756 8576 17759
rect 8628 17756 8634 17808
rect 8662 17756 8668 17808
rect 8720 17796 8726 17808
rect 10796 17796 10824 17836
rect 8720 17768 10824 17796
rect 13924 17796 13952 17836
rect 14182 17824 14188 17836
rect 14240 17824 14246 17876
rect 15470 17824 15476 17876
rect 15528 17864 15534 17876
rect 16390 17864 16396 17876
rect 15528 17836 16396 17864
rect 15528 17824 15534 17836
rect 16390 17824 16396 17836
rect 16448 17824 16454 17876
rect 17497 17867 17555 17873
rect 17497 17833 17509 17867
rect 17543 17864 17555 17867
rect 18230 17864 18236 17876
rect 17543 17836 18236 17864
rect 17543 17833 17555 17836
rect 17497 17827 17555 17833
rect 18230 17824 18236 17836
rect 18288 17824 18294 17876
rect 21634 17824 21640 17876
rect 21692 17864 21698 17876
rect 22649 17867 22707 17873
rect 22649 17864 22661 17867
rect 21692 17836 22661 17864
rect 21692 17824 21698 17836
rect 22649 17833 22661 17836
rect 22695 17833 22707 17867
rect 22649 17827 22707 17833
rect 26053 17867 26111 17873
rect 26053 17833 26065 17867
rect 26099 17864 26111 17867
rect 26510 17864 26516 17876
rect 26099 17836 26516 17864
rect 26099 17833 26111 17836
rect 26053 17827 26111 17833
rect 26510 17824 26516 17836
rect 26568 17824 26574 17876
rect 14645 17799 14703 17805
rect 14645 17796 14657 17799
rect 13924 17768 14657 17796
rect 8720 17756 8726 17768
rect 14200 17740 14228 17768
rect 14645 17765 14657 17768
rect 14691 17765 14703 17799
rect 23474 17796 23480 17808
rect 14645 17759 14703 17765
rect 22572 17768 23480 17796
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 1443 17700 2774 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 2746 17524 2774 17700
rect 3050 17688 3056 17740
rect 3108 17728 3114 17740
rect 3605 17731 3663 17737
rect 3605 17728 3617 17731
rect 3108 17700 3617 17728
rect 3108 17688 3114 17700
rect 3605 17697 3617 17700
rect 3651 17697 3663 17731
rect 3605 17691 3663 17697
rect 3697 17731 3755 17737
rect 3697 17697 3709 17731
rect 3743 17728 3755 17731
rect 4154 17728 4160 17740
rect 3743 17700 4160 17728
rect 3743 17697 3755 17700
rect 3697 17691 3755 17697
rect 4154 17688 4160 17700
rect 4212 17688 4218 17740
rect 4433 17731 4491 17737
rect 4433 17697 4445 17731
rect 4479 17697 4491 17731
rect 4433 17691 4491 17697
rect 7009 17731 7067 17737
rect 7009 17697 7021 17731
rect 7055 17728 7067 17731
rect 7374 17728 7380 17740
rect 7055 17700 7380 17728
rect 7055 17697 7067 17700
rect 7009 17691 7067 17697
rect 3878 17660 3884 17672
rect 3839 17632 3884 17660
rect 3878 17620 3884 17632
rect 3936 17620 3942 17672
rect 2958 17552 2964 17604
rect 3016 17592 3022 17604
rect 4448 17592 4476 17691
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 7466 17688 7472 17740
rect 7524 17728 7530 17740
rect 10597 17731 10655 17737
rect 10597 17728 10609 17731
rect 7524 17700 10609 17728
rect 7524 17688 7530 17700
rect 10597 17697 10609 17700
rect 10643 17697 10655 17731
rect 10597 17691 10655 17697
rect 12069 17731 12127 17737
rect 12069 17697 12081 17731
rect 12115 17728 12127 17731
rect 12710 17728 12716 17740
rect 12115 17700 12716 17728
rect 12115 17697 12127 17700
rect 12069 17691 12127 17697
rect 12710 17688 12716 17700
rect 12768 17688 12774 17740
rect 14182 17688 14188 17740
rect 14240 17688 14246 17740
rect 14550 17728 14556 17740
rect 14511 17700 14556 17728
rect 14550 17688 14556 17700
rect 14608 17688 14614 17740
rect 17586 17688 17592 17740
rect 17644 17728 17650 17740
rect 17773 17731 17831 17737
rect 17773 17728 17785 17731
rect 17644 17700 17785 17728
rect 17644 17688 17650 17700
rect 17773 17697 17785 17700
rect 17819 17697 17831 17731
rect 17954 17728 17960 17740
rect 17915 17700 17960 17728
rect 17773 17691 17831 17697
rect 17954 17688 17960 17700
rect 18012 17688 18018 17740
rect 22572 17737 22600 17768
rect 23474 17756 23480 17768
rect 23532 17756 23538 17808
rect 25038 17756 25044 17808
rect 25096 17796 25102 17808
rect 27985 17799 28043 17805
rect 27985 17796 27997 17799
rect 25096 17768 27997 17796
rect 25096 17756 25102 17768
rect 27985 17765 27997 17768
rect 28031 17765 28043 17799
rect 27985 17759 28043 17765
rect 22557 17731 22615 17737
rect 22557 17697 22569 17731
rect 22603 17697 22615 17731
rect 22557 17691 22615 17697
rect 22741 17731 22799 17737
rect 22741 17697 22753 17731
rect 22787 17728 22799 17731
rect 23014 17728 23020 17740
rect 22787 17700 23020 17728
rect 22787 17697 22799 17700
rect 22741 17691 22799 17697
rect 23014 17688 23020 17700
rect 23072 17688 23078 17740
rect 25961 17731 26019 17737
rect 25961 17697 25973 17731
rect 26007 17728 26019 17731
rect 26602 17728 26608 17740
rect 26007 17700 26608 17728
rect 26007 17697 26019 17700
rect 25961 17691 26019 17697
rect 26602 17688 26608 17700
rect 26660 17688 26666 17740
rect 26697 17731 26755 17737
rect 26697 17697 26709 17731
rect 26743 17697 26755 17731
rect 26878 17728 26884 17740
rect 26839 17700 26884 17728
rect 26697 17691 26755 17697
rect 5721 17663 5779 17669
rect 5721 17629 5733 17663
rect 5767 17629 5779 17663
rect 7101 17663 7159 17669
rect 7101 17660 7113 17663
rect 5721 17623 5779 17629
rect 7024 17632 7113 17660
rect 3016 17564 4476 17592
rect 5736 17592 5764 17623
rect 7024 17604 7052 17632
rect 7101 17629 7113 17632
rect 7147 17629 7159 17663
rect 8297 17663 8355 17669
rect 8297 17660 8309 17663
rect 7101 17623 7159 17629
rect 7208 17632 8309 17660
rect 5902 17592 5908 17604
rect 5736 17564 5908 17592
rect 3016 17552 3022 17564
rect 5902 17552 5908 17564
rect 5960 17552 5966 17604
rect 7006 17552 7012 17604
rect 7064 17552 7070 17604
rect 6730 17524 6736 17536
rect 2746 17496 6736 17524
rect 6730 17484 6736 17496
rect 6788 17524 6794 17536
rect 7208 17524 7236 17632
rect 8297 17629 8309 17632
rect 8343 17629 8355 17663
rect 8297 17623 8355 17629
rect 10873 17663 10931 17669
rect 10873 17629 10885 17663
rect 10919 17660 10931 17663
rect 11238 17660 11244 17672
rect 10919 17632 11244 17660
rect 10919 17629 10931 17632
rect 10873 17623 10931 17629
rect 6788 17496 7236 17524
rect 6788 17484 6794 17496
rect 7282 17484 7288 17536
rect 7340 17524 7346 17536
rect 7377 17527 7435 17533
rect 7377 17524 7389 17527
rect 7340 17496 7389 17524
rect 7340 17484 7346 17496
rect 7377 17493 7389 17496
rect 7423 17493 7435 17527
rect 8312 17524 8340 17623
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 12250 17620 12256 17672
rect 12308 17660 12314 17672
rect 12345 17663 12403 17669
rect 12345 17660 12357 17663
rect 12308 17632 12357 17660
rect 12308 17620 12314 17632
rect 12345 17629 12357 17632
rect 12391 17629 12403 17663
rect 12345 17623 12403 17629
rect 14642 17620 14648 17672
rect 14700 17660 14706 17672
rect 14737 17663 14795 17669
rect 14737 17660 14749 17663
rect 14700 17632 14749 17660
rect 14700 17620 14706 17632
rect 14737 17629 14749 17632
rect 14783 17629 14795 17663
rect 14737 17623 14795 17629
rect 17681 17663 17739 17669
rect 17681 17629 17693 17663
rect 17727 17629 17739 17663
rect 17862 17660 17868 17672
rect 17823 17632 17868 17660
rect 17681 17623 17739 17629
rect 17586 17552 17592 17604
rect 17644 17592 17650 17604
rect 17696 17592 17724 17623
rect 17862 17620 17868 17632
rect 17920 17620 17926 17672
rect 25682 17620 25688 17672
rect 25740 17660 25746 17672
rect 26712 17660 26740 17691
rect 26878 17688 26884 17700
rect 26936 17688 26942 17740
rect 25740 17632 26740 17660
rect 25740 17620 25746 17632
rect 28166 17592 28172 17604
rect 17644 17564 17724 17592
rect 28127 17564 28172 17592
rect 17644 17552 17650 17564
rect 28166 17552 28172 17564
rect 28224 17552 28230 17604
rect 8478 17524 8484 17536
rect 8312 17496 8484 17524
rect 7377 17487 7435 17493
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 11882 17484 11888 17536
rect 11940 17524 11946 17536
rect 13449 17527 13507 17533
rect 13449 17524 13461 17527
rect 11940 17496 13461 17524
rect 11940 17484 11946 17496
rect 13449 17493 13461 17496
rect 13495 17493 13507 17527
rect 13449 17487 13507 17493
rect 1104 17434 28888 17456
rect 1104 17382 5614 17434
rect 5666 17382 5678 17434
rect 5730 17382 5742 17434
rect 5794 17382 5806 17434
rect 5858 17382 14878 17434
rect 14930 17382 14942 17434
rect 14994 17382 15006 17434
rect 15058 17382 15070 17434
rect 15122 17382 24142 17434
rect 24194 17382 24206 17434
rect 24258 17382 24270 17434
rect 24322 17382 24334 17434
rect 24386 17382 28888 17434
rect 1104 17360 28888 17382
rect 3050 17320 3056 17332
rect 3011 17292 3056 17320
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 5166 17320 5172 17332
rect 5127 17292 5172 17320
rect 5166 17280 5172 17292
rect 5224 17280 5230 17332
rect 9677 17323 9735 17329
rect 9677 17289 9689 17323
rect 9723 17320 9735 17323
rect 9858 17320 9864 17332
rect 9723 17292 9864 17320
rect 9723 17289 9735 17292
rect 9677 17283 9735 17289
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 20530 17280 20536 17332
rect 20588 17320 20594 17332
rect 20898 17320 20904 17332
rect 20588 17292 20904 17320
rect 20588 17280 20594 17292
rect 20898 17280 20904 17292
rect 20956 17280 20962 17332
rect 26878 17320 26884 17332
rect 26839 17292 26884 17320
rect 26878 17280 26884 17292
rect 26936 17280 26942 17332
rect 1765 17255 1823 17261
rect 1765 17221 1777 17255
rect 1811 17252 1823 17255
rect 4982 17252 4988 17264
rect 1811 17224 4988 17252
rect 1811 17221 1823 17224
rect 1765 17215 1823 17221
rect 4982 17212 4988 17224
rect 5040 17212 5046 17264
rect 14550 17252 14556 17264
rect 5644 17224 14556 17252
rect 1670 17144 1676 17196
rect 1728 17184 1734 17196
rect 5644 17184 5672 17224
rect 14550 17212 14556 17224
rect 14608 17212 14614 17264
rect 19981 17255 20039 17261
rect 19981 17221 19993 17255
rect 20027 17252 20039 17255
rect 20990 17252 20996 17264
rect 20027 17224 20996 17252
rect 20027 17221 20039 17224
rect 19981 17215 20039 17221
rect 20990 17212 20996 17224
rect 21048 17252 21054 17264
rect 21358 17252 21364 17264
rect 21048 17224 21364 17252
rect 21048 17212 21054 17224
rect 21358 17212 21364 17224
rect 21416 17212 21422 17264
rect 21634 17252 21640 17264
rect 21595 17224 21640 17252
rect 21634 17212 21640 17224
rect 21692 17212 21698 17264
rect 1728 17156 5672 17184
rect 5813 17187 5871 17193
rect 1728 17144 1734 17156
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 6086 17184 6092 17196
rect 5859 17156 6092 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 6086 17144 6092 17156
rect 6144 17184 6150 17196
rect 6638 17184 6644 17196
rect 6144 17156 6644 17184
rect 6144 17144 6150 17156
rect 6638 17144 6644 17156
rect 6696 17144 6702 17196
rect 7558 17184 7564 17196
rect 7519 17156 7564 17184
rect 7558 17144 7564 17156
rect 7616 17144 7622 17196
rect 18969 17187 19027 17193
rect 18969 17153 18981 17187
rect 19015 17184 19027 17187
rect 19242 17184 19248 17196
rect 19015 17156 19248 17184
rect 19015 17153 19027 17156
rect 18969 17147 19027 17153
rect 19242 17144 19248 17156
rect 19300 17144 19306 17196
rect 20898 17144 20904 17196
rect 20956 17184 20962 17196
rect 21082 17184 21088 17196
rect 20956 17156 21088 17184
rect 20956 17144 20962 17156
rect 21082 17144 21088 17156
rect 21140 17184 21146 17196
rect 21269 17187 21327 17193
rect 21269 17184 21281 17187
rect 21140 17156 21281 17184
rect 21140 17144 21146 17156
rect 21269 17153 21281 17156
rect 21315 17153 21327 17187
rect 21269 17147 21327 17153
rect 28077 17187 28135 17193
rect 28077 17153 28089 17187
rect 28123 17184 28135 17187
rect 28350 17184 28356 17196
rect 28123 17156 28356 17184
rect 28123 17153 28135 17156
rect 28077 17147 28135 17153
rect 28350 17144 28356 17156
rect 28408 17144 28414 17196
rect 1946 17116 1952 17128
rect 1907 17088 1952 17116
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 2866 17076 2872 17128
rect 2924 17116 2930 17128
rect 2961 17119 3019 17125
rect 2961 17116 2973 17119
rect 2924 17088 2973 17116
rect 2924 17076 2930 17088
rect 2961 17085 2973 17088
rect 3007 17085 3019 17119
rect 2961 17079 3019 17085
rect 3970 17076 3976 17128
rect 4028 17116 4034 17128
rect 4982 17116 4988 17128
rect 4028 17088 4988 17116
rect 4028 17076 4034 17088
rect 4982 17076 4988 17088
rect 5040 17116 5046 17128
rect 5537 17119 5595 17125
rect 5537 17116 5549 17119
rect 5040 17088 5549 17116
rect 5040 17076 5046 17088
rect 5537 17085 5549 17088
rect 5583 17085 5595 17119
rect 7282 17116 7288 17128
rect 7243 17088 7288 17116
rect 5537 17079 5595 17085
rect 7282 17076 7288 17088
rect 7340 17076 7346 17128
rect 9582 17116 9588 17128
rect 9543 17088 9588 17116
rect 9582 17076 9588 17088
rect 9640 17076 9646 17128
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17085 11023 17119
rect 10965 17079 11023 17085
rect 2682 17008 2688 17060
rect 2740 17048 2746 17060
rect 5994 17048 6000 17060
rect 2740 17020 6000 17048
rect 2740 17008 2746 17020
rect 5994 17008 6000 17020
rect 6052 17008 6058 17060
rect 9398 17008 9404 17060
rect 9456 17048 9462 17060
rect 10980 17048 11008 17079
rect 11422 17076 11428 17128
rect 11480 17116 11486 17128
rect 11882 17116 11888 17128
rect 11480 17088 11888 17116
rect 11480 17076 11486 17088
rect 11882 17076 11888 17088
rect 11940 17076 11946 17128
rect 15194 17076 15200 17128
rect 15252 17116 15258 17128
rect 20165 17119 20223 17125
rect 20165 17116 20177 17119
rect 15252 17088 20177 17116
rect 15252 17076 15258 17088
rect 20165 17085 20177 17088
rect 20211 17085 20223 17119
rect 20165 17079 20223 17085
rect 26053 17119 26111 17125
rect 26053 17085 26065 17119
rect 26099 17116 26111 17119
rect 26099 17088 27936 17116
rect 26099 17085 26111 17088
rect 26053 17079 26111 17085
rect 9456 17020 11008 17048
rect 18785 17051 18843 17057
rect 9456 17008 9462 17020
rect 18785 17017 18797 17051
rect 18831 17048 18843 17051
rect 20070 17048 20076 17060
rect 18831 17020 20076 17048
rect 18831 17017 18843 17020
rect 18785 17011 18843 17017
rect 20070 17008 20076 17020
rect 20128 17008 20134 17060
rect 26234 17048 26240 17060
rect 26195 17020 26240 17048
rect 26234 17008 26240 17020
rect 26292 17008 26298 17060
rect 26326 17008 26332 17060
rect 26384 17048 26390 17060
rect 26789 17051 26847 17057
rect 26789 17048 26801 17051
rect 26384 17020 26801 17048
rect 26384 17008 26390 17020
rect 26789 17017 26801 17020
rect 26835 17017 26847 17051
rect 26789 17011 26847 17017
rect 27908 16992 27936 17088
rect 5626 16940 5632 16992
rect 5684 16980 5690 16992
rect 6914 16980 6920 16992
rect 5684 16952 5729 16980
rect 6875 16952 6920 16980
rect 5684 16940 5690 16952
rect 6914 16940 6920 16952
rect 6972 16940 6978 16992
rect 7377 16983 7435 16989
rect 7377 16949 7389 16983
rect 7423 16980 7435 16983
rect 8294 16980 8300 16992
rect 7423 16952 8300 16980
rect 7423 16949 7435 16952
rect 7377 16943 7435 16949
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 11146 16980 11152 16992
rect 11107 16952 11152 16980
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 18322 16980 18328 16992
rect 18283 16952 18328 16980
rect 18322 16940 18328 16952
rect 18380 16940 18386 16992
rect 18414 16940 18420 16992
rect 18472 16980 18478 16992
rect 18693 16983 18751 16989
rect 18693 16980 18705 16983
rect 18472 16952 18705 16980
rect 18472 16940 18478 16952
rect 18693 16949 18705 16952
rect 18739 16949 18751 16983
rect 18693 16943 18751 16949
rect 21174 16940 21180 16992
rect 21232 16980 21238 16992
rect 21729 16983 21787 16989
rect 21729 16980 21741 16983
rect 21232 16952 21741 16980
rect 21232 16940 21238 16952
rect 21729 16949 21741 16952
rect 21775 16949 21787 16983
rect 21729 16943 21787 16949
rect 24394 16940 24400 16992
rect 24452 16980 24458 16992
rect 24762 16980 24768 16992
rect 24452 16952 24768 16980
rect 24452 16940 24458 16952
rect 24762 16940 24768 16952
rect 24820 16940 24826 16992
rect 27430 16980 27436 16992
rect 27391 16952 27436 16980
rect 27430 16940 27436 16952
rect 27488 16940 27494 16992
rect 27798 16980 27804 16992
rect 27759 16952 27804 16980
rect 27798 16940 27804 16952
rect 27856 16940 27862 16992
rect 27890 16940 27896 16992
rect 27948 16980 27954 16992
rect 27948 16952 27993 16980
rect 27948 16940 27954 16952
rect 1104 16890 28888 16912
rect 1104 16838 10246 16890
rect 10298 16838 10310 16890
rect 10362 16838 10374 16890
rect 10426 16838 10438 16890
rect 10490 16838 19510 16890
rect 19562 16838 19574 16890
rect 19626 16838 19638 16890
rect 19690 16838 19702 16890
rect 19754 16838 28888 16890
rect 1104 16816 28888 16838
rect 1762 16776 1768 16788
rect 1723 16748 1768 16776
rect 1762 16736 1768 16748
rect 1820 16736 1826 16788
rect 3053 16779 3111 16785
rect 3053 16745 3065 16779
rect 3099 16745 3111 16779
rect 3053 16739 3111 16745
rect 3881 16779 3939 16785
rect 3881 16745 3893 16779
rect 3927 16776 3939 16779
rect 4614 16776 4620 16788
rect 3927 16748 4620 16776
rect 3927 16745 3939 16748
rect 3881 16739 3939 16745
rect 2682 16708 2688 16720
rect 2424 16680 2688 16708
rect 1946 16640 1952 16652
rect 1907 16612 1952 16640
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 2424 16513 2452 16680
rect 2682 16668 2688 16680
rect 2740 16668 2746 16720
rect 3068 16708 3096 16739
rect 4614 16736 4620 16748
rect 4672 16736 4678 16788
rect 5077 16779 5135 16785
rect 5077 16745 5089 16779
rect 5123 16776 5135 16779
rect 5626 16776 5632 16788
rect 5123 16748 5632 16776
rect 5123 16745 5135 16748
rect 5077 16739 5135 16745
rect 5626 16736 5632 16748
rect 5684 16736 5690 16788
rect 5721 16779 5779 16785
rect 5721 16745 5733 16779
rect 5767 16776 5779 16779
rect 5902 16776 5908 16788
rect 5767 16748 5908 16776
rect 5767 16745 5779 16748
rect 5721 16739 5779 16745
rect 5902 16736 5908 16748
rect 5960 16736 5966 16788
rect 7466 16776 7472 16788
rect 6840 16748 7472 16776
rect 6840 16708 6868 16748
rect 7466 16736 7472 16748
rect 7524 16736 7530 16788
rect 8294 16776 8300 16788
rect 8207 16748 8300 16776
rect 8294 16736 8300 16748
rect 8352 16776 8358 16788
rect 9490 16776 9496 16788
rect 8352 16748 9496 16776
rect 8352 16736 8358 16748
rect 9490 16736 9496 16748
rect 9548 16736 9554 16788
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 10505 16779 10563 16785
rect 10505 16776 10517 16779
rect 10100 16748 10517 16776
rect 10100 16736 10106 16748
rect 10505 16745 10517 16748
rect 10551 16745 10563 16779
rect 10505 16739 10563 16745
rect 16209 16779 16267 16785
rect 16209 16745 16221 16779
rect 16255 16776 16267 16779
rect 17126 16776 17132 16788
rect 16255 16748 17132 16776
rect 16255 16745 16267 16748
rect 16209 16739 16267 16745
rect 17126 16736 17132 16748
rect 17184 16736 17190 16788
rect 3068 16680 6868 16708
rect 6914 16668 6920 16720
rect 6972 16708 6978 16720
rect 7162 16711 7220 16717
rect 7162 16708 7174 16711
rect 6972 16680 7174 16708
rect 6972 16668 6978 16680
rect 7162 16677 7174 16680
rect 7208 16677 7220 16711
rect 7162 16671 7220 16677
rect 14458 16668 14464 16720
rect 14516 16708 14522 16720
rect 15074 16711 15132 16717
rect 15074 16708 15086 16711
rect 14516 16680 15086 16708
rect 14516 16668 14522 16680
rect 15074 16677 15086 16680
rect 15120 16677 15132 16711
rect 15074 16671 15132 16677
rect 15930 16668 15936 16720
rect 15988 16708 15994 16720
rect 17954 16708 17960 16720
rect 15988 16680 17960 16708
rect 15988 16668 15994 16680
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 18322 16668 18328 16720
rect 18380 16708 18386 16720
rect 18754 16711 18812 16717
rect 18754 16708 18766 16711
rect 18380 16680 18766 16708
rect 18380 16668 18386 16680
rect 18754 16677 18766 16680
rect 18800 16677 18812 16711
rect 18754 16671 18812 16677
rect 20806 16668 20812 16720
rect 20864 16708 20870 16720
rect 20864 16680 21128 16708
rect 20864 16668 20870 16680
rect 2593 16643 2651 16649
rect 2593 16609 2605 16643
rect 2639 16640 2651 16643
rect 2774 16640 2780 16652
rect 2639 16612 2780 16640
rect 2639 16609 2651 16612
rect 2593 16603 2651 16609
rect 2774 16600 2780 16612
rect 2832 16600 2838 16652
rect 3234 16640 3240 16652
rect 3195 16612 3240 16640
rect 3234 16600 3240 16612
rect 3292 16600 3298 16652
rect 3326 16600 3332 16652
rect 3384 16640 3390 16652
rect 3697 16643 3755 16649
rect 3697 16640 3709 16643
rect 3384 16612 3709 16640
rect 3384 16600 3390 16612
rect 3697 16609 3709 16612
rect 3743 16609 3755 16643
rect 3697 16603 3755 16609
rect 4985 16643 5043 16649
rect 4985 16609 4997 16643
rect 5031 16609 5043 16643
rect 4985 16603 5043 16609
rect 5629 16643 5687 16649
rect 5629 16609 5641 16643
rect 5675 16640 5687 16643
rect 6822 16640 6828 16652
rect 5675 16612 6828 16640
rect 5675 16609 5687 16612
rect 5629 16603 5687 16609
rect 2409 16507 2467 16513
rect 2409 16473 2421 16507
rect 2455 16473 2467 16507
rect 2409 16467 2467 16473
rect 2590 16464 2596 16516
rect 2648 16504 2654 16516
rect 5000 16504 5028 16603
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 9398 16600 9404 16652
rect 9456 16640 9462 16652
rect 10321 16643 10379 16649
rect 10321 16640 10333 16643
rect 9456 16612 10333 16640
rect 9456 16600 9462 16612
rect 10321 16609 10333 16612
rect 10367 16609 10379 16643
rect 10321 16603 10379 16609
rect 14274 16600 14280 16652
rect 14332 16640 14338 16652
rect 14829 16643 14887 16649
rect 14829 16640 14841 16643
rect 14332 16612 14841 16640
rect 14332 16600 14338 16612
rect 14829 16609 14841 16612
rect 14875 16609 14887 16643
rect 17586 16640 17592 16652
rect 14829 16603 14887 16609
rect 14936 16612 15884 16640
rect 17547 16612 17592 16640
rect 6730 16532 6736 16584
rect 6788 16572 6794 16584
rect 6917 16575 6975 16581
rect 6917 16572 6929 16575
rect 6788 16544 6929 16572
rect 6788 16532 6794 16544
rect 6917 16541 6929 16544
rect 6963 16541 6975 16575
rect 6917 16535 6975 16541
rect 13078 16532 13084 16584
rect 13136 16572 13142 16584
rect 14936 16572 14964 16612
rect 13136 16544 14964 16572
rect 15856 16572 15884 16612
rect 17586 16600 17592 16612
rect 17644 16600 17650 16652
rect 17862 16640 17868 16652
rect 17696 16612 17868 16640
rect 17696 16581 17724 16612
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 18414 16640 18420 16652
rect 17972 16612 18420 16640
rect 17972 16581 18000 16612
rect 18414 16600 18420 16612
rect 18472 16600 18478 16652
rect 18509 16643 18567 16649
rect 18509 16609 18521 16643
rect 18555 16640 18567 16643
rect 19978 16640 19984 16652
rect 18555 16612 19984 16640
rect 18555 16609 18567 16612
rect 18509 16603 18567 16609
rect 19978 16600 19984 16612
rect 20036 16600 20042 16652
rect 20990 16640 20996 16652
rect 20951 16612 20996 16640
rect 20990 16600 20996 16612
rect 21048 16600 21054 16652
rect 17681 16575 17739 16581
rect 15856 16544 17540 16572
rect 13136 16532 13142 16544
rect 17512 16504 17540 16544
rect 17681 16541 17693 16575
rect 17727 16541 17739 16575
rect 17681 16535 17739 16541
rect 17957 16575 18015 16581
rect 17957 16541 17969 16575
rect 18003 16541 18015 16575
rect 20162 16572 20168 16584
rect 17957 16535 18015 16541
rect 19536 16544 20168 16572
rect 2648 16476 5028 16504
rect 2648 16464 2654 16476
rect 5000 16436 5028 16476
rect 7852 16476 12434 16504
rect 17512 16476 18092 16504
rect 7852 16436 7880 16476
rect 5000 16408 7880 16436
rect 12406 16436 12434 16476
rect 17218 16436 17224 16448
rect 12406 16408 17224 16436
rect 17218 16396 17224 16408
rect 17276 16396 17282 16448
rect 18064 16436 18092 16476
rect 19536 16436 19564 16544
rect 20162 16532 20168 16544
rect 20220 16532 20226 16584
rect 20898 16572 20904 16584
rect 20859 16544 20904 16572
rect 20898 16532 20904 16544
rect 20956 16532 20962 16584
rect 21100 16581 21128 16680
rect 21174 16668 21180 16720
rect 21232 16668 21238 16720
rect 24670 16668 24676 16720
rect 24728 16668 24734 16720
rect 24762 16668 24768 16720
rect 24820 16708 24826 16720
rect 26697 16711 26755 16717
rect 26697 16708 26709 16711
rect 24820 16680 26709 16708
rect 24820 16668 24826 16680
rect 26697 16677 26709 16680
rect 26743 16677 26755 16711
rect 26697 16671 26755 16677
rect 27706 16668 27712 16720
rect 27764 16708 27770 16720
rect 27985 16711 28043 16717
rect 27985 16708 27997 16711
rect 27764 16680 27997 16708
rect 27764 16668 27770 16680
rect 27985 16677 27997 16680
rect 28031 16677 28043 16711
rect 27985 16671 28043 16677
rect 21192 16581 21220 16668
rect 23566 16600 23572 16652
rect 23624 16640 23630 16652
rect 23845 16643 23903 16649
rect 23845 16640 23857 16643
rect 23624 16612 23857 16640
rect 23624 16600 23630 16612
rect 23845 16609 23857 16612
rect 23891 16609 23903 16643
rect 24026 16640 24032 16652
rect 23845 16603 23903 16609
rect 23952 16612 24032 16640
rect 21085 16575 21143 16581
rect 21085 16541 21097 16575
rect 21131 16541 21143 16575
rect 21085 16535 21143 16541
rect 21177 16575 21235 16581
rect 21177 16541 21189 16575
rect 21223 16541 21235 16575
rect 21177 16535 21235 16541
rect 22646 16532 22652 16584
rect 22704 16572 22710 16584
rect 23106 16572 23112 16584
rect 22704 16544 23112 16572
rect 22704 16532 22710 16544
rect 23106 16532 23112 16544
rect 23164 16532 23170 16584
rect 23952 16581 23980 16612
rect 24026 16600 24032 16612
rect 24084 16640 24090 16652
rect 24688 16640 24716 16668
rect 24084 16612 24716 16640
rect 24940 16643 24998 16649
rect 24084 16600 24090 16612
rect 24940 16609 24952 16643
rect 24986 16640 24998 16643
rect 25222 16640 25228 16652
rect 24986 16612 25228 16640
rect 24986 16609 24998 16612
rect 24940 16603 24998 16609
rect 25222 16600 25228 16612
rect 25280 16600 25286 16652
rect 26878 16640 26884 16652
rect 26839 16612 26884 16640
rect 26878 16600 26884 16612
rect 26936 16600 26942 16652
rect 28166 16640 28172 16652
rect 28127 16612 28172 16640
rect 28166 16600 28172 16612
rect 28224 16600 28230 16652
rect 23937 16575 23995 16581
rect 23937 16541 23949 16575
rect 23983 16541 23995 16575
rect 24210 16572 24216 16584
rect 24171 16544 24216 16572
rect 23937 16535 23995 16541
rect 24210 16532 24216 16544
rect 24268 16532 24274 16584
rect 24673 16575 24731 16581
rect 24673 16541 24685 16575
rect 24719 16541 24731 16575
rect 24673 16535 24731 16541
rect 22278 16464 22284 16516
rect 22336 16504 22342 16516
rect 24394 16504 24400 16516
rect 22336 16476 24400 16504
rect 22336 16464 22342 16476
rect 24394 16464 24400 16476
rect 24452 16464 24458 16516
rect 18064 16408 19564 16436
rect 19889 16439 19947 16445
rect 19889 16405 19901 16439
rect 19935 16436 19947 16439
rect 20070 16436 20076 16448
rect 19935 16408 20076 16436
rect 19935 16405 19947 16408
rect 19889 16399 19947 16405
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 20714 16436 20720 16448
rect 20675 16408 20720 16436
rect 20714 16396 20720 16408
rect 20772 16396 20778 16448
rect 24688 16436 24716 16535
rect 24854 16436 24860 16448
rect 24688 16408 24860 16436
rect 24854 16396 24860 16408
rect 24912 16396 24918 16448
rect 25682 16396 25688 16448
rect 25740 16436 25746 16448
rect 26053 16439 26111 16445
rect 26053 16436 26065 16439
rect 25740 16408 26065 16436
rect 25740 16396 25746 16408
rect 26053 16405 26065 16408
rect 26099 16405 26111 16439
rect 26053 16399 26111 16405
rect 1104 16346 28888 16368
rect 1104 16294 5614 16346
rect 5666 16294 5678 16346
rect 5730 16294 5742 16346
rect 5794 16294 5806 16346
rect 5858 16294 14878 16346
rect 14930 16294 14942 16346
rect 14994 16294 15006 16346
rect 15058 16294 15070 16346
rect 15122 16294 24142 16346
rect 24194 16294 24206 16346
rect 24258 16294 24270 16346
rect 24322 16294 24334 16346
rect 24386 16294 28888 16346
rect 1104 16272 28888 16294
rect 4982 16232 4988 16244
rect 4943 16204 4988 16232
rect 4982 16192 4988 16204
rect 5040 16192 5046 16244
rect 12158 16192 12164 16244
rect 12216 16232 12222 16244
rect 15562 16232 15568 16244
rect 12216 16204 15568 16232
rect 12216 16192 12222 16204
rect 15562 16192 15568 16204
rect 15620 16192 15626 16244
rect 16945 16235 17003 16241
rect 16945 16201 16957 16235
rect 16991 16232 17003 16235
rect 17586 16232 17592 16244
rect 16991 16204 17592 16232
rect 16991 16201 17003 16204
rect 16945 16195 17003 16201
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 18414 16192 18420 16244
rect 18472 16232 18478 16244
rect 18966 16232 18972 16244
rect 18472 16204 18972 16232
rect 18472 16192 18478 16204
rect 18966 16192 18972 16204
rect 19024 16192 19030 16244
rect 19429 16235 19487 16241
rect 19429 16201 19441 16235
rect 19475 16232 19487 16235
rect 21634 16232 21640 16244
rect 19475 16204 21220 16232
rect 21595 16204 21640 16232
rect 19475 16201 19487 16204
rect 19429 16195 19487 16201
rect 3145 16167 3203 16173
rect 3145 16133 3157 16167
rect 3191 16164 3203 16167
rect 4246 16164 4252 16176
rect 3191 16136 4252 16164
rect 3191 16133 3203 16136
rect 3145 16127 3203 16133
rect 4246 16124 4252 16136
rect 4304 16124 4310 16176
rect 5902 16164 5908 16176
rect 4908 16136 5908 16164
rect 1854 16028 1860 16040
rect 1815 16000 1860 16028
rect 1854 15988 1860 16000
rect 1912 15988 1918 16040
rect 4908 16037 4936 16136
rect 5902 16124 5908 16136
rect 5960 16164 5966 16176
rect 15102 16164 15108 16176
rect 5960 16136 15108 16164
rect 5960 16124 5966 16136
rect 15102 16124 15108 16136
rect 15160 16124 15166 16176
rect 20162 16164 20168 16176
rect 16776 16136 20168 16164
rect 10796 16068 15424 16096
rect 4893 16031 4951 16037
rect 4893 15997 4905 16031
rect 4939 15997 4951 16031
rect 4893 15991 4951 15997
rect 5166 15988 5172 16040
rect 5224 16028 5230 16040
rect 10796 16037 10824 16068
rect 10781 16031 10839 16037
rect 10781 16028 10793 16031
rect 5224 16000 10793 16028
rect 5224 15988 5230 16000
rect 10781 15997 10793 16000
rect 10827 15997 10839 16031
rect 10781 15991 10839 15997
rect 13449 16031 13507 16037
rect 13449 15997 13461 16031
rect 13495 16028 13507 16031
rect 15194 16028 15200 16040
rect 13495 16000 15200 16028
rect 13495 15997 13507 16000
rect 13449 15991 13507 15997
rect 15194 15988 15200 16000
rect 15252 15988 15258 16040
rect 15396 16028 15424 16068
rect 15838 16056 15844 16108
rect 15896 16056 15902 16108
rect 16776 16028 16804 16136
rect 20162 16124 20168 16136
rect 20220 16124 20226 16176
rect 21192 16164 21220 16204
rect 21634 16192 21640 16204
rect 21692 16192 21698 16244
rect 22278 16232 22284 16244
rect 21744 16204 22284 16232
rect 21744 16164 21772 16204
rect 22278 16192 22284 16204
rect 22336 16192 22342 16244
rect 23566 16232 23572 16244
rect 23527 16204 23572 16232
rect 23566 16192 23572 16204
rect 23624 16192 23630 16244
rect 25222 16232 25228 16244
rect 25183 16204 25228 16232
rect 25222 16192 25228 16204
rect 25280 16192 25286 16244
rect 26786 16192 26792 16244
rect 26844 16232 26850 16244
rect 26881 16235 26939 16241
rect 26881 16232 26893 16235
rect 26844 16204 26893 16232
rect 26844 16192 26850 16204
rect 26881 16201 26893 16204
rect 26927 16201 26939 16235
rect 26881 16195 26939 16201
rect 27982 16164 27988 16176
rect 21192 16136 21772 16164
rect 24228 16136 27988 16164
rect 17218 16056 17224 16108
rect 17276 16096 17282 16108
rect 17276 16068 20392 16096
rect 17276 16056 17282 16068
rect 15396 16000 16804 16028
rect 17126 15988 17132 16040
rect 17184 16028 17190 16040
rect 17497 16031 17555 16037
rect 17497 16028 17509 16031
rect 17184 16000 17509 16028
rect 17184 15988 17190 16000
rect 17497 15997 17509 16000
rect 17543 15997 17555 16031
rect 17497 15991 17555 15997
rect 17589 16031 17647 16037
rect 17589 15997 17601 16031
rect 17635 16028 17647 16031
rect 17954 16028 17960 16040
rect 17635 16000 17960 16028
rect 17635 15997 17647 16000
rect 17589 15991 17647 15997
rect 17954 15988 17960 16000
rect 18012 15988 18018 16040
rect 18322 15988 18328 16040
rect 18380 16028 18386 16040
rect 19429 16031 19487 16037
rect 19429 16028 19441 16031
rect 18380 16000 19441 16028
rect 18380 15988 18386 16000
rect 19429 15997 19441 16000
rect 19475 15997 19487 16031
rect 19429 15991 19487 15997
rect 19978 15988 19984 16040
rect 20036 16028 20042 16040
rect 20257 16031 20315 16037
rect 20257 16028 20269 16031
rect 20036 16000 20269 16028
rect 20036 15988 20042 16000
rect 20257 15997 20269 16000
rect 20303 15997 20315 16031
rect 20364 16028 20392 16068
rect 22554 16056 22560 16108
rect 22612 16056 22618 16108
rect 22646 16028 22652 16040
rect 20364 16000 20852 16028
rect 22607 16000 22652 16028
rect 20257 15991 20315 15997
rect 2777 15963 2835 15969
rect 2777 15929 2789 15963
rect 2823 15960 2835 15963
rect 2958 15960 2964 15972
rect 2823 15932 2964 15960
rect 2823 15929 2835 15932
rect 2777 15923 2835 15929
rect 2958 15920 2964 15932
rect 3016 15920 3022 15972
rect 5074 15920 5080 15972
rect 5132 15960 5138 15972
rect 15930 15960 15936 15972
rect 5132 15932 15792 15960
rect 15891 15932 15936 15960
rect 5132 15920 5138 15932
rect 1946 15892 1952 15904
rect 1907 15864 1952 15892
rect 1946 15852 1952 15864
rect 2004 15852 2010 15904
rect 3237 15895 3295 15901
rect 3237 15861 3249 15895
rect 3283 15892 3295 15895
rect 3694 15892 3700 15904
rect 3283 15864 3700 15892
rect 3283 15861 3295 15864
rect 3237 15855 3295 15861
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 10870 15892 10876 15904
rect 10831 15864 10876 15892
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 11422 15852 11428 15904
rect 11480 15892 11486 15904
rect 13078 15892 13084 15904
rect 11480 15864 13084 15892
rect 11480 15852 11486 15864
rect 13078 15852 13084 15864
rect 13136 15852 13142 15904
rect 13262 15892 13268 15904
rect 13223 15864 13268 15892
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 15562 15852 15568 15904
rect 15620 15892 15626 15904
rect 15657 15895 15715 15901
rect 15657 15892 15669 15895
rect 15620 15864 15669 15892
rect 15620 15852 15626 15864
rect 15657 15861 15669 15864
rect 15703 15861 15715 15895
rect 15764 15892 15792 15932
rect 15930 15920 15936 15932
rect 15988 15920 15994 15972
rect 16025 15963 16083 15969
rect 16025 15929 16037 15963
rect 16071 15960 16083 15963
rect 16114 15960 16120 15972
rect 16071 15932 16120 15960
rect 16071 15929 16083 15932
rect 16025 15923 16083 15929
rect 16114 15920 16120 15932
rect 16172 15920 16178 15972
rect 16393 15963 16451 15969
rect 16393 15929 16405 15963
rect 16439 15960 16451 15963
rect 18966 15960 18972 15972
rect 16439 15932 18972 15960
rect 16439 15929 16451 15932
rect 16393 15923 16451 15929
rect 18966 15920 18972 15932
rect 19024 15920 19030 15972
rect 20524 15963 20582 15969
rect 20524 15929 20536 15963
rect 20570 15960 20582 15963
rect 20714 15960 20720 15972
rect 20570 15932 20720 15960
rect 20570 15929 20582 15932
rect 20524 15923 20582 15929
rect 20714 15920 20720 15932
rect 20772 15920 20778 15972
rect 20824 15960 20852 16000
rect 22646 15988 22652 16000
rect 22704 16028 22710 16040
rect 22922 16028 22928 16040
rect 22704 16000 22928 16028
rect 22704 15988 22710 16000
rect 22922 15988 22928 16000
rect 22980 15988 22986 16040
rect 23017 16031 23075 16037
rect 23017 15997 23029 16031
rect 23063 16028 23075 16031
rect 23106 16028 23112 16040
rect 23063 16000 23112 16028
rect 23063 15997 23075 16000
rect 23017 15991 23075 15997
rect 23106 15988 23112 16000
rect 23164 15988 23170 16040
rect 24228 16028 24256 16136
rect 27982 16124 27988 16136
rect 28040 16124 28046 16176
rect 25774 16096 25780 16108
rect 25735 16068 25780 16096
rect 25774 16056 25780 16068
rect 25832 16096 25838 16108
rect 25832 16068 26280 16096
rect 25832 16056 25838 16068
rect 26252 16040 26280 16068
rect 23308 16000 24256 16028
rect 22557 15963 22615 15969
rect 20824 15932 22508 15960
rect 16761 15895 16819 15901
rect 16761 15892 16773 15895
rect 15764 15864 16773 15892
rect 15657 15855 15715 15861
rect 16761 15861 16773 15864
rect 16807 15861 16819 15895
rect 16761 15855 16819 15861
rect 17218 15852 17224 15904
rect 17276 15892 17282 15904
rect 17494 15892 17500 15904
rect 17276 15864 17500 15892
rect 17276 15852 17282 15864
rect 17494 15852 17500 15864
rect 17552 15852 17558 15904
rect 17954 15852 17960 15904
rect 18012 15892 18018 15904
rect 20254 15892 20260 15904
rect 18012 15864 20260 15892
rect 18012 15852 18018 15864
rect 20254 15852 20260 15864
rect 20312 15852 20318 15904
rect 22278 15892 22284 15904
rect 22239 15864 22284 15892
rect 22278 15852 22284 15864
rect 22336 15852 22342 15904
rect 22480 15892 22508 15932
rect 22557 15929 22569 15963
rect 22603 15960 22615 15963
rect 22738 15960 22744 15972
rect 22603 15932 22744 15960
rect 22603 15929 22615 15932
rect 22557 15923 22615 15929
rect 22738 15920 22744 15932
rect 22796 15960 22802 15972
rect 23308 15960 23336 16000
rect 24946 15988 24952 16040
rect 25004 16028 25010 16040
rect 25593 16031 25651 16037
rect 25593 16028 25605 16031
rect 25004 16000 25605 16028
rect 25004 15988 25010 16000
rect 25593 15997 25605 16000
rect 25639 15997 25651 16031
rect 25593 15991 25651 15997
rect 25682 15988 25688 16040
rect 25740 16028 25746 16040
rect 25740 16000 25785 16028
rect 25740 15988 25746 16000
rect 26234 15988 26240 16040
rect 26292 15988 26298 16040
rect 26510 15988 26516 16040
rect 26568 16028 26574 16040
rect 26697 16031 26755 16037
rect 26697 16028 26709 16031
rect 26568 16000 26709 16028
rect 26568 15988 26574 16000
rect 26697 15997 26709 16000
rect 26743 15997 26755 16031
rect 27246 16028 27252 16040
rect 27207 16000 27252 16028
rect 26697 15991 26755 15997
rect 27246 15988 27252 16000
rect 27304 15988 27310 16040
rect 27522 16028 27528 16040
rect 27483 16000 27528 16028
rect 27522 15988 27528 16000
rect 27580 15988 27586 16040
rect 22796 15932 23336 15960
rect 22796 15920 22802 15932
rect 25498 15920 25504 15972
rect 25556 15960 25562 15972
rect 25866 15960 25872 15972
rect 25556 15932 25872 15960
rect 25556 15920 25562 15932
rect 25866 15920 25872 15932
rect 25924 15920 25930 15972
rect 23385 15895 23443 15901
rect 23385 15892 23397 15895
rect 22480 15864 23397 15892
rect 23385 15861 23397 15864
rect 23431 15861 23443 15895
rect 23385 15855 23443 15861
rect 1104 15802 28888 15824
rect 1104 15750 10246 15802
rect 10298 15750 10310 15802
rect 10362 15750 10374 15802
rect 10426 15750 10438 15802
rect 10490 15750 19510 15802
rect 19562 15750 19574 15802
rect 19626 15750 19638 15802
rect 19690 15750 19702 15802
rect 19754 15750 28888 15802
rect 1104 15728 28888 15750
rect 4985 15691 5043 15697
rect 4985 15657 4997 15691
rect 5031 15688 5043 15691
rect 5074 15688 5080 15700
rect 5031 15660 5080 15688
rect 5031 15657 5043 15660
rect 4985 15651 5043 15657
rect 5074 15648 5080 15660
rect 5132 15648 5138 15700
rect 5442 15648 5448 15700
rect 5500 15688 5506 15700
rect 20073 15691 20131 15697
rect 20073 15688 20085 15691
rect 5500 15660 20085 15688
rect 5500 15648 5506 15660
rect 20073 15657 20085 15660
rect 20119 15657 20131 15691
rect 20073 15651 20131 15657
rect 20162 15648 20168 15700
rect 20220 15688 20226 15700
rect 26237 15691 26295 15697
rect 26237 15688 26249 15691
rect 20220 15660 26249 15688
rect 20220 15648 20226 15660
rect 26237 15657 26249 15660
rect 26283 15657 26295 15691
rect 26418 15688 26424 15700
rect 26331 15660 26424 15688
rect 26237 15651 26295 15657
rect 26418 15648 26424 15660
rect 26476 15688 26482 15700
rect 27522 15688 27528 15700
rect 26476 15660 27528 15688
rect 26476 15648 26482 15660
rect 27522 15648 27528 15660
rect 27580 15648 27586 15700
rect 1854 15620 1860 15632
rect 1815 15592 1860 15620
rect 1854 15580 1860 15592
rect 1912 15580 1918 15632
rect 2041 15623 2099 15629
rect 2041 15589 2053 15623
rect 2087 15620 2099 15623
rect 2590 15620 2596 15632
rect 2087 15592 2596 15620
rect 2087 15589 2099 15592
rect 2041 15583 2099 15589
rect 1578 15512 1584 15564
rect 1636 15552 1642 15564
rect 2056 15552 2084 15583
rect 2590 15580 2596 15592
rect 2648 15580 2654 15632
rect 3878 15580 3884 15632
rect 3936 15620 3942 15632
rect 4065 15623 4123 15629
rect 4065 15620 4077 15623
rect 3936 15592 4077 15620
rect 3936 15580 3942 15592
rect 4065 15589 4077 15592
rect 4111 15589 4123 15623
rect 4065 15583 4123 15589
rect 4430 15580 4436 15632
rect 4488 15580 4494 15632
rect 4614 15580 4620 15632
rect 4672 15620 4678 15632
rect 5460 15620 5488 15648
rect 4672 15592 5488 15620
rect 4672 15580 4678 15592
rect 10686 15580 10692 15632
rect 10744 15620 10750 15632
rect 10965 15623 11023 15629
rect 10965 15620 10977 15623
rect 10744 15592 10977 15620
rect 10744 15580 10750 15592
rect 10965 15589 10977 15592
rect 11011 15589 11023 15623
rect 10965 15583 11023 15589
rect 11054 15580 11060 15632
rect 11112 15620 11118 15632
rect 11974 15620 11980 15632
rect 11112 15592 11980 15620
rect 11112 15580 11118 15592
rect 11974 15580 11980 15592
rect 12032 15580 12038 15632
rect 12084 15592 12480 15620
rect 2958 15552 2964 15564
rect 1636 15524 2084 15552
rect 2919 15524 2964 15552
rect 1636 15512 1642 15524
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 3970 15552 3976 15564
rect 3436 15524 3976 15552
rect 3436 15493 3464 15524
rect 3970 15512 3976 15524
rect 4028 15512 4034 15564
rect 4246 15552 4252 15564
rect 4080 15524 4252 15552
rect 3421 15487 3479 15493
rect 3421 15453 3433 15487
rect 3467 15453 3479 15487
rect 3421 15447 3479 15453
rect 3237 15351 3295 15357
rect 3237 15317 3249 15351
rect 3283 15348 3295 15351
rect 4080 15348 4108 15524
rect 4246 15512 4252 15524
rect 4304 15512 4310 15564
rect 4341 15555 4399 15561
rect 4341 15521 4353 15555
rect 4387 15552 4399 15555
rect 4448 15552 4476 15580
rect 4801 15555 4859 15561
rect 4387 15524 4660 15552
rect 4387 15521 4399 15524
rect 4341 15515 4399 15521
rect 4632 15496 4660 15524
rect 4801 15521 4813 15555
rect 4847 15521 4859 15555
rect 4801 15515 4859 15521
rect 8564 15555 8622 15561
rect 8564 15521 8576 15555
rect 8610 15552 8622 15555
rect 9490 15552 9496 15564
rect 8610 15524 9496 15552
rect 8610 15521 8622 15524
rect 8564 15515 8622 15521
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 4430 15484 4436 15496
rect 4203 15456 4436 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 4430 15444 4436 15456
rect 4488 15444 4494 15496
rect 4614 15444 4620 15496
rect 4672 15444 4678 15496
rect 4816 15416 4844 15515
rect 9490 15512 9496 15524
rect 9548 15512 9554 15564
rect 12084 15561 12112 15592
rect 12069 15555 12127 15561
rect 12069 15521 12081 15555
rect 12115 15521 12127 15555
rect 12069 15515 12127 15521
rect 12158 15512 12164 15564
rect 12216 15552 12222 15564
rect 12325 15555 12383 15561
rect 12325 15552 12337 15555
rect 12216 15524 12337 15552
rect 12216 15512 12222 15524
rect 12325 15521 12337 15524
rect 12371 15521 12383 15555
rect 12452 15552 12480 15592
rect 15562 15580 15568 15632
rect 15620 15620 15626 15632
rect 17954 15620 17960 15632
rect 15620 15592 17960 15620
rect 15620 15580 15626 15592
rect 17954 15580 17960 15592
rect 18012 15580 18018 15632
rect 18966 15620 18972 15632
rect 18927 15592 18972 15620
rect 18966 15580 18972 15592
rect 19024 15580 19030 15632
rect 19058 15580 19064 15632
rect 19116 15620 19122 15632
rect 19334 15629 19340 15632
rect 19224 15623 19282 15629
rect 19224 15620 19236 15623
rect 19116 15592 19236 15620
rect 19116 15580 19122 15592
rect 19224 15589 19236 15592
rect 19270 15589 19282 15623
rect 19224 15583 19282 15589
rect 19325 15623 19340 15629
rect 19325 15589 19337 15623
rect 19325 15583 19340 15589
rect 19334 15580 19340 15583
rect 19392 15580 19398 15632
rect 21634 15580 21640 15632
rect 21692 15620 21698 15632
rect 23106 15620 23112 15632
rect 21692 15592 23112 15620
rect 21692 15580 21698 15592
rect 23106 15580 23112 15592
rect 23164 15620 23170 15632
rect 24762 15620 24768 15632
rect 23164 15592 24768 15620
rect 23164 15580 23170 15592
rect 24762 15580 24768 15592
rect 24820 15620 24826 15632
rect 25133 15623 25191 15629
rect 25133 15620 25145 15623
rect 24820 15592 25145 15620
rect 24820 15580 24826 15592
rect 25133 15589 25145 15592
rect 25179 15589 25191 15623
rect 25133 15583 25191 15589
rect 25222 15580 25228 15632
rect 25280 15620 25286 15632
rect 25409 15623 25467 15629
rect 25409 15620 25421 15623
rect 25280 15592 25421 15620
rect 25280 15580 25286 15592
rect 25409 15589 25421 15592
rect 25455 15589 25467 15623
rect 25409 15583 25467 15589
rect 25501 15623 25559 15629
rect 25501 15589 25513 15623
rect 25547 15620 25559 15623
rect 25590 15620 25596 15632
rect 25547 15592 25596 15620
rect 25547 15589 25559 15592
rect 25501 15583 25559 15589
rect 12452 15524 13400 15552
rect 12325 15515 12383 15521
rect 8294 15484 8300 15496
rect 8255 15456 8300 15484
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 10962 15484 10968 15496
rect 10923 15456 10968 15484
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 13372 15484 13400 15524
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 14165 15555 14223 15561
rect 14165 15552 14177 15555
rect 13872 15524 14177 15552
rect 13872 15512 13878 15524
rect 14165 15521 14177 15524
rect 14211 15521 14223 15555
rect 14165 15515 14223 15521
rect 15470 15512 15476 15564
rect 15528 15552 15534 15564
rect 16025 15555 16083 15561
rect 16025 15552 16037 15555
rect 15528 15524 16037 15552
rect 15528 15512 15534 15524
rect 16025 15521 16037 15524
rect 16071 15552 16083 15555
rect 16298 15552 16304 15564
rect 16071 15524 16304 15552
rect 16071 15521 16083 15524
rect 16025 15515 16083 15521
rect 16298 15512 16304 15524
rect 16356 15512 16362 15564
rect 16666 15512 16672 15564
rect 16724 15552 16730 15564
rect 17126 15552 17132 15564
rect 16724 15524 17132 15552
rect 16724 15512 16730 15524
rect 17126 15512 17132 15524
rect 17184 15512 17190 15564
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15552 19763 15555
rect 20070 15552 20076 15564
rect 19751 15524 20076 15552
rect 19751 15521 19763 15524
rect 19705 15515 19763 15521
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 20254 15512 20260 15564
rect 20312 15552 20318 15564
rect 22738 15552 22744 15564
rect 20312 15524 22744 15552
rect 20312 15512 20318 15524
rect 22738 15512 22744 15524
rect 22796 15512 22802 15564
rect 25424 15552 25452 15583
rect 25590 15580 25596 15592
rect 25648 15580 25654 15632
rect 25682 15580 25688 15632
rect 25740 15620 25746 15632
rect 25869 15623 25927 15629
rect 25869 15620 25881 15623
rect 25740 15592 25881 15620
rect 25740 15580 25746 15592
rect 25869 15589 25881 15592
rect 25915 15589 25927 15623
rect 25869 15583 25927 15589
rect 27985 15555 28043 15561
rect 27985 15552 27997 15555
rect 25424 15524 27997 15552
rect 27985 15521 27997 15524
rect 28031 15521 28043 15555
rect 27985 15515 28043 15521
rect 13906 15484 13912 15496
rect 13372 15456 13912 15484
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 15194 15444 15200 15496
rect 15252 15484 15258 15496
rect 15930 15484 15936 15496
rect 15252 15456 15936 15484
rect 15252 15444 15258 15456
rect 15930 15444 15936 15456
rect 15988 15444 15994 15496
rect 18690 15444 18696 15496
rect 18748 15484 18754 15496
rect 20088 15484 20116 15512
rect 22278 15484 22284 15496
rect 18748 15470 18814 15484
rect 18748 15456 18828 15470
rect 20088 15456 22284 15484
rect 18748 15444 18754 15456
rect 4172 15388 4844 15416
rect 10505 15419 10563 15425
rect 4172 15360 4200 15388
rect 10505 15385 10517 15419
rect 10551 15416 10563 15419
rect 11422 15416 11428 15428
rect 10551 15388 11428 15416
rect 10551 15385 10563 15388
rect 10505 15379 10563 15385
rect 11422 15376 11428 15388
rect 11480 15376 11486 15428
rect 13078 15376 13084 15428
rect 13136 15416 13142 15428
rect 13136 15388 13581 15416
rect 13136 15376 13142 15388
rect 3283 15320 4108 15348
rect 3283 15317 3295 15320
rect 3237 15311 3295 15317
rect 4154 15308 4160 15360
rect 4212 15308 4218 15360
rect 4338 15348 4344 15360
rect 4299 15320 4344 15348
rect 4338 15308 4344 15320
rect 4396 15308 4402 15360
rect 9674 15348 9680 15360
rect 9635 15320 9680 15348
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 12342 15308 12348 15360
rect 12400 15348 12406 15360
rect 13449 15351 13507 15357
rect 13449 15348 13461 15351
rect 12400 15320 13461 15348
rect 12400 15308 12406 15320
rect 13449 15317 13461 15320
rect 13495 15317 13507 15351
rect 13553 15348 13581 15388
rect 14844 15388 15424 15416
rect 14844 15348 14872 15388
rect 13553 15320 14872 15348
rect 13449 15311 13507 15317
rect 15194 15308 15200 15360
rect 15252 15348 15258 15360
rect 15289 15351 15347 15357
rect 15289 15348 15301 15351
rect 15252 15320 15301 15348
rect 15252 15308 15258 15320
rect 15289 15317 15301 15320
rect 15335 15317 15347 15351
rect 15396 15348 15424 15388
rect 15562 15376 15568 15428
rect 15620 15416 15626 15428
rect 16114 15416 16120 15428
rect 15620 15388 16120 15416
rect 15620 15376 15626 15388
rect 16114 15376 16120 15388
rect 16172 15376 16178 15428
rect 16209 15419 16267 15425
rect 16209 15385 16221 15419
rect 16255 15416 16267 15419
rect 18322 15416 18328 15428
rect 16255 15388 18328 15416
rect 16255 15385 16267 15388
rect 16209 15379 16267 15385
rect 16224 15348 16252 15379
rect 18322 15376 18328 15388
rect 18380 15376 18386 15428
rect 15396 15320 16252 15348
rect 18800 15348 18828 15456
rect 22278 15444 22284 15456
rect 22336 15484 22342 15496
rect 23842 15484 23848 15496
rect 22336 15456 23848 15484
rect 22336 15444 22342 15456
rect 23842 15444 23848 15456
rect 23900 15444 23906 15496
rect 25498 15444 25504 15496
rect 25556 15444 25562 15496
rect 20257 15419 20315 15425
rect 20257 15385 20269 15419
rect 20303 15416 20315 15419
rect 20530 15416 20536 15428
rect 20303 15388 20536 15416
rect 20303 15385 20315 15388
rect 20257 15379 20315 15385
rect 20530 15376 20536 15388
rect 20588 15376 20594 15428
rect 23474 15376 23480 15428
rect 23532 15416 23538 15428
rect 24486 15416 24492 15428
rect 23532 15388 24492 15416
rect 23532 15376 23538 15388
rect 24486 15376 24492 15388
rect 24544 15376 24550 15428
rect 18966 15348 18972 15360
rect 18800 15320 18972 15348
rect 15289 15311 15347 15317
rect 18966 15308 18972 15320
rect 19024 15308 19030 15360
rect 27522 15308 27528 15360
rect 27580 15348 27586 15360
rect 28077 15351 28135 15357
rect 28077 15348 28089 15351
rect 27580 15320 28089 15348
rect 27580 15308 27586 15320
rect 28077 15317 28089 15320
rect 28123 15317 28135 15351
rect 28077 15311 28135 15317
rect 1104 15258 28888 15280
rect 1104 15206 5614 15258
rect 5666 15206 5678 15258
rect 5730 15206 5742 15258
rect 5794 15206 5806 15258
rect 5858 15206 14878 15258
rect 14930 15206 14942 15258
rect 14994 15206 15006 15258
rect 15058 15206 15070 15258
rect 15122 15206 24142 15258
rect 24194 15206 24206 15258
rect 24258 15206 24270 15258
rect 24322 15206 24334 15258
rect 24386 15206 28888 15258
rect 1104 15184 28888 15206
rect 2774 15104 2780 15156
rect 2832 15144 2838 15156
rect 2869 15147 2927 15153
rect 2869 15144 2881 15147
rect 2832 15116 2881 15144
rect 2832 15104 2838 15116
rect 2869 15113 2881 15116
rect 2915 15113 2927 15147
rect 2869 15107 2927 15113
rect 6822 15104 6828 15156
rect 6880 15144 6886 15156
rect 7009 15147 7067 15153
rect 7009 15144 7021 15147
rect 6880 15116 7021 15144
rect 6880 15104 6886 15116
rect 7009 15113 7021 15116
rect 7055 15113 7067 15147
rect 9490 15144 9496 15156
rect 9451 15116 9496 15144
rect 7009 15107 7067 15113
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 10686 15144 10692 15156
rect 10647 15116 10692 15144
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 12069 15147 12127 15153
rect 12069 15113 12081 15147
rect 12115 15144 12127 15147
rect 12158 15144 12164 15156
rect 12115 15116 12164 15144
rect 12115 15113 12127 15116
rect 12069 15107 12127 15113
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 13173 15147 13231 15153
rect 13173 15113 13185 15147
rect 13219 15144 13231 15147
rect 13814 15144 13820 15156
rect 13219 15116 13820 15144
rect 13219 15113 13231 15116
rect 13173 15107 13231 15113
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 15838 15104 15844 15156
rect 15896 15144 15902 15156
rect 16114 15144 16120 15156
rect 15896 15116 16120 15144
rect 15896 15104 15902 15116
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 17678 15144 17684 15156
rect 17639 15116 17684 15144
rect 17678 15104 17684 15116
rect 17736 15104 17742 15156
rect 21910 15144 21916 15156
rect 21871 15116 21916 15144
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 26329 15147 26387 15153
rect 26329 15113 26341 15147
rect 26375 15144 26387 15147
rect 27798 15144 27804 15156
rect 26375 15116 27804 15144
rect 26375 15113 26387 15116
rect 26329 15107 26387 15113
rect 27798 15104 27804 15116
rect 27856 15104 27862 15156
rect 27890 15104 27896 15156
rect 27948 15144 27954 15156
rect 28169 15147 28227 15153
rect 28169 15144 28181 15147
rect 27948 15116 28181 15144
rect 27948 15104 27954 15116
rect 28169 15113 28181 15116
rect 28215 15113 28227 15147
rect 28169 15107 28227 15113
rect 5074 15076 5080 15088
rect 2884 15048 5080 15076
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 1762 14900 1768 14952
rect 1820 14900 1826 14952
rect 1857 14943 1915 14949
rect 1857 14909 1869 14943
rect 1903 14940 1915 14943
rect 2317 14943 2375 14949
rect 1903 14912 2268 14940
rect 1903 14909 1915 14912
rect 1857 14903 1915 14909
rect 1578 14872 1584 14884
rect 1539 14844 1584 14872
rect 1578 14832 1584 14844
rect 1636 14832 1642 14884
rect 1780 14872 1808 14900
rect 1937 14875 1995 14881
rect 1937 14872 1949 14875
rect 1780 14844 1949 14872
rect 1937 14841 1949 14844
rect 1983 14841 1995 14875
rect 2240 14872 2268 14912
rect 2317 14909 2329 14943
rect 2363 14940 2375 14943
rect 2498 14940 2504 14952
rect 2363 14912 2504 14940
rect 2363 14909 2375 14912
rect 2317 14903 2375 14909
rect 2498 14900 2504 14912
rect 2556 14900 2562 14952
rect 2884 14940 2912 15048
rect 5074 15036 5080 15048
rect 5132 15036 5138 15088
rect 12526 15036 12532 15088
rect 12584 15076 12590 15088
rect 12584 15048 12756 15076
rect 12584 15036 12590 15048
rect 5092 14952 5120 14994
rect 6638 14968 6644 15020
rect 6696 15008 6702 15020
rect 7561 15011 7619 15017
rect 7561 15008 7573 15011
rect 6696 14980 7573 15008
rect 6696 14968 6702 14980
rect 7561 14977 7573 14980
rect 7607 14977 7619 15011
rect 10042 15008 10048 15020
rect 10003 14980 10048 15008
rect 7561 14971 7619 14977
rect 10042 14968 10048 14980
rect 10100 14968 10106 15020
rect 10870 14968 10876 15020
rect 10928 15008 10934 15020
rect 11149 15011 11207 15017
rect 11149 15008 11161 15011
rect 10928 14980 11161 15008
rect 10928 14968 10934 14980
rect 11149 14977 11161 14980
rect 11195 14977 11207 15011
rect 11149 14971 11207 14977
rect 11238 14968 11244 15020
rect 11296 15008 11302 15020
rect 11333 15011 11391 15017
rect 11333 15008 11345 15011
rect 11296 14980 11345 15008
rect 11296 14968 11302 14980
rect 11333 14977 11345 14980
rect 11379 15008 11391 15011
rect 11698 15008 11704 15020
rect 11379 14980 11704 15008
rect 11379 14977 11391 14980
rect 11333 14971 11391 14977
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 2792 14912 2912 14940
rect 2792 14872 2820 14912
rect 3694 14900 3700 14952
rect 3752 14940 3758 14952
rect 4249 14943 4307 14949
rect 4249 14940 4261 14943
rect 3752 14912 4261 14940
rect 3752 14900 3758 14912
rect 4249 14909 4261 14912
rect 4295 14909 4307 14943
rect 4249 14903 4307 14909
rect 5074 14900 5080 14952
rect 5132 14940 5138 14952
rect 5258 14940 5264 14952
rect 5132 14912 5264 14940
rect 5132 14900 5138 14912
rect 5258 14900 5264 14912
rect 5316 14900 5322 14952
rect 5442 14940 5448 14952
rect 5403 14912 5448 14940
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 5902 14940 5908 14952
rect 5863 14912 5908 14940
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 6270 14900 6276 14952
rect 6328 14900 6334 14952
rect 9674 14900 9680 14952
rect 9732 14940 9738 14952
rect 9861 14943 9919 14949
rect 9861 14940 9873 14943
rect 9732 14912 9873 14940
rect 9732 14900 9738 14912
rect 9861 14909 9873 14912
rect 9907 14909 9919 14943
rect 12342 14940 12348 14952
rect 12303 14912 12348 14940
rect 9861 14903 9919 14909
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 12728 14949 12756 15048
rect 13354 15036 13360 15088
rect 13412 15076 13418 15088
rect 13538 15076 13544 15088
rect 13412 15048 13544 15076
rect 13412 15036 13418 15048
rect 13538 15036 13544 15048
rect 13596 15036 13602 15088
rect 14642 15008 14648 15020
rect 13280 14980 14648 15008
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 12529 14943 12587 14949
rect 12529 14909 12541 14943
rect 12575 14909 12587 14943
rect 12529 14903 12587 14909
rect 12713 14943 12771 14949
rect 12713 14909 12725 14943
rect 12759 14909 12771 14943
rect 13280 14940 13308 14980
rect 14642 14968 14648 14980
rect 14700 15008 14706 15020
rect 15194 15008 15200 15020
rect 14700 14980 15200 15008
rect 14700 14968 14706 14980
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 17494 15008 17500 15020
rect 17328 14980 17500 15008
rect 13403 14943 13461 14949
rect 13403 14940 13415 14943
rect 13280 14912 13415 14940
rect 12713 14903 12771 14909
rect 13403 14909 13415 14912
rect 13449 14909 13461 14943
rect 13403 14903 13461 14909
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14909 13691 14943
rect 13814 14940 13820 14952
rect 13775 14912 13820 14940
rect 13633 14903 13691 14909
rect 2240 14844 2820 14872
rect 1937 14835 1995 14841
rect 2866 14832 2872 14884
rect 2924 14872 2930 14884
rect 5537 14875 5595 14881
rect 2924 14844 5304 14872
rect 2924 14832 2930 14844
rect 1762 14764 1768 14816
rect 1820 14804 1826 14816
rect 2685 14807 2743 14813
rect 2685 14804 2697 14807
rect 1820 14776 2697 14804
rect 1820 14764 1826 14776
rect 2685 14773 2697 14776
rect 2731 14773 2743 14807
rect 2685 14767 2743 14773
rect 3510 14764 3516 14816
rect 3568 14804 3574 14816
rect 4062 14804 4068 14816
rect 3568 14776 4068 14804
rect 3568 14764 3574 14776
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 4341 14807 4399 14813
rect 4341 14773 4353 14807
rect 4387 14804 4399 14807
rect 4430 14804 4436 14816
rect 4387 14776 4436 14804
rect 4387 14773 4399 14776
rect 4341 14767 4399 14773
rect 4430 14764 4436 14776
rect 4488 14804 4494 14816
rect 4798 14804 4804 14816
rect 4488 14776 4804 14804
rect 4488 14764 4494 14776
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 5166 14804 5172 14816
rect 5127 14776 5172 14804
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 5276 14804 5304 14844
rect 5537 14841 5549 14875
rect 5583 14872 5595 14875
rect 5810 14872 5816 14884
rect 5583 14844 5816 14872
rect 5583 14841 5595 14844
rect 5537 14835 5595 14841
rect 5810 14832 5816 14844
rect 5868 14872 5874 14884
rect 6288 14872 6316 14900
rect 5868 14844 6316 14872
rect 7469 14875 7527 14881
rect 5868 14832 5874 14844
rect 7469 14841 7481 14875
rect 7515 14872 7527 14875
rect 10594 14872 10600 14884
rect 7515 14844 10600 14872
rect 7515 14841 7527 14844
rect 7469 14835 7527 14841
rect 10594 14832 10600 14844
rect 10652 14832 10658 14884
rect 6273 14807 6331 14813
rect 6273 14804 6285 14807
rect 5276 14776 6285 14804
rect 6273 14773 6285 14776
rect 6319 14773 6331 14807
rect 6454 14804 6460 14816
rect 6415 14776 6460 14804
rect 6273 14767 6331 14773
rect 6454 14764 6460 14776
rect 6512 14764 6518 14816
rect 7374 14804 7380 14816
rect 7335 14776 7380 14804
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 9122 14764 9128 14816
rect 9180 14804 9186 14816
rect 9953 14807 10011 14813
rect 9953 14804 9965 14807
rect 9180 14776 9965 14804
rect 9180 14764 9186 14776
rect 9953 14773 9965 14776
rect 9999 14773 10011 14807
rect 9953 14767 10011 14773
rect 10134 14764 10140 14816
rect 10192 14804 10198 14816
rect 11057 14807 11115 14813
rect 11057 14804 11069 14807
rect 10192 14776 11069 14804
rect 10192 14764 10198 14776
rect 11057 14773 11069 14776
rect 11103 14773 11115 14807
rect 11057 14767 11115 14773
rect 12250 14764 12256 14816
rect 12308 14804 12314 14816
rect 12452 14804 12480 14903
rect 12544 14872 12572 14903
rect 12802 14872 12808 14884
rect 12544 14844 12808 14872
rect 12802 14832 12808 14844
rect 12860 14872 12866 14884
rect 13078 14872 13084 14884
rect 12860 14844 13084 14872
rect 12860 14832 12866 14844
rect 13078 14832 13084 14844
rect 13136 14832 13142 14884
rect 13556 14804 13584 14903
rect 13648 14872 13676 14903
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 17328 14949 17356 14980
rect 17494 14968 17500 14980
rect 17552 14968 17558 15020
rect 26050 15008 26056 15020
rect 26011 14980 26056 15008
rect 26050 14968 26056 14980
rect 26108 14968 26114 15020
rect 17313 14943 17371 14949
rect 17313 14909 17325 14943
rect 17359 14909 17371 14943
rect 17313 14903 17371 14909
rect 17405 14943 17463 14949
rect 17405 14909 17417 14943
rect 17451 14940 17463 14943
rect 17586 14940 17592 14952
rect 17451 14912 17592 14940
rect 17451 14909 17463 14912
rect 17405 14903 17463 14909
rect 17586 14900 17592 14912
rect 17644 14900 17650 14952
rect 21542 14900 21548 14952
rect 21600 14940 21606 14952
rect 21637 14943 21695 14949
rect 21637 14940 21649 14943
rect 21600 14912 21649 14940
rect 21600 14900 21606 14912
rect 21637 14909 21649 14912
rect 21683 14909 21695 14943
rect 21637 14903 21695 14909
rect 21726 14900 21732 14952
rect 21784 14949 21790 14952
rect 21784 14943 21833 14949
rect 21784 14909 21787 14943
rect 21821 14909 21833 14943
rect 21784 14903 21833 14909
rect 22097 14943 22155 14949
rect 22097 14909 22109 14943
rect 22143 14940 22155 14943
rect 22646 14940 22652 14952
rect 22143 14912 22652 14940
rect 22143 14909 22155 14912
rect 22097 14903 22155 14909
rect 21784 14900 21790 14903
rect 22646 14900 22652 14912
rect 22704 14900 22710 14952
rect 25961 14943 26019 14949
rect 25961 14909 25973 14943
rect 26007 14940 26019 14943
rect 26418 14940 26424 14952
rect 26007 14912 26424 14940
rect 26007 14909 26019 14912
rect 25961 14903 26019 14909
rect 26418 14900 26424 14912
rect 26476 14900 26482 14952
rect 26789 14943 26847 14949
rect 26789 14909 26801 14943
rect 26835 14909 26847 14943
rect 26789 14903 26847 14909
rect 27056 14943 27114 14949
rect 27056 14909 27068 14943
rect 27102 14940 27114 14943
rect 27430 14940 27436 14952
rect 27102 14912 27436 14940
rect 27102 14909 27114 14912
rect 27056 14903 27114 14909
rect 14274 14872 14280 14884
rect 13648 14844 14280 14872
rect 14274 14832 14280 14844
rect 14332 14832 14338 14884
rect 17126 14872 17132 14884
rect 17087 14844 17132 14872
rect 17126 14832 17132 14844
rect 17184 14832 17190 14884
rect 24854 14832 24860 14884
rect 24912 14872 24918 14884
rect 25866 14872 25872 14884
rect 24912 14844 25872 14872
rect 24912 14832 24918 14844
rect 25866 14832 25872 14844
rect 25924 14872 25930 14884
rect 26804 14872 26832 14903
rect 27430 14900 27436 14912
rect 27488 14900 27494 14952
rect 25924 14844 26832 14872
rect 25924 14832 25930 14844
rect 12308 14776 13584 14804
rect 17497 14807 17555 14813
rect 12308 14764 12314 14776
rect 17497 14773 17509 14807
rect 17543 14804 17555 14807
rect 17586 14804 17592 14816
rect 17543 14776 17592 14804
rect 17543 14773 17555 14776
rect 17497 14767 17555 14773
rect 17586 14764 17592 14776
rect 17644 14764 17650 14816
rect 22097 14807 22155 14813
rect 22097 14773 22109 14807
rect 22143 14804 22155 14807
rect 22462 14804 22468 14816
rect 22143 14776 22468 14804
rect 22143 14773 22155 14776
rect 22097 14767 22155 14773
rect 22462 14764 22468 14776
rect 22520 14764 22526 14816
rect 1104 14714 28888 14736
rect 1104 14662 10246 14714
rect 10298 14662 10310 14714
rect 10362 14662 10374 14714
rect 10426 14662 10438 14714
rect 10490 14662 19510 14714
rect 19562 14662 19574 14714
rect 19626 14662 19638 14714
rect 19690 14662 19702 14714
rect 19754 14662 28888 14714
rect 1104 14640 28888 14662
rect 1762 14600 1768 14612
rect 1723 14572 1768 14600
rect 1762 14560 1768 14572
rect 1820 14560 1826 14612
rect 2409 14603 2467 14609
rect 2409 14569 2421 14603
rect 2455 14600 2467 14603
rect 2498 14600 2504 14612
rect 2455 14572 2504 14600
rect 2455 14569 2467 14572
rect 2409 14563 2467 14569
rect 2498 14560 2504 14572
rect 2556 14560 2562 14612
rect 3878 14560 3884 14612
rect 3936 14600 3942 14612
rect 4430 14600 4436 14612
rect 3936 14572 4436 14600
rect 3936 14560 3942 14572
rect 4430 14560 4436 14572
rect 4488 14560 4494 14612
rect 4798 14560 4804 14612
rect 4856 14600 4862 14612
rect 5261 14603 5319 14609
rect 5261 14600 5273 14603
rect 4856 14572 5273 14600
rect 4856 14560 4862 14572
rect 5261 14569 5273 14572
rect 5307 14569 5319 14603
rect 10134 14600 10140 14612
rect 10095 14572 10140 14600
rect 5261 14563 5319 14569
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 10962 14600 10968 14612
rect 10923 14572 10968 14600
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 13541 14603 13599 14609
rect 13541 14569 13553 14603
rect 13587 14600 13599 14603
rect 13814 14600 13820 14612
rect 13587 14572 13820 14600
rect 13587 14569 13599 14572
rect 13541 14563 13599 14569
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 14182 14560 14188 14612
rect 14240 14600 14246 14612
rect 14642 14600 14648 14612
rect 14240 14572 14648 14600
rect 14240 14560 14246 14572
rect 14642 14560 14648 14572
rect 14700 14560 14706 14612
rect 17586 14560 17592 14612
rect 17644 14600 17650 14612
rect 17681 14603 17739 14609
rect 17681 14600 17693 14603
rect 17644 14572 17693 14600
rect 17644 14560 17650 14572
rect 17681 14569 17693 14572
rect 17727 14569 17739 14603
rect 17862 14600 17868 14612
rect 17823 14572 17868 14600
rect 17681 14563 17739 14569
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 19058 14560 19064 14612
rect 19116 14560 19122 14612
rect 21082 14600 21088 14612
rect 21043 14572 21088 14600
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 21361 14603 21419 14609
rect 21361 14569 21373 14603
rect 21407 14600 21419 14603
rect 21910 14600 21916 14612
rect 21407 14572 21916 14600
rect 21407 14569 21419 14572
rect 21361 14563 21419 14569
rect 21910 14560 21916 14572
rect 21968 14560 21974 14612
rect 22646 14600 22652 14612
rect 22607 14572 22652 14600
rect 22646 14560 22652 14572
rect 22704 14560 22710 14612
rect 26050 14560 26056 14612
rect 26108 14600 26114 14612
rect 26881 14603 26939 14609
rect 26881 14600 26893 14603
rect 26108 14572 26893 14600
rect 26108 14560 26114 14572
rect 26881 14569 26893 14572
rect 26927 14569 26939 14603
rect 26881 14563 26939 14569
rect 3786 14532 3792 14544
rect 3528 14504 3792 14532
rect 1946 14464 1952 14476
rect 1907 14436 1952 14464
rect 1946 14424 1952 14436
rect 2004 14424 2010 14476
rect 2593 14467 2651 14473
rect 2593 14433 2605 14467
rect 2639 14464 2651 14467
rect 2774 14464 2780 14476
rect 2639 14436 2780 14464
rect 2639 14433 2651 14436
rect 2593 14427 2651 14433
rect 2774 14424 2780 14436
rect 2832 14424 2838 14476
rect 3528 14473 3556 14504
rect 3786 14492 3792 14504
rect 3844 14532 3850 14544
rect 9674 14532 9680 14544
rect 3844 14504 5672 14532
rect 3844 14492 3850 14504
rect 3513 14467 3571 14473
rect 3513 14433 3525 14467
rect 3559 14433 3571 14467
rect 3694 14464 3700 14476
rect 3655 14436 3700 14464
rect 3513 14427 3571 14433
rect 3694 14424 3700 14436
rect 3752 14424 3758 14476
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 4249 14467 4307 14473
rect 4249 14464 4261 14467
rect 4028 14436 4261 14464
rect 4028 14424 4034 14436
rect 4249 14433 4261 14436
rect 4295 14433 4307 14467
rect 4249 14427 4307 14433
rect 4264 14396 4292 14427
rect 4430 14424 4436 14476
rect 4488 14464 4494 14476
rect 5077 14467 5135 14473
rect 5077 14464 5089 14467
rect 4488 14436 5089 14464
rect 4488 14424 4494 14436
rect 5077 14433 5089 14436
rect 5123 14433 5135 14467
rect 5077 14427 5135 14433
rect 5353 14467 5411 14473
rect 5353 14433 5365 14467
rect 5399 14433 5411 14467
rect 5353 14427 5411 14433
rect 5368 14396 5396 14427
rect 4264 14368 5396 14396
rect 4249 14331 4307 14337
rect 4249 14297 4261 14331
rect 4295 14328 4307 14331
rect 4798 14328 4804 14340
rect 4295 14300 4804 14328
rect 4295 14297 4307 14300
rect 4249 14291 4307 14297
rect 4798 14288 4804 14300
rect 4856 14288 4862 14340
rect 5644 14328 5672 14504
rect 9048 14504 9680 14532
rect 6454 14424 6460 14476
rect 6512 14464 6518 14476
rect 7098 14464 7104 14476
rect 6512 14436 7104 14464
rect 6512 14424 6518 14436
rect 7098 14424 7104 14436
rect 7156 14464 7162 14476
rect 9048 14473 9076 14504
rect 9674 14492 9680 14504
rect 9732 14492 9738 14544
rect 12434 14492 12440 14544
rect 12492 14532 12498 14544
rect 12621 14535 12679 14541
rect 12492 14504 12537 14532
rect 12492 14492 12498 14504
rect 12621 14501 12633 14535
rect 12667 14532 12679 14535
rect 13078 14532 13084 14544
rect 12667 14504 13084 14532
rect 12667 14501 12679 14504
rect 12621 14495 12679 14501
rect 13078 14492 13084 14504
rect 13136 14492 13142 14544
rect 7469 14467 7527 14473
rect 7469 14464 7481 14467
rect 7156 14436 7481 14464
rect 7156 14424 7162 14436
rect 7469 14433 7481 14436
rect 7515 14433 7527 14467
rect 7469 14427 7527 14433
rect 9033 14467 9091 14473
rect 9033 14433 9045 14467
rect 9079 14433 9091 14467
rect 9033 14427 9091 14433
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14464 9183 14467
rect 10045 14467 10103 14473
rect 10045 14464 10057 14467
rect 9171 14436 10057 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 10045 14433 10057 14436
rect 10091 14433 10103 14467
rect 10045 14427 10103 14433
rect 10873 14467 10931 14473
rect 10873 14433 10885 14467
rect 10919 14464 10931 14467
rect 10962 14464 10968 14476
rect 10919 14436 10968 14464
rect 10919 14433 10931 14436
rect 10873 14427 10931 14433
rect 10962 14424 10968 14436
rect 11020 14424 11026 14476
rect 12342 14424 12348 14476
rect 12400 14464 12406 14476
rect 12713 14467 12771 14473
rect 12713 14464 12725 14467
rect 12400 14436 12725 14464
rect 12400 14424 12406 14436
rect 12713 14433 12725 14436
rect 12759 14433 12771 14467
rect 13354 14464 13360 14476
rect 13315 14436 13360 14464
rect 12713 14427 12771 14433
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14464 13599 14467
rect 14182 14464 14188 14476
rect 13587 14436 14188 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 17494 14464 17500 14476
rect 17455 14436 17500 14464
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 17589 14467 17647 14473
rect 17589 14433 17601 14467
rect 17635 14433 17647 14467
rect 17589 14427 17647 14433
rect 9674 14356 9680 14408
rect 9732 14396 9738 14408
rect 9950 14396 9956 14408
rect 9732 14368 9956 14396
rect 9732 14356 9738 14368
rect 9950 14356 9956 14368
rect 10008 14396 10014 14408
rect 10229 14399 10287 14405
rect 10229 14396 10241 14399
rect 10008 14368 10241 14396
rect 10008 14356 10014 14368
rect 10229 14365 10241 14368
rect 10275 14365 10287 14399
rect 17604 14396 17632 14427
rect 17862 14396 17868 14408
rect 17604 14368 17868 14396
rect 10229 14359 10287 14365
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 12161 14331 12219 14337
rect 12161 14328 12173 14331
rect 5644 14300 12173 14328
rect 12161 14297 12173 14300
rect 12207 14297 12219 14331
rect 12161 14291 12219 14297
rect 17313 14331 17371 14337
rect 17313 14297 17325 14331
rect 17359 14328 17371 14331
rect 17678 14328 17684 14340
rect 17359 14300 17684 14328
rect 17359 14297 17371 14300
rect 17313 14291 17371 14297
rect 17678 14288 17684 14300
rect 17736 14288 17742 14340
rect 4893 14263 4951 14269
rect 4893 14229 4905 14263
rect 4939 14260 4951 14263
rect 4982 14260 4988 14272
rect 4939 14232 4988 14260
rect 4939 14229 4951 14232
rect 4893 14223 4951 14229
rect 4982 14220 4988 14232
rect 5040 14220 5046 14272
rect 7561 14263 7619 14269
rect 7561 14229 7573 14263
rect 7607 14260 7619 14263
rect 9122 14260 9128 14272
rect 7607 14232 9128 14260
rect 7607 14229 7619 14232
rect 7561 14223 7619 14229
rect 9122 14220 9128 14232
rect 9180 14220 9186 14272
rect 9677 14263 9735 14269
rect 9677 14229 9689 14263
rect 9723 14260 9735 14263
rect 9858 14260 9864 14272
rect 9723 14232 9864 14260
rect 9723 14229 9735 14232
rect 9677 14223 9735 14229
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 10594 14220 10600 14272
rect 10652 14260 10658 14272
rect 19076 14260 19104 14560
rect 25682 14492 25688 14544
rect 25740 14532 25746 14544
rect 25777 14535 25835 14541
rect 25777 14532 25789 14535
rect 25740 14504 25789 14532
rect 25740 14492 25746 14504
rect 25777 14501 25789 14504
rect 25823 14501 25835 14535
rect 25958 14532 25964 14544
rect 25919 14504 25964 14532
rect 25777 14495 25835 14501
rect 25958 14492 25964 14504
rect 26016 14492 26022 14544
rect 27982 14532 27988 14544
rect 27943 14504 27988 14532
rect 27982 14492 27988 14504
rect 28040 14492 28046 14544
rect 20714 14424 20720 14476
rect 20772 14464 20778 14476
rect 20993 14467 21051 14473
rect 20993 14464 21005 14467
rect 20772 14436 21005 14464
rect 20772 14424 20778 14436
rect 20993 14433 21005 14436
rect 21039 14433 21051 14467
rect 21174 14464 21180 14476
rect 21135 14436 21180 14464
rect 20993 14427 21051 14433
rect 21174 14424 21180 14436
rect 21232 14424 21238 14476
rect 22557 14467 22615 14473
rect 22557 14433 22569 14467
rect 22603 14464 22615 14467
rect 22646 14464 22652 14476
rect 22603 14436 22652 14464
rect 22603 14433 22615 14436
rect 22557 14427 22615 14433
rect 22646 14424 22652 14436
rect 22704 14424 22710 14476
rect 22741 14467 22799 14473
rect 22741 14433 22753 14467
rect 22787 14464 22799 14467
rect 23014 14464 23020 14476
rect 22787 14436 23020 14464
rect 22787 14433 22799 14436
rect 22741 14427 22799 14433
rect 23014 14424 23020 14436
rect 23072 14424 23078 14476
rect 20898 14356 20904 14408
rect 20956 14396 20962 14408
rect 21910 14396 21916 14408
rect 20956 14368 21916 14396
rect 20956 14356 20962 14368
rect 21910 14356 21916 14368
rect 21968 14356 21974 14408
rect 26418 14396 26424 14408
rect 26379 14368 26424 14396
rect 26418 14356 26424 14368
rect 26476 14356 26482 14408
rect 20806 14328 20812 14340
rect 20767 14300 20812 14328
rect 20806 14288 20812 14300
rect 20864 14288 20870 14340
rect 26694 14288 26700 14340
rect 26752 14328 26758 14340
rect 26789 14331 26847 14337
rect 26789 14328 26801 14331
rect 26752 14300 26801 14328
rect 26752 14288 26758 14300
rect 26789 14297 26801 14300
rect 26835 14328 26847 14331
rect 27246 14328 27252 14340
rect 26835 14300 27252 14328
rect 26835 14297 26847 14300
rect 26789 14291 26847 14297
rect 27246 14288 27252 14300
rect 27304 14288 27310 14340
rect 28166 14328 28172 14340
rect 28127 14300 28172 14328
rect 28166 14288 28172 14300
rect 28224 14288 28230 14340
rect 27982 14260 27988 14272
rect 10652 14232 27988 14260
rect 10652 14220 10658 14232
rect 27982 14220 27988 14232
rect 28040 14220 28046 14272
rect 1104 14170 28888 14192
rect 1104 14118 5614 14170
rect 5666 14118 5678 14170
rect 5730 14118 5742 14170
rect 5794 14118 5806 14170
rect 5858 14118 14878 14170
rect 14930 14118 14942 14170
rect 14994 14118 15006 14170
rect 15058 14118 15070 14170
rect 15122 14118 24142 14170
rect 24194 14118 24206 14170
rect 24258 14118 24270 14170
rect 24322 14118 24334 14170
rect 24386 14118 28888 14170
rect 1104 14096 28888 14118
rect 2314 14056 2320 14068
rect 2275 14028 2320 14056
rect 2314 14016 2320 14028
rect 2372 14016 2378 14068
rect 2866 14056 2872 14068
rect 2827 14028 2872 14056
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 4706 14056 4712 14068
rect 4667 14028 4712 14056
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 10962 14056 10968 14068
rect 10923 14028 10968 14056
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 17126 14056 17132 14068
rect 17087 14028 17132 14056
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 20533 14059 20591 14065
rect 20533 14025 20545 14059
rect 20579 14056 20591 14059
rect 20990 14056 20996 14068
rect 20579 14028 20996 14056
rect 20579 14025 20591 14028
rect 20533 14019 20591 14025
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 22646 14016 22652 14068
rect 22704 14056 22710 14068
rect 23290 14056 23296 14068
rect 22704 14028 23296 14056
rect 22704 14016 22710 14028
rect 23290 14016 23296 14028
rect 23348 14056 23354 14068
rect 23753 14059 23811 14065
rect 23753 14056 23765 14059
rect 23348 14028 23765 14056
rect 23348 14016 23354 14028
rect 23753 14025 23765 14028
rect 23799 14025 23811 14059
rect 23753 14019 23811 14025
rect 27341 14059 27399 14065
rect 27341 14025 27353 14059
rect 27387 14056 27399 14059
rect 27430 14056 27436 14068
rect 27387 14028 27436 14056
rect 27387 14025 27399 14028
rect 27341 14019 27399 14025
rect 27430 14016 27436 14028
rect 27488 14016 27494 14068
rect 2225 13991 2283 13997
rect 2225 13957 2237 13991
rect 2271 13988 2283 13991
rect 3326 13988 3332 14000
rect 2271 13960 3332 13988
rect 2271 13957 2283 13960
rect 2225 13951 2283 13957
rect 3326 13948 3332 13960
rect 3384 13948 3390 14000
rect 4614 13988 4620 14000
rect 4575 13960 4620 13988
rect 4614 13948 4620 13960
rect 4672 13948 4678 14000
rect 7190 13948 7196 14000
rect 7248 13988 7254 14000
rect 7929 13991 7987 13997
rect 7929 13988 7941 13991
rect 7248 13960 7941 13988
rect 7248 13948 7254 13960
rect 7929 13957 7941 13960
rect 7975 13957 7987 13991
rect 12066 13988 12072 14000
rect 7929 13951 7987 13957
rect 11440 13960 12072 13988
rect 2590 13920 2596 13932
rect 1872 13892 2596 13920
rect 1872 13861 1900 13892
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 4982 13920 4988 13932
rect 4264 13892 4988 13920
rect 1857 13855 1915 13861
rect 1857 13821 1869 13855
rect 1903 13821 1915 13855
rect 1857 13815 1915 13821
rect 2409 13855 2467 13861
rect 2409 13821 2421 13855
rect 2455 13852 2467 13855
rect 2498 13852 2504 13864
rect 2455 13824 2504 13852
rect 2455 13821 2467 13824
rect 2409 13815 2467 13821
rect 2498 13812 2504 13824
rect 2556 13812 2562 13864
rect 3050 13852 3056 13864
rect 3011 13824 3056 13852
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 4264 13861 4292 13892
rect 4982 13880 4988 13892
rect 5040 13880 5046 13932
rect 8202 13920 8208 13932
rect 8036 13892 8208 13920
rect 4249 13855 4307 13861
rect 4249 13821 4261 13855
rect 4295 13821 4307 13855
rect 4249 13815 4307 13821
rect 4801 13855 4859 13861
rect 4801 13821 4813 13855
rect 4847 13852 4859 13855
rect 4890 13852 4896 13864
rect 4847 13824 4896 13852
rect 4847 13821 4859 13824
rect 4801 13815 4859 13821
rect 4890 13812 4896 13824
rect 4948 13812 4954 13864
rect 7098 13852 7104 13864
rect 7059 13824 7104 13852
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 8036 13861 8064 13892
rect 8202 13880 8208 13892
rect 8260 13920 8266 13932
rect 11440 13929 11468 13960
rect 12066 13948 12072 13960
rect 12124 13948 12130 14000
rect 16574 13948 16580 14000
rect 16632 13988 16638 14000
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 16632 13960 17049 13988
rect 16632 13948 16638 13960
rect 17037 13957 17049 13960
rect 17083 13988 17095 13991
rect 17862 13988 17868 14000
rect 17083 13960 17868 13988
rect 17083 13957 17095 13960
rect 17037 13951 17095 13957
rect 17862 13948 17868 13960
rect 17920 13948 17926 14000
rect 23842 13948 23848 14000
rect 23900 13988 23906 14000
rect 23900 13960 27292 13988
rect 23900 13948 23906 13960
rect 10505 13923 10563 13929
rect 10505 13920 10517 13923
rect 8260 13892 10517 13920
rect 8260 13880 8266 13892
rect 10505 13889 10517 13892
rect 10551 13889 10563 13923
rect 10505 13883 10563 13889
rect 11425 13923 11483 13929
rect 11425 13889 11437 13923
rect 11471 13889 11483 13923
rect 11425 13883 11483 13889
rect 11609 13923 11667 13929
rect 11609 13889 11621 13923
rect 11655 13920 11667 13923
rect 11698 13920 11704 13932
rect 11655 13892 11704 13920
rect 11655 13889 11667 13892
rect 11609 13883 11667 13889
rect 11698 13880 11704 13892
rect 11756 13880 11762 13932
rect 18874 13920 18880 13932
rect 18835 13892 18880 13920
rect 18874 13880 18880 13892
rect 18932 13880 18938 13932
rect 20530 13880 20536 13932
rect 20588 13920 20594 13932
rect 20717 13923 20775 13929
rect 20717 13920 20729 13923
rect 20588 13892 20729 13920
rect 20588 13880 20594 13892
rect 20717 13889 20729 13892
rect 20763 13889 20775 13923
rect 21082 13920 21088 13932
rect 21043 13892 21088 13920
rect 20717 13883 20775 13889
rect 21082 13880 21088 13892
rect 21140 13880 21146 13932
rect 25792 13892 27200 13920
rect 8021 13855 8079 13861
rect 8021 13821 8033 13855
rect 8067 13821 8079 13855
rect 9766 13852 9772 13864
rect 9727 13824 9772 13852
rect 8021 13815 8079 13821
rect 9766 13812 9772 13824
rect 9824 13812 9830 13864
rect 9858 13812 9864 13864
rect 9916 13852 9922 13864
rect 9916 13824 9961 13852
rect 9916 13812 9922 13824
rect 11882 13812 11888 13864
rect 11940 13852 11946 13864
rect 12161 13855 12219 13861
rect 12161 13852 12173 13855
rect 11940 13824 12173 13852
rect 11940 13812 11946 13824
rect 12161 13821 12173 13824
rect 12207 13821 12219 13855
rect 12161 13815 12219 13821
rect 12345 13855 12403 13861
rect 12345 13821 12357 13855
rect 12391 13852 12403 13855
rect 14182 13852 14188 13864
rect 12391 13824 14188 13852
rect 12391 13821 12403 13824
rect 12345 13815 12403 13821
rect 14182 13812 14188 13824
rect 14240 13812 14246 13864
rect 16669 13855 16727 13861
rect 16669 13821 16681 13855
rect 16715 13852 16727 13855
rect 17034 13852 17040 13864
rect 16715 13824 17040 13852
rect 16715 13821 16727 13824
rect 16669 13815 16727 13821
rect 17034 13812 17040 13824
rect 17092 13852 17098 13864
rect 17589 13855 17647 13861
rect 17589 13852 17601 13855
rect 17092 13824 17601 13852
rect 17092 13812 17098 13824
rect 17589 13821 17601 13824
rect 17635 13821 17647 13855
rect 17589 13815 17647 13821
rect 17678 13812 17684 13864
rect 17736 13852 17742 13864
rect 18785 13855 18843 13861
rect 17736 13824 17781 13852
rect 17736 13812 17742 13824
rect 18785 13821 18797 13855
rect 18831 13852 18843 13855
rect 19978 13852 19984 13864
rect 18831 13824 19984 13852
rect 18831 13821 18843 13824
rect 18785 13815 18843 13821
rect 19978 13812 19984 13824
rect 20036 13812 20042 13864
rect 20806 13812 20812 13864
rect 20864 13852 20870 13864
rect 20864 13824 20909 13852
rect 20864 13812 20870 13824
rect 20990 13812 20996 13864
rect 21048 13852 21054 13864
rect 21174 13852 21180 13864
rect 21048 13824 21180 13852
rect 21048 13812 21054 13824
rect 21174 13812 21180 13824
rect 21232 13812 21238 13864
rect 22373 13855 22431 13861
rect 22373 13821 22385 13855
rect 22419 13821 22431 13855
rect 22373 13815 22431 13821
rect 1486 13744 1492 13796
rect 1544 13784 1550 13796
rect 1949 13787 2007 13793
rect 1949 13784 1961 13787
rect 1544 13756 1961 13784
rect 1544 13744 1550 13756
rect 1949 13753 1961 13756
rect 1995 13753 2007 13787
rect 4338 13784 4344 13796
rect 4299 13756 4344 13784
rect 1949 13747 2007 13753
rect 4338 13744 4344 13756
rect 4396 13744 4402 13796
rect 9214 13744 9220 13796
rect 9272 13784 9278 13796
rect 9490 13784 9496 13796
rect 9272 13756 9496 13784
rect 9272 13744 9278 13756
rect 9490 13744 9496 13756
rect 9548 13784 9554 13796
rect 9999 13787 10057 13793
rect 9999 13784 10011 13787
rect 9548 13756 10011 13784
rect 9548 13744 9554 13756
rect 9999 13753 10011 13756
rect 10045 13753 10057 13787
rect 9999 13747 10057 13753
rect 15930 13744 15936 13796
rect 15988 13784 15994 13796
rect 21542 13784 21548 13796
rect 15988 13756 21548 13784
rect 15988 13744 15994 13756
rect 21542 13744 21548 13756
rect 21600 13744 21606 13796
rect 22388 13784 22416 13815
rect 22462 13812 22468 13864
rect 22520 13852 22526 13864
rect 22629 13855 22687 13861
rect 22629 13852 22641 13855
rect 22520 13824 22641 13852
rect 22520 13812 22526 13824
rect 22629 13821 22641 13824
rect 22675 13821 22687 13855
rect 24854 13852 24860 13864
rect 22629 13815 22687 13821
rect 22756 13824 24860 13852
rect 22756 13784 22784 13824
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 25792 13861 25820 13892
rect 25777 13855 25835 13861
rect 25777 13821 25789 13855
rect 25823 13821 25835 13855
rect 25958 13852 25964 13864
rect 25919 13824 25964 13852
rect 25777 13815 25835 13821
rect 25958 13812 25964 13824
rect 26016 13812 26022 13864
rect 26697 13855 26755 13861
rect 26697 13821 26709 13855
rect 26743 13852 26755 13855
rect 26786 13852 26792 13864
rect 26743 13824 26792 13852
rect 26743 13821 26755 13824
rect 26697 13815 26755 13821
rect 26786 13812 26792 13824
rect 26844 13812 26850 13864
rect 22388 13756 22784 13784
rect 25222 13744 25228 13796
rect 25280 13784 25286 13796
rect 26513 13787 26571 13793
rect 26513 13784 26525 13787
rect 25280 13756 26525 13784
rect 25280 13744 25286 13756
rect 26513 13753 26525 13756
rect 26559 13753 26571 13787
rect 27172 13784 27200 13892
rect 27264 13861 27292 13960
rect 27249 13855 27307 13861
rect 27249 13821 27261 13855
rect 27295 13821 27307 13855
rect 27982 13852 27988 13864
rect 27943 13824 27988 13852
rect 27249 13815 27307 13821
rect 27982 13812 27988 13824
rect 28040 13812 28046 13864
rect 28166 13852 28172 13864
rect 28127 13824 28172 13852
rect 28166 13812 28172 13824
rect 28224 13812 28230 13864
rect 27890 13784 27896 13796
rect 27172 13756 27896 13784
rect 26513 13747 26571 13753
rect 27890 13744 27896 13756
rect 27948 13744 27954 13796
rect 3510 13676 3516 13728
rect 3568 13716 3574 13728
rect 11333 13719 11391 13725
rect 11333 13716 11345 13719
rect 3568 13688 11345 13716
rect 3568 13676 3574 13688
rect 11333 13685 11345 13688
rect 11379 13685 11391 13719
rect 12250 13716 12256 13728
rect 12211 13688 12256 13716
rect 11333 13679 11391 13685
rect 12250 13676 12256 13688
rect 12308 13676 12314 13728
rect 18322 13716 18328 13728
rect 18283 13688 18328 13716
rect 18322 13676 18328 13688
rect 18380 13676 18386 13728
rect 18690 13716 18696 13728
rect 18651 13688 18696 13716
rect 18690 13676 18696 13688
rect 18748 13676 18754 13728
rect 20714 13676 20720 13728
rect 20772 13716 20778 13728
rect 20901 13719 20959 13725
rect 20901 13716 20913 13719
rect 20772 13688 20913 13716
rect 20772 13676 20778 13688
rect 20901 13685 20913 13688
rect 20947 13685 20959 13719
rect 20901 13679 20959 13685
rect 1104 13626 28888 13648
rect 1104 13574 10246 13626
rect 10298 13574 10310 13626
rect 10362 13574 10374 13626
rect 10426 13574 10438 13626
rect 10490 13574 19510 13626
rect 19562 13574 19574 13626
rect 19626 13574 19638 13626
rect 19690 13574 19702 13626
rect 19754 13574 28888 13626
rect 1104 13552 28888 13574
rect 2314 13472 2320 13524
rect 2372 13512 2378 13524
rect 2685 13515 2743 13521
rect 2685 13512 2697 13515
rect 2372 13484 2697 13512
rect 2372 13472 2378 13484
rect 2685 13481 2697 13484
rect 2731 13481 2743 13515
rect 2685 13475 2743 13481
rect 3237 13515 3295 13521
rect 3237 13481 3249 13515
rect 3283 13512 3295 13515
rect 3510 13512 3516 13524
rect 3283 13484 3516 13512
rect 3283 13481 3295 13484
rect 3237 13475 3295 13481
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 3878 13472 3884 13524
rect 3936 13512 3942 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 3936 13484 4077 13512
rect 3936 13472 3942 13484
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4065 13475 4123 13481
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 5077 13515 5135 13521
rect 5077 13512 5089 13515
rect 4212 13484 5089 13512
rect 4212 13472 4218 13484
rect 5077 13481 5089 13484
rect 5123 13481 5135 13515
rect 5077 13475 5135 13481
rect 9125 13515 9183 13521
rect 9125 13481 9137 13515
rect 9171 13512 9183 13515
rect 9766 13512 9772 13524
rect 9171 13484 9772 13512
rect 9171 13481 9183 13484
rect 9125 13475 9183 13481
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 10505 13515 10563 13521
rect 10505 13512 10517 13515
rect 10192 13484 10517 13512
rect 10192 13472 10198 13484
rect 10505 13481 10517 13484
rect 10551 13481 10563 13515
rect 10505 13475 10563 13481
rect 12158 13472 12164 13524
rect 12216 13512 12222 13524
rect 12986 13512 12992 13524
rect 12216 13484 12992 13512
rect 12216 13472 12222 13484
rect 12986 13472 12992 13484
rect 13044 13472 13050 13524
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 13541 13515 13599 13521
rect 13541 13512 13553 13515
rect 13504 13484 13553 13512
rect 13504 13472 13510 13484
rect 13541 13481 13553 13484
rect 13587 13481 13599 13515
rect 13541 13475 13599 13481
rect 14090 13472 14096 13524
rect 14148 13512 14154 13524
rect 15473 13515 15531 13521
rect 15473 13512 15485 13515
rect 14148 13484 15485 13512
rect 14148 13472 14154 13484
rect 15473 13481 15485 13484
rect 15519 13481 15531 13515
rect 15473 13475 15531 13481
rect 16301 13515 16359 13521
rect 16301 13481 16313 13515
rect 16347 13512 16359 13515
rect 17678 13512 17684 13524
rect 16347 13484 17684 13512
rect 16347 13481 16359 13484
rect 16301 13475 16359 13481
rect 17678 13472 17684 13484
rect 17736 13472 17742 13524
rect 18141 13515 18199 13521
rect 18141 13481 18153 13515
rect 18187 13512 18199 13515
rect 18690 13512 18696 13524
rect 18187 13484 18696 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 18690 13472 18696 13484
rect 18748 13472 18754 13524
rect 19978 13512 19984 13524
rect 19939 13484 19984 13512
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 20714 13472 20720 13524
rect 20772 13512 20778 13524
rect 20809 13515 20867 13521
rect 20809 13512 20821 13515
rect 20772 13484 20821 13512
rect 20772 13472 20778 13484
rect 20809 13481 20821 13484
rect 20855 13481 20867 13515
rect 20809 13475 20867 13481
rect 20993 13515 21051 13521
rect 20993 13481 21005 13515
rect 21039 13512 21051 13515
rect 21726 13512 21732 13524
rect 21039 13484 21732 13512
rect 21039 13481 21051 13484
rect 20993 13475 21051 13481
rect 21726 13472 21732 13484
rect 21784 13472 21790 13524
rect 25406 13512 25412 13524
rect 21836 13484 25412 13512
rect 9030 13444 9036 13456
rect 8956 13416 9036 13444
rect 1854 13376 1860 13388
rect 1815 13348 1860 13376
rect 1854 13336 1860 13348
rect 1912 13336 1918 13388
rect 2590 13376 2596 13388
rect 2551 13348 2596 13376
rect 2590 13336 2596 13348
rect 2648 13336 2654 13388
rect 3418 13376 3424 13388
rect 3379 13348 3424 13376
rect 3418 13336 3424 13348
rect 3476 13336 3482 13388
rect 3786 13336 3792 13388
rect 3844 13376 3850 13388
rect 3973 13379 4031 13385
rect 3973 13376 3985 13379
rect 3844 13348 3985 13376
rect 3844 13336 3850 13348
rect 3973 13345 3985 13348
rect 4019 13345 4031 13379
rect 7650 13376 7656 13388
rect 7611 13348 7656 13376
rect 3973 13339 4031 13345
rect 7650 13336 7656 13348
rect 7708 13336 7714 13388
rect 7834 13336 7840 13388
rect 7892 13376 7898 13388
rect 8202 13376 8208 13388
rect 7892 13348 8208 13376
rect 7892 13336 7898 13348
rect 8202 13336 8208 13348
rect 8260 13376 8266 13388
rect 8956 13385 8984 13416
rect 9030 13404 9036 13416
rect 9088 13404 9094 13456
rect 11974 13404 11980 13456
rect 12032 13444 12038 13456
rect 12342 13444 12348 13456
rect 12032 13416 12348 13444
rect 12032 13404 12038 13416
rect 12342 13404 12348 13416
rect 12400 13404 12406 13456
rect 17586 13444 17592 13456
rect 16132 13416 17592 13444
rect 8297 13379 8355 13385
rect 8297 13376 8309 13379
rect 8260 13348 8309 13376
rect 8260 13336 8266 13348
rect 8297 13345 8309 13348
rect 8343 13345 8355 13379
rect 8297 13339 8355 13345
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13345 8999 13379
rect 9122 13376 9128 13388
rect 9083 13348 9128 13376
rect 8941 13339 8999 13345
rect 9122 13336 9128 13348
rect 9180 13336 9186 13388
rect 10413 13379 10471 13385
rect 10413 13345 10425 13379
rect 10459 13376 10471 13379
rect 10594 13376 10600 13388
rect 10459 13348 10600 13376
rect 10459 13345 10471 13348
rect 10413 13339 10471 13345
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 11238 13336 11244 13388
rect 11296 13376 11302 13388
rect 12428 13379 12486 13385
rect 12428 13376 12440 13379
rect 11296 13348 12440 13376
rect 11296 13336 11302 13348
rect 12428 13345 12440 13348
rect 12474 13345 12486 13379
rect 12428 13339 12486 13345
rect 13814 13336 13820 13388
rect 13872 13376 13878 13388
rect 16132 13385 16160 13416
rect 17586 13404 17592 13416
rect 17644 13404 17650 13456
rect 18322 13404 18328 13456
rect 18380 13444 18386 13456
rect 18846 13447 18904 13453
rect 18846 13444 18858 13447
rect 18380 13416 18858 13444
rect 18380 13404 18386 13416
rect 18846 13413 18858 13416
rect 18892 13413 18904 13447
rect 18846 13407 18904 13413
rect 19242 13404 19248 13456
rect 19300 13444 19306 13456
rect 21836 13444 21864 13484
rect 25406 13472 25412 13484
rect 25464 13512 25470 13524
rect 25682 13512 25688 13524
rect 25464 13484 25688 13512
rect 25464 13472 25470 13484
rect 25682 13472 25688 13484
rect 25740 13472 25746 13524
rect 27985 13447 28043 13453
rect 27985 13444 27997 13447
rect 19300 13416 21864 13444
rect 22066 13416 27997 13444
rect 19300 13404 19306 13416
rect 14349 13379 14407 13385
rect 14349 13376 14361 13379
rect 13872 13348 14361 13376
rect 13872 13336 13878 13348
rect 14349 13345 14361 13348
rect 14395 13345 14407 13379
rect 14349 13339 14407 13345
rect 16117 13379 16175 13385
rect 16117 13345 16129 13379
rect 16163 13345 16175 13379
rect 16117 13339 16175 13345
rect 16393 13379 16451 13385
rect 16393 13345 16405 13379
rect 16439 13376 16451 13379
rect 16574 13376 16580 13388
rect 16439 13348 16580 13376
rect 16439 13345 16451 13348
rect 16393 13339 16451 13345
rect 16574 13336 16580 13348
rect 16632 13336 16638 13388
rect 17494 13336 17500 13388
rect 17552 13376 17558 13388
rect 17773 13379 17831 13385
rect 17773 13376 17785 13379
rect 17552 13348 17785 13376
rect 17552 13336 17558 13348
rect 17773 13345 17785 13348
rect 17819 13345 17831 13379
rect 17773 13339 17831 13345
rect 18601 13379 18659 13385
rect 18601 13345 18613 13379
rect 18647 13376 18659 13379
rect 20162 13376 20168 13388
rect 18647 13348 20168 13376
rect 18647 13345 18659 13348
rect 18601 13339 18659 13345
rect 20162 13336 20168 13348
rect 20220 13336 20226 13388
rect 20717 13379 20775 13385
rect 20717 13345 20729 13379
rect 20763 13345 20775 13379
rect 21082 13376 21088 13388
rect 21043 13348 21088 13376
rect 20717 13339 20775 13345
rect 5166 13308 5172 13320
rect 5127 13280 5172 13308
rect 5166 13268 5172 13280
rect 5224 13268 5230 13320
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13308 5411 13311
rect 6454 13308 6460 13320
rect 5399 13280 6460 13308
rect 5399 13277 5411 13280
rect 5353 13271 5411 13277
rect 6454 13268 6460 13280
rect 6512 13308 6518 13320
rect 6638 13308 6644 13320
rect 6512 13280 6644 13308
rect 6512 13268 6518 13280
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 7745 13311 7803 13317
rect 7745 13277 7757 13311
rect 7791 13308 7803 13311
rect 7926 13308 7932 13320
rect 7791 13280 7932 13308
rect 7791 13277 7803 13280
rect 7745 13271 7803 13277
rect 7926 13268 7932 13280
rect 7984 13268 7990 13320
rect 8478 13308 8484 13320
rect 8391 13280 8484 13308
rect 8478 13268 8484 13280
rect 8536 13308 8542 13320
rect 9140 13308 9168 13336
rect 8536 13280 9168 13308
rect 12161 13311 12219 13317
rect 8536 13268 8542 13280
rect 12161 13277 12173 13311
rect 12207 13277 12219 13311
rect 12161 13271 12219 13277
rect 14093 13311 14151 13317
rect 14093 13277 14105 13311
rect 14139 13277 14151 13311
rect 17678 13308 17684 13320
rect 17639 13280 17684 13308
rect 14093 13271 14151 13277
rect 2041 13243 2099 13249
rect 2041 13209 2053 13243
rect 2087 13240 2099 13243
rect 2314 13240 2320 13252
rect 2087 13212 2320 13240
rect 2087 13209 2099 13212
rect 2041 13203 2099 13209
rect 2314 13200 2320 13212
rect 2372 13200 2378 13252
rect 8202 13240 8208 13252
rect 8163 13212 8208 13240
rect 8202 13200 8208 13212
rect 8260 13200 8266 13252
rect 4709 13175 4767 13181
rect 4709 13141 4721 13175
rect 4755 13172 4767 13175
rect 5994 13172 6000 13184
rect 4755 13144 6000 13172
rect 4755 13141 4767 13144
rect 4709 13135 4767 13141
rect 5994 13132 6000 13144
rect 6052 13132 6058 13184
rect 12176 13172 12204 13271
rect 13906 13172 13912 13184
rect 12176 13144 13912 13172
rect 13906 13132 13912 13144
rect 13964 13172 13970 13184
rect 14108 13172 14136 13271
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 15194 13200 15200 13252
rect 15252 13240 15258 13252
rect 15252 13212 18644 13240
rect 15252 13200 15258 13212
rect 14734 13172 14740 13184
rect 13964 13144 14740 13172
rect 13964 13132 13970 13144
rect 14734 13132 14740 13144
rect 14792 13132 14798 13184
rect 15933 13175 15991 13181
rect 15933 13141 15945 13175
rect 15979 13172 15991 13175
rect 18322 13172 18328 13184
rect 15979 13144 18328 13172
rect 15979 13141 15991 13144
rect 15933 13135 15991 13141
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 18616 13172 18644 13212
rect 20438 13172 20444 13184
rect 18616 13144 20444 13172
rect 20438 13132 20444 13144
rect 20496 13132 20502 13184
rect 20732 13172 20760 13339
rect 21082 13336 21088 13348
rect 21140 13336 21146 13388
rect 21542 13336 21548 13388
rect 21600 13376 21606 13388
rect 22066 13376 22094 13416
rect 27985 13413 27997 13416
rect 28031 13413 28043 13447
rect 27985 13407 28043 13413
rect 23842 13376 23848 13388
rect 21600 13348 22094 13376
rect 23803 13348 23848 13376
rect 21600 13336 21606 13348
rect 23842 13336 23848 13348
rect 23900 13336 23906 13388
rect 23937 13379 23995 13385
rect 23937 13345 23949 13379
rect 23983 13345 23995 13379
rect 23937 13339 23995 13345
rect 20901 13311 20959 13317
rect 20901 13277 20913 13311
rect 20947 13277 20959 13311
rect 20901 13271 20959 13277
rect 20806 13200 20812 13252
rect 20864 13240 20870 13252
rect 20916 13240 20944 13271
rect 21174 13268 21180 13320
rect 21232 13308 21238 13320
rect 21232 13280 22094 13308
rect 21232 13268 21238 13280
rect 20864 13212 20944 13240
rect 20864 13200 20870 13212
rect 20990 13172 20996 13184
rect 20732 13144 20996 13172
rect 20990 13132 20996 13144
rect 21048 13132 21054 13184
rect 22066 13172 22094 13280
rect 23566 13268 23572 13320
rect 23624 13308 23630 13320
rect 23952 13308 23980 13339
rect 24026 13336 24032 13388
rect 24084 13376 24090 13388
rect 24121 13379 24179 13385
rect 24121 13376 24133 13379
rect 24084 13348 24133 13376
rect 24084 13336 24090 13348
rect 24121 13345 24133 13348
rect 24167 13345 24179 13379
rect 24121 13339 24179 13345
rect 25038 13336 25044 13388
rect 25096 13376 25102 13388
rect 25205 13379 25263 13385
rect 25205 13376 25217 13379
rect 25096 13348 25217 13376
rect 25096 13336 25102 13348
rect 25205 13345 25217 13348
rect 25251 13345 25263 13379
rect 25205 13339 25263 13345
rect 23624 13280 23980 13308
rect 23624 13268 23630 13280
rect 24854 13268 24860 13320
rect 24912 13308 24918 13320
rect 24949 13311 25007 13317
rect 24949 13308 24961 13311
rect 24912 13280 24961 13308
rect 24912 13268 24918 13280
rect 24949 13277 24961 13280
rect 24995 13277 25007 13311
rect 24949 13271 25007 13277
rect 22922 13200 22928 13252
rect 22980 13240 22986 13252
rect 23106 13240 23112 13252
rect 22980 13212 23112 13240
rect 22980 13200 22986 13212
rect 23106 13200 23112 13212
rect 23164 13200 23170 13252
rect 23934 13240 23940 13252
rect 23895 13212 23940 13240
rect 23934 13200 23940 13212
rect 23992 13200 23998 13252
rect 24854 13172 24860 13184
rect 22066 13144 24860 13172
rect 24854 13132 24860 13144
rect 24912 13132 24918 13184
rect 24964 13172 24992 13271
rect 28166 13240 28172 13252
rect 28127 13212 28172 13240
rect 28166 13200 28172 13212
rect 28224 13200 28230 13252
rect 25866 13172 25872 13184
rect 24964 13144 25872 13172
rect 25866 13132 25872 13144
rect 25924 13132 25930 13184
rect 26142 13132 26148 13184
rect 26200 13172 26206 13184
rect 26329 13175 26387 13181
rect 26329 13172 26341 13175
rect 26200 13144 26341 13172
rect 26200 13132 26206 13144
rect 26329 13141 26341 13144
rect 26375 13141 26387 13175
rect 26329 13135 26387 13141
rect 1104 13082 28888 13104
rect 1104 13030 5614 13082
rect 5666 13030 5678 13082
rect 5730 13030 5742 13082
rect 5794 13030 5806 13082
rect 5858 13030 14878 13082
rect 14930 13030 14942 13082
rect 14994 13030 15006 13082
rect 15058 13030 15070 13082
rect 15122 13030 24142 13082
rect 24194 13030 24206 13082
rect 24258 13030 24270 13082
rect 24322 13030 24334 13082
rect 24386 13030 28888 13082
rect 1104 13008 28888 13030
rect 4154 12928 4160 12980
rect 4212 12968 4218 12980
rect 4341 12971 4399 12977
rect 4341 12968 4353 12971
rect 4212 12940 4353 12968
rect 4212 12928 4218 12940
rect 4341 12937 4353 12940
rect 4387 12937 4399 12971
rect 4341 12931 4399 12937
rect 5077 12971 5135 12977
rect 5077 12937 5089 12971
rect 5123 12968 5135 12971
rect 5166 12968 5172 12980
rect 5123 12940 5172 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 11606 12968 11612 12980
rect 5736 12940 11612 12968
rect 1578 12792 1584 12844
rect 1636 12832 1642 12844
rect 2041 12835 2099 12841
rect 2041 12832 2053 12835
rect 1636 12804 2053 12832
rect 1636 12792 1642 12804
rect 2041 12801 2053 12804
rect 2087 12832 2099 12835
rect 2087 12804 5028 12832
rect 2087 12801 2099 12804
rect 2041 12795 2099 12801
rect 2501 12767 2559 12773
rect 2501 12733 2513 12767
rect 2547 12764 2559 12767
rect 2774 12764 2780 12776
rect 2547 12736 2780 12764
rect 2547 12733 2559 12736
rect 2501 12727 2559 12733
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 2958 12724 2964 12776
rect 3016 12764 3022 12776
rect 4154 12764 4160 12776
rect 3016 12736 4160 12764
rect 3016 12724 3022 12736
rect 4154 12724 4160 12736
rect 4212 12724 4218 12776
rect 5000 12773 5028 12804
rect 4249 12767 4307 12773
rect 4249 12733 4261 12767
rect 4295 12733 4307 12767
rect 4249 12727 4307 12733
rect 4985 12767 5043 12773
rect 4985 12733 4997 12767
rect 5031 12764 5043 12767
rect 5736 12764 5764 12940
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 16761 12971 16819 12977
rect 11716 12940 15240 12968
rect 7006 12860 7012 12912
rect 7064 12900 7070 12912
rect 8481 12903 8539 12909
rect 8481 12900 8493 12903
rect 7064 12872 8493 12900
rect 7064 12860 7070 12872
rect 8481 12869 8493 12872
rect 8527 12869 8539 12903
rect 11716 12900 11744 12940
rect 8481 12863 8539 12869
rect 10980 12872 11744 12900
rect 11808 12872 13860 12900
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 8202 12832 8208 12844
rect 6687 12804 8064 12832
rect 8163 12804 8208 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 5902 12764 5908 12776
rect 5031 12736 5764 12764
rect 5863 12736 5908 12764
rect 5031 12733 5043 12736
rect 4985 12727 5043 12733
rect 1854 12696 1860 12708
rect 1815 12668 1860 12696
rect 1854 12656 1860 12668
rect 1912 12656 1918 12708
rect 4264 12696 4292 12727
rect 5902 12724 5908 12736
rect 5960 12724 5966 12776
rect 5994 12724 6000 12776
rect 6052 12764 6058 12776
rect 6178 12764 6184 12776
rect 6052 12736 6097 12764
rect 6139 12736 6184 12764
rect 6052 12724 6058 12736
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 7190 12764 7196 12776
rect 7151 12736 7196 12764
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 7466 12764 7472 12776
rect 7427 12736 7472 12764
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 7834 12764 7840 12776
rect 7795 12736 7840 12764
rect 7834 12724 7840 12736
rect 7892 12724 7898 12776
rect 8036 12764 8064 12804
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 10686 12764 10692 12776
rect 8036 12736 10692 12764
rect 10686 12724 10692 12736
rect 10744 12724 10750 12776
rect 4264 12668 5212 12696
rect 5184 12640 5212 12668
rect 7282 12656 7288 12708
rect 7340 12696 7346 12708
rect 7852 12696 7880 12724
rect 10980 12696 11008 12872
rect 11057 12835 11115 12841
rect 11057 12801 11069 12835
rect 11103 12832 11115 12835
rect 11808 12832 11836 12872
rect 11103 12804 11836 12832
rect 11103 12801 11115 12804
rect 11057 12795 11115 12801
rect 11974 12792 11980 12844
rect 12032 12832 12038 12844
rect 13832 12832 13860 12872
rect 13906 12860 13912 12912
rect 13964 12900 13970 12912
rect 14090 12900 14096 12912
rect 13964 12872 14096 12900
rect 13964 12860 13970 12872
rect 14090 12860 14096 12872
rect 14148 12860 14154 12912
rect 15102 12832 15108 12844
rect 12032 12804 12098 12832
rect 13832 12804 15108 12832
rect 12032 12792 12038 12804
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 11790 12724 11796 12776
rect 11848 12724 11854 12776
rect 13630 12764 13636 12776
rect 13591 12736 13636 12764
rect 13630 12724 13636 12736
rect 13688 12724 13694 12776
rect 13817 12767 13875 12773
rect 13817 12733 13829 12767
rect 13863 12764 13875 12767
rect 14182 12764 14188 12776
rect 13863 12736 14188 12764
rect 13863 12733 13875 12736
rect 13817 12727 13875 12733
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 15212 12764 15240 12940
rect 16761 12937 16773 12971
rect 16807 12968 16819 12971
rect 17494 12968 17500 12980
rect 16807 12940 17500 12968
rect 16807 12937 16819 12940
rect 16761 12931 16819 12937
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 17678 12968 17684 12980
rect 17639 12940 17684 12968
rect 17678 12928 17684 12940
rect 17736 12928 17742 12980
rect 18524 12940 18920 12968
rect 18524 12900 18552 12940
rect 16592 12872 18552 12900
rect 18785 12903 18843 12909
rect 16114 12792 16120 12844
rect 16172 12792 16178 12844
rect 15749 12767 15807 12773
rect 15749 12764 15761 12767
rect 15212 12736 15761 12764
rect 15749 12733 15761 12736
rect 15795 12764 15807 12767
rect 16592 12764 16620 12872
rect 18785 12869 18797 12903
rect 18831 12869 18843 12903
rect 18892 12900 18920 12940
rect 19150 12928 19156 12980
rect 19208 12968 19214 12980
rect 22278 12968 22284 12980
rect 19208 12940 22284 12968
rect 19208 12928 19214 12940
rect 22278 12928 22284 12940
rect 22336 12928 22342 12980
rect 23845 12971 23903 12977
rect 23845 12937 23857 12971
rect 23891 12968 23903 12971
rect 24026 12968 24032 12980
rect 23891 12940 24032 12968
rect 23891 12937 23903 12940
rect 23845 12931 23903 12937
rect 24026 12928 24032 12940
rect 24084 12928 24090 12980
rect 26694 12968 26700 12980
rect 26655 12940 26700 12968
rect 26694 12928 26700 12940
rect 26752 12928 26758 12980
rect 21174 12900 21180 12912
rect 18892 12872 21180 12900
rect 18785 12863 18843 12869
rect 17678 12792 17684 12844
rect 17736 12832 17742 12844
rect 17736 12804 18276 12832
rect 17736 12792 17742 12804
rect 15795 12736 16620 12764
rect 15795 12733 15807 12736
rect 15749 12727 15807 12733
rect 17034 12724 17040 12776
rect 17092 12764 17098 12776
rect 17405 12767 17463 12773
rect 17405 12764 17417 12767
rect 17092 12736 17417 12764
rect 17092 12724 17098 12736
rect 17405 12733 17417 12736
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 17494 12724 17500 12776
rect 17552 12764 17558 12776
rect 17862 12764 17868 12776
rect 17552 12736 17597 12764
rect 17823 12736 17868 12764
rect 17552 12724 17558 12736
rect 17862 12724 17868 12736
rect 17920 12724 17926 12776
rect 17954 12724 17960 12776
rect 18012 12764 18018 12776
rect 18138 12764 18144 12776
rect 18012 12736 18144 12764
rect 18012 12724 18018 12736
rect 18138 12724 18144 12736
rect 18196 12724 18202 12776
rect 18248 12764 18276 12804
rect 18322 12792 18328 12844
rect 18380 12832 18386 12844
rect 18800 12832 18828 12863
rect 21174 12860 21180 12872
rect 21232 12860 21238 12912
rect 22094 12860 22100 12912
rect 22152 12900 22158 12912
rect 22152 12872 22600 12900
rect 22152 12860 22158 12872
rect 22572 12844 22600 12872
rect 19150 12832 19156 12844
rect 18380 12804 18644 12832
rect 18800 12804 19156 12832
rect 18380 12792 18386 12804
rect 18509 12767 18567 12773
rect 18509 12764 18521 12767
rect 18248 12736 18521 12764
rect 18509 12733 18521 12736
rect 18555 12733 18567 12767
rect 18616 12764 18644 12804
rect 19150 12792 19156 12804
rect 19208 12792 19214 12844
rect 22554 12792 22560 12844
rect 22612 12792 22618 12844
rect 27890 12832 27896 12844
rect 25516 12776 25544 12818
rect 27851 12804 27896 12832
rect 27890 12792 27896 12804
rect 27948 12792 27954 12844
rect 28077 12835 28135 12841
rect 28077 12801 28089 12835
rect 28123 12832 28135 12835
rect 28350 12832 28356 12844
rect 28123 12804 28356 12832
rect 28123 12801 28135 12804
rect 28077 12795 28135 12801
rect 28350 12792 28356 12804
rect 28408 12792 28414 12844
rect 18797 12767 18855 12773
rect 18797 12764 18809 12767
rect 18616 12736 18809 12764
rect 18509 12727 18567 12733
rect 18797 12733 18809 12736
rect 18843 12733 18855 12767
rect 18797 12727 18855 12733
rect 21358 12724 21364 12776
rect 21416 12764 21422 12776
rect 21729 12767 21787 12773
rect 21729 12764 21741 12767
rect 21416 12736 21741 12764
rect 21416 12724 21422 12736
rect 21729 12733 21741 12736
rect 21775 12733 21787 12767
rect 22925 12767 22983 12773
rect 21729 12727 21787 12733
rect 21836 12736 22876 12764
rect 7340 12668 7880 12696
rect 9646 12668 11008 12696
rect 7340 12656 7346 12668
rect 2685 12631 2743 12637
rect 2685 12597 2697 12631
rect 2731 12628 2743 12631
rect 3970 12628 3976 12640
rect 2731 12600 3976 12628
rect 2731 12597 2743 12600
rect 2685 12591 2743 12597
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 5166 12588 5172 12640
rect 5224 12628 5230 12640
rect 9646 12628 9674 12668
rect 13722 12656 13728 12708
rect 13780 12696 13786 12708
rect 15473 12699 15531 12705
rect 15473 12696 15485 12699
rect 13780 12668 15485 12696
rect 13780 12656 13786 12668
rect 15473 12665 15485 12668
rect 15519 12665 15531 12699
rect 15473 12659 15531 12665
rect 12066 12628 12072 12640
rect 5224 12600 9674 12628
rect 12027 12600 12072 12628
rect 5224 12588 5230 12600
rect 12066 12588 12072 12600
rect 12124 12588 12130 12640
rect 12250 12588 12256 12640
rect 12308 12628 12314 12640
rect 13630 12628 13636 12640
rect 12308 12600 13636 12628
rect 12308 12588 12314 12600
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 13817 12631 13875 12637
rect 13817 12597 13829 12631
rect 13863 12628 13875 12631
rect 14458 12628 14464 12640
rect 13863 12600 14464 12628
rect 13863 12597 13875 12600
rect 13817 12591 13875 12597
rect 14458 12588 14464 12600
rect 14516 12588 14522 12640
rect 15488 12628 15516 12659
rect 15562 12656 15568 12708
rect 15620 12696 15626 12708
rect 15841 12699 15899 12705
rect 15841 12696 15853 12699
rect 15620 12668 15853 12696
rect 15620 12656 15626 12668
rect 15841 12665 15853 12668
rect 15887 12665 15899 12699
rect 15841 12659 15899 12665
rect 16209 12699 16267 12705
rect 16209 12665 16221 12699
rect 16255 12696 16267 12699
rect 18322 12696 18328 12708
rect 16255 12668 18328 12696
rect 16255 12665 16267 12668
rect 16209 12659 16267 12665
rect 18322 12656 18328 12668
rect 18380 12656 18386 12708
rect 18690 12696 18696 12708
rect 18651 12668 18696 12696
rect 18690 12656 18696 12668
rect 18748 12656 18754 12708
rect 21836 12696 21864 12736
rect 21192 12668 21864 12696
rect 16390 12628 16396 12640
rect 15488 12600 16396 12628
rect 16390 12588 16396 12600
rect 16448 12588 16454 12640
rect 16574 12628 16580 12640
rect 16535 12600 16580 12628
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 21192 12628 21220 12668
rect 22278 12656 22284 12708
rect 22336 12696 22342 12708
rect 22848 12705 22876 12736
rect 22925 12733 22937 12767
rect 22971 12764 22983 12767
rect 23106 12764 23112 12776
rect 22971 12736 23112 12764
rect 22971 12733 22983 12736
rect 22925 12727 22983 12733
rect 23106 12724 23112 12736
rect 23164 12724 23170 12776
rect 23290 12764 23296 12776
rect 23251 12736 23296 12764
rect 23290 12724 23296 12736
rect 23348 12764 23354 12776
rect 23348 12736 24440 12764
rect 23348 12724 23354 12736
rect 22833 12699 22891 12705
rect 22336 12668 22692 12696
rect 22336 12656 22342 12668
rect 17460 12600 21220 12628
rect 17460 12588 17466 12600
rect 21266 12588 21272 12640
rect 21324 12628 21330 12640
rect 21545 12631 21603 12637
rect 21545 12628 21557 12631
rect 21324 12600 21557 12628
rect 21324 12588 21330 12600
rect 21545 12597 21557 12600
rect 21591 12597 21603 12631
rect 22554 12628 22560 12640
rect 22515 12600 22560 12628
rect 21545 12591 21603 12597
rect 22554 12588 22560 12600
rect 22612 12588 22618 12640
rect 22664 12628 22692 12668
rect 22833 12665 22845 12699
rect 22879 12696 22891 12699
rect 23382 12696 23388 12708
rect 22879 12668 23388 12696
rect 22879 12665 22891 12668
rect 22833 12659 22891 12665
rect 23382 12656 23388 12668
rect 23440 12656 23446 12708
rect 24412 12696 24440 12736
rect 25498 12724 25504 12776
rect 25556 12724 25562 12776
rect 25590 12724 25596 12776
rect 25648 12764 25654 12776
rect 26142 12764 26148 12776
rect 25648 12736 25820 12764
rect 26103 12736 26148 12764
rect 25648 12724 25654 12736
rect 25222 12696 25228 12708
rect 24412 12668 25228 12696
rect 25222 12656 25228 12668
rect 25280 12696 25286 12708
rect 25409 12699 25467 12705
rect 25409 12696 25421 12699
rect 25280 12668 25421 12696
rect 25280 12656 25286 12668
rect 25409 12665 25421 12668
rect 25455 12665 25467 12699
rect 25682 12696 25688 12708
rect 25643 12668 25688 12696
rect 25409 12659 25467 12665
rect 25682 12656 25688 12668
rect 25740 12656 25746 12708
rect 25792 12705 25820 12736
rect 26142 12724 26148 12736
rect 26200 12724 26206 12776
rect 25777 12699 25835 12705
rect 25777 12665 25789 12699
rect 25823 12696 25835 12699
rect 26050 12696 26056 12708
rect 25823 12668 26056 12696
rect 25823 12665 25835 12668
rect 25777 12659 25835 12665
rect 26050 12656 26056 12668
rect 26108 12656 26114 12708
rect 23661 12631 23719 12637
rect 23661 12628 23673 12631
rect 22664 12600 23673 12628
rect 23661 12597 23673 12600
rect 23707 12597 23719 12631
rect 26510 12628 26516 12640
rect 26471 12600 26516 12628
rect 23661 12591 23719 12597
rect 26510 12588 26516 12600
rect 26568 12588 26574 12640
rect 27430 12628 27436 12640
rect 27391 12600 27436 12628
rect 27430 12588 27436 12600
rect 27488 12588 27494 12640
rect 27522 12588 27528 12640
rect 27580 12628 27586 12640
rect 27801 12631 27859 12637
rect 27801 12628 27813 12631
rect 27580 12600 27813 12628
rect 27580 12588 27586 12600
rect 27801 12597 27813 12600
rect 27847 12597 27859 12631
rect 27801 12591 27859 12597
rect 1104 12538 28888 12560
rect 1104 12486 10246 12538
rect 10298 12486 10310 12538
rect 10362 12486 10374 12538
rect 10426 12486 10438 12538
rect 10490 12486 19510 12538
rect 19562 12486 19574 12538
rect 19626 12486 19638 12538
rect 19690 12486 19702 12538
rect 19754 12486 28888 12538
rect 1104 12464 28888 12486
rect 1578 12424 1584 12436
rect 1539 12396 1584 12424
rect 1578 12384 1584 12396
rect 1636 12384 1642 12436
rect 2590 12384 2596 12436
rect 2648 12424 2654 12436
rect 2869 12427 2927 12433
rect 2869 12424 2881 12427
rect 2648 12396 2881 12424
rect 2648 12384 2654 12396
rect 2869 12393 2881 12396
rect 2915 12393 2927 12427
rect 2869 12387 2927 12393
rect 3234 12384 3240 12436
rect 3292 12424 3298 12436
rect 4798 12424 4804 12436
rect 3292 12396 4804 12424
rect 3292 12384 3298 12396
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 5813 12427 5871 12433
rect 5813 12393 5825 12427
rect 5859 12424 5871 12427
rect 5902 12424 5908 12436
rect 5859 12396 5908 12424
rect 5859 12393 5871 12396
rect 5813 12387 5871 12393
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 7193 12427 7251 12433
rect 7193 12393 7205 12427
rect 7239 12424 7251 12427
rect 8110 12424 8116 12436
rect 7239 12396 8116 12424
rect 7239 12393 7251 12396
rect 7193 12387 7251 12393
rect 8110 12384 8116 12396
rect 8168 12384 8174 12436
rect 13446 12424 13452 12436
rect 9324 12396 11008 12424
rect 1857 12359 1915 12365
rect 1857 12325 1869 12359
rect 1903 12356 1915 12359
rect 2682 12356 2688 12368
rect 1903 12328 2452 12356
rect 2643 12328 2688 12356
rect 1903 12325 1915 12328
rect 1857 12319 1915 12325
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 2038 12288 2044 12300
rect 1995 12260 2044 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 2314 12288 2320 12300
rect 2275 12260 2320 12288
rect 2314 12248 2320 12260
rect 2372 12248 2378 12300
rect 2424 12288 2452 12328
rect 2682 12316 2688 12328
rect 2740 12316 2746 12368
rect 4522 12316 4528 12368
rect 4580 12356 4586 12368
rect 9324 12356 9352 12396
rect 4580 12328 9352 12356
rect 9401 12359 9459 12365
rect 4580 12316 4586 12328
rect 9401 12325 9413 12359
rect 9447 12356 9459 12359
rect 9582 12356 9588 12368
rect 9447 12328 9588 12356
rect 9447 12325 9459 12328
rect 9401 12319 9459 12325
rect 9582 12316 9588 12328
rect 9640 12316 9646 12368
rect 2424 12260 2774 12288
rect 1400 12232 1452 12238
rect 2746 12220 2774 12260
rect 3326 12248 3332 12300
rect 3384 12288 3390 12300
rect 3421 12291 3479 12297
rect 3421 12288 3433 12291
rect 3384 12260 3433 12288
rect 3384 12248 3390 12260
rect 3421 12257 3433 12260
rect 3467 12257 3479 12291
rect 3421 12251 3479 12257
rect 3694 12248 3700 12300
rect 3752 12288 3758 12300
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 3752 12260 4077 12288
rect 3752 12248 3758 12260
rect 4065 12257 4077 12260
rect 4111 12257 4123 12291
rect 4065 12251 4123 12257
rect 5721 12291 5779 12297
rect 5721 12257 5733 12291
rect 5767 12288 5779 12291
rect 6362 12288 6368 12300
rect 5767 12260 6368 12288
rect 5767 12257 5779 12260
rect 5721 12251 5779 12257
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 7282 12248 7288 12300
rect 7340 12288 7346 12300
rect 7561 12291 7619 12297
rect 7561 12288 7573 12291
rect 7340 12260 7573 12288
rect 7340 12248 7346 12260
rect 7561 12257 7573 12260
rect 7607 12257 7619 12291
rect 7561 12251 7619 12257
rect 7653 12291 7711 12297
rect 7653 12257 7665 12291
rect 7699 12288 7711 12291
rect 8202 12288 8208 12300
rect 7699 12260 8208 12288
rect 7699 12257 7711 12260
rect 7653 12251 7711 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 9214 12288 9220 12300
rect 9175 12260 9220 12288
rect 9214 12248 9220 12260
rect 9272 12248 9278 12300
rect 9858 12248 9864 12300
rect 9916 12288 9922 12300
rect 10980 12297 11008 12396
rect 12636 12396 13452 12424
rect 11238 12316 11244 12368
rect 11296 12356 11302 12368
rect 11296 12328 12204 12356
rect 11296 12316 11302 12328
rect 10229 12291 10287 12297
rect 10229 12288 10241 12291
rect 9916 12260 10241 12288
rect 9916 12248 9922 12260
rect 10229 12257 10241 12260
rect 10275 12257 10287 12291
rect 10229 12251 10287 12257
rect 10965 12291 11023 12297
rect 10965 12257 10977 12291
rect 11011 12288 11023 12291
rect 11330 12288 11336 12300
rect 11011 12260 11336 12288
rect 11011 12257 11023 12260
rect 10965 12251 11023 12257
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 2866 12220 2872 12232
rect 2746 12192 2872 12220
rect 2866 12180 2872 12192
rect 2924 12220 2930 12232
rect 7374 12220 7380 12232
rect 2924 12192 4016 12220
rect 7335 12192 7380 12220
rect 2924 12180 2930 12192
rect 1400 12174 1452 12180
rect 3602 12152 3608 12164
rect 3563 12124 3608 12152
rect 3602 12112 3608 12124
rect 3660 12112 3666 12164
rect 3988 12152 4016 12192
rect 7374 12180 7380 12192
rect 7432 12180 7438 12232
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 7524 12192 7569 12220
rect 7524 12180 7530 12192
rect 9398 12180 9404 12232
rect 9456 12220 9462 12232
rect 9493 12223 9551 12229
rect 9493 12220 9505 12223
rect 9456 12192 9505 12220
rect 9456 12180 9462 12192
rect 9493 12189 9505 12192
rect 9539 12189 9551 12223
rect 11606 12220 11612 12232
rect 9493 12183 9551 12189
rect 9600 12192 11612 12220
rect 9600 12152 9628 12192
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 12176 12220 12204 12328
rect 12636 12297 12664 12396
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 13814 12424 13820 12436
rect 13775 12396 13820 12424
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 14274 12424 14280 12436
rect 14187 12396 14280 12424
rect 14274 12384 14280 12396
rect 14332 12424 14338 12436
rect 15746 12424 15752 12436
rect 14332 12396 15752 12424
rect 14332 12384 14338 12396
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 18322 12384 18328 12436
rect 18380 12424 18386 12436
rect 19153 12427 19211 12433
rect 19153 12424 19165 12427
rect 18380 12396 19165 12424
rect 18380 12384 18386 12396
rect 19153 12393 19165 12396
rect 19199 12424 19211 12427
rect 19242 12424 19248 12436
rect 19199 12396 19248 12424
rect 19199 12393 19211 12396
rect 19153 12387 19211 12393
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 19978 12424 19984 12436
rect 19904 12396 19984 12424
rect 13630 12356 13636 12368
rect 13004 12328 13636 12356
rect 12601 12291 12664 12297
rect 12601 12257 12613 12291
rect 12647 12260 12664 12291
rect 12713 12291 12771 12297
rect 12647 12257 12659 12260
rect 12601 12251 12659 12257
rect 12713 12257 12725 12291
rect 12759 12257 12771 12291
rect 12713 12251 12771 12257
rect 12345 12223 12403 12229
rect 12345 12220 12357 12223
rect 12176 12192 12357 12220
rect 12345 12189 12357 12192
rect 12391 12189 12403 12223
rect 12345 12183 12403 12189
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 12728 12220 12756 12251
rect 12802 12248 12808 12300
rect 12860 12288 12866 12300
rect 13004 12297 13032 12328
rect 13630 12316 13636 12328
rect 13688 12316 13694 12368
rect 12989 12291 13047 12297
rect 12860 12260 12905 12288
rect 12860 12248 12866 12260
rect 12989 12257 13001 12291
rect 13035 12257 13047 12291
rect 12989 12251 13047 12257
rect 13078 12248 13084 12300
rect 13136 12288 13142 12300
rect 13814 12288 13820 12300
rect 13136 12260 13820 12288
rect 13136 12248 13142 12260
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 14292 12297 14320 12384
rect 15286 12316 15292 12368
rect 15344 12356 15350 12368
rect 15838 12356 15844 12368
rect 15344 12328 15844 12356
rect 15344 12316 15350 12328
rect 15838 12316 15844 12328
rect 15896 12316 15902 12368
rect 16025 12359 16083 12365
rect 16025 12325 16037 12359
rect 16071 12356 16083 12359
rect 17218 12356 17224 12368
rect 16071 12328 17224 12356
rect 16071 12325 16083 12328
rect 16025 12319 16083 12325
rect 17218 12316 17224 12328
rect 17276 12316 17282 12368
rect 18598 12356 18604 12368
rect 17328 12328 18604 12356
rect 14093 12291 14151 12297
rect 14093 12288 14105 12291
rect 13964 12260 14105 12288
rect 13964 12248 13970 12260
rect 14093 12257 14105 12260
rect 14139 12257 14151 12291
rect 14093 12251 14151 12257
rect 14185 12291 14243 12297
rect 14185 12257 14197 12291
rect 14231 12257 14243 12291
rect 14185 12251 14243 12257
rect 14277 12291 14335 12297
rect 14277 12257 14289 12291
rect 14323 12257 14335 12291
rect 14458 12288 14464 12300
rect 14419 12260 14464 12288
rect 14277 12251 14335 12257
rect 13630 12220 13636 12232
rect 12492 12192 13636 12220
rect 12492 12180 12498 12192
rect 13630 12180 13636 12192
rect 13688 12220 13694 12232
rect 14200 12220 14228 12251
rect 14458 12248 14464 12260
rect 14516 12248 14522 12300
rect 15378 12288 15384 12300
rect 15339 12260 15384 12288
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 15565 12291 15623 12297
rect 15565 12257 15577 12291
rect 15611 12288 15623 12291
rect 15654 12288 15660 12300
rect 15611 12260 15660 12288
rect 15611 12257 15623 12260
rect 15565 12251 15623 12257
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 15286 12220 15292 12232
rect 13688 12192 14228 12220
rect 15247 12192 15292 12220
rect 13688 12180 13694 12192
rect 15286 12180 15292 12192
rect 15344 12220 15350 12232
rect 16206 12220 16212 12232
rect 15344 12192 16212 12220
rect 15344 12180 15350 12192
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 17328 12152 17356 12328
rect 18598 12316 18604 12328
rect 18656 12316 18662 12368
rect 19334 12316 19340 12368
rect 19392 12356 19398 12368
rect 19904 12365 19932 12396
rect 19978 12384 19984 12396
rect 20036 12424 20042 12436
rect 20441 12427 20499 12433
rect 20036 12396 20392 12424
rect 20036 12384 20042 12396
rect 19521 12359 19579 12365
rect 19521 12356 19533 12359
rect 19392 12328 19533 12356
rect 19392 12316 19398 12328
rect 19521 12325 19533 12328
rect 19567 12325 19579 12359
rect 19521 12319 19579 12325
rect 19889 12359 19947 12365
rect 19889 12325 19901 12359
rect 19935 12325 19947 12359
rect 20254 12356 20260 12368
rect 20215 12328 20260 12356
rect 19889 12319 19947 12325
rect 20254 12316 20260 12328
rect 20312 12316 20318 12368
rect 20364 12356 20392 12396
rect 20441 12393 20453 12427
rect 20487 12424 20499 12427
rect 21082 12424 21088 12436
rect 20487 12396 21088 12424
rect 20487 12393 20499 12396
rect 20441 12387 20499 12393
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 22554 12424 22560 12436
rect 21192 12396 22560 12424
rect 21192 12356 21220 12396
rect 22554 12384 22560 12396
rect 22612 12384 22618 12436
rect 24489 12427 24547 12433
rect 24489 12393 24501 12427
rect 24535 12424 24547 12427
rect 25317 12427 25375 12433
rect 25317 12424 25329 12427
rect 24535 12396 25329 12424
rect 24535 12393 24547 12396
rect 24489 12387 24547 12393
rect 25317 12393 25329 12396
rect 25363 12393 25375 12427
rect 25317 12387 25375 12393
rect 25406 12384 25412 12436
rect 25464 12424 25470 12436
rect 26142 12424 26148 12436
rect 25464 12396 26148 12424
rect 25464 12384 25470 12396
rect 26142 12384 26148 12396
rect 26200 12384 26206 12436
rect 26881 12427 26939 12433
rect 26881 12393 26893 12427
rect 26927 12424 26939 12427
rect 27522 12424 27528 12436
rect 26927 12396 27528 12424
rect 26927 12393 26939 12396
rect 26881 12387 26939 12393
rect 27522 12384 27528 12396
rect 27580 12384 27586 12436
rect 20364 12328 21220 12356
rect 21358 12316 21364 12368
rect 21416 12356 21422 12368
rect 21416 12328 22784 12356
rect 21416 12316 21422 12328
rect 19242 12248 19248 12300
rect 19300 12288 19306 12300
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 19300 12260 19441 12288
rect 19300 12248 19306 12260
rect 19429 12257 19441 12260
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 21269 12291 21327 12297
rect 21269 12257 21281 12291
rect 21315 12288 21327 12291
rect 21910 12288 21916 12300
rect 21315 12260 21916 12288
rect 21315 12257 21327 12260
rect 21269 12251 21327 12257
rect 21910 12248 21916 12260
rect 21968 12288 21974 12300
rect 22756 12297 22784 12328
rect 23382 12316 23388 12368
rect 23440 12356 23446 12368
rect 27985 12359 28043 12365
rect 27985 12356 27997 12359
rect 23440 12328 27997 12356
rect 23440 12316 23446 12328
rect 27985 12325 27997 12328
rect 28031 12325 28043 12359
rect 27985 12319 28043 12325
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 21968 12260 22017 12288
rect 21968 12248 21974 12260
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 22741 12291 22799 12297
rect 22741 12257 22753 12291
rect 22787 12257 22799 12291
rect 22741 12251 22799 12257
rect 23934 12248 23940 12300
rect 23992 12288 23998 12300
rect 24121 12291 24179 12297
rect 24121 12288 24133 12291
rect 23992 12260 24133 12288
rect 23992 12248 23998 12260
rect 24121 12257 24133 12260
rect 24167 12257 24179 12291
rect 24121 12251 24179 12257
rect 26513 12291 26571 12297
rect 26513 12257 26525 12291
rect 26559 12288 26571 12291
rect 26694 12288 26700 12300
rect 26559 12260 26700 12288
rect 26559 12257 26571 12260
rect 26513 12251 26571 12257
rect 26694 12248 26700 12260
rect 26752 12248 26758 12300
rect 18972 12232 19024 12238
rect 18598 12180 18604 12232
rect 18656 12220 18662 12232
rect 18656 12192 18972 12220
rect 18656 12180 18662 12192
rect 20806 12180 20812 12232
rect 20864 12220 20870 12232
rect 21174 12220 21180 12232
rect 20864 12192 21180 12220
rect 20864 12180 20870 12192
rect 21174 12180 21180 12192
rect 21232 12180 21238 12232
rect 21361 12223 21419 12229
rect 21361 12189 21373 12223
rect 21407 12189 21419 12223
rect 21361 12183 21419 12189
rect 21453 12223 21511 12229
rect 21453 12189 21465 12223
rect 21499 12220 21511 12223
rect 23382 12220 23388 12232
rect 21499 12192 23388 12220
rect 21499 12189 21511 12192
rect 21453 12183 21511 12189
rect 18972 12174 19024 12180
rect 3988 12124 9628 12152
rect 9876 12124 17356 12152
rect 3786 12044 3792 12096
rect 3844 12084 3850 12096
rect 4709 12087 4767 12093
rect 4709 12084 4721 12087
rect 3844 12056 4721 12084
rect 3844 12044 3850 12056
rect 4709 12053 4721 12056
rect 4755 12053 4767 12087
rect 4709 12047 4767 12053
rect 4982 12044 4988 12096
rect 5040 12084 5046 12096
rect 5902 12084 5908 12096
rect 5040 12056 5908 12084
rect 5040 12044 5046 12056
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 7282 12044 7288 12096
rect 7340 12084 7346 12096
rect 7466 12084 7472 12096
rect 7340 12056 7472 12084
rect 7340 12044 7346 12056
rect 7466 12044 7472 12056
rect 7524 12044 7530 12096
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 8110 12084 8116 12096
rect 7800 12056 8116 12084
rect 7800 12044 7806 12056
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8260 12056 8953 12084
rect 8260 12044 8266 12056
rect 8941 12053 8953 12056
rect 8987 12053 8999 12087
rect 8941 12047 8999 12053
rect 9122 12044 9128 12096
rect 9180 12084 9186 12096
rect 9876 12084 9904 12124
rect 20530 12112 20536 12164
rect 20588 12152 20594 12164
rect 21376 12152 21404 12183
rect 23382 12180 23388 12192
rect 23440 12180 23446 12232
rect 23842 12180 23848 12232
rect 23900 12220 23906 12232
rect 24213 12223 24271 12229
rect 24213 12220 24225 12223
rect 23900 12192 24225 12220
rect 23900 12180 23906 12192
rect 24213 12189 24225 12192
rect 24259 12220 24271 12223
rect 24762 12220 24768 12232
rect 24259 12192 24768 12220
rect 24259 12189 24271 12192
rect 24213 12183 24271 12189
rect 24762 12180 24768 12192
rect 24820 12180 24826 12232
rect 25593 12223 25651 12229
rect 25593 12189 25605 12223
rect 25639 12220 25651 12223
rect 26234 12220 26240 12232
rect 25639 12192 26240 12220
rect 25639 12189 25651 12192
rect 25593 12183 25651 12189
rect 20588 12124 21404 12152
rect 22005 12155 22063 12161
rect 20588 12112 20594 12124
rect 22005 12121 22017 12155
rect 22051 12152 22063 12155
rect 23290 12152 23296 12164
rect 22051 12124 23296 12152
rect 22051 12121 22063 12124
rect 22005 12115 22063 12121
rect 23290 12112 23296 12124
rect 23348 12112 23354 12164
rect 24949 12155 25007 12161
rect 24949 12121 24961 12155
rect 24995 12152 25007 12155
rect 25038 12152 25044 12164
rect 24995 12124 25044 12152
rect 24995 12121 25007 12124
rect 24949 12115 25007 12121
rect 25038 12112 25044 12124
rect 25096 12112 25102 12164
rect 25222 12112 25228 12164
rect 25280 12152 25286 12164
rect 25608 12152 25636 12183
rect 26234 12180 26240 12192
rect 26292 12180 26298 12232
rect 26418 12220 26424 12232
rect 26379 12192 26424 12220
rect 26418 12180 26424 12192
rect 26476 12180 26482 12232
rect 25280 12124 25636 12152
rect 28169 12155 28227 12161
rect 25280 12112 25286 12124
rect 28169 12121 28181 12155
rect 28215 12152 28227 12155
rect 28997 12155 29055 12161
rect 28997 12152 29009 12155
rect 28215 12124 29009 12152
rect 28215 12121 28227 12124
rect 28169 12115 28227 12121
rect 28997 12121 29009 12124
rect 29043 12121 29055 12155
rect 28997 12115 29055 12121
rect 9180 12056 9904 12084
rect 9180 12044 9186 12056
rect 9950 12044 9956 12096
rect 10008 12084 10014 12096
rect 10321 12087 10379 12093
rect 10321 12084 10333 12087
rect 10008 12056 10333 12084
rect 10008 12044 10014 12056
rect 10321 12053 10333 12056
rect 10367 12053 10379 12087
rect 10321 12047 10379 12053
rect 11057 12087 11115 12093
rect 11057 12053 11069 12087
rect 11103 12084 11115 12087
rect 11238 12084 11244 12096
rect 11103 12056 11244 12084
rect 11103 12053 11115 12056
rect 11057 12047 11115 12053
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 20993 12087 21051 12093
rect 20993 12053 21005 12087
rect 21039 12084 21051 12087
rect 21358 12084 21364 12096
rect 21039 12056 21364 12084
rect 21039 12053 21051 12056
rect 20993 12047 21051 12053
rect 21358 12044 21364 12056
rect 21416 12044 21422 12096
rect 21450 12044 21456 12096
rect 21508 12084 21514 12096
rect 22557 12087 22615 12093
rect 22557 12084 22569 12087
rect 21508 12056 22569 12084
rect 21508 12044 21514 12056
rect 22557 12053 22569 12056
rect 22603 12084 22615 12087
rect 25958 12084 25964 12096
rect 22603 12056 25964 12084
rect 22603 12053 22615 12056
rect 22557 12047 22615 12053
rect 25958 12044 25964 12056
rect 26016 12044 26022 12096
rect 1104 11994 28888 12016
rect 1104 11942 5614 11994
rect 5666 11942 5678 11994
rect 5730 11942 5742 11994
rect 5794 11942 5806 11994
rect 5858 11942 14878 11994
rect 14930 11942 14942 11994
rect 14994 11942 15006 11994
rect 15058 11942 15070 11994
rect 15122 11942 24142 11994
rect 24194 11942 24206 11994
rect 24258 11942 24270 11994
rect 24322 11942 24334 11994
rect 24386 11942 28888 11994
rect 1104 11920 28888 11942
rect 2593 11883 2651 11889
rect 2593 11849 2605 11883
rect 2639 11880 2651 11883
rect 2866 11880 2872 11892
rect 2639 11852 2872 11880
rect 2639 11849 2651 11852
rect 2593 11843 2651 11849
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 6362 11880 6368 11892
rect 6323 11852 6368 11880
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 7561 11883 7619 11889
rect 7561 11849 7573 11883
rect 7607 11880 7619 11883
rect 7650 11880 7656 11892
rect 7607 11852 7656 11880
rect 7607 11849 7619 11852
rect 7561 11843 7619 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 8297 11883 8355 11889
rect 8297 11849 8309 11883
rect 8343 11880 8355 11883
rect 9122 11880 9128 11892
rect 8343 11852 9128 11880
rect 8343 11849 8355 11852
rect 8297 11843 8355 11849
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 9582 11880 9588 11892
rect 9543 11852 9588 11880
rect 9582 11840 9588 11852
rect 9640 11840 9646 11892
rect 10781 11883 10839 11889
rect 10781 11849 10793 11883
rect 10827 11880 10839 11883
rect 11790 11880 11796 11892
rect 10827 11852 11796 11880
rect 10827 11849 10839 11852
rect 10781 11843 10839 11849
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 12066 11840 12072 11892
rect 12124 11880 12130 11892
rect 12989 11883 13047 11889
rect 12989 11880 13001 11883
rect 12124 11852 13001 11880
rect 12124 11840 12130 11852
rect 12989 11849 13001 11852
rect 13035 11849 13047 11883
rect 20530 11880 20536 11892
rect 20491 11852 20536 11880
rect 12989 11843 13047 11849
rect 20530 11840 20536 11852
rect 20588 11840 20594 11892
rect 23382 11840 23388 11892
rect 23440 11880 23446 11892
rect 23753 11883 23811 11889
rect 23753 11880 23765 11883
rect 23440 11852 23765 11880
rect 23440 11840 23446 11852
rect 23753 11849 23765 11852
rect 23799 11849 23811 11883
rect 23753 11843 23811 11849
rect 25038 11840 25044 11892
rect 25096 11880 25102 11892
rect 25222 11880 25228 11892
rect 25096 11852 25228 11880
rect 25096 11840 25102 11852
rect 25222 11840 25228 11852
rect 25280 11840 25286 11892
rect 27890 11840 27896 11892
rect 27948 11880 27954 11892
rect 28169 11883 28227 11889
rect 28169 11880 28181 11883
rect 27948 11852 28181 11880
rect 27948 11840 27954 11852
rect 28169 11849 28181 11852
rect 28215 11849 28227 11883
rect 28169 11843 28227 11849
rect 1765 11815 1823 11821
rect 1765 11781 1777 11815
rect 1811 11812 1823 11815
rect 5813 11815 5871 11821
rect 1811 11784 2774 11812
rect 1811 11781 1823 11784
rect 1765 11775 1823 11781
rect 1486 11636 1492 11688
rect 1544 11676 1550 11688
rect 1949 11679 2007 11685
rect 1949 11676 1961 11679
rect 1544 11648 1961 11676
rect 1544 11636 1550 11648
rect 1949 11645 1961 11648
rect 1995 11645 2007 11679
rect 2406 11676 2412 11688
rect 2367 11648 2412 11676
rect 1949 11639 2007 11645
rect 2406 11636 2412 11648
rect 2464 11636 2470 11688
rect 2746 11676 2774 11784
rect 5813 11781 5825 11815
rect 5859 11812 5871 11815
rect 7466 11812 7472 11824
rect 5859 11784 7472 11812
rect 5859 11781 5871 11784
rect 5813 11775 5871 11781
rect 7466 11772 7472 11784
rect 7524 11812 7530 11824
rect 7926 11812 7932 11824
rect 7524 11784 7932 11812
rect 7524 11772 7530 11784
rect 7926 11772 7932 11784
rect 7984 11812 7990 11824
rect 12345 11815 12403 11821
rect 7984 11784 8432 11812
rect 7984 11772 7990 11784
rect 5074 11704 5080 11756
rect 5132 11704 5138 11756
rect 6270 11704 6276 11756
rect 6328 11744 6334 11756
rect 6454 11744 6460 11756
rect 6328 11716 6460 11744
rect 6328 11704 6334 11716
rect 6454 11704 6460 11716
rect 6512 11744 6518 11756
rect 6917 11747 6975 11753
rect 6917 11744 6929 11747
rect 6512 11716 6929 11744
rect 6512 11704 6518 11716
rect 6917 11713 6929 11716
rect 6963 11713 6975 11747
rect 8202 11744 8208 11756
rect 6917 11707 6975 11713
rect 7576 11716 8208 11744
rect 7576 11685 7604 11716
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 6733 11679 6791 11685
rect 6733 11676 6745 11679
rect 2746 11648 6745 11676
rect 6733 11645 6745 11648
rect 6779 11645 6791 11679
rect 6733 11639 6791 11645
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 7561 11679 7619 11685
rect 6871 11648 7512 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 3970 11568 3976 11620
rect 4028 11608 4034 11620
rect 4801 11611 4859 11617
rect 4801 11608 4813 11611
rect 4028 11580 4813 11608
rect 4028 11568 4034 11580
rect 4801 11577 4813 11580
rect 4847 11577 4859 11611
rect 4801 11571 4859 11577
rect 4893 11611 4951 11617
rect 4893 11577 4905 11611
rect 4939 11608 4951 11611
rect 4982 11608 4988 11620
rect 4939 11580 4988 11608
rect 4939 11577 4951 11580
rect 4893 11571 4951 11577
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 4522 11540 4528 11552
rect 2372 11512 4528 11540
rect 2372 11500 2378 11512
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 4816 11540 4844 11571
rect 4982 11568 4988 11580
rect 5040 11568 5046 11620
rect 5166 11568 5172 11620
rect 5224 11608 5230 11620
rect 5261 11611 5319 11617
rect 5261 11608 5273 11611
rect 5224 11580 5273 11608
rect 5224 11568 5230 11580
rect 5261 11577 5273 11580
rect 5307 11577 5319 11611
rect 7484 11608 7512 11648
rect 7561 11645 7573 11679
rect 7607 11645 7619 11679
rect 7561 11639 7619 11645
rect 7837 11679 7895 11685
rect 7837 11645 7849 11679
rect 7883 11676 7895 11679
rect 8110 11676 8116 11688
rect 7883 11648 8116 11676
rect 7883 11645 7895 11648
rect 7837 11639 7895 11645
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 8404 11685 8432 11784
rect 12345 11781 12357 11815
rect 12391 11812 12403 11815
rect 12618 11812 12624 11824
rect 12391 11784 12624 11812
rect 12391 11781 12403 11784
rect 12345 11775 12403 11781
rect 12618 11772 12624 11784
rect 12676 11772 12682 11824
rect 14090 11772 14096 11824
rect 14148 11812 14154 11824
rect 14734 11812 14740 11824
rect 14148 11784 14740 11812
rect 14148 11772 14154 11784
rect 14734 11772 14740 11784
rect 14792 11772 14798 11824
rect 22738 11772 22744 11824
rect 22796 11812 22802 11824
rect 23569 11815 23627 11821
rect 23569 11812 23581 11815
rect 22796 11784 23581 11812
rect 22796 11772 22802 11784
rect 23569 11781 23581 11784
rect 23615 11781 23627 11815
rect 25590 11812 25596 11824
rect 25551 11784 25596 11812
rect 23569 11775 23627 11781
rect 25590 11772 25596 11784
rect 25648 11772 25654 11824
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 10137 11747 10195 11753
rect 10137 11744 10149 11747
rect 9732 11716 10149 11744
rect 9732 11704 9738 11716
rect 10137 11713 10149 11716
rect 10183 11713 10195 11747
rect 11238 11744 11244 11756
rect 11199 11716 11244 11744
rect 10137 11707 10195 11713
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 11425 11747 11483 11753
rect 11425 11713 11437 11747
rect 11471 11744 11483 11747
rect 11790 11744 11796 11756
rect 11471 11716 11796 11744
rect 11471 11713 11483 11716
rect 11425 11707 11483 11713
rect 11790 11704 11796 11716
rect 11848 11704 11854 11756
rect 13906 11744 13912 11756
rect 12452 11716 13912 11744
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11645 8447 11679
rect 8389 11639 8447 11645
rect 8478 11636 8484 11688
rect 8536 11636 8542 11688
rect 9950 11676 9956 11688
rect 9911 11648 9956 11676
rect 9950 11636 9956 11648
rect 10008 11636 10014 11688
rect 11514 11636 11520 11688
rect 11572 11676 11578 11688
rect 11974 11676 11980 11688
rect 11572 11648 11980 11676
rect 11572 11636 11578 11648
rect 11974 11636 11980 11648
rect 12032 11676 12038 11688
rect 12452 11685 12480 11716
rect 13906 11704 13912 11716
rect 13964 11704 13970 11756
rect 21450 11744 21456 11756
rect 21411 11716 21456 11744
rect 21450 11704 21456 11716
rect 21508 11704 21514 11756
rect 23290 11744 23296 11756
rect 23251 11716 23296 11744
rect 23290 11704 23296 11716
rect 23348 11704 23354 11756
rect 26142 11704 26148 11756
rect 26200 11744 26206 11756
rect 26329 11747 26387 11753
rect 26329 11744 26341 11747
rect 26200 11716 26341 11744
rect 26200 11704 26206 11716
rect 26329 11713 26341 11716
rect 26375 11713 26387 11747
rect 26329 11707 26387 11713
rect 27798 11704 27804 11756
rect 27856 11744 27862 11756
rect 28258 11744 28264 11756
rect 27856 11716 28264 11744
rect 27856 11704 27862 11716
rect 28258 11704 28264 11716
rect 28316 11704 28322 11756
rect 12253 11679 12311 11685
rect 12253 11676 12265 11679
rect 12032 11648 12265 11676
rect 12032 11636 12038 11648
rect 12253 11645 12265 11648
rect 12299 11645 12311 11679
rect 12253 11639 12311 11645
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11645 12495 11679
rect 12894 11676 12900 11688
rect 12855 11648 12900 11676
rect 12437 11639 12495 11645
rect 12894 11636 12900 11648
rect 12952 11636 12958 11688
rect 13262 11636 13268 11688
rect 13320 11676 13326 11688
rect 13725 11679 13783 11685
rect 13725 11676 13737 11679
rect 13320 11648 13737 11676
rect 13320 11636 13326 11648
rect 13725 11645 13737 11648
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11676 14243 11679
rect 14921 11679 14979 11685
rect 14921 11676 14933 11679
rect 14231 11648 14933 11676
rect 14231 11645 14243 11648
rect 14185 11639 14243 11645
rect 14921 11645 14933 11648
rect 14967 11645 14979 11679
rect 20714 11676 20720 11688
rect 20675 11648 20720 11676
rect 14921 11639 14979 11645
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 20990 11676 20996 11688
rect 20951 11648 20996 11676
rect 20990 11636 20996 11648
rect 21048 11636 21054 11688
rect 21358 11636 21364 11688
rect 21416 11676 21422 11688
rect 21709 11679 21767 11685
rect 21709 11676 21721 11679
rect 21416 11648 21721 11676
rect 21416 11636 21422 11648
rect 21709 11645 21721 11648
rect 21755 11645 21767 11679
rect 21709 11639 21767 11645
rect 22554 11636 22560 11688
rect 22612 11676 22618 11688
rect 25406 11676 25412 11688
rect 22612 11648 23060 11676
rect 25367 11648 25412 11676
rect 22612 11636 22618 11648
rect 7650 11608 7656 11620
rect 5261 11571 5319 11577
rect 5368 11580 7052 11608
rect 7484 11580 7656 11608
rect 5368 11540 5396 11580
rect 5626 11540 5632 11552
rect 4816 11512 5396 11540
rect 5587 11512 5632 11540
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 7024 11540 7052 11580
rect 7650 11568 7656 11580
rect 7708 11568 7714 11620
rect 7745 11611 7803 11617
rect 7745 11577 7757 11611
rect 7791 11608 7803 11611
rect 8496 11608 8524 11636
rect 7791 11580 8524 11608
rect 10045 11611 10103 11617
rect 7791 11577 7803 11580
rect 7745 11571 7803 11577
rect 10045 11577 10057 11611
rect 10091 11608 10103 11611
rect 10686 11608 10692 11620
rect 10091 11580 10692 11608
rect 10091 11577 10103 11580
rect 10045 11571 10103 11577
rect 10686 11568 10692 11580
rect 10744 11608 10750 11620
rect 11149 11611 11207 11617
rect 11149 11608 11161 11611
rect 10744 11580 11161 11608
rect 10744 11568 10750 11580
rect 11149 11577 11161 11580
rect 11195 11577 11207 11611
rect 11149 11571 11207 11577
rect 11330 11568 11336 11620
rect 11388 11608 11394 11620
rect 23032 11608 23060 11648
rect 25406 11636 25412 11648
rect 25464 11636 25470 11688
rect 25958 11636 25964 11688
rect 26016 11676 26022 11688
rect 26789 11679 26847 11685
rect 26789 11676 26801 11679
rect 26016 11648 26801 11676
rect 26016 11636 26022 11648
rect 26789 11645 26801 11648
rect 26835 11645 26847 11679
rect 26789 11639 26847 11645
rect 27056 11679 27114 11685
rect 27056 11645 27068 11679
rect 27102 11676 27114 11679
rect 27430 11676 27436 11688
rect 27102 11648 27436 11676
rect 27102 11645 27114 11648
rect 27056 11639 27114 11645
rect 27430 11636 27436 11648
rect 27488 11636 27494 11688
rect 26145 11611 26203 11617
rect 26145 11608 26157 11611
rect 11388 11580 21036 11608
rect 11388 11568 11394 11580
rect 8297 11543 8355 11549
rect 8297 11540 8309 11543
rect 7024 11512 8309 11540
rect 8297 11509 8309 11512
rect 8343 11509 8355 11543
rect 8478 11540 8484 11552
rect 8439 11512 8484 11540
rect 8297 11503 8355 11509
rect 8478 11500 8484 11512
rect 8536 11500 8542 11552
rect 9306 11500 9312 11552
rect 9364 11540 9370 11552
rect 9490 11540 9496 11552
rect 9364 11512 9496 11540
rect 9364 11500 9370 11512
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 13446 11500 13452 11552
rect 13504 11540 13510 11552
rect 13541 11543 13599 11549
rect 13541 11540 13553 11543
rect 13504 11512 13553 11540
rect 13504 11500 13510 11512
rect 13541 11509 13553 11512
rect 13587 11540 13599 11543
rect 14185 11543 14243 11549
rect 14185 11540 14197 11543
rect 13587 11512 14197 11540
rect 13587 11509 13599 11512
rect 13541 11503 13599 11509
rect 14185 11509 14197 11512
rect 14231 11509 14243 11543
rect 14185 11503 14243 11509
rect 14734 11500 14740 11552
rect 14792 11540 14798 11552
rect 19242 11540 19248 11552
rect 14792 11512 19248 11540
rect 14792 11500 14798 11512
rect 19242 11500 19248 11512
rect 19300 11540 19306 11552
rect 20622 11540 20628 11552
rect 19300 11512 20628 11540
rect 19300 11500 19306 11512
rect 20622 11500 20628 11512
rect 20680 11500 20686 11552
rect 20898 11540 20904 11552
rect 20859 11512 20904 11540
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 21008 11540 21036 11580
rect 22066 11580 22968 11608
rect 23032 11580 26157 11608
rect 22066 11540 22094 11580
rect 21008 11512 22094 11540
rect 22738 11500 22744 11552
rect 22796 11540 22802 11552
rect 22833 11543 22891 11549
rect 22833 11540 22845 11543
rect 22796 11512 22845 11540
rect 22796 11500 22802 11512
rect 22833 11509 22845 11512
rect 22879 11509 22891 11543
rect 22940 11540 22968 11580
rect 26145 11577 26157 11580
rect 26191 11577 26203 11611
rect 26145 11571 26203 11577
rect 26510 11540 26516 11552
rect 22940 11512 26516 11540
rect 22833 11503 22891 11509
rect 26510 11500 26516 11512
rect 26568 11500 26574 11552
rect 1104 11450 28888 11472
rect 1104 11398 10246 11450
rect 10298 11398 10310 11450
rect 10362 11398 10374 11450
rect 10426 11398 10438 11450
rect 10490 11398 19510 11450
rect 19562 11398 19574 11450
rect 19626 11398 19638 11450
rect 19690 11398 19702 11450
rect 19754 11398 28888 11450
rect 1104 11376 28888 11398
rect 1765 11339 1823 11345
rect 1765 11305 1777 11339
rect 1811 11305 1823 11339
rect 1765 11299 1823 11305
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11336 2467 11339
rect 2455 11308 7604 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 1780 11268 1808 11299
rect 5626 11268 5632 11280
rect 1780 11240 5632 11268
rect 5626 11228 5632 11240
rect 5684 11228 5690 11280
rect 7576 11268 7604 11308
rect 8220 11308 8432 11336
rect 8220 11268 8248 11308
rect 7576 11240 8248 11268
rect 8404 11268 8432 11308
rect 8478 11296 8484 11348
rect 8536 11336 8542 11348
rect 9306 11336 9312 11348
rect 8536 11308 9312 11336
rect 8536 11296 8542 11308
rect 9306 11296 9312 11308
rect 9364 11336 9370 11348
rect 9953 11339 10011 11345
rect 9953 11336 9965 11339
rect 9364 11308 9965 11336
rect 9364 11296 9370 11308
rect 9953 11305 9965 11308
rect 9999 11305 10011 11339
rect 9953 11299 10011 11305
rect 10686 11296 10692 11348
rect 10744 11336 10750 11348
rect 10781 11339 10839 11345
rect 10781 11336 10793 11339
rect 10744 11308 10793 11336
rect 10744 11296 10750 11308
rect 10781 11305 10793 11308
rect 10827 11305 10839 11339
rect 10781 11299 10839 11305
rect 12069 11339 12127 11345
rect 12069 11305 12081 11339
rect 12115 11336 12127 11339
rect 12894 11336 12900 11348
rect 12115 11308 12900 11336
rect 12115 11305 12127 11308
rect 12069 11299 12127 11305
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13630 11336 13636 11348
rect 13044 11308 13636 11336
rect 13044 11296 13050 11308
rect 13630 11296 13636 11308
rect 13688 11336 13694 11348
rect 18874 11336 18880 11348
rect 13688 11308 13860 11336
rect 13688 11296 13694 11308
rect 12437 11271 12495 11277
rect 12437 11268 12449 11271
rect 8404 11240 12449 11268
rect 12437 11237 12449 11240
rect 12483 11237 12495 11271
rect 12437 11231 12495 11237
rect 12529 11271 12587 11277
rect 12529 11237 12541 11271
rect 12575 11268 12587 11271
rect 13722 11268 13728 11280
rect 12575 11240 13728 11268
rect 12575 11237 12587 11240
rect 12529 11231 12587 11237
rect 13722 11228 13728 11240
rect 13780 11228 13786 11280
rect 13832 11277 13860 11308
rect 18524 11308 18880 11336
rect 13817 11271 13875 11277
rect 13817 11237 13829 11271
rect 13863 11237 13875 11271
rect 13817 11231 13875 11237
rect 1946 11200 1952 11212
rect 1907 11172 1952 11200
rect 1946 11160 1952 11172
rect 2004 11160 2010 11212
rect 2593 11203 2651 11209
rect 2593 11169 2605 11203
rect 2639 11200 2651 11203
rect 2774 11200 2780 11212
rect 2639 11172 2780 11200
rect 2639 11169 2651 11172
rect 2593 11163 2651 11169
rect 2774 11160 2780 11172
rect 2832 11160 2838 11212
rect 3234 11200 3240 11212
rect 3195 11172 3240 11200
rect 3234 11160 3240 11172
rect 3292 11160 3298 11212
rect 3421 11203 3479 11209
rect 3421 11169 3433 11203
rect 3467 11169 3479 11203
rect 3421 11163 3479 11169
rect 3142 11092 3148 11144
rect 3200 11132 3206 11144
rect 3436 11132 3464 11163
rect 3510 11160 3516 11212
rect 3568 11200 3574 11212
rect 3970 11200 3976 11212
rect 3568 11172 3613 11200
rect 3931 11172 3976 11200
rect 3568 11160 3574 11172
rect 3970 11160 3976 11172
rect 4028 11160 4034 11212
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 5350 11200 5356 11212
rect 5123 11172 5356 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 3200 11104 4077 11132
rect 3200 11092 3206 11104
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 5000 11132 5028 11163
rect 5350 11160 5356 11172
rect 5408 11160 5414 11212
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 7524 11172 7573 11200
rect 7524 11160 7530 11172
rect 7561 11169 7573 11172
rect 7607 11169 7619 11203
rect 8202 11200 8208 11212
rect 8163 11172 8208 11200
rect 7561 11163 7619 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 9858 11200 9864 11212
rect 9819 11172 9864 11200
rect 9858 11160 9864 11172
rect 9916 11160 9922 11212
rect 10689 11203 10747 11209
rect 10689 11200 10701 11203
rect 10612 11172 10701 11200
rect 5258 11132 5264 11144
rect 5000 11104 5264 11132
rect 4065 11095 4123 11101
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 10042 11132 10048 11144
rect 10003 11104 10048 11132
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 3050 11064 3056 11076
rect 3011 11036 3056 11064
rect 3050 11024 3056 11036
rect 3108 11024 3114 11076
rect 5074 11024 5080 11076
rect 5132 11064 5138 11076
rect 5994 11064 6000 11076
rect 5132 11036 6000 11064
rect 5132 11024 5138 11036
rect 5994 11024 6000 11036
rect 6052 11024 6058 11076
rect 8389 11067 8447 11073
rect 8389 11064 8401 11067
rect 7300 11036 8401 11064
rect 7300 11008 7328 11036
rect 8389 11033 8401 11036
rect 8435 11033 8447 11067
rect 10612 11064 10640 11172
rect 10689 11169 10701 11172
rect 10735 11200 10747 11203
rect 13633 11203 13691 11209
rect 10735 11172 13584 11200
rect 10735 11169 10747 11172
rect 10689 11163 10747 11169
rect 11790 11092 11796 11144
rect 11848 11132 11854 11144
rect 12621 11135 12679 11141
rect 12621 11132 12633 11135
rect 11848 11104 12633 11132
rect 11848 11092 11854 11104
rect 12621 11101 12633 11104
rect 12667 11101 12679 11135
rect 13556 11132 13584 11172
rect 13633 11169 13645 11203
rect 13679 11200 13691 11203
rect 13906 11200 13912 11212
rect 13679 11172 13912 11200
rect 13679 11169 13691 11172
rect 13633 11163 13691 11169
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 18046 11200 18052 11212
rect 18007 11172 18052 11200
rect 18046 11160 18052 11172
rect 18104 11160 18110 11212
rect 14734 11132 14740 11144
rect 13556 11104 14740 11132
rect 12621 11095 12679 11101
rect 14734 11092 14740 11104
rect 14792 11092 14798 11144
rect 18141 11135 18199 11141
rect 18141 11101 18153 11135
rect 18187 11101 18199 11135
rect 18141 11095 18199 11101
rect 18325 11135 18383 11141
rect 18325 11101 18337 11135
rect 18371 11132 18383 11135
rect 18524 11132 18552 11308
rect 18874 11296 18880 11308
rect 18932 11336 18938 11348
rect 19705 11339 19763 11345
rect 19705 11336 19717 11339
rect 18932 11308 19717 11336
rect 18932 11296 18938 11308
rect 19705 11305 19717 11308
rect 19751 11305 19763 11339
rect 19705 11299 19763 11305
rect 20162 11296 20168 11348
rect 20220 11336 20226 11348
rect 20257 11339 20315 11345
rect 20257 11336 20269 11339
rect 20220 11308 20269 11336
rect 20220 11296 20226 11308
rect 20257 11305 20269 11308
rect 20303 11305 20315 11339
rect 20257 11299 20315 11305
rect 24854 11296 24860 11348
rect 24912 11336 24918 11348
rect 24912 11308 28028 11336
rect 24912 11296 24918 11308
rect 19794 11268 19800 11280
rect 18371 11104 18552 11132
rect 18616 11240 19800 11268
rect 18616 11132 18644 11240
rect 19794 11228 19800 11240
rect 19852 11228 19858 11280
rect 20622 11228 20628 11280
rect 20680 11268 20686 11280
rect 28000 11277 28028 11308
rect 26697 11271 26755 11277
rect 26697 11268 26709 11271
rect 20680 11240 26709 11268
rect 20680 11228 20686 11240
rect 26697 11237 26709 11240
rect 26743 11237 26755 11271
rect 26697 11231 26755 11237
rect 27985 11271 28043 11277
rect 27985 11237 27997 11271
rect 28031 11237 28043 11271
rect 27985 11231 28043 11237
rect 18690 11160 18696 11212
rect 18748 11200 18754 11212
rect 18877 11203 18935 11209
rect 18877 11200 18889 11203
rect 18748 11172 18889 11200
rect 18748 11160 18754 11172
rect 18877 11169 18889 11172
rect 18923 11200 18935 11203
rect 19613 11203 19671 11209
rect 19613 11200 19625 11203
rect 18923 11172 19625 11200
rect 18923 11169 18935 11172
rect 18877 11163 18935 11169
rect 19613 11169 19625 11172
rect 19659 11169 19671 11203
rect 19613 11163 19671 11169
rect 20441 11203 20499 11209
rect 20441 11169 20453 11203
rect 20487 11200 20499 11203
rect 21266 11200 21272 11212
rect 20487 11172 21272 11200
rect 20487 11169 20499 11172
rect 20441 11163 20499 11169
rect 21266 11160 21272 11172
rect 21324 11160 21330 11212
rect 24213 11203 24271 11209
rect 24213 11169 24225 11203
rect 24259 11200 24271 11203
rect 25041 11203 25099 11209
rect 25041 11200 25053 11203
rect 24259 11172 25053 11200
rect 24259 11169 24271 11172
rect 24213 11163 24271 11169
rect 25041 11169 25053 11172
rect 25087 11169 25099 11203
rect 25041 11163 25099 11169
rect 25682 11160 25688 11212
rect 25740 11200 25746 11212
rect 25961 11203 26019 11209
rect 25961 11200 25973 11203
rect 25740 11172 25973 11200
rect 25740 11160 25746 11172
rect 25961 11169 25973 11172
rect 26007 11169 26019 11203
rect 26142 11200 26148 11212
rect 26103 11172 26148 11200
rect 25961 11163 26019 11169
rect 26142 11160 26148 11172
rect 26200 11160 26206 11212
rect 18969 11135 19027 11141
rect 18969 11132 18981 11135
rect 18616 11104 18981 11132
rect 18371 11101 18383 11104
rect 18325 11095 18383 11101
rect 18969 11101 18981 11104
rect 19015 11101 19027 11135
rect 19150 11132 19156 11144
rect 19111 11104 19156 11132
rect 18969 11095 19027 11101
rect 8389 11027 8447 11033
rect 8496 11036 10640 11064
rect 13648 11036 13860 11064
rect 7282 10956 7288 11008
rect 7340 10956 7346 11008
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 8496 10996 8524 11036
rect 7708 10968 8524 10996
rect 9493 10999 9551 11005
rect 7708 10956 7714 10968
rect 9493 10965 9505 10999
rect 9539 10996 9551 10999
rect 9582 10996 9588 11008
rect 9539 10968 9588 10996
rect 9539 10965 9551 10968
rect 9493 10959 9551 10965
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 9766 10956 9772 11008
rect 9824 10996 9830 11008
rect 13648 10996 13676 11036
rect 9824 10968 13676 10996
rect 13832 10996 13860 11036
rect 17586 11024 17592 11076
rect 17644 11064 17650 11076
rect 17681 11067 17739 11073
rect 17681 11064 17693 11067
rect 17644 11036 17693 11064
rect 17644 11024 17650 11036
rect 17681 11033 17693 11036
rect 17727 11033 17739 11067
rect 18156 11064 18184 11095
rect 19150 11092 19156 11104
rect 19208 11092 19214 11144
rect 19886 11092 19892 11144
rect 19944 11132 19950 11144
rect 20162 11132 20168 11144
rect 19944 11104 20168 11132
rect 19944 11092 19950 11104
rect 20162 11092 20168 11104
rect 20220 11092 20226 11144
rect 23566 11132 23572 11144
rect 23527 11104 23572 11132
rect 23566 11092 23572 11104
rect 23624 11092 23630 11144
rect 23842 11092 23848 11144
rect 23900 11132 23906 11144
rect 23937 11135 23995 11141
rect 23937 11132 23949 11135
rect 23900 11104 23949 11132
rect 23900 11092 23906 11104
rect 23937 11101 23949 11104
rect 23983 11101 23995 11135
rect 23937 11095 23995 11101
rect 24026 11092 24032 11144
rect 24084 11132 24090 11144
rect 24084 11104 24129 11132
rect 24084 11092 24090 11104
rect 24762 11092 24768 11144
rect 24820 11132 24826 11144
rect 24857 11135 24915 11141
rect 24857 11132 24869 11135
rect 24820 11104 24869 11132
rect 24820 11092 24826 11104
rect 24857 11101 24869 11104
rect 24903 11101 24915 11135
rect 24857 11095 24915 11101
rect 24949 11135 25007 11141
rect 24949 11101 24961 11135
rect 24995 11101 25007 11135
rect 24949 11095 25007 11101
rect 18690 11064 18696 11076
rect 18156 11036 18696 11064
rect 17681 11027 17739 11033
rect 18690 11024 18696 11036
rect 18748 11024 18754 11076
rect 19058 11064 19064 11076
rect 19019 11036 19064 11064
rect 19058 11024 19064 11036
rect 19116 11024 19122 11076
rect 24964 11064 24992 11095
rect 25130 11092 25136 11144
rect 25188 11132 25194 11144
rect 25188 11104 25233 11132
rect 25188 11092 25194 11104
rect 25314 11064 25320 11076
rect 19628 11036 20392 11064
rect 24964 11036 25320 11064
rect 19628 10996 19656 11036
rect 13832 10968 19656 10996
rect 20364 10996 20392 11036
rect 25314 11024 25320 11036
rect 25372 11024 25378 11076
rect 26878 11064 26884 11076
rect 26839 11036 26884 11064
rect 26878 11024 26884 11036
rect 26936 11024 26942 11076
rect 27522 11024 27528 11076
rect 27580 11064 27586 11076
rect 28169 11067 28227 11073
rect 28169 11064 28181 11067
rect 27580 11036 28181 11064
rect 27580 11024 27586 11036
rect 28169 11033 28181 11036
rect 28215 11033 28227 11067
rect 28994 11064 29000 11076
rect 28955 11036 29000 11064
rect 28169 11027 28227 11033
rect 28994 11024 29000 11036
rect 29052 11024 29058 11076
rect 22554 10996 22560 11008
rect 20364 10968 22560 10996
rect 9824 10956 9830 10968
rect 22554 10956 22560 10968
rect 22612 10956 22618 11008
rect 24670 10996 24676 11008
rect 24631 10968 24676 10996
rect 24670 10956 24676 10968
rect 24728 10956 24734 11008
rect 1104 10906 28888 10928
rect 1104 10854 5614 10906
rect 5666 10854 5678 10906
rect 5730 10854 5742 10906
rect 5794 10854 5806 10906
rect 5858 10854 14878 10906
rect 14930 10854 14942 10906
rect 14994 10854 15006 10906
rect 15058 10854 15070 10906
rect 15122 10854 24142 10906
rect 24194 10854 24206 10906
rect 24258 10854 24270 10906
rect 24322 10854 24334 10906
rect 24386 10854 28888 10906
rect 1104 10832 28888 10854
rect 2041 10795 2099 10801
rect 2041 10761 2053 10795
rect 2087 10792 2099 10795
rect 2222 10792 2228 10804
rect 2087 10764 2228 10792
rect 2087 10761 2099 10764
rect 2041 10755 2099 10761
rect 2222 10752 2228 10764
rect 2280 10752 2286 10804
rect 2958 10752 2964 10804
rect 3016 10792 3022 10804
rect 3053 10795 3111 10801
rect 3053 10792 3065 10795
rect 3016 10764 3065 10792
rect 3016 10752 3022 10764
rect 3053 10761 3065 10764
rect 3099 10792 3111 10795
rect 3970 10792 3976 10804
rect 3099 10764 3976 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 9766 10792 9772 10804
rect 5276 10764 9772 10792
rect 2866 10724 2872 10736
rect 2827 10696 2872 10724
rect 2866 10684 2872 10696
rect 2924 10684 2930 10736
rect 2130 10616 2136 10668
rect 2188 10656 2194 10668
rect 2593 10659 2651 10665
rect 2593 10656 2605 10659
rect 2188 10628 2605 10656
rect 2188 10616 2194 10628
rect 2593 10625 2605 10628
rect 2639 10625 2651 10659
rect 2593 10619 2651 10625
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 5276 10665 5304 10764
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 10873 10795 10931 10801
rect 10873 10792 10885 10795
rect 9916 10764 10885 10792
rect 9916 10752 9922 10764
rect 10873 10761 10885 10764
rect 10919 10761 10931 10795
rect 13446 10792 13452 10804
rect 10873 10755 10931 10761
rect 12406 10764 13452 10792
rect 5261 10659 5319 10665
rect 5261 10656 5273 10659
rect 4396 10628 5273 10656
rect 4396 10616 4402 10628
rect 5261 10625 5273 10628
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 5445 10659 5503 10665
rect 5445 10625 5457 10659
rect 5491 10656 5503 10659
rect 6270 10656 6276 10668
rect 5491 10628 6276 10656
rect 5491 10625 5503 10628
rect 5445 10619 5503 10625
rect 6270 10616 6276 10628
rect 6328 10616 6334 10668
rect 9416 10628 9628 10656
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10588 2007 10591
rect 2866 10588 2872 10600
rect 1995 10560 2872 10588
rect 1995 10557 2007 10560
rect 1949 10551 2007 10557
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 4706 10548 4712 10600
rect 4764 10588 4770 10600
rect 9416 10588 9444 10628
rect 4764 10560 9444 10588
rect 9493 10591 9551 10597
rect 4764 10548 4770 10560
rect 9493 10557 9505 10591
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 5169 10523 5227 10529
rect 5169 10489 5181 10523
rect 5215 10520 5227 10523
rect 5350 10520 5356 10532
rect 5215 10492 5356 10520
rect 5215 10489 5227 10492
rect 5169 10483 5227 10489
rect 5350 10480 5356 10492
rect 5408 10480 5414 10532
rect 8294 10480 8300 10532
rect 8352 10520 8358 10532
rect 9508 10520 9536 10551
rect 8352 10492 9536 10520
rect 9600 10520 9628 10628
rect 9766 10597 9772 10600
rect 9760 10588 9772 10597
rect 9727 10560 9772 10588
rect 9760 10551 9772 10560
rect 9766 10548 9772 10551
rect 9824 10548 9830 10600
rect 11517 10591 11575 10597
rect 11517 10557 11529 10591
rect 11563 10588 11575 10591
rect 12406 10588 12434 10764
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 16393 10795 16451 10801
rect 16393 10761 16405 10795
rect 16439 10792 16451 10795
rect 17034 10792 17040 10804
rect 16439 10764 17040 10792
rect 16439 10761 16451 10764
rect 16393 10755 16451 10761
rect 17034 10752 17040 10764
rect 17092 10752 17098 10804
rect 18966 10752 18972 10804
rect 19024 10792 19030 10804
rect 19150 10792 19156 10804
rect 19024 10764 19156 10792
rect 19024 10752 19030 10764
rect 19150 10752 19156 10764
rect 19208 10752 19214 10804
rect 24026 10752 24032 10804
rect 24084 10752 24090 10804
rect 24213 10795 24271 10801
rect 24213 10761 24225 10795
rect 24259 10792 24271 10795
rect 24486 10792 24492 10804
rect 24259 10764 24492 10792
rect 24259 10761 24271 10764
rect 24213 10755 24271 10761
rect 24486 10752 24492 10764
rect 24544 10752 24550 10804
rect 25130 10752 25136 10804
rect 25188 10792 25194 10804
rect 25685 10795 25743 10801
rect 25685 10792 25697 10795
rect 25188 10764 25697 10792
rect 25188 10752 25194 10764
rect 25685 10761 25697 10764
rect 25731 10761 25743 10795
rect 25685 10755 25743 10761
rect 12986 10684 12992 10736
rect 13044 10684 13050 10736
rect 18417 10727 18475 10733
rect 18417 10724 18429 10727
rect 18248 10696 18429 10724
rect 13004 10656 13032 10684
rect 12912 10628 13032 10656
rect 11563 10560 12434 10588
rect 11563 10557 11575 10560
rect 11517 10551 11575 10557
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 12912 10597 12940 10628
rect 16114 10616 16120 10668
rect 16172 10656 16178 10668
rect 16172 10628 16974 10656
rect 16172 10616 16178 10628
rect 12759 10591 12817 10597
rect 12759 10588 12771 10591
rect 12676 10560 12771 10588
rect 12676 10548 12682 10560
rect 12759 10557 12771 10560
rect 12805 10557 12817 10591
rect 12759 10551 12817 10557
rect 12878 10591 12940 10597
rect 12878 10557 12890 10591
rect 12924 10560 12940 10591
rect 12924 10557 12936 10560
rect 12878 10551 12936 10557
rect 12986 10548 12992 10600
rect 13044 10588 13050 10600
rect 13185 10591 13243 10597
rect 13044 10560 13089 10588
rect 13044 10548 13050 10560
rect 13185 10557 13197 10591
rect 13231 10588 13243 10591
rect 13446 10588 13452 10600
rect 13231 10560 13452 10588
rect 13231 10557 13243 10560
rect 13185 10551 13243 10557
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 15473 10591 15531 10597
rect 15473 10557 15485 10591
rect 15519 10588 15531 10591
rect 15562 10588 15568 10600
rect 15519 10560 15568 10588
rect 15519 10557 15531 10560
rect 15473 10551 15531 10557
rect 15562 10548 15568 10560
rect 15620 10588 15626 10600
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 15620 10560 17509 10588
rect 15620 10548 15626 10560
rect 17497 10557 17509 10560
rect 17543 10557 17555 10591
rect 17497 10551 17555 10557
rect 17678 10548 17684 10600
rect 17736 10588 17742 10600
rect 18248 10588 18276 10696
rect 18417 10693 18429 10696
rect 18463 10693 18475 10727
rect 18417 10687 18475 10693
rect 22741 10727 22799 10733
rect 22741 10693 22753 10727
rect 22787 10693 22799 10727
rect 22741 10687 22799 10693
rect 22094 10616 22100 10668
rect 22152 10616 22158 10668
rect 22756 10656 22784 10687
rect 23566 10656 23572 10668
rect 22756 10628 23572 10656
rect 23566 10616 23572 10628
rect 23624 10616 23630 10668
rect 23934 10656 23940 10668
rect 23895 10628 23940 10656
rect 23934 10616 23940 10628
rect 23992 10616 23998 10668
rect 17736 10560 18276 10588
rect 17736 10548 17742 10560
rect 18414 10548 18420 10600
rect 18472 10588 18478 10600
rect 21729 10591 21787 10597
rect 21729 10588 21741 10591
rect 18472 10560 21741 10588
rect 18472 10548 18478 10560
rect 21729 10557 21741 10560
rect 21775 10557 21787 10591
rect 22278 10588 22284 10600
rect 21729 10551 21787 10557
rect 22112 10560 22284 10588
rect 12066 10520 12072 10532
rect 9600 10492 12072 10520
rect 8352 10480 8358 10492
rect 4798 10452 4804 10464
rect 4759 10424 4804 10452
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 9416 10452 9444 10492
rect 12066 10480 12072 10492
rect 12124 10480 12130 10532
rect 15194 10480 15200 10532
rect 15252 10520 15258 10532
rect 15930 10529 15936 10532
rect 15381 10523 15439 10529
rect 15381 10520 15393 10523
rect 15252 10492 15393 10520
rect 15252 10480 15258 10492
rect 15381 10489 15393 10492
rect 15427 10489 15439 10523
rect 15381 10483 15439 10489
rect 15887 10523 15936 10529
rect 15887 10489 15899 10523
rect 15933 10489 15936 10523
rect 15887 10483 15936 10489
rect 15930 10480 15936 10483
rect 15988 10480 15994 10532
rect 17126 10520 17132 10532
rect 17087 10492 17132 10520
rect 17126 10480 17132 10492
rect 17184 10480 17190 10532
rect 17405 10523 17463 10529
rect 17405 10489 17417 10523
rect 17451 10520 17463 10523
rect 17865 10523 17923 10529
rect 17451 10492 17724 10520
rect 17451 10489 17463 10492
rect 17405 10483 17463 10489
rect 17696 10464 17724 10492
rect 17865 10489 17877 10523
rect 17911 10520 17923 10523
rect 21174 10520 21180 10532
rect 17911 10492 21180 10520
rect 17911 10489 17923 10492
rect 17865 10483 17923 10489
rect 21174 10480 21180 10492
rect 21232 10520 21238 10532
rect 21542 10520 21548 10532
rect 21232 10492 21548 10520
rect 21232 10480 21238 10492
rect 21542 10480 21548 10492
rect 21600 10480 21606 10532
rect 21821 10523 21879 10529
rect 21821 10489 21833 10523
rect 21867 10520 21879 10523
rect 22112 10520 22140 10560
rect 22278 10548 22284 10560
rect 22336 10588 22342 10600
rect 22922 10588 22928 10600
rect 22336 10560 22928 10588
rect 22336 10548 22342 10560
rect 22922 10548 22928 10560
rect 22980 10548 22986 10600
rect 21867 10492 22140 10520
rect 22189 10523 22247 10529
rect 21867 10489 21879 10492
rect 21821 10483 21879 10489
rect 22189 10489 22201 10523
rect 22235 10520 22247 10523
rect 22646 10520 22652 10532
rect 22235 10492 22652 10520
rect 22235 10489 22247 10492
rect 22189 10483 22247 10489
rect 22646 10480 22652 10492
rect 22704 10480 22710 10532
rect 23934 10480 23940 10532
rect 23992 10520 23998 10532
rect 24044 10529 24072 10752
rect 25593 10727 25651 10733
rect 25593 10693 25605 10727
rect 25639 10724 25651 10727
rect 25866 10724 25872 10736
rect 25639 10696 25872 10724
rect 25639 10693 25651 10696
rect 25593 10687 25651 10693
rect 25866 10684 25872 10696
rect 25924 10684 25930 10736
rect 25225 10659 25283 10665
rect 25225 10625 25237 10659
rect 25271 10656 25283 10659
rect 25314 10656 25320 10668
rect 25271 10628 25320 10656
rect 25271 10625 25283 10628
rect 25225 10619 25283 10625
rect 25314 10616 25320 10628
rect 25372 10616 25378 10668
rect 25498 10616 25504 10668
rect 25556 10656 25562 10668
rect 25958 10656 25964 10668
rect 25556 10628 25964 10656
rect 25556 10616 25562 10628
rect 25958 10616 25964 10628
rect 26016 10656 26022 10668
rect 26789 10659 26847 10665
rect 26789 10656 26801 10659
rect 26016 10628 26801 10656
rect 26016 10616 26022 10628
rect 26789 10625 26801 10628
rect 26835 10625 26847 10659
rect 26789 10619 26847 10625
rect 25406 10548 25412 10600
rect 25464 10588 25470 10600
rect 26145 10591 26203 10597
rect 26145 10588 26157 10591
rect 25464 10560 26157 10588
rect 25464 10548 25470 10560
rect 26145 10557 26157 10560
rect 26191 10557 26203 10591
rect 26145 10551 26203 10557
rect 24044 10523 24112 10529
rect 24044 10520 24066 10523
rect 23992 10492 24066 10520
rect 23992 10480 23998 10492
rect 24054 10489 24066 10492
rect 24100 10489 24112 10523
rect 24054 10483 24112 10489
rect 27056 10523 27114 10529
rect 27056 10489 27068 10523
rect 27102 10520 27114 10523
rect 27982 10520 27988 10532
rect 27102 10492 27988 10520
rect 27102 10489 27114 10492
rect 27056 10483 27114 10489
rect 27982 10480 27988 10492
rect 28040 10480 28046 10532
rect 11333 10455 11391 10461
rect 11333 10452 11345 10455
rect 9416 10424 11345 10452
rect 11333 10421 11345 10424
rect 11379 10421 11391 10455
rect 12526 10452 12532 10464
rect 12487 10424 12532 10452
rect 11333 10415 11391 10421
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 15105 10455 15163 10461
rect 15105 10421 15117 10455
rect 15151 10452 15163 10455
rect 15562 10452 15568 10464
rect 15151 10424 15568 10452
rect 15151 10421 15163 10424
rect 15105 10415 15163 10421
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 16206 10452 16212 10464
rect 16167 10424 16212 10452
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 17678 10412 17684 10464
rect 17736 10412 17742 10464
rect 18230 10452 18236 10464
rect 18191 10424 18236 10452
rect 18230 10412 18236 10424
rect 18288 10412 18294 10464
rect 19794 10412 19800 10464
rect 19852 10452 19858 10464
rect 21453 10455 21511 10461
rect 21453 10452 21465 10455
rect 19852 10424 21465 10452
rect 19852 10412 19858 10424
rect 21453 10421 21465 10424
rect 21499 10452 21511 10455
rect 21910 10452 21916 10464
rect 21499 10424 21916 10452
rect 21499 10421 21511 10424
rect 21453 10415 21511 10421
rect 21910 10412 21916 10424
rect 21968 10412 21974 10464
rect 22554 10452 22560 10464
rect 22515 10424 22560 10452
rect 22554 10412 22560 10424
rect 22612 10412 22618 10464
rect 23842 10452 23848 10464
rect 23803 10424 23848 10452
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 26234 10412 26240 10464
rect 26292 10452 26298 10464
rect 28169 10455 28227 10461
rect 26292 10424 26337 10452
rect 26292 10412 26298 10424
rect 28169 10421 28181 10455
rect 28215 10452 28227 10455
rect 28258 10452 28264 10464
rect 28215 10424 28264 10452
rect 28215 10421 28227 10424
rect 28169 10415 28227 10421
rect 28258 10412 28264 10424
rect 28316 10412 28322 10464
rect 1104 10362 28888 10384
rect 1104 10310 10246 10362
rect 10298 10310 10310 10362
rect 10362 10310 10374 10362
rect 10426 10310 10438 10362
rect 10490 10310 19510 10362
rect 19562 10310 19574 10362
rect 19626 10310 19638 10362
rect 19690 10310 19702 10362
rect 19754 10310 28888 10362
rect 1104 10288 28888 10310
rect 1397 10251 1455 10257
rect 1397 10217 1409 10251
rect 1443 10248 1455 10251
rect 2682 10248 2688 10260
rect 1443 10220 2688 10248
rect 1443 10217 1455 10220
rect 1397 10211 1455 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 2961 10251 3019 10257
rect 2961 10248 2973 10251
rect 2832 10220 2973 10248
rect 2832 10208 2838 10220
rect 2961 10217 2973 10220
rect 3007 10248 3019 10251
rect 3694 10248 3700 10260
rect 3007 10220 3700 10248
rect 3007 10217 3019 10220
rect 2961 10211 3019 10217
rect 3694 10208 3700 10220
rect 3752 10208 3758 10260
rect 8113 10251 8171 10257
rect 8113 10248 8125 10251
rect 6932 10220 8125 10248
rect 2130 10180 2136 10192
rect 2056 10152 2136 10180
rect 1578 10112 1584 10124
rect 1539 10084 1584 10112
rect 1578 10072 1584 10084
rect 1636 10072 1642 10124
rect 2056 10121 2084 10152
rect 2130 10140 2136 10152
rect 2188 10140 2194 10192
rect 6932 10189 6960 10220
rect 8113 10217 8125 10220
rect 8159 10217 8171 10251
rect 9214 10248 9220 10260
rect 9175 10220 9220 10248
rect 8113 10211 8171 10217
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 15194 10248 15200 10260
rect 12124 10220 15200 10248
rect 12124 10208 12130 10220
rect 15194 10208 15200 10220
rect 15252 10208 15258 10260
rect 15562 10208 15568 10260
rect 15620 10248 15626 10260
rect 16022 10248 16028 10260
rect 15620 10220 16028 10248
rect 15620 10208 15626 10220
rect 16022 10208 16028 10220
rect 16080 10248 16086 10260
rect 16574 10248 16580 10260
rect 16080 10220 16580 10248
rect 16080 10208 16086 10220
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 17865 10251 17923 10257
rect 17865 10217 17877 10251
rect 17911 10248 17923 10251
rect 18046 10248 18052 10260
rect 17911 10220 18052 10248
rect 17911 10217 17923 10220
rect 17865 10211 17923 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 18138 10208 18144 10260
rect 18196 10248 18202 10260
rect 19705 10251 19763 10257
rect 19705 10248 19717 10251
rect 18196 10220 19717 10248
rect 18196 10208 18202 10220
rect 19705 10217 19717 10220
rect 19751 10217 19763 10251
rect 19705 10211 19763 10217
rect 25866 10208 25872 10260
rect 25924 10248 25930 10260
rect 26789 10251 26847 10257
rect 26789 10248 26801 10251
rect 25924 10220 26801 10248
rect 25924 10208 25930 10220
rect 26789 10217 26801 10220
rect 26835 10217 26847 10251
rect 28074 10248 28080 10260
rect 28035 10220 28080 10248
rect 26789 10211 26847 10217
rect 28074 10208 28080 10220
rect 28132 10208 28138 10260
rect 6917 10183 6975 10189
rect 6917 10149 6929 10183
rect 6963 10149 6975 10183
rect 7098 10180 7104 10192
rect 7011 10152 7104 10180
rect 6917 10143 6975 10149
rect 7098 10140 7104 10152
rect 7156 10180 7162 10192
rect 7653 10183 7711 10189
rect 7156 10152 7604 10180
rect 7156 10140 7162 10152
rect 2041 10115 2099 10121
rect 2041 10081 2053 10115
rect 2087 10081 2099 10115
rect 2222 10112 2228 10124
rect 2183 10084 2228 10112
rect 2041 10075 2099 10081
rect 2222 10072 2228 10084
rect 2280 10072 2286 10124
rect 2958 10112 2964 10124
rect 2919 10084 2964 10112
rect 2958 10072 2964 10084
rect 3016 10072 3022 10124
rect 3234 10072 3240 10124
rect 3292 10112 3298 10124
rect 3421 10115 3479 10121
rect 3421 10112 3433 10115
rect 3292 10084 3433 10112
rect 3292 10072 3298 10084
rect 3421 10081 3433 10084
rect 3467 10081 3479 10115
rect 3421 10075 3479 10081
rect 3510 10072 3516 10124
rect 3568 10112 3574 10124
rect 3697 10115 3755 10121
rect 3697 10112 3709 10115
rect 3568 10084 3709 10112
rect 3568 10072 3574 10084
rect 3697 10081 3709 10084
rect 3743 10081 3755 10115
rect 3697 10075 3755 10081
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 5169 10115 5227 10121
rect 5169 10112 5181 10115
rect 4856 10084 5181 10112
rect 4856 10072 4862 10084
rect 5169 10081 5181 10084
rect 5215 10081 5227 10115
rect 5169 10075 5227 10081
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10112 5411 10115
rect 6178 10112 6184 10124
rect 5399 10084 6184 10112
rect 5399 10081 5411 10084
rect 5353 10075 5411 10081
rect 6178 10072 6184 10084
rect 6236 10072 6242 10124
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10112 7251 10115
rect 7282 10112 7288 10124
rect 7239 10084 7288 10112
rect 7239 10081 7251 10084
rect 7193 10075 7251 10081
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 7576 10112 7604 10152
rect 7653 10149 7665 10183
rect 7699 10180 7711 10183
rect 8202 10180 8208 10192
rect 7699 10152 8208 10180
rect 7699 10149 7711 10152
rect 7653 10143 7711 10149
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 12526 10140 12532 10192
rect 12584 10180 12590 10192
rect 12682 10183 12740 10189
rect 12682 10180 12694 10183
rect 12584 10152 12694 10180
rect 12584 10140 12590 10152
rect 12682 10149 12694 10152
rect 12728 10149 12740 10183
rect 18414 10180 18420 10192
rect 12682 10143 12740 10149
rect 18340 10152 18420 10180
rect 7834 10112 7840 10124
rect 7576 10084 7840 10112
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 9030 10112 9036 10124
rect 8991 10084 9036 10112
rect 9030 10072 9036 10084
rect 9088 10072 9094 10124
rect 9217 10115 9275 10121
rect 9217 10081 9229 10115
rect 9263 10112 9275 10115
rect 9306 10112 9312 10124
rect 9263 10084 9312 10112
rect 9263 10081 9275 10084
rect 9217 10075 9275 10081
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10112 12495 10115
rect 14090 10112 14096 10124
rect 12483 10084 14096 10112
rect 12483 10081 12495 10084
rect 12437 10075 12495 10081
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 17034 10072 17040 10124
rect 17092 10112 17098 10124
rect 17497 10115 17555 10121
rect 17497 10112 17509 10115
rect 17092 10084 17509 10112
rect 17092 10072 17098 10084
rect 17497 10081 17509 10084
rect 17543 10081 17555 10115
rect 17497 10075 17555 10081
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 3528 10044 3556 10072
rect 2455 10016 3556 10044
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 4246 10004 4252 10056
rect 4304 10044 4310 10056
rect 5077 10047 5135 10053
rect 5077 10044 5089 10047
rect 4304 10016 5089 10044
rect 4304 10004 4310 10016
rect 5077 10013 5089 10016
rect 5123 10013 5135 10047
rect 5077 10007 5135 10013
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10044 5871 10047
rect 12158 10044 12164 10056
rect 5859 10016 12164 10044
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 12158 10004 12164 10016
rect 12216 10004 12222 10056
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10044 17647 10047
rect 17862 10044 17868 10056
rect 17635 10016 17868 10044
rect 17635 10013 17647 10016
rect 17589 10007 17647 10013
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 7466 9936 7472 9988
rect 7524 9976 7530 9988
rect 7929 9979 7987 9985
rect 7929 9976 7941 9979
rect 7524 9948 7941 9976
rect 7524 9936 7530 9948
rect 7929 9945 7941 9948
rect 7975 9945 7987 9979
rect 7929 9939 7987 9945
rect 15102 9936 15108 9988
rect 15160 9976 15166 9988
rect 18340 9976 18368 10152
rect 18414 10140 18420 10152
rect 18472 10140 18478 10192
rect 18601 10183 18659 10189
rect 18601 10149 18613 10183
rect 18647 10180 18659 10183
rect 19150 10180 19156 10192
rect 18647 10152 19156 10180
rect 18647 10149 18659 10152
rect 18601 10143 18659 10149
rect 19150 10140 19156 10152
rect 19208 10180 19214 10192
rect 22833 10183 22891 10189
rect 22833 10180 22845 10183
rect 19208 10152 22845 10180
rect 19208 10140 19214 10152
rect 22833 10149 22845 10152
rect 22879 10180 22891 10183
rect 23382 10180 23388 10192
rect 22879 10152 23388 10180
rect 22879 10149 22891 10152
rect 22833 10143 22891 10149
rect 23382 10140 23388 10152
rect 23440 10140 23446 10192
rect 23934 10140 23940 10192
rect 23992 10180 23998 10192
rect 23992 10152 24532 10180
rect 23992 10140 23998 10152
rect 18874 10112 18880 10124
rect 18835 10084 18880 10112
rect 18874 10072 18880 10084
rect 18932 10072 18938 10124
rect 18969 10115 19027 10121
rect 18969 10081 18981 10115
rect 19015 10112 19027 10115
rect 19242 10112 19248 10124
rect 19015 10084 19248 10112
rect 19015 10081 19027 10084
rect 18969 10075 19027 10081
rect 19242 10072 19248 10084
rect 19300 10072 19306 10124
rect 19383 10115 19441 10121
rect 19383 10081 19395 10115
rect 19429 10112 19441 10115
rect 19794 10112 19800 10124
rect 19429 10084 19800 10112
rect 19429 10081 19441 10084
rect 19383 10075 19441 10081
rect 19794 10072 19800 10084
rect 19852 10072 19858 10124
rect 20441 10115 20499 10121
rect 20441 10081 20453 10115
rect 20487 10081 20499 10115
rect 20714 10112 20720 10124
rect 20675 10084 20720 10112
rect 20441 10075 20499 10081
rect 18598 10004 18604 10056
rect 18656 10004 18662 10056
rect 15160 9948 18368 9976
rect 20456 9976 20484 10075
rect 20714 10072 20720 10084
rect 20772 10072 20778 10124
rect 21082 10112 21088 10124
rect 21043 10084 21088 10112
rect 21082 10072 21088 10084
rect 21140 10072 21146 10124
rect 21174 10072 21180 10124
rect 21232 10112 21238 10124
rect 22741 10115 22799 10121
rect 22741 10112 22753 10115
rect 21232 10084 22753 10112
rect 21232 10072 21238 10084
rect 22741 10081 22753 10084
rect 22787 10081 22799 10115
rect 22741 10075 22799 10081
rect 20806 10044 20812 10056
rect 20767 10016 20812 10044
rect 20806 10004 20812 10016
rect 20864 10004 20870 10056
rect 20456 9948 20852 9976
rect 15160 9936 15166 9948
rect 20824 9920 20852 9948
rect 6917 9911 6975 9917
rect 6917 9877 6929 9911
rect 6963 9908 6975 9911
rect 7650 9908 7656 9920
rect 6963 9880 7656 9908
rect 6963 9877 6975 9880
rect 6917 9871 6975 9877
rect 7650 9868 7656 9880
rect 7708 9868 7714 9920
rect 12618 9868 12624 9920
rect 12676 9908 12682 9920
rect 13817 9911 13875 9917
rect 13817 9908 13829 9911
rect 12676 9880 13829 9908
rect 12676 9868 12682 9880
rect 13817 9877 13829 9880
rect 13863 9877 13875 9911
rect 13817 9871 13875 9877
rect 19889 9911 19947 9917
rect 19889 9877 19901 9911
rect 19935 9908 19947 9911
rect 20438 9908 20444 9920
rect 19935 9880 20444 9908
rect 19935 9877 19947 9880
rect 19889 9871 19947 9877
rect 20438 9868 20444 9880
rect 20496 9868 20502 9920
rect 20806 9868 20812 9920
rect 20864 9868 20870 9920
rect 22756 9908 22784 10075
rect 23566 10072 23572 10124
rect 23624 10112 23630 10124
rect 23661 10115 23719 10121
rect 23661 10112 23673 10115
rect 23624 10084 23673 10112
rect 23624 10072 23630 10084
rect 23661 10081 23673 10084
rect 23707 10081 23719 10115
rect 23661 10075 23719 10081
rect 23842 10072 23848 10124
rect 23900 10112 23906 10124
rect 24504 10121 24532 10152
rect 24670 10140 24676 10192
rect 24728 10180 24734 10192
rect 25654 10183 25712 10189
rect 25654 10180 25666 10183
rect 24728 10152 25666 10180
rect 24728 10140 24734 10152
rect 25654 10149 25666 10152
rect 25700 10149 25712 10183
rect 25654 10143 25712 10149
rect 24213 10115 24271 10121
rect 24213 10112 24225 10115
rect 23900 10084 24225 10112
rect 23900 10072 23906 10084
rect 24213 10081 24225 10084
rect 24259 10081 24271 10115
rect 24213 10075 24271 10081
rect 24489 10115 24547 10121
rect 24489 10081 24501 10115
rect 24535 10081 24547 10115
rect 24489 10075 24547 10081
rect 25409 10115 25467 10121
rect 25409 10081 25421 10115
rect 25455 10112 25467 10115
rect 25498 10112 25504 10124
rect 25455 10084 25504 10112
rect 25455 10081 25467 10084
rect 25409 10075 25467 10081
rect 25498 10072 25504 10084
rect 25556 10072 25562 10124
rect 27893 10115 27951 10121
rect 27893 10081 27905 10115
rect 27939 10112 27951 10115
rect 28350 10112 28356 10124
rect 27939 10084 28356 10112
rect 27939 10081 27951 10084
rect 27893 10075 27951 10081
rect 28350 10072 28356 10084
rect 28408 10072 28414 10124
rect 24762 10044 24768 10056
rect 24723 10016 24768 10044
rect 24762 10004 24768 10016
rect 24820 10004 24826 10056
rect 27890 9908 27896 9920
rect 22756 9880 27896 9908
rect 27890 9868 27896 9880
rect 27948 9868 27954 9920
rect 1104 9818 28888 9840
rect 1104 9766 5614 9818
rect 5666 9766 5678 9818
rect 5730 9766 5742 9818
rect 5794 9766 5806 9818
rect 5858 9766 14878 9818
rect 14930 9766 14942 9818
rect 14994 9766 15006 9818
rect 15058 9766 15070 9818
rect 15122 9766 24142 9818
rect 24194 9766 24206 9818
rect 24258 9766 24270 9818
rect 24322 9766 24334 9818
rect 24386 9766 28888 9818
rect 1104 9744 28888 9766
rect 2866 9704 2872 9716
rect 2827 9676 2872 9704
rect 2866 9664 2872 9676
rect 2924 9664 2930 9716
rect 4709 9707 4767 9713
rect 4709 9673 4721 9707
rect 4755 9704 4767 9707
rect 5350 9704 5356 9716
rect 4755 9676 5356 9704
rect 4755 9673 4767 9676
rect 4709 9667 4767 9673
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 12437 9707 12495 9713
rect 12437 9673 12449 9707
rect 12483 9704 12495 9707
rect 13446 9704 13452 9716
rect 12483 9676 13452 9704
rect 12483 9673 12495 9676
rect 12437 9667 12495 9673
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 15562 9664 15568 9716
rect 15620 9704 15626 9716
rect 16206 9704 16212 9716
rect 15620 9676 16212 9704
rect 15620 9664 15626 9676
rect 16206 9664 16212 9676
rect 16264 9664 16270 9716
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 21910 9704 21916 9716
rect 16632 9676 20024 9704
rect 21871 9676 21916 9704
rect 16632 9664 16638 9676
rect 7009 9639 7067 9645
rect 7009 9605 7021 9639
rect 7055 9636 7067 9639
rect 7466 9636 7472 9648
rect 7055 9608 7472 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 7466 9596 7472 9608
rect 7524 9636 7530 9648
rect 10594 9636 10600 9648
rect 7524 9608 10600 9636
rect 7524 9596 7530 9608
rect 10594 9596 10600 9608
rect 10652 9596 10658 9648
rect 11149 9639 11207 9645
rect 11149 9605 11161 9639
rect 11195 9636 11207 9639
rect 11195 9608 15148 9636
rect 11195 9605 11207 9608
rect 11149 9599 11207 9605
rect 1400 9580 1452 9586
rect 7650 9568 7656 9580
rect 7611 9540 7656 9568
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 11790 9568 11796 9580
rect 11751 9540 11796 9568
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 12250 9528 12256 9580
rect 12308 9568 12314 9580
rect 12308 9540 14688 9568
rect 12308 9528 12314 9540
rect 1400 9522 1452 9528
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9500 1915 9503
rect 2406 9500 2412 9512
rect 1903 9472 2412 9500
rect 1903 9469 1915 9472
rect 1857 9463 1915 9469
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 3050 9460 3056 9512
rect 3108 9500 3114 9512
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 3108 9472 4261 9500
rect 3108 9460 3114 9472
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4801 9503 4859 9509
rect 4801 9469 4813 9503
rect 4847 9500 4859 9503
rect 4890 9500 4896 9512
rect 4847 9472 4896 9500
rect 4847 9469 4859 9472
rect 4801 9463 4859 9469
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 1949 9435 2007 9441
rect 1949 9401 1961 9435
rect 1995 9432 2007 9435
rect 2038 9432 2044 9444
rect 1995 9404 2044 9432
rect 1995 9401 2007 9404
rect 1949 9395 2007 9401
rect 2038 9392 2044 9404
rect 2096 9392 2102 9444
rect 2314 9432 2320 9444
rect 2275 9404 2320 9432
rect 2314 9392 2320 9404
rect 2372 9392 2378 9444
rect 2958 9432 2964 9444
rect 2424 9404 2964 9432
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 2424 9364 2452 9404
rect 2958 9392 2964 9404
rect 3016 9432 3022 9444
rect 3694 9432 3700 9444
rect 3016 9404 3700 9432
rect 3016 9392 3022 9404
rect 3694 9392 3700 9404
rect 3752 9392 3758 9444
rect 2682 9364 2688 9376
rect 1627 9336 2452 9364
rect 2643 9336 2688 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 4341 9367 4399 9373
rect 4341 9364 4353 9367
rect 3476 9336 4353 9364
rect 3476 9324 3482 9336
rect 4341 9333 4353 9336
rect 4387 9333 4399 9367
rect 4522 9364 4528 9376
rect 4483 9336 4528 9364
rect 4341 9327 4399 9333
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 4890 9324 4896 9376
rect 4948 9364 4954 9376
rect 5644 9364 5672 9463
rect 6178 9460 6184 9512
rect 6236 9500 6242 9512
rect 6236 9472 6960 9500
rect 6236 9460 6242 9472
rect 5896 9435 5954 9441
rect 5896 9401 5908 9435
rect 5942 9432 5954 9435
rect 6822 9432 6828 9444
rect 5942 9404 6828 9432
rect 5942 9401 5954 9404
rect 5896 9395 5954 9401
rect 6822 9392 6828 9404
rect 6880 9392 6886 9444
rect 6932 9432 6960 9472
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7432 9472 7757 9500
rect 7432 9460 7438 9472
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 10778 9460 10784 9512
rect 10836 9500 10842 9512
rect 11698 9500 11704 9512
rect 10836 9472 11704 9500
rect 10836 9460 10842 9472
rect 11698 9460 11704 9472
rect 11756 9500 11762 9512
rect 12345 9503 12403 9509
rect 12345 9500 12357 9503
rect 11756 9472 12357 9500
rect 11756 9460 11762 9472
rect 12345 9469 12357 9472
rect 12391 9469 12403 9503
rect 12345 9463 12403 9469
rect 12529 9503 12587 9509
rect 12529 9469 12541 9503
rect 12575 9500 12587 9503
rect 14182 9500 14188 9512
rect 12575 9472 14188 9500
rect 12575 9469 12587 9472
rect 12529 9463 12587 9469
rect 14182 9460 14188 9472
rect 14240 9460 14246 9512
rect 11514 9432 11520 9444
rect 6932 9404 8248 9432
rect 11475 9404 11520 9432
rect 6914 9364 6920 9376
rect 4948 9336 6920 9364
rect 4948 9324 4954 9336
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 8113 9367 8171 9373
rect 8113 9364 8125 9367
rect 7248 9336 8125 9364
rect 7248 9324 7254 9336
rect 8113 9333 8125 9336
rect 8159 9333 8171 9367
rect 8220 9364 8248 9404
rect 11514 9392 11520 9404
rect 11572 9392 11578 9444
rect 12066 9392 12072 9444
rect 12124 9432 12130 9444
rect 14458 9432 14464 9444
rect 12124 9404 14464 9432
rect 12124 9392 12130 9404
rect 14458 9392 14464 9404
rect 14516 9392 14522 9444
rect 14660 9432 14688 9540
rect 14734 9460 14740 9512
rect 14792 9500 14798 9512
rect 15120 9509 15148 9608
rect 15749 9571 15807 9577
rect 15749 9537 15761 9571
rect 15795 9568 15807 9571
rect 16758 9568 16764 9580
rect 15795 9540 16764 9568
rect 15795 9537 15807 9540
rect 15749 9531 15807 9537
rect 16758 9528 16764 9540
rect 16816 9528 16822 9580
rect 19996 9568 20024 9676
rect 21910 9664 21916 9676
rect 21968 9664 21974 9716
rect 22925 9639 22983 9645
rect 22925 9605 22937 9639
rect 22971 9636 22983 9639
rect 22971 9608 25820 9636
rect 22971 9605 22983 9608
rect 22925 9599 22983 9605
rect 23382 9568 23388 9580
rect 19996 9540 20116 9568
rect 23343 9540 23388 9568
rect 17586 9509 17592 9512
rect 15013 9503 15071 9509
rect 15013 9500 15025 9503
rect 14792 9472 15025 9500
rect 14792 9460 14798 9472
rect 15013 9469 15025 9472
rect 15059 9469 15071 9503
rect 15013 9463 15071 9469
rect 15105 9503 15163 9509
rect 15105 9469 15117 9503
rect 15151 9469 15163 9503
rect 15105 9463 15163 9469
rect 15289 9503 15347 9509
rect 15289 9469 15301 9503
rect 15335 9469 15347 9503
rect 15289 9463 15347 9469
rect 17313 9503 17371 9509
rect 17313 9469 17325 9503
rect 17359 9469 17371 9503
rect 17580 9500 17592 9509
rect 17547 9472 17592 9500
rect 17313 9463 17371 9469
rect 17580 9463 17592 9472
rect 15304 9432 15332 9463
rect 16390 9432 16396 9444
rect 14660 9404 16396 9432
rect 16390 9392 16396 9404
rect 16448 9392 16454 9444
rect 17126 9392 17132 9444
rect 17184 9432 17190 9444
rect 17328 9432 17356 9463
rect 17586 9460 17592 9463
rect 17644 9460 17650 9512
rect 19886 9500 19892 9512
rect 17696 9472 19892 9500
rect 17696 9432 17724 9472
rect 19886 9460 19892 9472
rect 19944 9500 19950 9512
rect 19981 9503 20039 9509
rect 19981 9500 19993 9503
rect 19944 9472 19993 9500
rect 19944 9460 19950 9472
rect 19981 9469 19993 9472
rect 20027 9469 20039 9503
rect 20088 9500 20116 9540
rect 23382 9528 23388 9540
rect 23440 9528 23446 9580
rect 23566 9568 23572 9580
rect 23527 9540 23572 9568
rect 23566 9528 23572 9540
rect 23624 9568 23630 9580
rect 25590 9568 25596 9580
rect 23624 9540 25596 9568
rect 23624 9528 23630 9540
rect 25590 9528 25596 9540
rect 25648 9528 25654 9580
rect 25792 9577 25820 9608
rect 26418 9596 26424 9648
rect 26476 9636 26482 9648
rect 26789 9639 26847 9645
rect 26789 9636 26801 9639
rect 26476 9608 26801 9636
rect 26476 9596 26482 9608
rect 26789 9605 26801 9608
rect 26835 9605 26847 9639
rect 26789 9599 26847 9605
rect 25777 9571 25835 9577
rect 25777 9537 25789 9571
rect 25823 9537 25835 9571
rect 25777 9531 25835 9537
rect 25961 9571 26019 9577
rect 25961 9537 25973 9571
rect 26007 9568 26019 9571
rect 26050 9568 26056 9580
rect 26007 9540 26056 9568
rect 26007 9537 26019 9540
rect 25961 9531 26019 9537
rect 26050 9528 26056 9540
rect 26108 9528 26114 9580
rect 21818 9500 21824 9512
rect 20088 9472 20944 9500
rect 21779 9472 21824 9500
rect 19981 9463 20039 9469
rect 20916 9444 20944 9472
rect 21818 9460 21824 9472
rect 21876 9460 21882 9512
rect 22646 9460 22652 9512
rect 22704 9500 22710 9512
rect 23293 9503 23351 9509
rect 23293 9500 23305 9503
rect 22704 9472 23305 9500
rect 22704 9460 22710 9472
rect 23293 9469 23305 9472
rect 23339 9469 23351 9503
rect 23293 9463 23351 9469
rect 25685 9503 25743 9509
rect 25685 9469 25697 9503
rect 25731 9500 25743 9503
rect 26234 9500 26240 9512
rect 25731 9472 26240 9500
rect 25731 9469 25743 9472
rect 25685 9463 25743 9469
rect 26234 9460 26240 9472
rect 26292 9460 26298 9512
rect 26602 9500 26608 9512
rect 26563 9472 26608 9500
rect 26602 9460 26608 9472
rect 26660 9460 26666 9512
rect 27154 9460 27160 9512
rect 27212 9500 27218 9512
rect 27430 9500 27436 9512
rect 27212 9472 27257 9500
rect 27391 9472 27436 9500
rect 27212 9460 27218 9472
rect 27430 9460 27436 9472
rect 27488 9460 27494 9512
rect 17184 9404 17724 9432
rect 17184 9392 17190 9404
rect 19058 9392 19064 9444
rect 19116 9432 19122 9444
rect 20226 9435 20284 9441
rect 20226 9432 20238 9435
rect 19116 9404 20238 9432
rect 19116 9392 19122 9404
rect 20226 9401 20238 9404
rect 20272 9401 20284 9435
rect 20226 9395 20284 9401
rect 20898 9392 20904 9444
rect 20956 9392 20962 9444
rect 26620 9432 26648 9460
rect 25332 9404 26648 9432
rect 11054 9364 11060 9376
rect 8220 9336 11060 9364
rect 8113 9327 8171 9333
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 11606 9364 11612 9376
rect 11567 9336 11612 9364
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 11790 9324 11796 9376
rect 11848 9364 11854 9376
rect 14274 9364 14280 9376
rect 11848 9336 14280 9364
rect 11848 9324 11854 9336
rect 14274 9324 14280 9336
rect 14332 9324 14338 9376
rect 15470 9324 15476 9376
rect 15528 9364 15534 9376
rect 15930 9364 15936 9376
rect 15528 9336 15936 9364
rect 15528 9324 15534 9336
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 18690 9364 18696 9376
rect 18603 9336 18696 9364
rect 18690 9324 18696 9336
rect 18748 9364 18754 9376
rect 19334 9364 19340 9376
rect 18748 9336 19340 9364
rect 18748 9324 18754 9336
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 21361 9367 21419 9373
rect 21361 9333 21373 9367
rect 21407 9364 21419 9367
rect 21818 9364 21824 9376
rect 21407 9336 21824 9364
rect 21407 9333 21419 9336
rect 21361 9327 21419 9333
rect 21818 9324 21824 9336
rect 21876 9324 21882 9376
rect 25332 9373 25360 9404
rect 25317 9367 25375 9373
rect 25317 9333 25329 9367
rect 25363 9333 25375 9367
rect 25317 9327 25375 9333
rect 1104 9274 28888 9296
rect 1104 9222 10246 9274
rect 10298 9222 10310 9274
rect 10362 9222 10374 9274
rect 10426 9222 10438 9274
rect 10490 9222 19510 9274
rect 19562 9222 19574 9274
rect 19626 9222 19638 9274
rect 19690 9222 19702 9274
rect 19754 9222 28888 9274
rect 1104 9200 28888 9222
rect 3142 9120 3148 9172
rect 3200 9160 3206 9172
rect 3237 9163 3295 9169
rect 3237 9160 3249 9163
rect 3200 9132 3249 9160
rect 3200 9120 3206 9132
rect 3237 9129 3249 9132
rect 3283 9129 3295 9163
rect 3418 9160 3424 9172
rect 3379 9132 3424 9160
rect 3237 9123 3295 9129
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 4430 9160 4436 9172
rect 3528 9132 4436 9160
rect 1854 9092 1860 9104
rect 1815 9064 1860 9092
rect 1854 9052 1860 9064
rect 1912 9052 1918 9104
rect 2501 9027 2559 9033
rect 2501 8993 2513 9027
rect 2547 9024 2559 9027
rect 3050 9024 3056 9036
rect 2547 8996 3056 9024
rect 2547 8993 2559 8996
rect 2501 8987 2559 8993
rect 3050 8984 3056 8996
rect 3108 8984 3114 9036
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 9024 3203 9027
rect 3418 9024 3424 9036
rect 3191 8996 3424 9024
rect 3191 8993 3203 8996
rect 3145 8987 3203 8993
rect 3418 8984 3424 8996
rect 3476 8984 3482 9036
rect 3528 9033 3556 9132
rect 4430 9120 4436 9132
rect 4488 9120 4494 9172
rect 6822 9160 6828 9172
rect 6783 9132 6828 9160
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7190 9160 7196 9172
rect 7151 9132 7196 9160
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 7285 9163 7343 9169
rect 7285 9129 7297 9163
rect 7331 9160 7343 9163
rect 7466 9160 7472 9172
rect 7331 9132 7472 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 8941 9163 8999 9169
rect 8941 9129 8953 9163
rect 8987 9160 8999 9163
rect 10413 9163 10471 9169
rect 10413 9160 10425 9163
rect 8987 9132 10425 9160
rect 8987 9129 8999 9132
rect 8941 9123 8999 9129
rect 10413 9129 10425 9132
rect 10459 9129 10471 9163
rect 10413 9123 10471 9129
rect 10781 9163 10839 9169
rect 10781 9129 10793 9163
rect 10827 9160 10839 9163
rect 11606 9160 11612 9172
rect 10827 9132 11612 9160
rect 10827 9129 10839 9132
rect 10781 9123 10839 9129
rect 11606 9120 11612 9132
rect 11664 9160 11670 9172
rect 12161 9163 12219 9169
rect 12161 9160 12173 9163
rect 11664 9132 12173 9160
rect 11664 9120 11670 9132
rect 12161 9129 12173 9132
rect 12207 9129 12219 9163
rect 25777 9163 25835 9169
rect 25777 9160 25789 9163
rect 12161 9123 12219 9129
rect 12268 9132 25789 9160
rect 4338 9052 4344 9104
rect 4396 9092 4402 9104
rect 12268 9092 12296 9132
rect 25777 9129 25789 9132
rect 25823 9129 25835 9163
rect 25777 9123 25835 9129
rect 25866 9120 25872 9172
rect 25924 9160 25930 9172
rect 28258 9160 28264 9172
rect 25924 9132 25969 9160
rect 26206 9132 28264 9160
rect 25924 9120 25930 9132
rect 14366 9092 14372 9104
rect 4396 9064 4441 9092
rect 6840 9064 12296 9092
rect 12406 9064 13952 9092
rect 14327 9064 14372 9092
rect 4396 9052 4402 9064
rect 3513 9027 3571 9033
rect 3513 8993 3525 9027
rect 3559 8993 3571 9027
rect 3513 8987 3571 8993
rect 3694 8984 3700 9036
rect 3752 9024 3758 9036
rect 4249 9027 4307 9033
rect 4249 9024 4261 9027
rect 3752 8996 4261 9024
rect 3752 8984 3758 8996
rect 4249 8993 4261 8996
rect 4295 8993 4307 9027
rect 4249 8987 4307 8993
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3329 8959 3387 8965
rect 3329 8956 3341 8959
rect 3292 8928 3341 8956
rect 3292 8916 3298 8928
rect 3329 8925 3341 8928
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 6840 8956 6868 9064
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 8294 9024 8300 9036
rect 6972 8996 8300 9024
rect 6972 8984 6978 8996
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 8754 9024 8760 9036
rect 8715 8996 8760 9024
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 9585 9027 9643 9033
rect 9585 8993 9597 9027
rect 9631 9024 9643 9027
rect 9858 9024 9864 9036
rect 9631 8996 9864 9024
rect 9631 8993 9643 8996
rect 9585 8987 9643 8993
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 12084 9033 12112 9064
rect 12069 9027 12127 9033
rect 10796 8996 11008 9024
rect 4203 8928 6868 8956
rect 7469 8959 7527 8965
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 7469 8925 7481 8959
rect 7515 8956 7527 8959
rect 7558 8956 7564 8968
rect 7515 8928 7564 8956
rect 7515 8925 7527 8928
rect 7469 8919 7527 8925
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 7834 8916 7840 8968
rect 7892 8956 7898 8968
rect 9033 8959 9091 8965
rect 9033 8956 9045 8959
rect 7892 8928 9045 8956
rect 7892 8916 7898 8928
rect 9033 8925 9045 8928
rect 9079 8925 9091 8959
rect 9033 8919 9091 8925
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 10796 8956 10824 8996
rect 10980 8965 11008 8996
rect 12069 8993 12081 9027
rect 12115 8993 12127 9027
rect 12069 8987 12127 8993
rect 9548 8928 10824 8956
rect 10873 8959 10931 8965
rect 9548 8916 9554 8928
rect 10873 8925 10885 8959
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 2593 8891 2651 8897
rect 2593 8857 2605 8891
rect 2639 8888 2651 8891
rect 10888 8888 10916 8919
rect 11054 8916 11060 8968
rect 11112 8956 11118 8968
rect 12406 8956 12434 9064
rect 12618 8984 12624 9036
rect 12676 9024 12682 9036
rect 12713 9027 12771 9033
rect 12713 9024 12725 9027
rect 12676 8996 12725 9024
rect 12676 8984 12682 8996
rect 12713 8993 12725 8996
rect 12759 8993 12771 9027
rect 12713 8987 12771 8993
rect 12805 9027 12863 9033
rect 12805 8993 12817 9027
rect 12851 9024 12863 9027
rect 13078 9024 13084 9036
rect 12851 8996 13084 9024
rect 12851 8993 12863 8996
rect 12805 8987 12863 8993
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 13924 9033 13952 9064
rect 14366 9052 14372 9064
rect 14424 9052 14430 9104
rect 15194 9092 15200 9104
rect 15155 9064 15200 9092
rect 15194 9052 15200 9064
rect 15252 9052 15258 9104
rect 20533 9095 20591 9101
rect 20533 9061 20545 9095
rect 20579 9092 20591 9095
rect 20714 9092 20720 9104
rect 20579 9064 20720 9092
rect 20579 9061 20591 9064
rect 20533 9055 20591 9061
rect 20714 9052 20720 9064
rect 20772 9052 20778 9104
rect 22646 9092 22652 9104
rect 22607 9064 22652 9092
rect 22646 9052 22652 9064
rect 22704 9052 22710 9104
rect 24029 9095 24087 9101
rect 24029 9061 24041 9095
rect 24075 9092 24087 9095
rect 26206 9092 26234 9132
rect 28258 9120 28264 9132
rect 28316 9120 28322 9172
rect 24075 9064 26234 9092
rect 24075 9061 24087 9064
rect 24029 9055 24087 9061
rect 26418 9052 26424 9104
rect 26476 9092 26482 9104
rect 26605 9095 26663 9101
rect 26605 9092 26617 9095
rect 26476 9064 26617 9092
rect 26476 9052 26482 9064
rect 26605 9061 26617 9064
rect 26651 9061 26663 9095
rect 26786 9092 26792 9104
rect 26747 9064 26792 9092
rect 26605 9055 26663 9061
rect 26786 9052 26792 9064
rect 26844 9052 26850 9104
rect 27890 9052 27896 9104
rect 27948 9092 27954 9104
rect 27985 9095 28043 9101
rect 27985 9092 27997 9095
rect 27948 9064 27997 9092
rect 27948 9052 27954 9064
rect 27985 9061 27997 9064
rect 28031 9061 28043 9095
rect 27985 9055 28043 9061
rect 13725 9027 13783 9033
rect 13725 8993 13737 9027
rect 13771 8993 13783 9027
rect 13725 8987 13783 8993
rect 13909 9027 13967 9033
rect 13909 8993 13921 9027
rect 13955 8993 13967 9027
rect 13909 8987 13967 8993
rect 11112 8928 12434 8956
rect 11112 8916 11118 8928
rect 13354 8916 13360 8968
rect 13412 8956 13418 8968
rect 13633 8959 13691 8965
rect 13633 8956 13645 8959
rect 13412 8928 13645 8956
rect 13412 8916 13418 8928
rect 13633 8925 13645 8928
rect 13679 8925 13691 8959
rect 13740 8956 13768 8987
rect 14458 8984 14464 9036
rect 14516 9024 14522 9036
rect 16022 9024 16028 9036
rect 14516 8996 15608 9024
rect 15983 8996 16028 9024
rect 14516 8984 14522 8996
rect 13740 8928 14872 8956
rect 13633 8919 13691 8925
rect 14844 8897 14872 8928
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 15160 8928 15301 8956
rect 15160 8916 15166 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 15470 8956 15476 8968
rect 15431 8928 15476 8956
rect 15289 8919 15347 8925
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 15580 8956 15608 8996
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 20438 9024 20444 9036
rect 20399 8996 20444 9024
rect 20438 8984 20444 8996
rect 20496 8984 20502 9036
rect 22557 9027 22615 9033
rect 22557 8993 22569 9027
rect 22603 8993 22615 9027
rect 22557 8987 22615 8993
rect 23293 9027 23351 9033
rect 23293 8993 23305 9027
rect 23339 9024 23351 9027
rect 23382 9024 23388 9036
rect 23339 8996 23388 9024
rect 23339 8993 23351 8996
rect 23293 8987 23351 8993
rect 17678 8956 17684 8968
rect 15580 8928 17684 8956
rect 17678 8916 17684 8928
rect 17736 8916 17742 8968
rect 22572 8956 22600 8987
rect 23382 8984 23388 8996
rect 23440 8984 23446 9036
rect 24765 9027 24823 9033
rect 24765 9024 24777 9027
rect 23492 8996 24777 9024
rect 22738 8956 22744 8968
rect 22572 8928 22744 8956
rect 22738 8916 22744 8928
rect 22796 8956 22802 8968
rect 23492 8956 23520 8996
rect 24765 8993 24777 8996
rect 24811 8993 24823 9027
rect 24765 8987 24823 8993
rect 26881 9027 26939 9033
rect 26881 8993 26893 9027
rect 26927 9024 26939 9027
rect 26970 9024 26976 9036
rect 26927 8996 26976 9024
rect 26927 8993 26939 8996
rect 26881 8987 26939 8993
rect 26970 8984 26976 8996
rect 27028 8984 27034 9036
rect 22796 8928 23520 8956
rect 24213 8959 24271 8965
rect 22796 8916 22802 8928
rect 24213 8925 24225 8959
rect 24259 8956 24271 8959
rect 24854 8956 24860 8968
rect 24259 8928 24860 8956
rect 24259 8925 24271 8928
rect 24213 8919 24271 8925
rect 24854 8916 24860 8928
rect 24912 8916 24918 8968
rect 25590 8916 25596 8968
rect 25648 8956 25654 8968
rect 25961 8959 26019 8965
rect 25961 8956 25973 8959
rect 25648 8928 25973 8956
rect 25648 8916 25654 8928
rect 25961 8925 25973 8928
rect 26007 8925 26019 8959
rect 25961 8919 26019 8925
rect 14829 8891 14887 8897
rect 2639 8860 12434 8888
rect 2639 8857 2651 8860
rect 2593 8851 2651 8857
rect 1949 8823 2007 8829
rect 1949 8789 1961 8823
rect 1995 8820 2007 8823
rect 2314 8820 2320 8832
rect 1995 8792 2320 8820
rect 1995 8789 2007 8792
rect 1949 8783 2007 8789
rect 2314 8780 2320 8792
rect 2372 8820 2378 8832
rect 4157 8823 4215 8829
rect 4157 8820 4169 8823
rect 2372 8792 4169 8820
rect 2372 8780 2378 8792
rect 4157 8789 4169 8792
rect 4203 8789 4215 8823
rect 4157 8783 4215 8789
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 7834 8820 7840 8832
rect 5960 8792 7840 8820
rect 5960 8780 5966 8792
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 8481 8823 8539 8829
rect 8481 8820 8493 8823
rect 8444 8792 8493 8820
rect 8444 8780 8450 8792
rect 8481 8789 8493 8792
rect 8527 8789 8539 8823
rect 8481 8783 8539 8789
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 9769 8823 9827 8829
rect 9769 8820 9781 8823
rect 8628 8792 9781 8820
rect 8628 8780 8634 8792
rect 9769 8789 9781 8792
rect 9815 8820 9827 8823
rect 10134 8820 10140 8832
rect 9815 8792 10140 8820
rect 9815 8789 9827 8792
rect 9769 8783 9827 8789
rect 10134 8780 10140 8792
rect 10192 8780 10198 8832
rect 12406 8820 12434 8860
rect 14829 8857 14841 8891
rect 14875 8857 14887 8891
rect 18138 8888 18144 8900
rect 14829 8851 14887 8857
rect 15948 8860 18144 8888
rect 15948 8820 15976 8860
rect 18138 8848 18144 8860
rect 18196 8848 18202 8900
rect 23385 8891 23443 8897
rect 23385 8857 23397 8891
rect 23431 8888 23443 8891
rect 23842 8888 23848 8900
rect 23431 8860 23848 8888
rect 23431 8857 23443 8860
rect 23385 8851 23443 8857
rect 23842 8848 23848 8860
rect 23900 8848 23906 8900
rect 24946 8888 24952 8900
rect 24907 8860 24952 8888
rect 24946 8848 24952 8860
rect 25004 8848 25010 8900
rect 25406 8888 25412 8900
rect 25367 8860 25412 8888
rect 25406 8848 25412 8860
rect 25464 8848 25470 8900
rect 16114 8820 16120 8832
rect 12406 8792 15976 8820
rect 16075 8792 16120 8820
rect 16114 8780 16120 8792
rect 16172 8780 16178 8832
rect 24854 8780 24860 8832
rect 24912 8820 24918 8832
rect 26050 8820 26056 8832
rect 24912 8792 26056 8820
rect 24912 8780 24918 8792
rect 26050 8780 26056 8792
rect 26108 8780 26114 8832
rect 26881 8823 26939 8829
rect 26881 8789 26893 8823
rect 26927 8820 26939 8823
rect 27522 8820 27528 8832
rect 26927 8792 27528 8820
rect 26927 8789 26939 8792
rect 26881 8783 26939 8789
rect 27522 8780 27528 8792
rect 27580 8780 27586 8832
rect 28074 8820 28080 8832
rect 28035 8792 28080 8820
rect 28074 8780 28080 8792
rect 28132 8780 28138 8832
rect 1104 8730 28888 8752
rect 1104 8678 5614 8730
rect 5666 8678 5678 8730
rect 5730 8678 5742 8730
rect 5794 8678 5806 8730
rect 5858 8678 14878 8730
rect 14930 8678 14942 8730
rect 14994 8678 15006 8730
rect 15058 8678 15070 8730
rect 15122 8678 24142 8730
rect 24194 8678 24206 8730
rect 24258 8678 24270 8730
rect 24322 8678 24334 8730
rect 24386 8678 28888 8730
rect 1104 8656 28888 8678
rect 2406 8576 2412 8628
rect 2464 8616 2470 8628
rect 2593 8619 2651 8625
rect 2593 8616 2605 8619
rect 2464 8588 2605 8616
rect 2464 8576 2470 8588
rect 2593 8585 2605 8588
rect 2639 8585 2651 8619
rect 3050 8616 3056 8628
rect 3011 8588 3056 8616
rect 2593 8579 2651 8585
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 4890 8616 4896 8628
rect 4264 8588 4896 8616
rect 1765 8551 1823 8557
rect 1765 8517 1777 8551
rect 1811 8548 1823 8551
rect 4062 8548 4068 8560
rect 1811 8520 4068 8548
rect 1811 8517 1823 8520
rect 1765 8511 1823 8517
rect 4062 8508 4068 8520
rect 4120 8508 4126 8560
rect 4264 8489 4292 8588
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5258 8576 5264 8628
rect 5316 8616 5322 8628
rect 5629 8619 5687 8625
rect 5629 8616 5641 8619
rect 5316 8588 5641 8616
rect 5316 8576 5322 8588
rect 5629 8585 5641 8588
rect 5675 8616 5687 8619
rect 12066 8616 12072 8628
rect 5675 8588 12072 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 12342 8576 12348 8628
rect 12400 8616 12406 8628
rect 13170 8616 13176 8628
rect 12400 8588 13176 8616
rect 12400 8576 12406 8588
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13354 8616 13360 8628
rect 13315 8588 13360 8616
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 14829 8619 14887 8625
rect 14829 8616 14841 8619
rect 14792 8588 14841 8616
rect 14792 8576 14798 8588
rect 14829 8585 14841 8588
rect 14875 8585 14887 8619
rect 26970 8616 26976 8628
rect 26931 8588 26976 8616
rect 14829 8579 14887 8585
rect 26970 8576 26976 8588
rect 27028 8576 27034 8628
rect 27982 8576 27988 8628
rect 28040 8616 28046 8628
rect 28169 8619 28227 8625
rect 28169 8616 28181 8619
rect 28040 8588 28181 8616
rect 28040 8576 28046 8588
rect 28169 8585 28181 8588
rect 28215 8585 28227 8619
rect 28169 8579 28227 8585
rect 5994 8508 6000 8560
rect 6052 8548 6058 8560
rect 9490 8548 9496 8560
rect 6052 8520 9496 8548
rect 6052 8508 6058 8520
rect 9490 8508 9496 8520
rect 9548 8508 9554 8560
rect 9858 8508 9864 8560
rect 9916 8548 9922 8560
rect 9916 8520 10088 8548
rect 9916 8508 9922 8520
rect 10060 8489 10088 8520
rect 10870 8508 10876 8560
rect 10928 8548 10934 8560
rect 11793 8551 11851 8557
rect 11793 8548 11805 8551
rect 10928 8520 11805 8548
rect 10928 8508 10934 8520
rect 11793 8517 11805 8520
rect 11839 8517 11851 8551
rect 18230 8548 18236 8560
rect 11793 8511 11851 8517
rect 11992 8520 18236 8548
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 10045 8483 10103 8489
rect 10045 8449 10057 8483
rect 10091 8480 10103 8483
rect 10962 8480 10968 8492
rect 10091 8452 10968 8480
rect 10091 8449 10103 8452
rect 10045 8443 10103 8449
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 1946 8412 1952 8424
rect 1907 8384 1952 8412
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 2406 8412 2412 8424
rect 2367 8384 2412 8412
rect 2406 8372 2412 8384
rect 2464 8372 2470 8424
rect 3234 8412 3240 8424
rect 3195 8384 3240 8412
rect 3234 8372 3240 8384
rect 3292 8372 3298 8424
rect 4522 8421 4528 8424
rect 4516 8412 4528 8421
rect 4483 8384 4528 8412
rect 4516 8375 4528 8384
rect 4522 8372 4528 8375
rect 4580 8372 4586 8424
rect 9953 8415 10011 8421
rect 9953 8381 9965 8415
rect 9999 8412 10011 8415
rect 11514 8412 11520 8424
rect 9999 8384 11520 8412
rect 9999 8381 10011 8384
rect 9953 8375 10011 8381
rect 11514 8372 11520 8384
rect 11572 8372 11578 8424
rect 2314 8304 2320 8356
rect 2372 8344 2378 8356
rect 11992 8344 12020 8520
rect 18230 8508 18236 8520
rect 18288 8508 18294 8560
rect 24213 8551 24271 8557
rect 24213 8517 24225 8551
rect 24259 8548 24271 8551
rect 24259 8520 26740 8548
rect 24259 8517 24271 8520
rect 24213 8511 24271 8517
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8480 12311 8483
rect 13078 8480 13084 8492
rect 12299 8452 13084 8480
rect 12299 8449 12311 8452
rect 12253 8443 12311 8449
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 16114 8480 16120 8492
rect 16075 8452 16120 8480
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16850 8480 16856 8492
rect 16811 8452 16856 8480
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 21818 8440 21824 8492
rect 21876 8480 21882 8492
rect 26329 8483 26387 8489
rect 21876 8452 25728 8480
rect 21876 8440 21882 8452
rect 12894 8372 12900 8424
rect 12952 8412 12958 8424
rect 13265 8415 13323 8421
rect 13265 8412 13277 8415
rect 12952 8384 13277 8412
rect 12952 8372 12958 8384
rect 13265 8381 13277 8384
rect 13311 8381 13323 8415
rect 14734 8412 14740 8424
rect 14695 8384 14740 8412
rect 13265 8375 13323 8381
rect 14734 8372 14740 8384
rect 14792 8372 14798 8424
rect 16206 8412 16212 8424
rect 16167 8384 16212 8412
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 16390 8412 16396 8424
rect 16351 8384 16396 8412
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 24121 8415 24179 8421
rect 24121 8381 24133 8415
rect 24167 8412 24179 8415
rect 24762 8412 24768 8424
rect 24167 8384 24768 8412
rect 24167 8381 24179 8384
rect 24121 8375 24179 8381
rect 24762 8372 24768 8384
rect 24820 8372 24826 8424
rect 25700 8421 25728 8452
rect 26329 8449 26341 8483
rect 26375 8480 26387 8483
rect 26602 8480 26608 8492
rect 26375 8452 26608 8480
rect 26375 8449 26387 8452
rect 26329 8443 26387 8449
rect 26602 8440 26608 8452
rect 26660 8440 26666 8492
rect 26712 8489 26740 8520
rect 26697 8483 26755 8489
rect 26697 8449 26709 8483
rect 26743 8480 26755 8483
rect 27154 8480 27160 8492
rect 26743 8452 27160 8480
rect 26743 8449 26755 8452
rect 26697 8443 26755 8449
rect 27154 8440 27160 8452
rect 27212 8440 27218 8492
rect 27522 8480 27528 8492
rect 27483 8452 27528 8480
rect 27522 8440 27528 8452
rect 27580 8440 27586 8492
rect 27893 8483 27951 8489
rect 27893 8449 27905 8483
rect 27939 8480 27951 8483
rect 28166 8480 28172 8492
rect 27939 8452 28172 8480
rect 27939 8449 27951 8452
rect 27893 8443 27951 8449
rect 28166 8440 28172 8452
rect 28224 8440 28230 8492
rect 25685 8415 25743 8421
rect 25685 8381 25697 8415
rect 25731 8381 25743 8415
rect 25866 8412 25872 8424
rect 25827 8384 25872 8412
rect 25685 8375 25743 8381
rect 25866 8372 25872 8384
rect 25924 8372 25930 8424
rect 26234 8372 26240 8424
rect 26292 8412 26298 8424
rect 26789 8415 26847 8421
rect 26789 8412 26801 8415
rect 26292 8384 26801 8412
rect 26292 8372 26298 8384
rect 26789 8381 26801 8384
rect 26835 8412 26847 8415
rect 27430 8412 27436 8424
rect 26835 8384 27436 8412
rect 26835 8381 26847 8384
rect 26789 8375 26847 8381
rect 27430 8372 27436 8384
rect 27488 8372 27494 8424
rect 27985 8415 28043 8421
rect 27985 8381 27997 8415
rect 28031 8412 28043 8415
rect 28258 8412 28264 8424
rect 28031 8384 28264 8412
rect 28031 8381 28043 8384
rect 27985 8375 28043 8381
rect 28258 8372 28264 8384
rect 28316 8372 28322 8424
rect 2372 8316 12020 8344
rect 2372 8304 2378 8316
rect 12066 8304 12072 8356
rect 12124 8344 12130 8356
rect 12207 8347 12265 8353
rect 12207 8344 12219 8347
rect 12124 8316 12219 8344
rect 12124 8304 12130 8316
rect 12207 8313 12219 8316
rect 12253 8313 12265 8347
rect 12342 8344 12348 8356
rect 12303 8316 12348 8344
rect 12207 8307 12265 8313
rect 12342 8304 12348 8316
rect 12400 8304 12406 8356
rect 15470 8344 15476 8356
rect 13740 8316 15476 8344
rect 13740 8288 13768 8316
rect 15470 8304 15476 8316
rect 15528 8304 15534 8356
rect 6546 8236 6552 8288
rect 6604 8276 6610 8288
rect 9306 8276 9312 8288
rect 6604 8248 9312 8276
rect 6604 8236 6610 8248
rect 9306 8236 9312 8248
rect 9364 8236 9370 8288
rect 9490 8276 9496 8288
rect 9451 8248 9496 8276
rect 9490 8236 9496 8248
rect 9548 8236 9554 8288
rect 9858 8276 9864 8288
rect 9819 8248 9864 8276
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 13722 8276 13728 8288
rect 10008 8248 13728 8276
rect 10008 8236 10014 8248
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 19886 8236 19892 8288
rect 19944 8276 19950 8288
rect 20162 8276 20168 8288
rect 19944 8248 20168 8276
rect 19944 8236 19950 8248
rect 20162 8236 20168 8248
rect 20220 8236 20226 8288
rect 25590 8236 25596 8288
rect 25648 8276 25654 8288
rect 26786 8276 26792 8288
rect 25648 8248 26792 8276
rect 25648 8236 25654 8248
rect 26786 8236 26792 8248
rect 26844 8236 26850 8288
rect 1104 8186 28888 8208
rect 1104 8134 10246 8186
rect 10298 8134 10310 8186
rect 10362 8134 10374 8186
rect 10426 8134 10438 8186
rect 10490 8134 19510 8186
rect 19562 8134 19574 8186
rect 19626 8134 19638 8186
rect 19690 8134 19702 8186
rect 19754 8134 28888 8186
rect 1104 8112 28888 8134
rect 1765 8075 1823 8081
rect 1765 8041 1777 8075
rect 1811 8072 1823 8075
rect 2682 8072 2688 8084
rect 1811 8044 2688 8072
rect 1811 8041 1823 8044
rect 1765 8035 1823 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 2958 8032 2964 8084
rect 3016 8072 3022 8084
rect 3237 8075 3295 8081
rect 3237 8072 3249 8075
rect 3016 8044 3249 8072
rect 3016 8032 3022 8044
rect 3237 8041 3249 8044
rect 3283 8041 3295 8075
rect 3237 8035 3295 8041
rect 4062 8032 4068 8084
rect 4120 8072 4126 8084
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 4120 8044 5181 8072
rect 4120 8032 4126 8044
rect 5169 8041 5181 8044
rect 5215 8041 5227 8075
rect 5169 8035 5227 8041
rect 6917 8075 6975 8081
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 8754 8072 8760 8084
rect 6963 8044 8760 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 9125 8075 9183 8081
rect 9125 8041 9137 8075
rect 9171 8072 9183 8075
rect 9490 8072 9496 8084
rect 9171 8044 9496 8072
rect 9171 8041 9183 8044
rect 9125 8035 9183 8041
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 12124 8044 12169 8072
rect 12124 8032 12130 8044
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 13078 8072 13084 8084
rect 12676 8044 13084 8072
rect 12676 8032 12682 8044
rect 13078 8032 13084 8044
rect 13136 8032 13142 8084
rect 14461 8075 14519 8081
rect 14461 8041 14473 8075
rect 14507 8072 14519 8075
rect 14734 8072 14740 8084
rect 14507 8044 14740 8072
rect 14507 8041 14519 8044
rect 14461 8035 14519 8041
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 15657 8075 15715 8081
rect 15657 8041 15669 8075
rect 15703 8072 15715 8075
rect 16022 8072 16028 8084
rect 15703 8044 16028 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 16022 8032 16028 8044
rect 16080 8032 16086 8084
rect 16117 8075 16175 8081
rect 16117 8041 16129 8075
rect 16163 8072 16175 8075
rect 16666 8072 16672 8084
rect 16163 8044 16672 8072
rect 16163 8041 16175 8044
rect 16117 8035 16175 8041
rect 16666 8032 16672 8044
rect 16724 8072 16730 8084
rect 16850 8072 16856 8084
rect 16724 8044 16856 8072
rect 16724 8032 16730 8044
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 17218 8072 17224 8084
rect 16960 8044 17224 8072
rect 4246 8004 4252 8016
rect 4207 7976 4252 8004
rect 4246 7964 4252 7976
rect 4304 7964 4310 8016
rect 5261 8007 5319 8013
rect 5261 7973 5273 8007
rect 5307 8004 5319 8007
rect 5902 8004 5908 8016
rect 5307 7976 5908 8004
rect 5307 7973 5319 7976
rect 5261 7967 5319 7973
rect 5902 7964 5908 7976
rect 5960 7964 5966 8016
rect 8021 8007 8079 8013
rect 8021 7973 8033 8007
rect 8067 8004 8079 8007
rect 8941 8007 8999 8013
rect 8941 8004 8953 8007
rect 8067 7976 8953 8004
rect 8067 7973 8079 7976
rect 8021 7967 8079 7973
rect 8941 7973 8953 7976
rect 8987 7973 8999 8007
rect 8941 7967 8999 7973
rect 9306 7964 9312 8016
rect 9364 8004 9370 8016
rect 10226 8004 10232 8016
rect 9364 7976 10232 8004
rect 9364 7964 9370 7976
rect 10226 7964 10232 7976
rect 10284 7964 10290 8016
rect 10410 8004 10416 8016
rect 10371 7976 10416 8004
rect 10410 7964 10416 7976
rect 10468 7964 10474 8016
rect 14829 8007 14887 8013
rect 14829 8004 14841 8007
rect 10520 7976 14841 8004
rect 1486 7896 1492 7948
rect 1544 7936 1550 7948
rect 1949 7939 2007 7945
rect 1949 7936 1961 7939
rect 1544 7908 1961 7936
rect 1544 7896 1550 7908
rect 1949 7905 1961 7908
rect 1995 7905 2007 7939
rect 2406 7936 2412 7948
rect 2367 7908 2412 7936
rect 1949 7899 2007 7905
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 2866 7896 2872 7948
rect 2924 7936 2930 7948
rect 3053 7939 3111 7945
rect 3053 7936 3065 7939
rect 2924 7908 3065 7936
rect 2924 7896 2930 7908
rect 3053 7905 3065 7908
rect 3099 7905 3111 7939
rect 3053 7899 3111 7905
rect 4157 7939 4215 7945
rect 4157 7905 4169 7939
rect 4203 7936 4215 7939
rect 6822 7936 6828 7948
rect 4203 7908 4844 7936
rect 4203 7905 4215 7908
rect 4157 7899 4215 7905
rect 4816 7809 4844 7908
rect 5184 7908 5488 7936
rect 6783 7908 6828 7936
rect 2593 7803 2651 7809
rect 2593 7769 2605 7803
rect 2639 7800 2651 7803
rect 4801 7803 4859 7809
rect 2639 7772 2774 7800
rect 2639 7769 2651 7772
rect 2593 7763 2651 7769
rect 2746 7732 2774 7772
rect 4801 7769 4813 7803
rect 4847 7769 4859 7803
rect 4801 7763 4859 7769
rect 5184 7732 5212 7908
rect 5353 7871 5411 7877
rect 5353 7837 5365 7871
rect 5399 7837 5411 7871
rect 5460 7868 5488 7908
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 7926 7936 7932 7948
rect 7887 7908 7932 7936
rect 7926 7896 7932 7908
rect 7984 7896 7990 7948
rect 8110 7936 8116 7948
rect 8071 7908 8116 7936
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 10520 7936 10548 7976
rect 14829 7973 14841 7976
rect 14875 7973 14887 8007
rect 14829 7967 14887 7973
rect 14921 8007 14979 8013
rect 14921 7973 14933 8007
rect 14967 8004 14979 8007
rect 16960 8004 16988 8044
rect 17218 8032 17224 8044
rect 17276 8072 17282 8084
rect 17276 8044 18644 8072
rect 17276 8032 17282 8044
rect 14967 7976 16988 8004
rect 14967 7973 14979 7976
rect 14921 7967 14979 7973
rect 17034 7964 17040 8016
rect 17092 8004 17098 8016
rect 17865 8007 17923 8013
rect 17865 8004 17877 8007
rect 17092 7976 17877 8004
rect 17092 7964 17098 7976
rect 17865 7973 17877 7976
rect 17911 7973 17923 8007
rect 17865 7967 17923 7973
rect 17957 8007 18015 8013
rect 17957 7973 17969 8007
rect 18003 8004 18015 8007
rect 18506 8004 18512 8016
rect 18003 7976 18512 8004
rect 18003 7973 18015 7976
rect 17957 7967 18015 7973
rect 18506 7964 18512 7976
rect 18564 7964 18570 8016
rect 18616 8004 18644 8044
rect 18690 8032 18696 8084
rect 18748 8072 18754 8084
rect 18748 8044 28028 8072
rect 18748 8032 18754 8044
rect 25958 8004 25964 8016
rect 18616 7976 25728 8004
rect 25919 7976 25964 8004
rect 8220 7908 10548 7936
rect 8220 7868 8248 7908
rect 10686 7896 10692 7948
rect 10744 7936 10750 7948
rect 12437 7939 12495 7945
rect 12437 7936 12449 7939
rect 10744 7908 12449 7936
rect 10744 7896 10750 7908
rect 12437 7905 12449 7908
rect 12483 7905 12495 7939
rect 12437 7899 12495 7905
rect 12526 7896 12532 7948
rect 12584 7936 12590 7948
rect 16022 7936 16028 7948
rect 12584 7908 12629 7936
rect 15983 7908 16028 7936
rect 12584 7896 12590 7908
rect 16022 7896 16028 7908
rect 16080 7896 16086 7948
rect 18690 7936 18696 7948
rect 18651 7908 18696 7936
rect 18690 7896 18696 7908
rect 18748 7896 18754 7948
rect 19334 7936 19340 7948
rect 19247 7908 19340 7936
rect 19334 7896 19340 7908
rect 19392 7936 19398 7948
rect 19886 7936 19892 7948
rect 19392 7908 19892 7936
rect 19392 7896 19398 7908
rect 19886 7896 19892 7908
rect 19944 7896 19950 7948
rect 20714 7936 20720 7948
rect 20675 7908 20720 7936
rect 20714 7896 20720 7908
rect 20772 7936 20778 7948
rect 21082 7936 21088 7948
rect 20772 7908 21088 7936
rect 20772 7896 20778 7908
rect 21082 7896 21088 7908
rect 21140 7896 21146 7948
rect 22922 7936 22928 7948
rect 22883 7908 22928 7936
rect 22922 7896 22928 7908
rect 22980 7896 22986 7948
rect 23382 7896 23388 7948
rect 23440 7936 23446 7948
rect 23937 7939 23995 7945
rect 23937 7936 23949 7939
rect 23440 7908 23949 7936
rect 23440 7896 23446 7908
rect 23937 7905 23949 7908
rect 23983 7905 23995 7939
rect 23937 7899 23995 7905
rect 25225 7939 25283 7945
rect 25225 7905 25237 7939
rect 25271 7936 25283 7939
rect 25590 7936 25596 7948
rect 25271 7908 25596 7936
rect 25271 7905 25283 7908
rect 25225 7899 25283 7905
rect 25590 7896 25596 7908
rect 25648 7896 25654 7948
rect 25700 7936 25728 7976
rect 25958 7964 25964 7976
rect 26016 7964 26022 8016
rect 26142 8004 26148 8016
rect 26103 7976 26148 8004
rect 26142 7964 26148 7976
rect 26200 7964 26206 8016
rect 28000 8013 28028 8044
rect 27985 8007 28043 8013
rect 27985 7973 27997 8007
rect 28031 7973 28043 8007
rect 27985 7967 28043 7973
rect 26697 7939 26755 7945
rect 26697 7936 26709 7939
rect 25700 7908 26709 7936
rect 26697 7905 26709 7908
rect 26743 7905 26755 7939
rect 26697 7899 26755 7905
rect 5460 7840 8248 7868
rect 9217 7871 9275 7877
rect 5353 7831 5411 7837
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9398 7868 9404 7880
rect 9263 7840 9404 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 2746 7704 5212 7732
rect 5368 7732 5396 7831
rect 9398 7828 9404 7840
rect 9456 7868 9462 7880
rect 10318 7868 10324 7880
rect 9456 7840 10180 7868
rect 10279 7840 10324 7868
rect 9456 7828 9462 7840
rect 5534 7760 5540 7812
rect 5592 7800 5598 7812
rect 10152 7800 10180 7840
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7868 12771 7871
rect 13078 7868 13084 7880
rect 12759 7840 13084 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 10520 7800 10548 7831
rect 13078 7828 13084 7840
rect 13136 7828 13142 7880
rect 14274 7828 14280 7880
rect 14332 7868 14338 7880
rect 15013 7871 15071 7877
rect 15013 7868 15025 7871
rect 14332 7840 15025 7868
rect 14332 7828 14338 7840
rect 15013 7837 15025 7840
rect 15059 7868 15071 7871
rect 16209 7871 16267 7877
rect 16209 7868 16221 7871
rect 15059 7840 16221 7868
rect 15059 7837 15071 7840
rect 15013 7831 15071 7837
rect 16209 7837 16221 7840
rect 16255 7868 16267 7871
rect 16482 7868 16488 7880
rect 16255 7840 16488 7868
rect 16255 7837 16267 7840
rect 16209 7831 16267 7837
rect 16482 7828 16488 7840
rect 16540 7828 16546 7880
rect 17770 7868 17776 7880
rect 17731 7840 17776 7868
rect 17770 7828 17776 7840
rect 17828 7828 17834 7880
rect 18966 7828 18972 7880
rect 19024 7868 19030 7880
rect 23014 7868 23020 7880
rect 19024 7840 22094 7868
rect 22975 7840 23020 7868
rect 19024 7828 19030 7840
rect 15562 7800 15568 7812
rect 5592 7772 10088 7800
rect 10152 7772 10548 7800
rect 10704 7772 15568 7800
rect 5592 7760 5598 7772
rect 6270 7732 6276 7744
rect 5368 7704 6276 7732
rect 6270 7692 6276 7704
rect 6328 7732 6334 7744
rect 7374 7732 7380 7744
rect 6328 7704 7380 7732
rect 6328 7692 6334 7704
rect 7374 7692 7380 7704
rect 7432 7692 7438 7744
rect 8202 7692 8208 7744
rect 8260 7732 8266 7744
rect 8665 7735 8723 7741
rect 8665 7732 8677 7735
rect 8260 7704 8677 7732
rect 8260 7692 8266 7704
rect 8665 7701 8677 7704
rect 8711 7701 8723 7735
rect 8665 7695 8723 7701
rect 9674 7692 9680 7744
rect 9732 7732 9738 7744
rect 9953 7735 10011 7741
rect 9953 7732 9965 7735
rect 9732 7704 9965 7732
rect 9732 7692 9738 7704
rect 9953 7701 9965 7704
rect 9999 7701 10011 7735
rect 10060 7732 10088 7772
rect 10704 7732 10732 7772
rect 15562 7760 15568 7772
rect 15620 7760 15626 7812
rect 17405 7803 17463 7809
rect 17405 7769 17417 7803
rect 17451 7800 17463 7803
rect 17862 7800 17868 7812
rect 17451 7772 17868 7800
rect 17451 7769 17463 7772
rect 17405 7763 17463 7769
rect 17862 7760 17868 7772
rect 17920 7760 17926 7812
rect 20901 7803 20959 7809
rect 20901 7769 20913 7803
rect 20947 7800 20959 7803
rect 20990 7800 20996 7812
rect 20947 7772 20996 7800
rect 20947 7769 20959 7772
rect 20901 7763 20959 7769
rect 20990 7760 20996 7772
rect 21048 7760 21054 7812
rect 22066 7800 22094 7840
rect 23014 7828 23020 7840
rect 23072 7828 23078 7880
rect 23106 7828 23112 7880
rect 23164 7868 23170 7880
rect 23842 7868 23848 7880
rect 23164 7840 23209 7868
rect 23803 7840 23848 7868
rect 23164 7828 23170 7840
rect 23842 7828 23848 7840
rect 23900 7828 23906 7880
rect 28350 7868 28356 7880
rect 26206 7840 28356 7868
rect 22462 7800 22468 7812
rect 22066 7772 22468 7800
rect 22462 7760 22468 7772
rect 22520 7760 22526 7812
rect 25317 7803 25375 7809
rect 25317 7769 25329 7803
rect 25363 7800 25375 7803
rect 26206 7800 26234 7840
rect 28350 7828 28356 7840
rect 28408 7828 28414 7880
rect 28166 7800 28172 7812
rect 25363 7772 26234 7800
rect 28127 7772 28172 7800
rect 25363 7769 25375 7772
rect 25317 7763 25375 7769
rect 28166 7760 28172 7772
rect 28224 7760 28230 7812
rect 10060 7704 10732 7732
rect 9953 7695 10011 7701
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 18690 7732 18696 7744
rect 10836 7704 18696 7732
rect 10836 7692 10842 7704
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 18785 7735 18843 7741
rect 18785 7701 18797 7735
rect 18831 7732 18843 7735
rect 18874 7732 18880 7744
rect 18831 7704 18880 7732
rect 18831 7701 18843 7704
rect 18785 7695 18843 7701
rect 18874 7692 18880 7704
rect 18932 7692 18938 7744
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 19429 7735 19487 7741
rect 19429 7732 19441 7735
rect 19392 7704 19441 7732
rect 19392 7692 19398 7704
rect 19429 7701 19441 7704
rect 19475 7701 19487 7735
rect 22554 7732 22560 7744
rect 22515 7704 22560 7732
rect 19429 7695 19487 7701
rect 22554 7692 22560 7704
rect 22612 7692 22618 7744
rect 24213 7735 24271 7741
rect 24213 7701 24225 7735
rect 24259 7732 24271 7735
rect 25958 7732 25964 7744
rect 24259 7704 25964 7732
rect 24259 7701 24271 7704
rect 24213 7695 24271 7701
rect 25958 7692 25964 7704
rect 26016 7692 26022 7744
rect 26786 7732 26792 7744
rect 26747 7704 26792 7732
rect 26786 7692 26792 7704
rect 26844 7692 26850 7744
rect 1104 7642 28888 7664
rect 1104 7590 5614 7642
rect 5666 7590 5678 7642
rect 5730 7590 5742 7642
rect 5794 7590 5806 7642
rect 5858 7590 14878 7642
rect 14930 7590 14942 7642
rect 14994 7590 15006 7642
rect 15058 7590 15070 7642
rect 15122 7590 24142 7642
rect 24194 7590 24206 7642
rect 24258 7590 24270 7642
rect 24322 7590 24334 7642
rect 24386 7590 28888 7642
rect 1104 7568 28888 7590
rect 4985 7531 5043 7537
rect 4985 7497 4997 7531
rect 5031 7528 5043 7531
rect 6822 7528 6828 7540
rect 5031 7500 6828 7528
rect 5031 7497 5043 7500
rect 4985 7491 5043 7497
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7926 7488 7932 7540
rect 7984 7528 7990 7540
rect 8386 7528 8392 7540
rect 7984 7500 8392 7528
rect 7984 7488 7990 7500
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 9585 7531 9643 7537
rect 9585 7497 9597 7531
rect 9631 7528 9643 7531
rect 9858 7528 9864 7540
rect 9631 7500 9864 7528
rect 9631 7497 9643 7500
rect 9585 7491 9643 7497
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 10410 7528 10416 7540
rect 10371 7500 10416 7528
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 13633 7531 13691 7537
rect 13633 7497 13645 7531
rect 13679 7528 13691 7531
rect 13998 7528 14004 7540
rect 13679 7500 14004 7528
rect 13679 7497 13691 7500
rect 13633 7491 13691 7497
rect 13998 7488 14004 7500
rect 14056 7488 14062 7540
rect 14185 7531 14243 7537
rect 14185 7497 14197 7531
rect 14231 7528 14243 7531
rect 15841 7531 15899 7537
rect 15841 7528 15853 7531
rect 14231 7500 15853 7528
rect 14231 7497 14243 7500
rect 14185 7491 14243 7497
rect 15841 7497 15853 7500
rect 15887 7497 15899 7531
rect 15841 7491 15899 7497
rect 15933 7531 15991 7537
rect 15933 7497 15945 7531
rect 15979 7528 15991 7531
rect 16206 7528 16212 7540
rect 15979 7500 16212 7528
rect 15979 7497 15991 7500
rect 15933 7491 15991 7497
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 18506 7528 18512 7540
rect 18467 7500 18512 7528
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 20625 7531 20683 7537
rect 20625 7497 20637 7531
rect 20671 7528 20683 7531
rect 20806 7528 20812 7540
rect 20671 7500 20812 7528
rect 20671 7497 20683 7500
rect 20625 7491 20683 7497
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 22649 7531 22707 7537
rect 22649 7497 22661 7531
rect 22695 7528 22707 7531
rect 23382 7528 23388 7540
rect 22695 7500 23388 7528
rect 22695 7497 22707 7500
rect 22649 7491 22707 7497
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 1673 7463 1731 7469
rect 1673 7429 1685 7463
rect 1719 7460 1731 7463
rect 5350 7460 5356 7472
rect 1719 7432 5356 7460
rect 1719 7429 1731 7432
rect 1673 7423 1731 7429
rect 5350 7420 5356 7432
rect 5408 7420 5414 7472
rect 11606 7460 11612 7472
rect 5460 7432 11612 7460
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 5460 7392 5488 7432
rect 11606 7420 11612 7432
rect 11664 7420 11670 7472
rect 15746 7460 15752 7472
rect 15212 7432 15752 7460
rect 2363 7364 5488 7392
rect 5629 7395 5687 7401
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 5629 7361 5641 7395
rect 5675 7392 5687 7395
rect 5810 7392 5816 7404
rect 5675 7364 5816 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 5810 7352 5816 7364
rect 5868 7392 5874 7404
rect 5994 7392 6000 7404
rect 5868 7364 6000 7392
rect 5868 7352 5874 7364
rect 5994 7352 6000 7364
rect 6052 7392 6058 7404
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 6052 7364 7297 7392
rect 6052 7352 6058 7364
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 10778 7392 10784 7404
rect 7285 7355 7343 7361
rect 7392 7364 10784 7392
rect 1581 7327 1639 7333
rect 1581 7293 1593 7327
rect 1627 7324 1639 7327
rect 1854 7324 1860 7336
rect 1627 7296 1860 7324
rect 1627 7293 1639 7296
rect 1581 7287 1639 7293
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7293 2283 7327
rect 3050 7324 3056 7336
rect 3011 7296 3056 7324
rect 2225 7287 2283 7293
rect 2240 7256 2268 7287
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 5258 7284 5264 7336
rect 5316 7324 5322 7336
rect 5445 7327 5503 7333
rect 5445 7324 5457 7327
rect 5316 7296 5457 7324
rect 5316 7284 5322 7296
rect 5445 7293 5457 7296
rect 5491 7293 5503 7327
rect 5445 7287 5503 7293
rect 5902 7284 5908 7336
rect 5960 7324 5966 7336
rect 6638 7324 6644 7336
rect 5960 7296 6644 7324
rect 5960 7284 5966 7296
rect 6638 7284 6644 7296
rect 6696 7324 6702 7336
rect 7392 7324 7420 7364
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 10962 7392 10968 7404
rect 10923 7364 10968 7392
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 14185 7395 14243 7401
rect 14185 7392 14197 7395
rect 11072 7364 14197 7392
rect 9490 7324 9496 7336
rect 6696 7296 7420 7324
rect 9451 7296 9496 7324
rect 6696 7284 6702 7296
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 11072 7324 11100 7364
rect 14185 7361 14197 7364
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 11606 7324 11612 7336
rect 9600 7296 11100 7324
rect 11567 7296 11612 7324
rect 5353 7259 5411 7265
rect 5353 7256 5365 7259
rect 1596 7228 2268 7256
rect 2884 7228 5365 7256
rect 1596 7200 1624 7228
rect 1578 7148 1584 7200
rect 1636 7148 1642 7200
rect 2884 7197 2912 7228
rect 5353 7225 5365 7228
rect 5399 7225 5411 7259
rect 5353 7219 5411 7225
rect 5534 7216 5540 7268
rect 5592 7256 5598 7268
rect 7101 7259 7159 7265
rect 7101 7256 7113 7259
rect 5592 7228 7113 7256
rect 5592 7216 5598 7228
rect 7101 7225 7113 7228
rect 7147 7256 7159 7259
rect 9600 7256 9628 7296
rect 11606 7284 11612 7296
rect 11664 7284 11670 7336
rect 13446 7324 13452 7336
rect 13407 7296 13452 7324
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 15010 7324 15016 7336
rect 14971 7296 15016 7324
rect 15010 7284 15016 7296
rect 15068 7284 15074 7336
rect 15212 7333 15240 7432
rect 15746 7420 15752 7432
rect 15804 7420 15810 7472
rect 16482 7392 16488 7404
rect 16443 7364 16488 7392
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 17126 7392 17132 7404
rect 17087 7364 17132 7392
rect 17126 7352 17132 7364
rect 17184 7352 17190 7404
rect 22094 7352 22100 7404
rect 22152 7352 22158 7404
rect 28077 7395 28135 7401
rect 28077 7361 28089 7395
rect 28123 7392 28135 7395
rect 28350 7392 28356 7404
rect 28123 7364 28356 7392
rect 28123 7361 28135 7364
rect 28077 7355 28135 7361
rect 28350 7352 28356 7364
rect 28408 7352 28414 7404
rect 15102 7327 15160 7333
rect 15102 7293 15114 7327
rect 15148 7293 15160 7327
rect 15102 7287 15160 7293
rect 15197 7327 15255 7333
rect 15197 7293 15209 7327
rect 15243 7293 15255 7327
rect 15197 7287 15255 7293
rect 7147 7228 9628 7256
rect 10781 7259 10839 7265
rect 7147 7225 7159 7228
rect 7101 7219 7159 7225
rect 10781 7225 10793 7259
rect 10827 7256 10839 7259
rect 11701 7259 11759 7265
rect 11701 7256 11713 7259
rect 10827 7228 11713 7256
rect 10827 7225 10839 7228
rect 10781 7219 10839 7225
rect 11701 7225 11713 7228
rect 11747 7225 11759 7259
rect 11701 7219 11759 7225
rect 2869 7191 2927 7197
rect 2869 7157 2881 7191
rect 2915 7157 2927 7191
rect 6730 7188 6736 7200
rect 6691 7160 6736 7188
rect 2869 7151 2927 7157
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 7374 7148 7380 7200
rect 7432 7188 7438 7200
rect 9950 7188 9956 7200
rect 7432 7160 9956 7188
rect 7432 7148 7438 7160
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 10873 7191 10931 7197
rect 10873 7157 10885 7191
rect 10919 7188 10931 7191
rect 11330 7188 11336 7200
rect 10919 7160 11336 7188
rect 10919 7157 10931 7160
rect 10873 7151 10931 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 14734 7188 14740 7200
rect 14695 7160 14740 7188
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 14826 7148 14832 7200
rect 14884 7188 14890 7200
rect 15120 7188 15148 7287
rect 15378 7284 15384 7336
rect 15436 7324 15442 7336
rect 20530 7324 20536 7336
rect 15436 7296 15481 7324
rect 20491 7296 20536 7324
rect 15436 7284 15442 7296
rect 20530 7284 20536 7296
rect 20588 7284 20594 7336
rect 20898 7284 20904 7336
rect 20956 7324 20962 7336
rect 21637 7327 21695 7333
rect 21637 7324 21649 7327
rect 20956 7296 21649 7324
rect 20956 7284 20962 7296
rect 21637 7293 21649 7296
rect 21683 7293 21695 7327
rect 21637 7287 21695 7293
rect 21729 7327 21787 7333
rect 21729 7293 21741 7327
rect 21775 7324 21787 7327
rect 22278 7324 22284 7336
rect 21775 7296 22284 7324
rect 21775 7293 21787 7296
rect 21729 7287 21787 7293
rect 22278 7284 22284 7296
rect 22336 7284 22342 7336
rect 24213 7327 24271 7333
rect 24213 7293 24225 7327
rect 24259 7324 24271 7327
rect 24486 7324 24492 7336
rect 24259 7296 24492 7324
rect 24259 7293 24271 7296
rect 24213 7287 24271 7293
rect 24486 7284 24492 7296
rect 24544 7284 24550 7336
rect 25317 7327 25375 7333
rect 25317 7293 25329 7327
rect 25363 7324 25375 7327
rect 25406 7324 25412 7336
rect 25363 7296 25412 7324
rect 25363 7293 25375 7296
rect 25317 7287 25375 7293
rect 25406 7284 25412 7296
rect 25464 7284 25470 7336
rect 15841 7259 15899 7265
rect 15841 7225 15853 7259
rect 15887 7256 15899 7259
rect 15887 7228 16436 7256
rect 15887 7225 15899 7228
rect 15841 7219 15899 7225
rect 14884 7160 15148 7188
rect 14884 7148 14890 7160
rect 15470 7148 15476 7200
rect 15528 7188 15534 7200
rect 16408 7197 16436 7228
rect 17310 7216 17316 7268
rect 17368 7265 17374 7268
rect 17368 7259 17432 7265
rect 17368 7225 17386 7259
rect 17420 7225 17432 7259
rect 17368 7219 17432 7225
rect 17368 7216 17374 7219
rect 19334 7216 19340 7268
rect 19392 7256 19398 7268
rect 21361 7259 21419 7265
rect 21361 7256 21373 7259
rect 19392 7228 21373 7256
rect 19392 7216 19398 7228
rect 21361 7225 21373 7228
rect 21407 7225 21419 7259
rect 21361 7219 21419 7225
rect 22097 7259 22155 7265
rect 22097 7225 22109 7259
rect 22143 7256 22155 7259
rect 23106 7256 23112 7268
rect 22143 7228 23112 7256
rect 22143 7225 22155 7228
rect 22097 7219 22155 7225
rect 23106 7216 23112 7228
rect 23164 7216 23170 7268
rect 25584 7259 25642 7265
rect 25584 7225 25596 7259
rect 25630 7256 25642 7259
rect 25682 7256 25688 7268
rect 25630 7228 25688 7256
rect 25630 7225 25642 7228
rect 25584 7219 25642 7225
rect 25682 7216 25688 7228
rect 25740 7216 25746 7268
rect 16301 7191 16359 7197
rect 16301 7188 16313 7191
rect 15528 7160 16313 7188
rect 15528 7148 15534 7160
rect 16301 7157 16313 7160
rect 16347 7157 16359 7191
rect 16301 7151 16359 7157
rect 16393 7191 16451 7197
rect 16393 7157 16405 7191
rect 16439 7188 16451 7191
rect 20070 7188 20076 7200
rect 16439 7160 20076 7188
rect 16439 7157 16451 7160
rect 16393 7151 16451 7157
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 22462 7188 22468 7200
rect 22423 7160 22468 7188
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 23934 7188 23940 7200
rect 23895 7160 23940 7188
rect 23934 7148 23940 7160
rect 23992 7148 23998 7200
rect 26142 7148 26148 7200
rect 26200 7188 26206 7200
rect 26697 7191 26755 7197
rect 26697 7188 26709 7191
rect 26200 7160 26709 7188
rect 26200 7148 26206 7160
rect 26697 7157 26709 7160
rect 26743 7157 26755 7191
rect 27430 7188 27436 7200
rect 27391 7160 27436 7188
rect 26697 7151 26755 7157
rect 27430 7148 27436 7160
rect 27488 7148 27494 7200
rect 27522 7148 27528 7200
rect 27580 7188 27586 7200
rect 27801 7191 27859 7197
rect 27801 7188 27813 7191
rect 27580 7160 27813 7188
rect 27580 7148 27586 7160
rect 27801 7157 27813 7160
rect 27847 7157 27859 7191
rect 27801 7151 27859 7157
rect 27893 7191 27951 7197
rect 27893 7157 27905 7191
rect 27939 7188 27951 7191
rect 28074 7188 28080 7200
rect 27939 7160 28080 7188
rect 27939 7157 27951 7160
rect 27893 7151 27951 7157
rect 28074 7148 28080 7160
rect 28132 7148 28138 7200
rect 1104 7098 28888 7120
rect 1104 7046 10246 7098
rect 10298 7046 10310 7098
rect 10362 7046 10374 7098
rect 10426 7046 10438 7098
rect 10490 7046 19510 7098
rect 19562 7046 19574 7098
rect 19626 7046 19638 7098
rect 19690 7046 19702 7098
rect 19754 7046 28888 7098
rect 1104 7024 28888 7046
rect 2685 6987 2743 6993
rect 2685 6953 2697 6987
rect 2731 6953 2743 6987
rect 2685 6947 2743 6953
rect 1489 6851 1547 6857
rect 1489 6817 1501 6851
rect 1535 6848 1547 6851
rect 2130 6848 2136 6860
rect 1535 6820 2136 6848
rect 1535 6817 1547 6820
rect 1489 6811 1547 6817
rect 2130 6808 2136 6820
rect 2188 6808 2194 6860
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6848 2375 6851
rect 2498 6848 2504 6860
rect 2363 6820 2504 6848
rect 2363 6817 2375 6820
rect 2317 6811 2375 6817
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 2700 6848 2728 6947
rect 4522 6944 4528 6996
rect 4580 6984 4586 6996
rect 8662 6984 8668 6996
rect 4580 6956 8668 6984
rect 4580 6944 4586 6956
rect 8662 6944 8668 6956
rect 8720 6944 8726 6996
rect 8757 6987 8815 6993
rect 8757 6953 8769 6987
rect 8803 6984 8815 6987
rect 9490 6984 9496 6996
rect 8803 6956 9496 6984
rect 8803 6953 8815 6956
rect 8757 6947 8815 6953
rect 9490 6944 9496 6956
rect 9548 6984 9554 6996
rect 9585 6987 9643 6993
rect 9585 6984 9597 6987
rect 9548 6956 9597 6984
rect 9548 6944 9554 6956
rect 9585 6953 9597 6956
rect 9631 6953 9643 6987
rect 10594 6984 10600 6996
rect 10555 6956 10600 6984
rect 9585 6947 9643 6953
rect 10594 6944 10600 6956
rect 10652 6944 10658 6996
rect 11330 6944 11336 6996
rect 11388 6984 11394 6996
rect 15470 6984 15476 6996
rect 11388 6956 15476 6984
rect 11388 6944 11394 6956
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 15654 6984 15660 6996
rect 15615 6956 15660 6984
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 17310 6984 17316 6996
rect 17271 6956 17316 6984
rect 17310 6944 17316 6956
rect 17368 6944 17374 6996
rect 18506 6984 18512 6996
rect 17972 6956 18512 6984
rect 5537 6919 5595 6925
rect 5537 6885 5549 6919
rect 5583 6916 5595 6919
rect 5902 6916 5908 6928
rect 5583 6888 5908 6916
rect 5583 6885 5595 6888
rect 5537 6879 5595 6885
rect 5902 6876 5908 6888
rect 5960 6876 5966 6928
rect 8386 6876 8392 6928
rect 8444 6916 8450 6928
rect 9677 6919 9735 6925
rect 9677 6916 9689 6919
rect 8444 6888 9689 6916
rect 8444 6876 8450 6888
rect 9677 6885 9689 6888
rect 9723 6885 9735 6919
rect 9677 6879 9735 6885
rect 10134 6876 10140 6928
rect 10192 6916 10198 6928
rect 10192 6888 10640 6916
rect 10192 6876 10198 6888
rect 3145 6851 3203 6857
rect 3145 6848 3157 6851
rect 2700 6820 3157 6848
rect 3145 6817 3157 6820
rect 3191 6817 3203 6851
rect 3145 6811 3203 6817
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 3786 6848 3792 6860
rect 3292 6820 3792 6848
rect 3292 6808 3298 6820
rect 3786 6808 3792 6820
rect 3844 6808 3850 6860
rect 3970 6848 3976 6860
rect 3931 6820 3976 6848
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 4433 6851 4491 6857
rect 4433 6848 4445 6851
rect 4120 6820 4445 6848
rect 4120 6808 4126 6820
rect 4433 6817 4445 6820
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 5994 6848 6000 6860
rect 5675 6820 6000 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 5994 6808 6000 6820
rect 6052 6808 6058 6860
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7377 6851 7435 6857
rect 7377 6848 7389 6851
rect 6972 6820 7389 6848
rect 6972 6808 6978 6820
rect 7377 6817 7389 6820
rect 7423 6817 7435 6851
rect 7377 6811 7435 6817
rect 7644 6851 7702 6857
rect 7644 6817 7656 6851
rect 7690 6848 7702 6851
rect 7690 6820 9260 6848
rect 7690 6817 7702 6820
rect 7644 6811 7702 6817
rect 2222 6780 2228 6792
rect 2183 6752 2228 6780
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 5534 6780 5540 6792
rect 2332 6752 5540 6780
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 2332 6712 2360 6752
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 5810 6780 5816 6792
rect 5771 6752 5816 6780
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 9232 6721 9260 6820
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 10612 6857 10640 6888
rect 12618 6876 12624 6928
rect 12676 6916 12682 6928
rect 13630 6916 13636 6928
rect 12676 6888 13636 6916
rect 12676 6876 12682 6888
rect 13630 6876 13636 6888
rect 13688 6876 13694 6928
rect 14544 6919 14602 6925
rect 14544 6885 14556 6919
rect 14590 6916 14602 6919
rect 14734 6916 14740 6928
rect 14590 6888 14740 6916
rect 14590 6885 14602 6888
rect 14544 6879 14602 6885
rect 14734 6876 14740 6888
rect 14792 6876 14798 6928
rect 10413 6851 10471 6857
rect 10413 6848 10425 6851
rect 9916 6820 10425 6848
rect 9916 6808 9922 6820
rect 10413 6817 10425 6820
rect 10459 6817 10471 6851
rect 10413 6811 10471 6817
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 11882 6808 11888 6860
rect 11940 6848 11946 6860
rect 12253 6851 12311 6857
rect 12253 6848 12265 6851
rect 11940 6820 12265 6848
rect 11940 6808 11946 6820
rect 12253 6817 12265 6820
rect 12299 6848 12311 6851
rect 12802 6848 12808 6860
rect 12299 6820 12808 6848
rect 12299 6817 12311 6820
rect 12253 6811 12311 6817
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 13262 6848 13268 6860
rect 13223 6820 13268 6848
rect 13262 6808 13268 6820
rect 13320 6808 13326 6860
rect 14090 6808 14096 6860
rect 14148 6848 14154 6860
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 14148 6820 14289 6848
rect 14148 6808 14154 6820
rect 14277 6817 14289 6820
rect 14323 6817 14335 6851
rect 14277 6811 14335 6817
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6780 9827 6783
rect 10042 6780 10048 6792
rect 9815 6752 10048 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 10042 6740 10048 6752
rect 10100 6780 10106 6792
rect 10686 6780 10692 6792
rect 10100 6752 10692 6780
rect 10100 6740 10106 6752
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6749 13415 6783
rect 13357 6743 13415 6749
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6780 13599 6783
rect 13722 6780 13728 6792
rect 13587 6752 13728 6780
rect 13587 6749 13599 6752
rect 13541 6743 13599 6749
rect 1627 6684 2360 6712
rect 9217 6715 9275 6721
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 9217 6681 9229 6715
rect 9263 6681 9275 6715
rect 12894 6712 12900 6724
rect 12855 6684 12900 6712
rect 9217 6675 9275 6681
rect 12894 6672 12900 6684
rect 12952 6672 12958 6724
rect 13372 6712 13400 6743
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 13630 6712 13636 6724
rect 13372 6684 13636 6712
rect 13630 6672 13636 6684
rect 13688 6672 13694 6724
rect 3786 6644 3792 6656
rect 3747 6616 3792 6644
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 3878 6604 3884 6656
rect 3936 6644 3942 6656
rect 4617 6647 4675 6653
rect 4617 6644 4629 6647
rect 3936 6616 4629 6644
rect 3936 6604 3942 6616
rect 4617 6613 4629 6616
rect 4663 6613 4675 6647
rect 5166 6644 5172 6656
rect 5127 6616 5172 6644
rect 4617 6607 4675 6613
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 12345 6647 12403 6653
rect 12345 6613 12357 6647
rect 12391 6644 12403 6647
rect 13446 6644 13452 6656
rect 12391 6616 13452 6644
rect 12391 6613 12403 6616
rect 12345 6607 12403 6613
rect 13446 6604 13452 6616
rect 13504 6604 13510 6656
rect 15488 6644 15516 6944
rect 17972 6916 18000 6956
rect 18506 6944 18512 6956
rect 18564 6944 18570 6996
rect 19981 6987 20039 6993
rect 19981 6953 19993 6987
rect 20027 6953 20039 6987
rect 23106 6984 23112 6996
rect 23067 6956 23112 6984
rect 19981 6947 20039 6953
rect 17604 6888 18000 6916
rect 17604 6857 17632 6888
rect 18414 6876 18420 6928
rect 18472 6916 18478 6928
rect 18693 6919 18751 6925
rect 18693 6916 18705 6919
rect 18472 6888 18705 6916
rect 18472 6876 18478 6888
rect 18693 6885 18705 6888
rect 18739 6916 18751 6919
rect 18739 6888 19288 6916
rect 18739 6885 18751 6888
rect 18693 6879 18751 6885
rect 17589 6851 17647 6857
rect 17589 6817 17601 6851
rect 17635 6817 17647 6851
rect 17589 6811 17647 6817
rect 17681 6851 17739 6857
rect 17681 6817 17693 6851
rect 17727 6817 17739 6851
rect 17681 6811 17739 6817
rect 17773 6851 17831 6857
rect 17773 6817 17785 6851
rect 17819 6817 17831 6851
rect 17954 6848 17960 6860
rect 17915 6820 17960 6848
rect 17773 6811 17831 6817
rect 16574 6740 16580 6792
rect 16632 6780 16638 6792
rect 17696 6780 17724 6811
rect 16632 6752 17724 6780
rect 16632 6740 16638 6752
rect 17788 6712 17816 6811
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 18782 6848 18788 6860
rect 18156 6820 18788 6848
rect 18046 6712 18052 6724
rect 17788 6684 18052 6712
rect 18046 6672 18052 6684
rect 18104 6672 18110 6724
rect 18156 6644 18184 6820
rect 18782 6808 18788 6820
rect 18840 6848 18846 6860
rect 18969 6851 19027 6857
rect 18969 6848 18981 6851
rect 18840 6820 18981 6848
rect 18840 6808 18846 6820
rect 18969 6817 18981 6820
rect 19015 6817 19027 6851
rect 18969 6811 19027 6817
rect 19058 6808 19064 6860
rect 19116 6848 19122 6860
rect 19260 6848 19288 6888
rect 19334 6876 19340 6928
rect 19392 6916 19398 6928
rect 19429 6919 19487 6925
rect 19429 6916 19441 6919
rect 19392 6888 19441 6916
rect 19392 6876 19398 6888
rect 19429 6885 19441 6888
rect 19475 6885 19487 6919
rect 19794 6916 19800 6928
rect 19755 6888 19800 6916
rect 19429 6879 19487 6885
rect 19794 6876 19800 6888
rect 19852 6876 19858 6928
rect 19996 6848 20024 6947
rect 23106 6944 23112 6956
rect 23164 6984 23170 6996
rect 23845 6987 23903 6993
rect 23845 6984 23857 6987
rect 23164 6956 23857 6984
rect 23164 6944 23170 6956
rect 23845 6953 23857 6956
rect 23891 6953 23903 6987
rect 24949 6987 25007 6993
rect 24949 6984 24961 6987
rect 23845 6947 23903 6953
rect 23952 6956 24961 6984
rect 20070 6876 20076 6928
rect 20128 6916 20134 6928
rect 23952 6916 23980 6956
rect 24949 6953 24961 6956
rect 24995 6953 25007 6987
rect 25682 6984 25688 6996
rect 25643 6956 25688 6984
rect 24949 6947 25007 6953
rect 25682 6944 25688 6956
rect 25740 6944 25746 6996
rect 25958 6944 25964 6996
rect 26016 6984 26022 6996
rect 26053 6987 26111 6993
rect 26053 6984 26065 6987
rect 26016 6956 26065 6984
rect 26016 6944 26022 6956
rect 26053 6953 26065 6956
rect 26099 6953 26111 6987
rect 26053 6947 26111 6953
rect 24854 6916 24860 6928
rect 20128 6888 23980 6916
rect 24412 6888 24860 6916
rect 20128 6876 20134 6888
rect 20530 6848 20536 6860
rect 19116 6820 19161 6848
rect 19260 6820 19840 6848
rect 19996 6820 20536 6848
rect 19116 6808 19122 6820
rect 18598 6740 18604 6792
rect 18656 6740 18662 6792
rect 19812 6712 19840 6820
rect 20530 6808 20536 6820
rect 20588 6848 20594 6860
rect 20809 6851 20867 6857
rect 20809 6848 20821 6851
rect 20588 6820 20821 6848
rect 20588 6808 20594 6820
rect 20809 6817 20821 6820
rect 20855 6817 20867 6851
rect 23014 6848 23020 6860
rect 22975 6820 23020 6848
rect 20809 6811 20867 6817
rect 23014 6808 23020 6820
rect 23072 6808 23078 6860
rect 23934 6808 23940 6860
rect 23992 6848 23998 6860
rect 24121 6851 24179 6857
rect 24121 6848 24133 6851
rect 23992 6820 24133 6848
rect 23992 6808 23998 6820
rect 24121 6817 24133 6820
rect 24167 6817 24179 6851
rect 24121 6811 24179 6817
rect 24213 6851 24271 6857
rect 24213 6817 24225 6851
rect 24259 6848 24271 6851
rect 24412 6848 24440 6888
rect 24854 6876 24860 6888
rect 24912 6876 24918 6928
rect 24578 6848 24584 6860
rect 24259 6820 24440 6848
rect 24539 6820 24584 6848
rect 24259 6817 24271 6820
rect 24213 6811 24271 6817
rect 24578 6808 24584 6820
rect 24636 6808 24642 6860
rect 24670 6808 24676 6860
rect 24728 6848 24734 6860
rect 27985 6851 28043 6857
rect 27985 6848 27997 6851
rect 24728 6820 27997 6848
rect 24728 6808 24734 6820
rect 27985 6817 27997 6820
rect 28031 6817 28043 6851
rect 27985 6811 28043 6817
rect 20901 6783 20959 6789
rect 20901 6749 20913 6783
rect 20947 6780 20959 6783
rect 20990 6780 20996 6792
rect 20947 6752 20996 6780
rect 20947 6749 20959 6752
rect 20901 6743 20959 6749
rect 20990 6740 20996 6752
rect 21048 6740 21054 6792
rect 23566 6740 23572 6792
rect 23624 6780 23630 6792
rect 23624 6752 23690 6780
rect 23624 6740 23630 6752
rect 25866 6740 25872 6792
rect 25924 6780 25930 6792
rect 26142 6780 26148 6792
rect 25924 6752 26148 6780
rect 25924 6740 25930 6752
rect 26142 6740 26148 6752
rect 26200 6740 26206 6792
rect 26237 6783 26295 6789
rect 26237 6749 26249 6783
rect 26283 6749 26295 6783
rect 26237 6743 26295 6749
rect 21082 6712 21088 6724
rect 19812 6684 21088 6712
rect 21082 6672 21088 6684
rect 21140 6672 21146 6724
rect 21177 6715 21235 6721
rect 21177 6681 21189 6715
rect 21223 6712 21235 6715
rect 22922 6712 22928 6724
rect 21223 6684 22928 6712
rect 21223 6681 21235 6684
rect 21177 6675 21235 6681
rect 22922 6672 22928 6684
rect 22980 6672 22986 6724
rect 25038 6672 25044 6724
rect 25096 6712 25102 6724
rect 26252 6712 26280 6743
rect 28166 6712 28172 6724
rect 25096 6684 26280 6712
rect 28127 6684 28172 6712
rect 25096 6672 25102 6684
rect 28166 6672 28172 6684
rect 28224 6672 28230 6724
rect 25130 6644 25136 6656
rect 15488 6616 18184 6644
rect 25091 6616 25136 6644
rect 25130 6604 25136 6616
rect 25188 6604 25194 6656
rect 1104 6554 28888 6576
rect 1104 6502 5614 6554
rect 5666 6502 5678 6554
rect 5730 6502 5742 6554
rect 5794 6502 5806 6554
rect 5858 6502 14878 6554
rect 14930 6502 14942 6554
rect 14994 6502 15006 6554
rect 15058 6502 15070 6554
rect 15122 6502 24142 6554
rect 24194 6502 24206 6554
rect 24258 6502 24270 6554
rect 24322 6502 24334 6554
rect 24386 6502 28888 6554
rect 1104 6480 28888 6502
rect 2869 6443 2927 6449
rect 2869 6409 2881 6443
rect 2915 6440 2927 6443
rect 4154 6440 4160 6452
rect 2915 6412 4160 6440
rect 2915 6409 2927 6412
rect 2869 6403 2927 6409
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 11238 6440 11244 6452
rect 11199 6412 11244 6440
rect 11238 6400 11244 6412
rect 11296 6400 11302 6452
rect 11330 6400 11336 6452
rect 11388 6440 11394 6452
rect 12158 6440 12164 6452
rect 11388 6412 11433 6440
rect 12119 6412 12164 6440
rect 11388 6400 11394 6412
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 14921 6443 14979 6449
rect 14921 6409 14933 6443
rect 14967 6440 14979 6443
rect 15378 6440 15384 6452
rect 14967 6412 15384 6440
rect 14967 6409 14979 6412
rect 14921 6403 14979 6409
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 15746 6400 15752 6452
rect 15804 6440 15810 6452
rect 16025 6443 16083 6449
rect 16025 6440 16037 6443
rect 15804 6412 16037 6440
rect 15804 6400 15810 6412
rect 16025 6409 16037 6412
rect 16071 6440 16083 6443
rect 16206 6440 16212 6452
rect 16071 6412 16212 6440
rect 16071 6409 16083 6412
rect 16025 6403 16083 6409
rect 16206 6400 16212 6412
rect 16264 6400 16270 6452
rect 16482 6400 16488 6452
rect 16540 6440 16546 6452
rect 16761 6443 16819 6449
rect 16761 6440 16773 6443
rect 16540 6412 16773 6440
rect 16540 6400 16546 6412
rect 16761 6409 16773 6412
rect 16807 6440 16819 6443
rect 18598 6440 18604 6452
rect 16807 6412 18604 6440
rect 16807 6409 16819 6412
rect 16761 6403 16819 6409
rect 18598 6400 18604 6412
rect 18656 6400 18662 6452
rect 18782 6440 18788 6452
rect 18743 6412 18788 6440
rect 18782 6400 18788 6412
rect 18840 6400 18846 6452
rect 18892 6412 21036 6440
rect 6549 6375 6607 6381
rect 6549 6341 6561 6375
rect 6595 6372 6607 6375
rect 9858 6372 9864 6384
rect 6595 6344 9864 6372
rect 6595 6341 6607 6344
rect 6549 6335 6607 6341
rect 9858 6332 9864 6344
rect 9916 6332 9922 6384
rect 15838 6372 15844 6384
rect 9968 6344 12112 6372
rect 1400 6316 1452 6322
rect 3418 6264 3424 6316
rect 3476 6304 3482 6316
rect 3476 6276 4936 6304
rect 3476 6264 3482 6276
rect 1400 6258 1452 6264
rect 1854 6236 1860 6248
rect 1815 6208 1860 6236
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 1949 6239 2007 6245
rect 1949 6205 1961 6239
rect 1995 6236 2007 6239
rect 2038 6236 2044 6248
rect 1995 6208 2044 6236
rect 1995 6205 2007 6208
rect 1949 6199 2007 6205
rect 2038 6196 2044 6208
rect 2096 6196 2102 6248
rect 2130 6196 2136 6248
rect 2188 6236 2194 6248
rect 2317 6239 2375 6245
rect 2317 6236 2329 6239
rect 2188 6208 2329 6236
rect 2188 6196 2194 6208
rect 2317 6205 2329 6208
rect 2363 6236 2375 6239
rect 3878 6236 3884 6248
rect 2363 6208 3884 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 4154 6196 4160 6248
rect 4212 6236 4218 6248
rect 4908 6245 4936 6276
rect 5994 6264 6000 6316
rect 6052 6304 6058 6316
rect 9968 6304 9996 6344
rect 6052 6276 9996 6304
rect 6052 6264 6058 6276
rect 10962 6264 10968 6316
rect 11020 6304 11026 6316
rect 11241 6307 11299 6313
rect 11241 6304 11253 6307
rect 11020 6276 11253 6304
rect 11020 6264 11026 6276
rect 11241 6273 11253 6276
rect 11287 6273 11299 6307
rect 11241 6267 11299 6273
rect 4249 6239 4307 6245
rect 4249 6236 4261 6239
rect 4212 6208 4261 6236
rect 4212 6196 4218 6208
rect 4249 6205 4261 6208
rect 4295 6205 4307 6239
rect 4249 6199 4307 6205
rect 4893 6239 4951 6245
rect 4893 6205 4905 6239
rect 4939 6205 4951 6239
rect 4893 6199 4951 6205
rect 5166 6196 5172 6248
rect 5224 6236 5230 6248
rect 5813 6239 5871 6245
rect 5813 6236 5825 6239
rect 5224 6208 5825 6236
rect 5224 6196 5230 6208
rect 5813 6205 5825 6208
rect 5859 6205 5871 6239
rect 5813 6199 5871 6205
rect 7101 6239 7159 6245
rect 7101 6205 7113 6239
rect 7147 6236 7159 6239
rect 7834 6236 7840 6248
rect 7147 6208 7840 6236
rect 7147 6205 7159 6208
rect 7101 6199 7159 6205
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 11146 6196 11152 6248
rect 11204 6236 11210 6248
rect 12084 6245 12112 6344
rect 14844 6344 15844 6372
rect 12342 6264 12348 6316
rect 12400 6304 12406 6316
rect 13446 6304 13452 6316
rect 12400 6276 12848 6304
rect 13407 6276 13452 6304
rect 12400 6264 12406 6276
rect 11425 6239 11483 6245
rect 11425 6236 11437 6239
rect 11204 6208 11437 6236
rect 11204 6196 11210 6208
rect 11425 6205 11437 6208
rect 11471 6205 11483 6239
rect 11425 6199 11483 6205
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6236 12127 6239
rect 12250 6236 12256 6248
rect 12115 6208 12256 6236
rect 12115 6205 12127 6208
rect 12069 6199 12127 6205
rect 12250 6196 12256 6208
rect 12308 6196 12314 6248
rect 12710 6236 12716 6248
rect 12671 6208 12716 6236
rect 12710 6196 12716 6208
rect 12768 6196 12774 6248
rect 12820 6236 12848 6276
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 13541 6239 13599 6245
rect 13541 6236 13553 6239
rect 12820 6208 13553 6236
rect 13541 6205 13553 6208
rect 13587 6236 13599 6239
rect 14550 6236 14556 6248
rect 13587 6208 14556 6236
rect 13587 6205 13599 6208
rect 13541 6199 13599 6205
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 14844 6245 14872 6344
rect 15838 6332 15844 6344
rect 15896 6332 15902 6384
rect 17678 6332 17684 6384
rect 17736 6372 17742 6384
rect 18892 6372 18920 6412
rect 17736 6344 18920 6372
rect 17736 6332 17742 6344
rect 19794 6304 19800 6316
rect 15856 6276 19800 6304
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6205 14887 6239
rect 15010 6236 15016 6248
rect 14971 6208 15016 6236
rect 14829 6199 14887 6205
rect 15010 6196 15016 6208
rect 15068 6196 15074 6248
rect 1872 6168 1900 6196
rect 5905 6171 5963 6177
rect 1872 6140 4476 6168
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 1762 6060 1768 6112
rect 1820 6100 1826 6112
rect 4448 6109 4476 6140
rect 5905 6137 5917 6171
rect 5951 6168 5963 6171
rect 6825 6171 6883 6177
rect 6825 6168 6837 6171
rect 5951 6140 6837 6168
rect 5951 6137 5963 6140
rect 5905 6131 5963 6137
rect 6825 6137 6837 6140
rect 6871 6137 6883 6171
rect 11054 6168 11060 6180
rect 11015 6140 11060 6168
rect 6825 6131 6883 6137
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 15856 6168 15884 6276
rect 19794 6264 19800 6276
rect 19852 6264 19858 6316
rect 21008 6304 21036 6412
rect 21082 6400 21088 6452
rect 21140 6440 21146 6452
rect 23934 6440 23940 6452
rect 21140 6412 23940 6440
rect 21140 6400 21146 6412
rect 23934 6400 23940 6412
rect 23992 6400 23998 6452
rect 24213 6443 24271 6449
rect 24213 6409 24225 6443
rect 24259 6440 24271 6443
rect 24578 6440 24584 6452
rect 24259 6412 24584 6440
rect 24259 6409 24271 6412
rect 24213 6403 24271 6409
rect 24578 6400 24584 6412
rect 24636 6400 24642 6452
rect 26237 6443 26295 6449
rect 26237 6409 26249 6443
rect 26283 6440 26295 6443
rect 27522 6440 27528 6452
rect 26283 6412 27528 6440
rect 26283 6409 26295 6412
rect 26237 6403 26295 6409
rect 27522 6400 27528 6412
rect 27580 6400 27586 6452
rect 25498 6332 25504 6384
rect 25556 6372 25562 6384
rect 25958 6372 25964 6384
rect 25556 6344 25964 6372
rect 25556 6332 25562 6344
rect 25958 6332 25964 6344
rect 26016 6372 26022 6384
rect 26016 6344 26832 6372
rect 26016 6332 26022 6344
rect 24670 6304 24676 6316
rect 21008 6276 22140 6304
rect 15930 6196 15936 6248
rect 15988 6236 15994 6248
rect 16669 6239 16727 6245
rect 16669 6236 16681 6239
rect 15988 6208 16681 6236
rect 15988 6196 15994 6208
rect 16669 6205 16681 6208
rect 16715 6236 16727 6239
rect 17589 6239 17647 6245
rect 17589 6236 17601 6239
rect 16715 6208 17601 6236
rect 16715 6205 16727 6208
rect 16669 6199 16727 6205
rect 17589 6205 17601 6208
rect 17635 6205 17647 6239
rect 18690 6236 18696 6248
rect 18651 6208 18696 6236
rect 17589 6199 17647 6205
rect 18690 6196 18696 6208
rect 18748 6196 18754 6248
rect 19981 6239 20039 6245
rect 19981 6205 19993 6239
rect 20027 6236 20039 6239
rect 20070 6236 20076 6248
rect 20027 6208 20076 6236
rect 20027 6205 20039 6208
rect 19981 6199 20039 6205
rect 20070 6196 20076 6208
rect 20128 6196 20134 6248
rect 22005 6239 22063 6245
rect 22005 6205 22017 6239
rect 22051 6205 22063 6239
rect 22005 6199 22063 6205
rect 11164 6140 15884 6168
rect 2685 6103 2743 6109
rect 2685 6100 2697 6103
rect 1820 6072 2697 6100
rect 1820 6060 1826 6072
rect 2685 6069 2697 6072
rect 2731 6069 2743 6103
rect 2685 6063 2743 6069
rect 4433 6103 4491 6109
rect 4433 6069 4445 6103
rect 4479 6069 4491 6103
rect 4433 6063 4491 6069
rect 5077 6103 5135 6109
rect 5077 6069 5089 6103
rect 5123 6100 5135 6103
rect 5442 6100 5448 6112
rect 5123 6072 5448 6100
rect 5123 6069 5135 6072
rect 5077 6063 5135 6069
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 7009 6103 7067 6109
rect 7009 6100 7021 6103
rect 6788 6072 7021 6100
rect 6788 6060 6794 6072
rect 7009 6069 7021 6072
rect 7055 6069 7067 6103
rect 7009 6063 7067 6069
rect 7190 6060 7196 6112
rect 7248 6100 7254 6112
rect 11164 6100 11192 6140
rect 18322 6128 18328 6180
rect 18380 6168 18386 6180
rect 20226 6171 20284 6177
rect 20226 6168 20238 6171
rect 18380 6140 20238 6168
rect 18380 6128 18386 6140
rect 20226 6137 20238 6140
rect 20272 6137 20284 6171
rect 20226 6131 20284 6137
rect 7248 6072 11192 6100
rect 7248 6060 7254 6072
rect 12986 6060 12992 6112
rect 13044 6100 13050 6112
rect 13446 6100 13452 6112
rect 13044 6072 13452 6100
rect 13044 6060 13050 6072
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 13814 6100 13820 6112
rect 13775 6072 13820 6100
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 17681 6103 17739 6109
rect 17681 6069 17693 6103
rect 17727 6100 17739 6103
rect 18046 6100 18052 6112
rect 17727 6072 18052 6100
rect 17727 6069 17739 6072
rect 17681 6063 17739 6069
rect 18046 6060 18052 6072
rect 18104 6100 18110 6112
rect 18414 6100 18420 6112
rect 18104 6072 18420 6100
rect 18104 6060 18110 6072
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 21358 6100 21364 6112
rect 21319 6072 21364 6100
rect 21358 6060 21364 6072
rect 21416 6060 21422 6112
rect 22020 6100 22048 6199
rect 22112 6168 22140 6276
rect 23032 6276 24676 6304
rect 22272 6239 22330 6245
rect 22272 6205 22284 6239
rect 22318 6236 22330 6239
rect 22554 6236 22560 6248
rect 22318 6208 22560 6236
rect 22318 6205 22330 6208
rect 22272 6199 22330 6205
rect 22554 6196 22560 6208
rect 22612 6196 22618 6248
rect 23032 6168 23060 6276
rect 24670 6264 24676 6276
rect 24728 6264 24734 6316
rect 26053 6307 26111 6313
rect 26053 6273 26065 6307
rect 26099 6304 26111 6307
rect 26234 6304 26240 6316
rect 26099 6276 26240 6304
rect 26099 6273 26111 6276
rect 26053 6267 26111 6273
rect 26234 6264 26240 6276
rect 26292 6304 26298 6316
rect 26510 6304 26516 6316
rect 26292 6276 26516 6304
rect 26292 6264 26298 6276
rect 26510 6264 26516 6276
rect 26568 6264 26574 6316
rect 26804 6313 26832 6344
rect 26789 6307 26847 6313
rect 26789 6273 26801 6307
rect 26835 6273 26847 6307
rect 26789 6267 26847 6273
rect 24121 6239 24179 6245
rect 24121 6205 24133 6239
rect 24167 6205 24179 6239
rect 24121 6199 24179 6205
rect 22112 6140 23060 6168
rect 24136 6168 24164 6199
rect 24762 6196 24768 6248
rect 24820 6236 24826 6248
rect 25130 6236 25136 6248
rect 24820 6208 25136 6236
rect 24820 6196 24826 6208
rect 25130 6196 25136 6208
rect 25188 6236 25194 6248
rect 25961 6239 26019 6245
rect 25961 6236 25973 6239
rect 25188 6208 25973 6236
rect 25188 6196 25194 6208
rect 25961 6205 25973 6208
rect 26007 6205 26019 6239
rect 25961 6199 26019 6205
rect 27056 6239 27114 6245
rect 27056 6205 27068 6239
rect 27102 6236 27114 6239
rect 27430 6236 27436 6248
rect 27102 6208 27436 6236
rect 27102 6205 27114 6208
rect 27056 6199 27114 6205
rect 27430 6196 27436 6208
rect 27488 6196 27494 6248
rect 25866 6168 25872 6180
rect 24136 6140 25872 6168
rect 25866 6128 25872 6140
rect 25924 6128 25930 6180
rect 22738 6100 22744 6112
rect 22020 6072 22744 6100
rect 22738 6060 22744 6072
rect 22796 6060 22802 6112
rect 23014 6060 23020 6112
rect 23072 6100 23078 6112
rect 23385 6103 23443 6109
rect 23385 6100 23397 6103
rect 23072 6072 23397 6100
rect 23072 6060 23078 6072
rect 23385 6069 23397 6072
rect 23431 6100 23443 6103
rect 26142 6100 26148 6112
rect 23431 6072 26148 6100
rect 23431 6069 23443 6072
rect 23385 6063 23443 6069
rect 26142 6060 26148 6072
rect 26200 6060 26206 6112
rect 28166 6100 28172 6112
rect 28127 6072 28172 6100
rect 28166 6060 28172 6072
rect 28224 6060 28230 6112
rect 1104 6010 28888 6032
rect 1104 5958 10246 6010
rect 10298 5958 10310 6010
rect 10362 5958 10374 6010
rect 10426 5958 10438 6010
rect 10490 5958 19510 6010
rect 19562 5958 19574 6010
rect 19626 5958 19638 6010
rect 19690 5958 19702 6010
rect 19754 5958 28888 6010
rect 1104 5936 28888 5958
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 6362 5896 6368 5908
rect 3752 5868 6368 5896
rect 3752 5856 3758 5868
rect 6362 5856 6368 5868
rect 6420 5856 6426 5908
rect 8573 5899 8631 5905
rect 8573 5865 8585 5899
rect 8619 5896 8631 5899
rect 10962 5896 10968 5908
rect 8619 5868 10824 5896
rect 10923 5868 10968 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 2222 5828 2228 5840
rect 2183 5800 2228 5828
rect 2222 5788 2228 5800
rect 2280 5788 2286 5840
rect 3786 5828 3792 5840
rect 2746 5800 3792 5828
rect 1581 5763 1639 5769
rect 1581 5729 1593 5763
rect 1627 5760 1639 5763
rect 2746 5760 2774 5800
rect 3786 5788 3792 5800
rect 3844 5788 3850 5840
rect 7190 5828 7196 5840
rect 4080 5800 7196 5828
rect 1627 5732 2774 5760
rect 3421 5763 3479 5769
rect 1627 5729 1639 5732
rect 1581 5723 1639 5729
rect 3421 5729 3433 5763
rect 3467 5760 3479 5763
rect 3602 5760 3608 5772
rect 3467 5732 3608 5760
rect 3467 5729 3479 5732
rect 3421 5723 3479 5729
rect 3602 5720 3608 5732
rect 3660 5720 3666 5772
rect 3326 5692 3332 5704
rect 2332 5664 2774 5692
rect 3287 5664 3332 5692
rect 1673 5627 1731 5633
rect 1673 5593 1685 5627
rect 1719 5624 1731 5627
rect 2332 5624 2360 5664
rect 2498 5624 2504 5636
rect 1719 5596 2360 5624
rect 2459 5596 2504 5624
rect 1719 5593 1731 5596
rect 1673 5587 1731 5593
rect 2498 5584 2504 5596
rect 2556 5584 2562 5636
rect 2746 5624 2774 5664
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 4080 5624 4108 5800
rect 7190 5788 7196 5800
rect 7248 5788 7254 5840
rect 10796 5828 10824 5868
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 17497 5899 17555 5905
rect 17497 5865 17509 5899
rect 17543 5896 17555 5899
rect 17954 5896 17960 5908
rect 17543 5868 17960 5896
rect 17543 5865 17555 5868
rect 17497 5859 17555 5865
rect 17954 5856 17960 5868
rect 18012 5856 18018 5908
rect 21358 5856 21364 5908
rect 21416 5896 21422 5908
rect 24486 5896 24492 5908
rect 21416 5868 24492 5896
rect 21416 5856 21422 5868
rect 24486 5856 24492 5868
rect 24544 5856 24550 5908
rect 25314 5896 25320 5908
rect 25275 5868 25320 5896
rect 25314 5856 25320 5868
rect 25372 5856 25378 5908
rect 26050 5896 26056 5908
rect 26011 5868 26056 5896
rect 26050 5856 26056 5868
rect 26108 5856 26114 5908
rect 10796 5800 11192 5828
rect 4246 5760 4252 5772
rect 4207 5732 4252 5760
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 4338 5720 4344 5772
rect 4396 5760 4402 5772
rect 5353 5763 5411 5769
rect 5353 5760 5365 5763
rect 4396 5732 5365 5760
rect 4396 5720 4402 5732
rect 5353 5729 5365 5732
rect 5399 5729 5411 5763
rect 6546 5760 6552 5772
rect 5353 5723 5411 5729
rect 5460 5732 6552 5760
rect 2746 5596 4108 5624
rect 4433 5627 4491 5633
rect 4433 5593 4445 5627
rect 4479 5624 4491 5627
rect 5460 5624 5488 5732
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 6822 5760 6828 5772
rect 6783 5732 6828 5760
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 7650 5720 7656 5772
rect 7708 5760 7714 5772
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 7708 5732 8401 5760
rect 7708 5720 7714 5732
rect 8389 5729 8401 5732
rect 8435 5729 8447 5763
rect 9674 5760 9680 5772
rect 9635 5732 9680 5760
rect 8389 5723 8447 5729
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 9858 5760 9864 5772
rect 9819 5732 9864 5760
rect 9858 5720 9864 5732
rect 9916 5720 9922 5772
rect 10505 5763 10563 5769
rect 10505 5729 10517 5763
rect 10551 5760 10563 5763
rect 10551 5732 10732 5760
rect 10551 5729 10563 5732
rect 10505 5723 10563 5729
rect 9950 5692 9956 5704
rect 4479 5596 5488 5624
rect 6472 5664 9956 5692
rect 4479 5593 4491 5596
rect 4433 5587 4491 5593
rect 2682 5556 2688 5568
rect 2643 5528 2688 5556
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 3786 5556 3792 5568
rect 3747 5528 3792 5556
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 5537 5559 5595 5565
rect 5537 5525 5549 5559
rect 5583 5556 5595 5559
rect 6472 5556 6500 5664
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10045 5695 10103 5701
rect 10045 5661 10057 5695
rect 10091 5692 10103 5695
rect 10594 5692 10600 5704
rect 10091 5664 10600 5692
rect 10091 5661 10103 5664
rect 10045 5655 10103 5661
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 10704 5692 10732 5732
rect 10778 5720 10784 5772
rect 10836 5760 10842 5772
rect 10962 5760 10968 5772
rect 10836 5732 10968 5760
rect 10836 5720 10842 5732
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 11164 5760 11192 5800
rect 11238 5788 11244 5840
rect 11296 5828 11302 5840
rect 12314 5831 12372 5837
rect 12314 5828 12326 5831
rect 11296 5800 12326 5828
rect 11296 5788 11302 5800
rect 12314 5797 12326 5800
rect 12360 5797 12372 5831
rect 12314 5791 12372 5797
rect 13814 5788 13820 5840
rect 13872 5828 13878 5840
rect 14001 5831 14059 5837
rect 14001 5828 14013 5831
rect 13872 5800 14013 5828
rect 13872 5788 13878 5800
rect 14001 5797 14013 5800
rect 14047 5828 14059 5831
rect 14737 5831 14795 5837
rect 14737 5828 14749 5831
rect 14047 5800 14749 5828
rect 14047 5797 14059 5800
rect 14001 5791 14059 5797
rect 14737 5797 14749 5800
rect 14783 5797 14795 5831
rect 14737 5791 14795 5797
rect 14921 5831 14979 5837
rect 14921 5797 14933 5831
rect 14967 5828 14979 5831
rect 15010 5828 15016 5840
rect 14967 5800 15016 5828
rect 14967 5797 14979 5800
rect 14921 5791 14979 5797
rect 15010 5788 15016 5800
rect 15068 5828 15074 5840
rect 25225 5831 25283 5837
rect 15068 5800 17540 5828
rect 15068 5788 15074 5800
rect 17126 5760 17132 5772
rect 11164 5732 17132 5760
rect 17126 5720 17132 5732
rect 17184 5720 17190 5772
rect 17313 5763 17371 5769
rect 17313 5729 17325 5763
rect 17359 5760 17371 5763
rect 17402 5760 17408 5772
rect 17359 5732 17408 5760
rect 17359 5729 17371 5732
rect 17313 5723 17371 5729
rect 17402 5720 17408 5732
rect 17460 5720 17466 5772
rect 17512 5769 17540 5800
rect 19306 5800 25176 5828
rect 17497 5763 17555 5769
rect 17497 5729 17509 5763
rect 17543 5760 17555 5763
rect 17862 5760 17868 5772
rect 17543 5732 17868 5760
rect 17543 5729 17555 5732
rect 17497 5723 17555 5729
rect 17862 5720 17868 5732
rect 17920 5720 17926 5772
rect 18322 5720 18328 5772
rect 18380 5760 18386 5772
rect 18509 5763 18567 5769
rect 18509 5760 18521 5763
rect 18380 5732 18521 5760
rect 18380 5720 18386 5732
rect 18509 5729 18521 5732
rect 18555 5729 18567 5763
rect 18509 5723 18567 5729
rect 10870 5692 10876 5704
rect 10704 5664 10876 5692
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 12066 5692 12072 5704
rect 12027 5664 12072 5692
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14185 5695 14243 5701
rect 14185 5692 14197 5695
rect 13964 5664 14197 5692
rect 13964 5652 13970 5664
rect 14185 5661 14197 5664
rect 14231 5661 14243 5695
rect 17420 5692 17448 5720
rect 18230 5692 18236 5704
rect 17420 5664 18236 5692
rect 14185 5655 14243 5661
rect 18230 5652 18236 5664
rect 18288 5652 18294 5704
rect 18598 5652 18604 5704
rect 18656 5692 18662 5704
rect 19306 5692 19334 5800
rect 24029 5763 24087 5769
rect 24029 5729 24041 5763
rect 24075 5729 24087 5763
rect 24029 5723 24087 5729
rect 24673 5763 24731 5769
rect 24673 5729 24685 5763
rect 24719 5760 24731 5763
rect 24762 5760 24768 5772
rect 24719 5732 24768 5760
rect 24719 5729 24731 5732
rect 24673 5723 24731 5729
rect 18656 5664 19334 5692
rect 24044 5692 24072 5723
rect 24762 5720 24768 5732
rect 24820 5720 24826 5772
rect 25148 5760 25176 5800
rect 25225 5797 25237 5831
rect 25271 5828 25283 5831
rect 28166 5828 28172 5840
rect 25271 5800 28172 5828
rect 25271 5797 25283 5800
rect 25225 5791 25283 5797
rect 28166 5788 28172 5800
rect 28224 5788 28230 5840
rect 25774 5760 25780 5772
rect 25148 5732 25780 5760
rect 25774 5720 25780 5732
rect 25832 5720 25838 5772
rect 25866 5720 25872 5772
rect 25924 5760 25930 5772
rect 25961 5763 26019 5769
rect 25961 5760 25973 5763
rect 25924 5732 25973 5760
rect 25924 5720 25930 5732
rect 25961 5729 25973 5732
rect 26007 5729 26019 5763
rect 26418 5760 26424 5772
rect 25961 5723 26019 5729
rect 26068 5732 26424 5760
rect 26068 5692 26096 5732
rect 26418 5720 26424 5732
rect 26476 5720 26482 5772
rect 26697 5763 26755 5769
rect 26697 5729 26709 5763
rect 26743 5729 26755 5763
rect 26697 5723 26755 5729
rect 27985 5763 28043 5769
rect 27985 5729 27997 5763
rect 28031 5729 28043 5763
rect 27985 5723 28043 5729
rect 24044 5664 26096 5692
rect 18656 5652 18662 5664
rect 26142 5652 26148 5704
rect 26200 5692 26206 5704
rect 26712 5692 26740 5723
rect 26200 5664 26740 5692
rect 26200 5652 26206 5664
rect 6546 5584 6552 5636
rect 6604 5624 6610 5636
rect 13449 5627 13507 5633
rect 6604 5596 11008 5624
rect 6604 5584 6610 5596
rect 7006 5556 7012 5568
rect 5583 5528 6500 5556
rect 6967 5528 7012 5556
rect 5583 5525 5595 5528
rect 5537 5519 5595 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 10686 5565 10692 5568
rect 10643 5559 10692 5565
rect 10643 5525 10655 5559
rect 10689 5525 10692 5559
rect 10643 5519 10692 5525
rect 10686 5516 10692 5519
rect 10744 5516 10750 5568
rect 10778 5516 10784 5568
rect 10836 5556 10842 5568
rect 10980 5556 11008 5596
rect 13449 5593 13461 5627
rect 13495 5624 13507 5627
rect 13630 5624 13636 5636
rect 13495 5596 13636 5624
rect 13495 5593 13507 5596
rect 13449 5587 13507 5593
rect 13630 5584 13636 5596
rect 13688 5624 13694 5636
rect 23845 5627 23903 5633
rect 13688 5596 18736 5624
rect 13688 5584 13694 5596
rect 18708 5568 18736 5596
rect 23845 5593 23857 5627
rect 23891 5624 23903 5627
rect 26694 5624 26700 5636
rect 23891 5596 26700 5624
rect 23891 5593 23903 5596
rect 23845 5587 23903 5593
rect 26694 5584 26700 5596
rect 26752 5584 26758 5636
rect 26878 5624 26884 5636
rect 26839 5596 26884 5624
rect 26878 5584 26884 5596
rect 26936 5584 26942 5636
rect 28000 5624 28028 5723
rect 27080 5596 28028 5624
rect 13262 5556 13268 5568
rect 10836 5528 10881 5556
rect 10980 5528 13268 5556
rect 10836 5516 10842 5528
rect 13262 5516 13268 5528
rect 13320 5516 13326 5568
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 18325 5559 18383 5565
rect 18325 5556 18337 5559
rect 18012 5528 18337 5556
rect 18012 5516 18018 5528
rect 18325 5525 18337 5528
rect 18371 5525 18383 5559
rect 18325 5519 18383 5525
rect 18690 5516 18696 5568
rect 18748 5556 18754 5568
rect 23934 5556 23940 5568
rect 18748 5528 23940 5556
rect 18748 5516 18754 5528
rect 23934 5516 23940 5528
rect 23992 5516 23998 5568
rect 24486 5556 24492 5568
rect 24447 5528 24492 5556
rect 24486 5516 24492 5528
rect 24544 5516 24550 5568
rect 24578 5516 24584 5568
rect 24636 5556 24642 5568
rect 27080 5556 27108 5596
rect 24636 5528 27108 5556
rect 24636 5516 24642 5528
rect 27430 5516 27436 5568
rect 27488 5556 27494 5568
rect 28077 5559 28135 5565
rect 28077 5556 28089 5559
rect 27488 5528 28089 5556
rect 27488 5516 27494 5528
rect 28077 5525 28089 5528
rect 28123 5525 28135 5559
rect 28077 5519 28135 5525
rect 1104 5466 28888 5488
rect 1104 5414 5614 5466
rect 5666 5414 5678 5466
rect 5730 5414 5742 5466
rect 5794 5414 5806 5466
rect 5858 5414 14878 5466
rect 14930 5414 14942 5466
rect 14994 5414 15006 5466
rect 15058 5414 15070 5466
rect 15122 5414 24142 5466
rect 24194 5414 24206 5466
rect 24258 5414 24270 5466
rect 24322 5414 24334 5466
rect 24386 5414 28888 5466
rect 1104 5392 28888 5414
rect 1762 5352 1768 5364
rect 1723 5324 1768 5352
rect 1762 5312 1768 5324
rect 1820 5312 1826 5364
rect 2682 5352 2688 5364
rect 2643 5324 2688 5352
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 2961 5355 3019 5361
rect 2961 5321 2973 5355
rect 3007 5352 3019 5355
rect 3326 5352 3332 5364
rect 3007 5324 3332 5352
rect 3007 5321 3019 5324
rect 2961 5315 3019 5321
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 6549 5355 6607 5361
rect 6549 5352 6561 5355
rect 4448 5324 6561 5352
rect 1578 5244 1584 5296
rect 1636 5284 1642 5296
rect 4448 5284 4476 5324
rect 6549 5321 6561 5324
rect 6595 5321 6607 5355
rect 6549 5315 6607 5321
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 11149 5355 11207 5361
rect 11149 5352 11161 5355
rect 11112 5324 11161 5352
rect 11112 5312 11118 5324
rect 11149 5321 11161 5324
rect 11195 5321 11207 5355
rect 11149 5315 11207 5321
rect 14734 5312 14740 5364
rect 14792 5352 14798 5364
rect 16485 5355 16543 5361
rect 16485 5352 16497 5355
rect 14792 5324 16497 5352
rect 14792 5312 14798 5324
rect 16485 5321 16497 5324
rect 16531 5352 16543 5355
rect 16574 5352 16580 5364
rect 16531 5324 16580 5352
rect 16531 5321 16543 5324
rect 16485 5315 16543 5321
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 22830 5312 22836 5364
rect 22888 5352 22894 5364
rect 25777 5355 25835 5361
rect 25777 5352 25789 5355
rect 22888 5324 25789 5352
rect 22888 5312 22894 5324
rect 25777 5321 25789 5324
rect 25823 5321 25835 5355
rect 25777 5315 25835 5321
rect 26510 5312 26516 5364
rect 26568 5352 26574 5364
rect 27157 5355 27215 5361
rect 27157 5352 27169 5355
rect 26568 5324 27169 5352
rect 26568 5312 26574 5324
rect 27157 5321 27169 5324
rect 27203 5321 27215 5355
rect 27157 5315 27215 5321
rect 27338 5312 27344 5364
rect 27396 5312 27402 5364
rect 1636 5256 4476 5284
rect 5813 5287 5871 5293
rect 1636 5244 1642 5256
rect 5813 5253 5825 5287
rect 5859 5284 5871 5287
rect 5994 5284 6000 5296
rect 5859 5256 6000 5284
rect 5859 5253 5871 5256
rect 5813 5247 5871 5253
rect 5994 5244 6000 5256
rect 6052 5244 6058 5296
rect 10778 5244 10784 5296
rect 10836 5284 10842 5296
rect 11517 5287 11575 5293
rect 11517 5284 11529 5287
rect 10836 5256 11529 5284
rect 10836 5244 10842 5256
rect 11517 5253 11529 5256
rect 11563 5284 11575 5287
rect 12161 5287 12219 5293
rect 12161 5284 12173 5287
rect 11563 5256 12173 5284
rect 11563 5253 11575 5256
rect 11517 5247 11575 5253
rect 12161 5253 12173 5256
rect 12207 5253 12219 5287
rect 12161 5247 12219 5253
rect 13817 5287 13875 5293
rect 13817 5253 13829 5287
rect 13863 5284 13875 5287
rect 14182 5284 14188 5296
rect 13863 5256 14188 5284
rect 13863 5253 13875 5256
rect 13817 5247 13875 5253
rect 14182 5244 14188 5256
rect 14240 5244 14246 5296
rect 19886 5244 19892 5296
rect 19944 5284 19950 5296
rect 25593 5287 25651 5293
rect 25593 5284 25605 5287
rect 19944 5256 25605 5284
rect 19944 5244 19950 5256
rect 25593 5253 25605 5256
rect 25639 5253 25651 5287
rect 27356 5284 27384 5312
rect 27356 5256 27568 5284
rect 25593 5247 25651 5253
rect 6914 5216 6920 5228
rect 5460 5188 6920 5216
rect 1946 5148 1952 5160
rect 1907 5120 1952 5148
rect 1946 5108 1952 5120
rect 2004 5108 2010 5160
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 2958 5148 2964 5160
rect 2832 5120 2964 5148
rect 2832 5108 2838 5120
rect 2958 5108 2964 5120
rect 3016 5108 3022 5160
rect 3145 5151 3203 5157
rect 3145 5117 3157 5151
rect 3191 5148 3203 5151
rect 3234 5148 3240 5160
rect 3191 5120 3240 5148
rect 3191 5117 3203 5120
rect 3145 5111 3203 5117
rect 3234 5108 3240 5120
rect 3292 5108 3298 5160
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 4982 5148 4988 5160
rect 4479 5120 4988 5148
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 4982 5108 4988 5120
rect 5040 5148 5046 5160
rect 5460 5148 5488 5188
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 9674 5176 9680 5228
rect 9732 5216 9738 5228
rect 10686 5216 10692 5228
rect 9732 5188 10456 5216
rect 10599 5188 10692 5216
rect 9732 5176 9738 5188
rect 6362 5148 6368 5160
rect 5040 5120 5488 5148
rect 6323 5120 6368 5148
rect 5040 5108 5046 5120
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 6454 5108 6460 5160
rect 6512 5148 6518 5160
rect 7009 5151 7067 5157
rect 7009 5148 7021 5151
rect 6512 5120 7021 5148
rect 6512 5108 6518 5120
rect 7009 5117 7021 5120
rect 7055 5117 7067 5151
rect 8202 5148 8208 5160
rect 8163 5120 8208 5148
rect 7009 5111 7067 5117
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 8386 5148 8392 5160
rect 8347 5120 8392 5148
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 9858 5108 9864 5160
rect 9916 5148 9922 5160
rect 10428 5157 10456 5188
rect 10686 5176 10692 5188
rect 10744 5216 10750 5228
rect 11609 5219 11667 5225
rect 11609 5216 11621 5219
rect 10744 5188 11621 5216
rect 10744 5176 10750 5188
rect 11609 5185 11621 5188
rect 11655 5185 11667 5219
rect 21726 5216 21732 5228
rect 11609 5179 11667 5185
rect 17604 5188 21732 5216
rect 9953 5151 10011 5157
rect 9953 5148 9965 5151
rect 9916 5120 9965 5148
rect 9916 5108 9922 5120
rect 9953 5117 9965 5120
rect 9999 5117 10011 5151
rect 9953 5111 10011 5117
rect 10413 5151 10471 5157
rect 10413 5117 10425 5151
rect 10459 5117 10471 5151
rect 10413 5111 10471 5117
rect 10870 5108 10876 5160
rect 10928 5148 10934 5160
rect 11333 5151 11391 5157
rect 11333 5148 11345 5151
rect 10928 5120 11345 5148
rect 10928 5108 10934 5120
rect 11333 5117 11345 5120
rect 11379 5117 11391 5151
rect 11333 5111 11391 5117
rect 12069 5151 12127 5157
rect 12069 5117 12081 5151
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 13633 5151 13691 5157
rect 13633 5117 13645 5151
rect 13679 5148 13691 5151
rect 13814 5148 13820 5160
rect 13679 5120 13820 5148
rect 13679 5117 13691 5120
rect 13633 5111 13691 5117
rect 4614 5040 4620 5092
rect 4672 5089 4678 5092
rect 4672 5083 4736 5089
rect 4672 5049 4690 5083
rect 4724 5049 4736 5083
rect 4672 5043 4736 5049
rect 4672 5040 4678 5043
rect 10594 5040 10600 5092
rect 10652 5080 10658 5092
rect 12084 5080 12112 5111
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 13906 5108 13912 5160
rect 13964 5148 13970 5160
rect 16393 5151 16451 5157
rect 16393 5148 16405 5151
rect 13964 5120 16405 5148
rect 13964 5108 13970 5120
rect 16393 5117 16405 5120
rect 16439 5117 16451 5151
rect 16393 5111 16451 5117
rect 10652 5052 12112 5080
rect 16408 5080 16436 5111
rect 16942 5108 16948 5160
rect 17000 5148 17006 5160
rect 17604 5157 17632 5188
rect 21726 5176 21732 5188
rect 21784 5176 21790 5228
rect 27338 5216 27344 5228
rect 23676 5188 27344 5216
rect 17589 5151 17647 5157
rect 17589 5148 17601 5151
rect 17000 5120 17601 5148
rect 17000 5108 17006 5120
rect 17589 5117 17601 5120
rect 17635 5117 17647 5151
rect 17589 5111 17647 5117
rect 17773 5151 17831 5157
rect 17773 5117 17785 5151
rect 17819 5148 17831 5151
rect 17862 5148 17868 5160
rect 17819 5120 17868 5148
rect 17819 5117 17831 5120
rect 17773 5111 17831 5117
rect 17862 5108 17868 5120
rect 17920 5108 17926 5160
rect 19794 5108 19800 5160
rect 19852 5148 19858 5160
rect 20165 5151 20223 5157
rect 20165 5148 20177 5151
rect 19852 5120 20177 5148
rect 19852 5108 19858 5120
rect 20165 5117 20177 5120
rect 20211 5117 20223 5151
rect 20165 5111 20223 5117
rect 21174 5108 21180 5160
rect 21232 5148 21238 5160
rect 23676 5157 23704 5188
rect 27338 5176 27344 5188
rect 27396 5176 27402 5228
rect 27540 5225 27568 5256
rect 27525 5219 27583 5225
rect 27525 5185 27537 5219
rect 27571 5185 27583 5219
rect 27525 5179 27583 5185
rect 21269 5151 21327 5157
rect 21269 5148 21281 5151
rect 21232 5120 21281 5148
rect 21232 5108 21238 5120
rect 21269 5117 21281 5120
rect 21315 5117 21327 5151
rect 21269 5111 21327 5117
rect 23661 5151 23719 5157
rect 23661 5117 23673 5151
rect 23707 5117 23719 5151
rect 23661 5111 23719 5117
rect 23750 5108 23756 5160
rect 23808 5148 23814 5160
rect 24121 5151 24179 5157
rect 24121 5148 24133 5151
rect 23808 5120 24133 5148
rect 23808 5108 23814 5120
rect 24121 5117 24133 5120
rect 24167 5117 24179 5151
rect 24121 5111 24179 5117
rect 24305 5151 24363 5157
rect 24305 5117 24317 5151
rect 24351 5117 24363 5151
rect 24305 5111 24363 5117
rect 18325 5083 18383 5089
rect 18325 5080 18337 5083
rect 16408 5052 18337 5080
rect 10652 5040 10658 5052
rect 18325 5049 18337 5052
rect 18371 5049 18383 5083
rect 18325 5043 18383 5049
rect 18509 5083 18567 5089
rect 18509 5049 18521 5083
rect 18555 5080 18567 5083
rect 18782 5080 18788 5092
rect 18555 5052 18788 5080
rect 18555 5049 18567 5052
rect 18509 5043 18567 5049
rect 18782 5040 18788 5052
rect 18840 5040 18846 5092
rect 22462 5040 22468 5092
rect 22520 5080 22526 5092
rect 24320 5080 24348 5111
rect 25222 5108 25228 5160
rect 25280 5148 25286 5160
rect 25685 5151 25743 5157
rect 25685 5148 25697 5151
rect 25280 5120 25697 5148
rect 25280 5108 25286 5120
rect 25685 5117 25697 5120
rect 25731 5117 25743 5151
rect 25685 5111 25743 5117
rect 22520 5052 24348 5080
rect 26421 5083 26479 5089
rect 22520 5040 22526 5052
rect 26421 5049 26433 5083
rect 26467 5049 26479 5083
rect 26602 5080 26608 5092
rect 26563 5052 26608 5080
rect 26421 5043 26479 5049
rect 6270 4972 6276 5024
rect 6328 5012 6334 5024
rect 7193 5015 7251 5021
rect 7193 5012 7205 5015
rect 6328 4984 7205 5012
rect 6328 4972 6334 4984
rect 7193 4981 7205 4984
rect 7239 4981 7251 5015
rect 7193 4975 7251 4981
rect 8110 4972 8116 5024
rect 8168 5012 8174 5024
rect 8297 5015 8355 5021
rect 8297 5012 8309 5015
rect 8168 4984 8309 5012
rect 8168 4972 8174 4984
rect 8297 4981 8309 4984
rect 8343 4981 8355 5015
rect 8297 4975 8355 4981
rect 9582 4972 9588 5024
rect 9640 5012 9646 5024
rect 15378 5012 15384 5024
rect 9640 4984 15384 5012
rect 9640 4972 9646 4984
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 18138 4972 18144 5024
rect 18196 5012 18202 5024
rect 19242 5012 19248 5024
rect 18196 4984 19248 5012
rect 18196 4972 18202 4984
rect 19242 4972 19248 4984
rect 19300 4972 19306 5024
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 19981 5015 20039 5021
rect 19981 5012 19993 5015
rect 19392 4984 19993 5012
rect 19392 4972 19398 4984
rect 19981 4981 19993 4984
rect 20027 4981 20039 5015
rect 19981 4975 20039 4981
rect 20162 4972 20168 5024
rect 20220 5012 20226 5024
rect 21085 5015 21143 5021
rect 21085 5012 21097 5015
rect 20220 4984 21097 5012
rect 20220 4972 20226 4984
rect 21085 4981 21097 4984
rect 21131 4981 21143 5015
rect 23474 5012 23480 5024
rect 23435 4984 23480 5012
rect 21085 4975 21143 4981
rect 23474 4972 23480 4984
rect 23532 4972 23538 5024
rect 24305 5015 24363 5021
rect 24305 4981 24317 5015
rect 24351 5012 24363 5015
rect 25038 5012 25044 5024
rect 24351 4984 25044 5012
rect 24351 4981 24363 4984
rect 24305 4975 24363 4981
rect 25038 4972 25044 4984
rect 25096 4972 25102 5024
rect 25593 5015 25651 5021
rect 25593 4981 25605 5015
rect 25639 5012 25651 5015
rect 26436 5012 26464 5043
rect 26602 5040 26608 5052
rect 26660 5040 26666 5092
rect 27706 5080 27712 5092
rect 27667 5052 27712 5080
rect 27706 5040 27712 5052
rect 27764 5040 27770 5092
rect 25639 4984 26464 5012
rect 25639 4981 25651 4984
rect 25593 4975 25651 4981
rect 27522 4972 27528 5024
rect 27580 5012 27586 5024
rect 27617 5015 27675 5021
rect 27617 5012 27629 5015
rect 27580 4984 27629 5012
rect 27580 4972 27586 4984
rect 27617 4981 27629 4984
rect 27663 4981 27675 5015
rect 27617 4975 27675 4981
rect 1104 4922 28888 4944
rect 1104 4870 10246 4922
rect 10298 4870 10310 4922
rect 10362 4870 10374 4922
rect 10426 4870 10438 4922
rect 10490 4870 19510 4922
rect 19562 4870 19574 4922
rect 19626 4870 19638 4922
rect 19690 4870 19702 4922
rect 19754 4870 28888 4922
rect 1104 4848 28888 4870
rect 2409 4811 2467 4817
rect 2409 4777 2421 4811
rect 2455 4808 2467 4811
rect 2455 4780 2774 4808
rect 2455 4777 2467 4780
rect 2409 4771 2467 4777
rect 2746 4740 2774 4780
rect 3786 4768 3792 4820
rect 3844 4808 3850 4820
rect 4525 4811 4583 4817
rect 4525 4808 4537 4811
rect 3844 4780 4537 4808
rect 3844 4768 3850 4780
rect 4525 4777 4537 4780
rect 4571 4777 4583 4811
rect 4525 4771 4583 4777
rect 5902 4768 5908 4820
rect 5960 4768 5966 4820
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 15194 4808 15200 4820
rect 12492 4780 12537 4808
rect 15155 4780 15200 4808
rect 12492 4768 12498 4780
rect 15194 4768 15200 4780
rect 15252 4768 15258 4820
rect 16298 4808 16304 4820
rect 15304 4780 16304 4808
rect 5920 4740 5948 4768
rect 10686 4740 10692 4752
rect 2746 4712 5948 4740
rect 10152 4712 10692 4740
rect 1394 4632 1400 4684
rect 1452 4672 1458 4684
rect 1949 4675 2007 4681
rect 1949 4672 1961 4675
rect 1452 4644 1961 4672
rect 1452 4632 1458 4644
rect 1949 4641 1961 4644
rect 1995 4641 2007 4675
rect 1949 4635 2007 4641
rect 2593 4675 2651 4681
rect 2593 4641 2605 4675
rect 2639 4672 2651 4675
rect 2774 4672 2780 4684
rect 2639 4644 2780 4672
rect 2639 4641 2651 4644
rect 2593 4635 2651 4641
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 3234 4672 3240 4684
rect 3195 4644 3240 4672
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 4430 4632 4436 4684
rect 4488 4672 4494 4684
rect 5537 4675 5595 4681
rect 4488 4644 4752 4672
rect 4488 4632 4494 4644
rect 4724 4613 4752 4644
rect 5537 4641 5549 4675
rect 5583 4672 5595 4675
rect 5902 4672 5908 4684
rect 5583 4644 5908 4672
rect 5583 4641 5595 4644
rect 5537 4635 5595 4641
rect 5902 4632 5908 4644
rect 5960 4632 5966 4684
rect 7009 4675 7067 4681
rect 7009 4641 7021 4675
rect 7055 4672 7067 4675
rect 7282 4672 7288 4684
rect 7055 4644 7288 4672
rect 7055 4641 7067 4644
rect 7009 4635 7067 4641
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 8110 4672 8116 4684
rect 8071 4644 8116 4672
rect 8110 4632 8116 4644
rect 8168 4632 8174 4684
rect 8754 4672 8760 4684
rect 8715 4644 8760 4672
rect 8754 4632 8760 4644
rect 8812 4632 8818 4684
rect 9030 4672 9036 4684
rect 8991 4644 9036 4672
rect 9030 4632 9036 4644
rect 9088 4632 9094 4684
rect 10152 4681 10180 4712
rect 10686 4700 10692 4712
rect 10744 4700 10750 4752
rect 13814 4740 13820 4752
rect 13775 4712 13820 4740
rect 13814 4700 13820 4712
rect 13872 4700 13878 4752
rect 14182 4700 14188 4752
rect 14240 4740 14246 4752
rect 14240 4712 14688 4740
rect 14240 4700 14246 4712
rect 10137 4675 10195 4681
rect 10137 4641 10149 4675
rect 10183 4641 10195 4675
rect 10594 4672 10600 4684
rect 10555 4644 10600 4672
rect 10137 4635 10195 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 12158 4632 12164 4684
rect 12216 4672 12222 4684
rect 14660 4681 14688 4712
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 12216 4644 12357 4672
rect 12216 4632 12222 4644
rect 12345 4641 12357 4644
rect 12391 4641 12403 4675
rect 12345 4635 12403 4641
rect 14461 4675 14519 4681
rect 14461 4641 14473 4675
rect 14507 4641 14519 4675
rect 14461 4635 14519 4641
rect 14645 4675 14703 4681
rect 14645 4641 14657 4675
rect 14691 4641 14703 4675
rect 14645 4635 14703 4641
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4573 4675 4607
rect 4617 4567 4675 4573
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 7098 4604 7104 4616
rect 7059 4576 7104 4604
rect 4709 4567 4767 4573
rect 1765 4539 1823 4545
rect 1765 4505 1777 4539
rect 1811 4536 1823 4539
rect 3510 4536 3516 4548
rect 1811 4508 3516 4536
rect 1811 4505 1823 4508
rect 1765 4499 1823 4505
rect 3510 4496 3516 4508
rect 3568 4496 3574 4548
rect 4632 4536 4660 4567
rect 7098 4564 7104 4576
rect 7156 4604 7162 4616
rect 10870 4604 10876 4616
rect 7156 4576 8340 4604
rect 10831 4576 10876 4604
rect 7156 4564 7162 4576
rect 6086 4536 6092 4548
rect 4632 4508 6092 4536
rect 6086 4496 6092 4508
rect 6144 4496 6150 4548
rect 8312 4545 8340 4576
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 14476 4604 14504 4635
rect 14734 4632 14740 4684
rect 14792 4672 14798 4684
rect 15105 4675 15163 4681
rect 15105 4672 15117 4675
rect 14792 4644 15117 4672
rect 14792 4632 14798 4644
rect 15105 4641 15117 4644
rect 15151 4641 15163 4675
rect 15105 4635 15163 4641
rect 15304 4604 15332 4780
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 16666 4768 16672 4820
rect 16724 4808 16730 4820
rect 17862 4808 17868 4820
rect 16724 4780 17868 4808
rect 16724 4768 16730 4780
rect 17862 4768 17868 4780
rect 17920 4808 17926 4820
rect 19613 4811 19671 4817
rect 17920 4780 19196 4808
rect 17920 4768 17926 4780
rect 16574 4740 16580 4752
rect 16132 4712 16580 4740
rect 16132 4681 16160 4712
rect 16574 4700 16580 4712
rect 16632 4700 16638 4752
rect 17770 4700 17776 4752
rect 17828 4740 17834 4752
rect 17828 4712 18552 4740
rect 17828 4700 17834 4712
rect 16025 4675 16083 4681
rect 16025 4641 16037 4675
rect 16071 4641 16083 4675
rect 16025 4635 16083 4641
rect 16117 4675 16175 4681
rect 16117 4641 16129 4675
rect 16163 4641 16175 4675
rect 16117 4635 16175 4641
rect 14476 4576 15332 4604
rect 16040 4604 16068 4635
rect 16206 4632 16212 4684
rect 16264 4672 16270 4684
rect 16390 4672 16396 4684
rect 16264 4644 16309 4672
rect 16351 4644 16396 4672
rect 16264 4632 16270 4644
rect 16390 4632 16396 4644
rect 16448 4632 16454 4684
rect 18138 4672 18144 4684
rect 18099 4644 18144 4672
rect 18138 4632 18144 4644
rect 18196 4632 18202 4684
rect 18524 4681 18552 4712
rect 18233 4675 18291 4681
rect 18233 4641 18245 4675
rect 18279 4641 18291 4675
rect 18233 4635 18291 4641
rect 18325 4675 18383 4681
rect 18325 4641 18337 4675
rect 18371 4641 18383 4675
rect 18325 4635 18383 4641
rect 18509 4675 18567 4681
rect 18509 4641 18521 4675
rect 18555 4641 18567 4675
rect 18509 4635 18567 4641
rect 16040 4576 16160 4604
rect 8297 4539 8355 4545
rect 8297 4505 8309 4539
rect 8343 4505 8355 4539
rect 8297 4499 8355 4505
rect 9030 4496 9036 4548
rect 9088 4536 9094 4548
rect 10045 4539 10103 4545
rect 10045 4536 10057 4539
rect 9088 4508 10057 4536
rect 9088 4496 9094 4508
rect 10045 4505 10057 4508
rect 10091 4505 10103 4539
rect 10045 4499 10103 4505
rect 13262 4496 13268 4548
rect 13320 4536 13326 4548
rect 14001 4539 14059 4545
rect 14001 4536 14013 4539
rect 13320 4508 14013 4536
rect 13320 4496 13326 4508
rect 14001 4505 14013 4508
rect 14047 4536 14059 4539
rect 15654 4536 15660 4548
rect 14047 4508 15660 4536
rect 14047 4505 14059 4508
rect 14001 4499 14059 4505
rect 15654 4496 15660 4508
rect 15712 4496 15718 4548
rect 16132 4536 16160 4576
rect 16574 4564 16580 4616
rect 16632 4604 16638 4616
rect 18248 4604 18276 4635
rect 18340 4604 18368 4635
rect 18874 4632 18880 4684
rect 18932 4672 18938 4684
rect 19168 4681 19196 4780
rect 19613 4777 19625 4811
rect 19659 4808 19671 4811
rect 20714 4808 20720 4820
rect 19659 4780 20720 4808
rect 19659 4777 19671 4780
rect 19613 4771 19671 4777
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 23934 4768 23940 4820
rect 23992 4808 23998 4820
rect 23992 4780 28028 4808
rect 23992 4768 23998 4780
rect 19242 4700 19248 4752
rect 19300 4740 19306 4752
rect 19981 4743 20039 4749
rect 19981 4740 19993 4743
rect 19300 4712 19993 4740
rect 19300 4700 19306 4712
rect 19981 4709 19993 4712
rect 20027 4709 20039 4743
rect 19981 4703 20039 4709
rect 20070 4700 20076 4752
rect 20128 4700 20134 4752
rect 22002 4740 22008 4752
rect 21284 4712 22008 4740
rect 18969 4675 19027 4681
rect 18969 4672 18981 4675
rect 18932 4644 18981 4672
rect 18932 4632 18938 4644
rect 18969 4641 18981 4644
rect 19015 4641 19027 4675
rect 18969 4635 19027 4641
rect 19153 4675 19211 4681
rect 19153 4641 19165 4675
rect 19199 4641 19211 4675
rect 19153 4635 19211 4641
rect 18414 4604 18420 4616
rect 16632 4576 18276 4604
rect 18327 4576 18420 4604
rect 16632 4564 16638 4576
rect 18414 4564 18420 4576
rect 18472 4604 18478 4616
rect 18984 4604 19012 4635
rect 19702 4632 19708 4684
rect 19760 4672 19766 4684
rect 20088 4672 20116 4700
rect 21284 4681 21312 4712
rect 22002 4700 22008 4712
rect 22060 4740 22066 4752
rect 22370 4740 22376 4752
rect 22060 4712 22376 4740
rect 22060 4700 22066 4712
rect 22370 4700 22376 4712
rect 22428 4740 22434 4752
rect 23106 4740 23112 4752
rect 22428 4712 23112 4740
rect 22428 4700 22434 4712
rect 23106 4700 23112 4712
rect 23164 4740 23170 4752
rect 23385 4743 23443 4749
rect 23385 4740 23397 4743
rect 23164 4712 23397 4740
rect 23164 4700 23170 4712
rect 23385 4709 23397 4712
rect 23431 4709 23443 4743
rect 23566 4740 23572 4752
rect 23527 4712 23572 4740
rect 23385 4703 23443 4709
rect 23566 4700 23572 4712
rect 23624 4700 23630 4752
rect 23658 4700 23664 4752
rect 23716 4740 23722 4752
rect 24578 4740 24584 4752
rect 23716 4712 24584 4740
rect 23716 4700 23722 4712
rect 24578 4700 24584 4712
rect 24636 4700 24642 4752
rect 25406 4700 25412 4752
rect 25464 4740 25470 4752
rect 28000 4749 28028 4780
rect 27985 4743 28043 4749
rect 25464 4712 26464 4740
rect 25464 4700 25470 4712
rect 19760 4644 20116 4672
rect 21269 4675 21327 4681
rect 19760 4632 19766 4644
rect 21269 4641 21281 4675
rect 21315 4641 21327 4675
rect 21269 4635 21327 4641
rect 21358 4675 21416 4681
rect 21358 4641 21370 4675
rect 21404 4641 21416 4675
rect 21358 4635 21416 4641
rect 21453 4675 21511 4681
rect 21453 4641 21465 4675
rect 21499 4641 21511 4675
rect 21634 4672 21640 4684
rect 21595 4644 21640 4672
rect 21453 4635 21511 4641
rect 19886 4604 19892 4616
rect 18472 4576 18920 4604
rect 18984 4576 19892 4604
rect 18472 4564 18478 4576
rect 18892 4548 18920 4576
rect 19886 4564 19892 4576
rect 19944 4564 19950 4616
rect 20070 4604 20076 4616
rect 20031 4576 20076 4604
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 20165 4607 20223 4613
rect 20165 4573 20177 4607
rect 20211 4573 20223 4607
rect 20165 4567 20223 4573
rect 17678 4536 17684 4548
rect 16132 4508 17684 4536
rect 17678 4496 17684 4508
rect 17736 4496 17742 4548
rect 18874 4496 18880 4548
rect 18932 4496 18938 4548
rect 19978 4496 19984 4548
rect 20036 4536 20042 4548
rect 20180 4536 20208 4567
rect 20990 4564 20996 4616
rect 21048 4604 21054 4616
rect 21376 4604 21404 4635
rect 21048 4576 21404 4604
rect 21468 4604 21496 4635
rect 21634 4632 21640 4644
rect 21692 4632 21698 4684
rect 22738 4632 22744 4684
rect 22796 4672 22802 4684
rect 24486 4672 24492 4684
rect 22796 4644 24072 4672
rect 24447 4644 24492 4672
rect 22796 4632 22802 4644
rect 21542 4604 21548 4616
rect 21468 4576 21548 4604
rect 21048 4564 21054 4576
rect 20622 4536 20628 4548
rect 20036 4508 20628 4536
rect 20036 4496 20042 4508
rect 20622 4496 20628 4508
rect 20680 4496 20686 4548
rect 21376 4536 21404 4576
rect 21542 4564 21548 4576
rect 21600 4564 21606 4616
rect 23382 4564 23388 4616
rect 23440 4604 23446 4616
rect 23934 4604 23940 4616
rect 23440 4576 23940 4604
rect 23440 4564 23446 4576
rect 23934 4564 23940 4576
rect 23992 4564 23998 4616
rect 24044 4604 24072 4644
rect 24486 4632 24492 4644
rect 24544 4632 24550 4684
rect 25314 4632 25320 4684
rect 25372 4672 25378 4684
rect 25665 4675 25723 4681
rect 25665 4672 25677 4675
rect 25372 4644 25677 4672
rect 25372 4632 25378 4644
rect 25665 4641 25677 4644
rect 25711 4641 25723 4675
rect 25665 4635 25723 4641
rect 25409 4607 25467 4613
rect 25409 4604 25421 4607
rect 24044 4576 25421 4604
rect 25409 4573 25421 4576
rect 25455 4573 25467 4607
rect 25409 4567 25467 4573
rect 23014 4536 23020 4548
rect 21376 4508 23020 4536
rect 23014 4496 23020 4508
rect 23072 4496 23078 4548
rect 23109 4539 23167 4545
rect 23109 4505 23121 4539
rect 23155 4536 23167 4539
rect 23842 4536 23848 4548
rect 23155 4508 23848 4536
rect 23155 4505 23167 4508
rect 23109 4499 23167 4505
rect 23842 4496 23848 4508
rect 23900 4496 23906 4548
rect 3050 4468 3056 4480
rect 3011 4440 3056 4468
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 4157 4471 4215 4477
rect 4157 4437 4169 4471
rect 4203 4468 4215 4471
rect 4338 4468 4344 4480
rect 4203 4440 4344 4468
rect 4203 4437 4215 4440
rect 4157 4431 4215 4437
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 4430 4428 4436 4480
rect 4488 4468 4494 4480
rect 5353 4471 5411 4477
rect 5353 4468 5365 4471
rect 4488 4440 5365 4468
rect 4488 4428 4494 4440
rect 5353 4437 5365 4440
rect 5399 4437 5411 4471
rect 7374 4468 7380 4480
rect 7335 4440 7380 4468
rect 5353 4431 5411 4437
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 14553 4471 14611 4477
rect 14553 4437 14565 4471
rect 14599 4468 14611 4471
rect 15562 4468 15568 4480
rect 14599 4440 15568 4468
rect 14599 4437 14611 4440
rect 14553 4431 14611 4437
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 15749 4471 15807 4477
rect 15749 4437 15761 4471
rect 15795 4468 15807 4471
rect 16022 4468 16028 4480
rect 15795 4440 16028 4468
rect 15795 4437 15807 4440
rect 15749 4431 15807 4437
rect 16022 4428 16028 4440
rect 16080 4428 16086 4480
rect 17862 4468 17868 4480
rect 17823 4440 17868 4468
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 19058 4468 19064 4480
rect 19019 4440 19064 4468
rect 19058 4428 19064 4440
rect 19116 4428 19122 4480
rect 20993 4471 21051 4477
rect 20993 4437 21005 4471
rect 21039 4468 21051 4471
rect 21082 4468 21088 4480
rect 21039 4440 21088 4468
rect 21039 4437 21051 4440
rect 20993 4431 21051 4437
rect 21082 4428 21088 4440
rect 21140 4428 21146 4480
rect 21910 4428 21916 4480
rect 21968 4468 21974 4480
rect 24581 4471 24639 4477
rect 24581 4468 24593 4471
rect 21968 4440 24593 4468
rect 21968 4428 21974 4440
rect 24581 4437 24593 4440
rect 24627 4437 24639 4471
rect 25424 4468 25452 4567
rect 26436 4536 26464 4712
rect 27985 4709 27997 4743
rect 28031 4709 28043 4743
rect 27985 4703 28043 4709
rect 26789 4539 26847 4545
rect 26789 4536 26801 4539
rect 26436 4508 26801 4536
rect 26789 4505 26801 4508
rect 26835 4536 26847 4539
rect 27706 4536 27712 4548
rect 26835 4508 27712 4536
rect 26835 4505 26847 4508
rect 26789 4499 26847 4505
rect 27706 4496 27712 4508
rect 27764 4496 27770 4548
rect 26050 4468 26056 4480
rect 25424 4440 26056 4468
rect 24581 4431 24639 4437
rect 26050 4428 26056 4440
rect 26108 4428 26114 4480
rect 28074 4468 28080 4480
rect 28035 4440 28080 4468
rect 28074 4428 28080 4440
rect 28132 4428 28138 4480
rect 1104 4378 28888 4400
rect 1104 4326 5614 4378
rect 5666 4326 5678 4378
rect 5730 4326 5742 4378
rect 5794 4326 5806 4378
rect 5858 4326 14878 4378
rect 14930 4326 14942 4378
rect 14994 4326 15006 4378
rect 15058 4326 15070 4378
rect 15122 4326 24142 4378
rect 24194 4326 24206 4378
rect 24258 4326 24270 4378
rect 24322 4326 24334 4378
rect 24386 4326 28888 4378
rect 1104 4304 28888 4326
rect 4154 4224 4160 4276
rect 4212 4264 4218 4276
rect 4982 4264 4988 4276
rect 4212 4236 4988 4264
rect 4212 4224 4218 4236
rect 4982 4224 4988 4236
rect 5040 4224 5046 4276
rect 5629 4267 5687 4273
rect 5629 4233 5641 4267
rect 5675 4264 5687 4267
rect 6086 4264 6092 4276
rect 5675 4236 6092 4264
rect 5675 4233 5687 4236
rect 5629 4227 5687 4233
rect 6086 4224 6092 4236
rect 6144 4224 6150 4276
rect 10870 4264 10876 4276
rect 10831 4236 10876 4264
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 12894 4224 12900 4276
rect 12952 4264 12958 4276
rect 13906 4264 13912 4276
rect 12952 4236 13912 4264
rect 12952 4224 12958 4236
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 16574 4264 16580 4276
rect 15120 4236 16580 4264
rect 4246 4196 4252 4208
rect 3252 4168 4252 4196
rect 1670 4128 1676 4140
rect 1631 4100 1676 4128
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 3252 4137 3280 4168
rect 4246 4156 4252 4168
rect 4304 4156 4310 4208
rect 10962 4196 10968 4208
rect 10244 4168 10968 4196
rect 3237 4131 3295 4137
rect 3237 4097 3249 4131
rect 3283 4097 3295 4131
rect 6638 4128 6644 4140
rect 6599 4100 6644 4128
rect 3237 4091 3295 4097
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4128 6883 4131
rect 7558 4128 7564 4140
rect 6871 4100 7564 4128
rect 6871 4097 6883 4100
rect 6825 4091 6883 4097
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 8386 4128 8392 4140
rect 7944 4100 8392 4128
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4060 1639 4063
rect 3050 4060 3056 4072
rect 1627 4032 3056 4060
rect 1627 4029 1639 4032
rect 1581 4023 1639 4029
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 4212 4032 4261 4060
rect 4212 4020 4218 4032
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 4338 4020 4344 4072
rect 4396 4060 4402 4072
rect 4505 4063 4563 4069
rect 4505 4060 4517 4063
rect 4396 4032 4517 4060
rect 4396 4020 4402 4032
rect 4505 4029 4517 4032
rect 4551 4029 4563 4063
rect 7466 4060 7472 4072
rect 4505 4023 4563 4029
rect 4632 4032 7472 4060
rect 1670 3952 1676 4004
rect 1728 3992 1734 4004
rect 4632 3992 4660 4032
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 7944 4069 7972 4100
rect 8386 4088 8392 4100
rect 8444 4088 8450 4140
rect 8478 4088 8484 4140
rect 8536 4128 8542 4140
rect 8573 4131 8631 4137
rect 8573 4128 8585 4131
rect 8536 4100 8585 4128
rect 8536 4088 8542 4100
rect 8573 4097 8585 4100
rect 8619 4128 8631 4131
rect 8754 4128 8760 4140
rect 8619 4100 8760 4128
rect 8619 4097 8631 4100
rect 8573 4091 8631 4097
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 9858 4088 9864 4140
rect 9916 4128 9922 4140
rect 10244 4137 10272 4168
rect 10962 4156 10968 4168
rect 11020 4156 11026 4208
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9916 4100 10057 4128
rect 9916 4088 9922 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4097 10287 4131
rect 11606 4128 11612 4140
rect 10229 4091 10287 4097
rect 10612 4100 11612 4128
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4029 7987 4063
rect 8202 4060 8208 4072
rect 8163 4032 8208 4060
rect 7929 4023 7987 4029
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 9953 4063 10011 4069
rect 9953 4029 9965 4063
rect 9999 4060 10011 4063
rect 10612 4060 10640 4100
rect 11606 4088 11612 4100
rect 11664 4088 11670 4140
rect 12158 4088 12164 4140
rect 12216 4128 12222 4140
rect 12216 4100 13032 4128
rect 12216 4088 12222 4100
rect 10778 4060 10784 4072
rect 9999 4032 10640 4060
rect 10739 4032 10784 4060
rect 9999 4029 10011 4032
rect 9953 4023 10011 4029
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 11514 4020 11520 4072
rect 11572 4060 11578 4072
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 11572 4032 11713 4060
rect 11572 4020 11578 4032
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 11701 4023 11759 4029
rect 12253 4063 12311 4069
rect 12253 4029 12265 4063
rect 12299 4029 12311 4063
rect 12253 4023 12311 4029
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4060 12495 4063
rect 12894 4060 12900 4072
rect 12483 4032 12900 4060
rect 12483 4029 12495 4032
rect 12437 4023 12495 4029
rect 1728 3964 4660 3992
rect 1728 3952 1734 3964
rect 4706 3952 4712 4004
rect 4764 3992 4770 4004
rect 6454 3992 6460 4004
rect 4764 3964 6460 3992
rect 4764 3952 4770 3964
rect 6454 3952 6460 3964
rect 6512 3952 6518 4004
rect 7006 3952 7012 4004
rect 7064 3992 7070 4004
rect 11330 3992 11336 4004
rect 7064 3964 11336 3992
rect 7064 3952 7070 3964
rect 11330 3952 11336 3964
rect 11388 3952 11394 4004
rect 11422 3952 11428 4004
rect 11480 3992 11486 4004
rect 12268 3992 12296 4023
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 13004 4060 13032 4100
rect 13078 4060 13084 4072
rect 12991 4032 13084 4060
rect 13078 4020 13084 4032
rect 13136 4069 13142 4072
rect 13136 4063 13185 4069
rect 13136 4029 13139 4063
rect 13173 4029 13185 4063
rect 13262 4060 13268 4072
rect 13223 4032 13268 4060
rect 13136 4023 13185 4029
rect 13136 4020 13142 4023
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 13357 4063 13415 4069
rect 13357 4029 13369 4063
rect 13403 4060 13415 4063
rect 13446 4060 13452 4072
rect 13403 4032 13452 4060
rect 13403 4029 13415 4032
rect 13357 4023 13415 4029
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 13541 4063 13599 4069
rect 13541 4029 13553 4063
rect 13587 4029 13599 4063
rect 13541 4023 13599 4029
rect 11480 3964 12296 3992
rect 12345 3995 12403 4001
rect 11480 3952 11486 3964
rect 12345 3961 12357 3995
rect 12391 3992 12403 3995
rect 13556 3992 13584 4023
rect 14734 4020 14740 4072
rect 14792 4060 14798 4072
rect 15010 4060 15016 4072
rect 14792 4032 15016 4060
rect 14792 4020 14798 4032
rect 15010 4020 15016 4032
rect 15068 4020 15074 4072
rect 15120 4069 15148 4236
rect 16574 4224 16580 4236
rect 16632 4224 16638 4276
rect 17313 4267 17371 4273
rect 17313 4233 17325 4267
rect 17359 4264 17371 4267
rect 17678 4264 17684 4276
rect 17359 4236 17684 4264
rect 17359 4233 17371 4236
rect 17313 4227 17371 4233
rect 17678 4224 17684 4236
rect 17736 4224 17742 4276
rect 18874 4224 18880 4276
rect 18932 4264 18938 4276
rect 21542 4264 21548 4276
rect 18932 4236 21548 4264
rect 18932 4224 18938 4236
rect 21542 4224 21548 4236
rect 21600 4224 21606 4276
rect 22830 4264 22836 4276
rect 21928 4236 22836 4264
rect 15930 4196 15936 4208
rect 15212 4168 15936 4196
rect 15212 4069 15240 4168
rect 15930 4156 15936 4168
rect 15988 4156 15994 4208
rect 18598 4156 18604 4208
rect 18656 4196 18662 4208
rect 19978 4196 19984 4208
rect 18656 4168 19984 4196
rect 18656 4156 18662 4168
rect 19978 4156 19984 4168
rect 20036 4156 20042 4208
rect 15562 4128 15568 4140
rect 15396 4100 15568 4128
rect 15396 4069 15424 4100
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 18230 4088 18236 4140
rect 18288 4128 18294 4140
rect 18414 4128 18420 4140
rect 18288 4100 18420 4128
rect 18288 4088 18294 4100
rect 18414 4088 18420 4100
rect 18472 4088 18478 4140
rect 18800 4100 20116 4128
rect 18800 4072 18828 4100
rect 15102 4063 15160 4069
rect 15102 4029 15114 4063
rect 15148 4029 15160 4063
rect 15102 4023 15160 4029
rect 15197 4063 15255 4069
rect 15197 4029 15209 4063
rect 15243 4029 15255 4063
rect 15197 4023 15255 4029
rect 15381 4063 15439 4069
rect 15381 4029 15393 4063
rect 15427 4029 15439 4063
rect 15381 4023 15439 4029
rect 15470 4020 15476 4072
rect 15528 4060 15534 4072
rect 15933 4063 15991 4069
rect 15933 4060 15945 4063
rect 15528 4032 15945 4060
rect 15528 4020 15534 4032
rect 15933 4029 15945 4032
rect 15979 4029 15991 4063
rect 15933 4023 15991 4029
rect 16022 4020 16028 4072
rect 16080 4060 16086 4072
rect 16189 4063 16247 4069
rect 16189 4060 16201 4063
rect 16080 4032 16201 4060
rect 16080 4020 16086 4032
rect 16189 4029 16201 4032
rect 16235 4029 16247 4063
rect 16189 4023 16247 4029
rect 16482 4020 16488 4072
rect 16540 4060 16546 4072
rect 18506 4060 18512 4072
rect 16540 4032 18512 4060
rect 16540 4020 16546 4032
rect 18506 4020 18512 4032
rect 18564 4020 18570 4072
rect 18598 4020 18604 4072
rect 18656 4069 18662 4072
rect 18656 4063 18705 4069
rect 18656 4029 18659 4063
rect 18693 4029 18705 4063
rect 18782 4060 18788 4072
rect 18743 4032 18788 4060
rect 18656 4023 18705 4029
rect 18656 4020 18662 4023
rect 18782 4020 18788 4032
rect 18840 4020 18846 4072
rect 18874 4020 18880 4072
rect 18932 4060 18938 4072
rect 19058 4060 19064 4072
rect 18932 4032 18977 4060
rect 19019 4032 19064 4060
rect 18932 4020 18938 4032
rect 19058 4020 19064 4032
rect 19116 4020 19122 4072
rect 19702 4020 19708 4072
rect 19760 4060 19766 4072
rect 19978 4060 19984 4072
rect 19760 4032 19984 4060
rect 19760 4020 19766 4032
rect 19978 4020 19984 4032
rect 20036 4020 20042 4072
rect 20088 4060 20116 4100
rect 20990 4060 20996 4072
rect 20088 4032 20996 4060
rect 20990 4020 20996 4032
rect 21048 4020 21054 4072
rect 21928 4069 21956 4236
rect 22830 4224 22836 4236
rect 22888 4224 22894 4276
rect 23750 4224 23756 4276
rect 23808 4264 23814 4276
rect 24213 4267 24271 4273
rect 24213 4264 24225 4267
rect 23808 4236 24225 4264
rect 23808 4224 23814 4236
rect 24213 4233 24225 4236
rect 24259 4233 24271 4267
rect 24213 4227 24271 4233
rect 26068 4236 27016 4264
rect 22005 4199 22063 4205
rect 22005 4165 22017 4199
rect 22051 4196 22063 4199
rect 23658 4196 23664 4208
rect 22051 4168 23664 4196
rect 22051 4165 22063 4168
rect 22005 4159 22063 4165
rect 23658 4156 23664 4168
rect 23716 4156 23722 4208
rect 25038 4156 25044 4208
rect 25096 4196 25102 4208
rect 25958 4196 25964 4208
rect 25096 4168 25964 4196
rect 25096 4156 25102 4168
rect 25958 4156 25964 4168
rect 26016 4156 26022 4208
rect 22186 4088 22192 4140
rect 22244 4128 22250 4140
rect 23017 4131 23075 4137
rect 23017 4128 23029 4131
rect 22244 4100 23029 4128
rect 22244 4088 22250 4100
rect 23017 4097 23029 4100
rect 23063 4097 23075 4131
rect 23017 4091 23075 4097
rect 21913 4063 21971 4069
rect 21913 4029 21925 4063
rect 21959 4029 21971 4063
rect 21913 4023 21971 4029
rect 22097 4063 22155 4069
rect 22097 4029 22109 4063
rect 22143 4060 22155 4063
rect 22281 4063 22339 4069
rect 22281 4060 22293 4063
rect 22143 4032 22293 4060
rect 22143 4029 22155 4032
rect 22097 4023 22155 4029
rect 22281 4029 22293 4032
rect 22327 4029 22339 4063
rect 22925 4063 22983 4069
rect 22925 4060 22937 4063
rect 22281 4023 22339 4029
rect 22388 4032 22937 4060
rect 22388 4001 22416 4032
rect 22925 4029 22937 4032
rect 22971 4029 22983 4063
rect 23032 4060 23060 4091
rect 23106 4088 23112 4140
rect 23164 4128 23170 4140
rect 23164 4100 23209 4128
rect 23164 4088 23170 4100
rect 23290 4088 23296 4140
rect 23348 4128 23354 4140
rect 26068 4128 26096 4236
rect 26988 4196 27016 4236
rect 27246 4224 27252 4276
rect 27304 4264 27310 4276
rect 27433 4267 27491 4273
rect 27433 4264 27445 4267
rect 27304 4236 27445 4264
rect 27304 4224 27310 4236
rect 27433 4233 27445 4236
rect 27479 4233 27491 4267
rect 27433 4227 27491 4233
rect 26988 4168 27108 4196
rect 23348 4100 26096 4128
rect 27080 4128 27108 4168
rect 28077 4131 28135 4137
rect 28077 4128 28089 4131
rect 27080 4100 28089 4128
rect 23348 4088 23354 4100
rect 28077 4097 28089 4100
rect 28123 4097 28135 4131
rect 28077 4091 28135 4097
rect 23382 4060 23388 4072
rect 23032 4032 23388 4060
rect 22925 4023 22983 4029
rect 23382 4020 23388 4032
rect 23440 4020 23446 4072
rect 23474 4020 23480 4072
rect 23532 4060 23538 4072
rect 24121 4063 24179 4069
rect 24121 4060 24133 4063
rect 23532 4032 24133 4060
rect 23532 4020 23538 4032
rect 24121 4029 24133 4032
rect 24167 4029 24179 4063
rect 26050 4060 26056 4072
rect 26011 4032 26056 4060
rect 24121 4023 24179 4029
rect 26050 4020 26056 4032
rect 26108 4020 26114 4072
rect 26694 4020 26700 4072
rect 26752 4060 26758 4072
rect 27985 4063 28043 4069
rect 27985 4060 27997 4063
rect 26752 4032 27997 4060
rect 26752 4020 26758 4032
rect 27985 4029 27997 4032
rect 28031 4029 28043 4063
rect 27985 4023 28043 4029
rect 12391 3964 13584 3992
rect 18417 3995 18475 4001
rect 12391 3961 12403 3964
rect 12345 3955 12403 3961
rect 18417 3961 18429 3995
rect 18463 3992 18475 3995
rect 20226 3995 20284 4001
rect 20226 3992 20238 3995
rect 18463 3964 20238 3992
rect 18463 3961 18475 3964
rect 18417 3955 18475 3961
rect 20226 3961 20238 3964
rect 20272 3961 20284 3995
rect 22373 3995 22431 4001
rect 22373 3992 22385 3995
rect 20226 3955 20284 3961
rect 20364 3964 22385 3992
rect 2590 3924 2596 3936
rect 2551 3896 2596 3924
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 2866 3884 2872 3936
rect 2924 3924 2930 3936
rect 2961 3927 3019 3933
rect 2961 3924 2973 3927
rect 2924 3896 2973 3924
rect 2924 3884 2930 3896
rect 2961 3893 2973 3896
rect 3007 3893 3019 3927
rect 2961 3887 3019 3893
rect 3053 3927 3111 3933
rect 3053 3893 3065 3927
rect 3099 3924 3111 3927
rect 4154 3924 4160 3936
rect 3099 3896 4160 3924
rect 3099 3893 3111 3896
rect 3053 3887 3111 3893
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 6178 3924 6184 3936
rect 6139 3896 6184 3924
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 6549 3927 6607 3933
rect 6549 3893 6561 3927
rect 6595 3924 6607 3927
rect 8662 3924 8668 3936
rect 6595 3896 8668 3924
rect 6595 3893 6607 3896
rect 6549 3887 6607 3893
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 9582 3924 9588 3936
rect 9543 3896 9588 3924
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 11517 3927 11575 3933
rect 11517 3893 11529 3927
rect 11563 3924 11575 3927
rect 12250 3924 12256 3936
rect 11563 3896 12256 3924
rect 11563 3893 11575 3896
rect 11517 3887 11575 3893
rect 12250 3884 12256 3896
rect 12308 3884 12314 3936
rect 12894 3924 12900 3936
rect 12855 3896 12900 3924
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 14734 3924 14740 3936
rect 14695 3896 14740 3924
rect 14734 3884 14740 3896
rect 14792 3884 14798 3936
rect 14826 3884 14832 3936
rect 14884 3924 14890 3936
rect 20364 3924 20392 3964
rect 22373 3961 22385 3964
rect 22419 3961 22431 3995
rect 23566 3992 23572 4004
rect 22373 3955 22431 3961
rect 22572 3964 23572 3992
rect 14884 3896 20392 3924
rect 14884 3884 14890 3896
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 21361 3927 21419 3933
rect 21361 3924 21373 3927
rect 20680 3896 21373 3924
rect 20680 3884 20686 3896
rect 21361 3893 21373 3896
rect 21407 3893 21419 3927
rect 21361 3887 21419 3893
rect 22281 3927 22339 3933
rect 22281 3893 22293 3927
rect 22327 3924 22339 3927
rect 22462 3924 22468 3936
rect 22327 3896 22468 3924
rect 22327 3893 22339 3896
rect 22281 3887 22339 3893
rect 22462 3884 22468 3896
rect 22520 3884 22526 3936
rect 22572 3933 22600 3964
rect 23566 3952 23572 3964
rect 23624 3952 23630 4004
rect 25409 3995 25467 4001
rect 25409 3961 25421 3995
rect 25455 3992 25467 3995
rect 25455 3964 25820 3992
rect 25455 3961 25467 3964
rect 25409 3955 25467 3961
rect 22557 3927 22615 3933
rect 22557 3893 22569 3927
rect 22603 3893 22615 3927
rect 22557 3887 22615 3893
rect 22646 3884 22652 3936
rect 22704 3924 22710 3936
rect 23198 3924 23204 3936
rect 22704 3896 23204 3924
rect 22704 3884 22710 3896
rect 23198 3884 23204 3896
rect 23256 3884 23262 3936
rect 25498 3924 25504 3936
rect 25459 3896 25504 3924
rect 25498 3884 25504 3896
rect 25556 3884 25562 3936
rect 25792 3924 25820 3964
rect 25866 3952 25872 4004
rect 25924 3992 25930 4004
rect 26298 3995 26356 4001
rect 26298 3992 26310 3995
rect 25924 3964 26310 3992
rect 25924 3952 25930 3964
rect 26298 3961 26310 3964
rect 26344 3961 26356 3995
rect 27890 3992 27896 4004
rect 26298 3955 26356 3961
rect 27080 3964 27896 3992
rect 27080 3924 27108 3964
rect 27890 3952 27896 3964
rect 27948 3952 27954 4004
rect 25792 3896 27108 3924
rect 1104 3834 28888 3856
rect 1104 3782 10246 3834
rect 10298 3782 10310 3834
rect 10362 3782 10374 3834
rect 10426 3782 10438 3834
rect 10490 3782 19510 3834
rect 19562 3782 19574 3834
rect 19626 3782 19638 3834
rect 19690 3782 19702 3834
rect 19754 3782 28888 3834
rect 1104 3760 28888 3782
rect 1670 3720 1676 3732
rect 1631 3692 1676 3720
rect 1670 3680 1676 3692
rect 1728 3680 1734 3732
rect 4154 3720 4160 3732
rect 4067 3692 4160 3720
rect 4154 3680 4160 3692
rect 4212 3720 4218 3732
rect 5074 3720 5080 3732
rect 4212 3692 5080 3720
rect 4212 3680 4218 3692
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 7193 3723 7251 3729
rect 7193 3689 7205 3723
rect 7239 3720 7251 3723
rect 7374 3720 7380 3732
rect 7239 3692 7380 3720
rect 7239 3689 7251 3692
rect 7193 3683 7251 3689
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 10042 3720 10048 3732
rect 7524 3692 10048 3720
rect 7524 3680 7530 3692
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 10689 3723 10747 3729
rect 10689 3689 10701 3723
rect 10735 3720 10747 3723
rect 11974 3720 11980 3732
rect 10735 3692 11980 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 13078 3680 13084 3732
rect 13136 3720 13142 3732
rect 13817 3723 13875 3729
rect 13817 3720 13829 3723
rect 13136 3692 13829 3720
rect 13136 3680 13142 3692
rect 13817 3689 13829 3692
rect 13863 3689 13875 3723
rect 13817 3683 13875 3689
rect 15010 3680 15016 3732
rect 15068 3720 15074 3732
rect 15749 3723 15807 3729
rect 15749 3720 15761 3723
rect 15068 3692 15761 3720
rect 15068 3680 15074 3692
rect 15749 3689 15761 3692
rect 15795 3689 15807 3723
rect 16390 3720 16396 3732
rect 16351 3692 16396 3720
rect 15749 3683 15807 3689
rect 16390 3680 16396 3692
rect 16448 3680 16454 3732
rect 19705 3723 19763 3729
rect 19705 3720 19717 3723
rect 16500 3692 19717 3720
rect 2590 3612 2596 3664
rect 2648 3652 2654 3664
rect 3022 3655 3080 3661
rect 3022 3652 3034 3655
rect 2648 3624 3034 3652
rect 2648 3612 2654 3624
rect 3022 3621 3034 3624
rect 3068 3621 3080 3655
rect 3022 3615 3080 3621
rect 5092 3624 11284 3652
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 4430 3584 4436 3596
rect 1627 3556 4436 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 4430 3544 4436 3556
rect 4488 3544 4494 3596
rect 4982 3584 4988 3596
rect 4943 3556 4988 3584
rect 4982 3544 4988 3556
rect 5040 3544 5046 3596
rect 5092 3593 5120 3624
rect 5077 3587 5135 3593
rect 5077 3553 5089 3587
rect 5123 3553 5135 3587
rect 5077 3547 5135 3553
rect 5445 3587 5503 3593
rect 5445 3553 5457 3587
rect 5491 3584 5503 3587
rect 6270 3584 6276 3596
rect 5491 3556 6276 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 7285 3587 7343 3593
rect 7285 3553 7297 3587
rect 7331 3584 7343 3587
rect 7742 3584 7748 3596
rect 7331 3556 7748 3584
rect 7331 3553 7343 3556
rect 7285 3547 7343 3553
rect 7742 3544 7748 3556
rect 7800 3544 7806 3596
rect 8389 3587 8447 3593
rect 8389 3553 8401 3587
rect 8435 3584 8447 3587
rect 9030 3584 9036 3596
rect 8435 3556 9036 3584
rect 8435 3553 8447 3556
rect 8389 3547 8447 3553
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 9398 3584 9404 3596
rect 9359 3556 9404 3584
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 10594 3584 10600 3596
rect 10555 3556 10600 3584
rect 10594 3544 10600 3556
rect 10652 3544 10658 3596
rect 11256 3584 11284 3624
rect 11330 3612 11336 3664
rect 11388 3652 11394 3664
rect 12704 3655 12762 3661
rect 11388 3624 12480 3652
rect 11388 3612 11394 3624
rect 12342 3584 12348 3596
rect 11256 3556 12348 3584
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 12452 3584 12480 3624
rect 12704 3621 12716 3655
rect 12750 3652 12762 3655
rect 12894 3652 12900 3664
rect 12750 3624 12900 3652
rect 12750 3621 12762 3624
rect 12704 3615 12762 3621
rect 12894 3612 12900 3624
rect 12952 3612 12958 3664
rect 14636 3655 14694 3661
rect 14636 3621 14648 3655
rect 14682 3652 14694 3655
rect 14734 3652 14740 3664
rect 14682 3624 14740 3652
rect 14682 3621 14694 3624
rect 14636 3615 14694 3621
rect 14734 3612 14740 3624
rect 14792 3612 14798 3664
rect 16500 3652 16528 3692
rect 19705 3689 19717 3692
rect 19751 3689 19763 3723
rect 19705 3683 19763 3689
rect 19889 3723 19947 3729
rect 19889 3689 19901 3723
rect 19935 3720 19947 3723
rect 20070 3720 20076 3732
rect 19935 3692 20076 3720
rect 19935 3689 19947 3692
rect 19889 3683 19947 3689
rect 14844 3624 16528 3652
rect 14844 3584 14872 3624
rect 17862 3612 17868 3664
rect 17920 3652 17926 3664
rect 18202 3655 18260 3661
rect 18202 3652 18214 3655
rect 17920 3624 18214 3652
rect 17920 3612 17926 3624
rect 18202 3621 18214 3624
rect 18248 3621 18260 3655
rect 18202 3615 18260 3621
rect 18506 3612 18512 3664
rect 18564 3652 18570 3664
rect 19521 3655 19579 3661
rect 19521 3652 19533 3655
rect 18564 3624 19533 3652
rect 18564 3612 18570 3624
rect 19521 3621 19533 3624
rect 19567 3621 19579 3655
rect 19720 3652 19748 3683
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 20346 3720 20352 3732
rect 20307 3692 20352 3720
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 21269 3723 21327 3729
rect 21269 3689 21281 3723
rect 21315 3720 21327 3723
rect 21634 3720 21640 3732
rect 21315 3692 21640 3720
rect 21315 3689 21327 3692
rect 21269 3683 21327 3689
rect 21634 3680 21640 3692
rect 21692 3680 21698 3732
rect 23198 3680 23204 3732
rect 23256 3720 23262 3732
rect 24578 3720 24584 3732
rect 23256 3692 24584 3720
rect 23256 3680 23262 3692
rect 24578 3680 24584 3692
rect 24636 3680 24642 3732
rect 25314 3720 25320 3732
rect 25275 3692 25320 3720
rect 25314 3680 25320 3692
rect 25372 3680 25378 3732
rect 26786 3720 26792 3732
rect 25608 3692 26004 3720
rect 26747 3692 26792 3720
rect 20257 3655 20315 3661
rect 20257 3652 20269 3655
rect 19720 3624 20269 3652
rect 19521 3615 19579 3621
rect 20257 3621 20269 3624
rect 20303 3621 20315 3655
rect 21910 3652 21916 3664
rect 20257 3615 20315 3621
rect 21100 3624 21916 3652
rect 16206 3584 16212 3596
rect 12452 3556 14872 3584
rect 16167 3556 16212 3584
rect 16206 3544 16212 3556
rect 16264 3544 16270 3596
rect 16393 3587 16451 3593
rect 16393 3553 16405 3587
rect 16439 3584 16451 3587
rect 16666 3584 16672 3596
rect 16439 3556 16672 3584
rect 16439 3553 16451 3556
rect 16393 3547 16451 3553
rect 16666 3544 16672 3556
rect 16724 3544 16730 3596
rect 17313 3587 17371 3593
rect 17313 3553 17325 3587
rect 17359 3584 17371 3587
rect 19978 3584 19984 3596
rect 17359 3556 17908 3584
rect 17359 3553 17371 3556
rect 17313 3547 17371 3553
rect 17880 3528 17908 3556
rect 18064 3556 19984 3584
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3485 2835 3519
rect 2777 3479 2835 3485
rect 7469 3519 7527 3525
rect 7469 3485 7481 3519
rect 7515 3516 7527 3519
rect 7558 3516 7564 3528
rect 7515 3488 7564 3516
rect 7515 3485 7527 3488
rect 7469 3479 7527 3485
rect 2792 3380 2820 3479
rect 7558 3476 7564 3488
rect 7616 3476 7622 3528
rect 8478 3516 8484 3528
rect 8439 3488 8484 3516
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 11330 3516 11336 3528
rect 8588 3488 11336 3516
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 8588 3448 8616 3488
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 11698 3476 11704 3528
rect 11756 3516 11762 3528
rect 11974 3516 11980 3528
rect 11756 3488 11980 3516
rect 11756 3476 11762 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 12066 3476 12072 3528
rect 12124 3516 12130 3528
rect 12434 3516 12440 3528
rect 12124 3488 12440 3516
rect 12124 3476 12130 3488
rect 12434 3476 12440 3488
rect 12492 3516 12498 3528
rect 12492 3488 12537 3516
rect 12492 3476 12498 3488
rect 14090 3476 14096 3528
rect 14148 3516 14154 3528
rect 14369 3519 14427 3525
rect 14369 3516 14381 3519
rect 14148 3488 14381 3516
rect 14148 3476 14154 3488
rect 14369 3485 14381 3488
rect 14415 3485 14427 3519
rect 14369 3479 14427 3485
rect 15654 3476 15660 3528
rect 15712 3516 15718 3528
rect 15712 3488 17540 3516
rect 15712 3476 15718 3488
rect 5500 3420 8616 3448
rect 5500 3408 5506 3420
rect 8662 3408 8668 3460
rect 8720 3448 8726 3460
rect 8757 3451 8815 3457
rect 8757 3448 8769 3451
rect 8720 3420 8769 3448
rect 8720 3408 8726 3420
rect 8757 3417 8769 3420
rect 8803 3417 8815 3451
rect 8757 3411 8815 3417
rect 9493 3451 9551 3457
rect 9493 3417 9505 3451
rect 9539 3448 9551 3451
rect 11422 3448 11428 3460
rect 9539 3420 11428 3448
rect 9539 3417 9551 3420
rect 9493 3411 9551 3417
rect 11422 3408 11428 3420
rect 11480 3408 11486 3460
rect 15838 3408 15844 3460
rect 15896 3448 15902 3460
rect 17405 3451 17463 3457
rect 17405 3448 17417 3451
rect 15896 3420 17417 3448
rect 15896 3408 15902 3420
rect 17405 3417 17417 3420
rect 17451 3417 17463 3451
rect 17405 3411 17463 3417
rect 4890 3380 4896 3392
rect 2792 3352 4896 3380
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 6825 3383 6883 3389
rect 6825 3349 6837 3383
rect 6871 3380 6883 3383
rect 7098 3380 7104 3392
rect 6871 3352 7104 3380
rect 6871 3349 6883 3352
rect 6825 3343 6883 3349
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 17218 3380 17224 3392
rect 11204 3352 17224 3380
rect 11204 3340 11210 3352
rect 17218 3340 17224 3352
rect 17276 3340 17282 3392
rect 17512 3380 17540 3488
rect 17862 3476 17868 3528
rect 17920 3476 17926 3528
rect 17957 3519 18015 3525
rect 17957 3485 17969 3519
rect 18003 3516 18015 3519
rect 18064 3516 18092 3556
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 21100 3593 21128 3624
rect 21910 3612 21916 3624
rect 21968 3612 21974 3664
rect 22649 3655 22707 3661
rect 22649 3621 22661 3655
rect 22695 3652 22707 3655
rect 25608 3652 25636 3692
rect 22695 3624 25636 3652
rect 22695 3621 22707 3624
rect 22649 3615 22707 3621
rect 21085 3587 21143 3593
rect 21085 3553 21097 3587
rect 21131 3553 21143 3587
rect 21269 3587 21327 3593
rect 21269 3584 21281 3587
rect 21085 3547 21143 3553
rect 21264 3553 21281 3584
rect 21315 3584 21327 3587
rect 21315 3556 22508 3584
rect 21315 3553 21327 3556
rect 21264 3547 21327 3553
rect 18003 3488 18092 3516
rect 18003 3485 18015 3488
rect 17957 3479 18015 3485
rect 19242 3476 19248 3528
rect 19300 3516 19306 3528
rect 20441 3519 20499 3525
rect 20441 3516 20453 3519
rect 19300 3488 20453 3516
rect 19300 3476 19306 3488
rect 20441 3485 20453 3488
rect 20487 3485 20499 3519
rect 20441 3479 20499 3485
rect 21264 3448 21292 3547
rect 22480 3528 22508 3556
rect 22554 3544 22560 3596
rect 22612 3584 22618 3596
rect 22741 3587 22799 3593
rect 22612 3556 22657 3584
rect 22612 3544 22618 3556
rect 22741 3553 22753 3587
rect 22787 3553 22799 3587
rect 22741 3547 22799 3553
rect 22462 3476 22468 3528
rect 22520 3516 22526 3528
rect 22756 3516 22784 3547
rect 22922 3544 22928 3596
rect 22980 3584 22986 3596
rect 23457 3587 23515 3593
rect 23457 3584 23469 3587
rect 22980 3556 23469 3584
rect 22980 3544 22986 3556
rect 23457 3553 23469 3556
rect 23503 3553 23515 3587
rect 23457 3547 23515 3553
rect 25406 3544 25412 3596
rect 25464 3584 25470 3596
rect 25547 3587 25605 3593
rect 25547 3584 25559 3587
rect 25464 3556 25559 3584
rect 25464 3544 25470 3556
rect 25547 3553 25559 3556
rect 25593 3553 25605 3587
rect 25547 3547 25605 3553
rect 25666 3587 25724 3593
rect 25666 3553 25678 3587
rect 25712 3553 25724 3587
rect 25666 3547 25724 3553
rect 22520 3488 22784 3516
rect 22520 3476 22526 3488
rect 22830 3476 22836 3528
rect 22888 3516 22894 3528
rect 23201 3519 23259 3525
rect 23201 3516 23213 3519
rect 22888 3488 23213 3516
rect 22888 3476 22894 3488
rect 23201 3485 23213 3488
rect 23247 3485 23259 3519
rect 23201 3479 23259 3485
rect 25130 3476 25136 3528
rect 25188 3516 25194 3528
rect 25680 3516 25708 3547
rect 25774 3544 25780 3596
rect 25832 3593 25838 3596
rect 25976 3593 26004 3692
rect 26786 3680 26792 3692
rect 26844 3680 26850 3732
rect 27985 3655 28043 3661
rect 27985 3652 27997 3655
rect 26206 3624 27997 3652
rect 25832 3584 25840 3593
rect 25961 3587 26019 3593
rect 25832 3556 25877 3584
rect 25832 3547 25840 3556
rect 25961 3553 25973 3587
rect 26007 3553 26019 3587
rect 26206 3584 26234 3624
rect 27985 3621 27997 3624
rect 28031 3621 28043 3655
rect 27985 3615 28043 3621
rect 25961 3547 26019 3553
rect 26068 3556 26234 3584
rect 26697 3587 26755 3593
rect 25832 3544 25838 3547
rect 25188 3488 25708 3516
rect 25188 3476 25194 3488
rect 26068 3448 26096 3556
rect 26697 3553 26709 3587
rect 26743 3553 26755 3587
rect 26697 3547 26755 3553
rect 26142 3476 26148 3528
rect 26200 3516 26206 3528
rect 26712 3516 26740 3547
rect 26200 3488 26740 3516
rect 26200 3476 26206 3488
rect 18892 3420 21292 3448
rect 24136 3420 26096 3448
rect 18892 3380 18920 3420
rect 17512 3352 18920 3380
rect 19242 3340 19248 3392
rect 19300 3380 19306 3392
rect 19337 3383 19395 3389
rect 19337 3380 19349 3383
rect 19300 3352 19349 3380
rect 19300 3340 19306 3352
rect 19337 3349 19349 3352
rect 19383 3349 19395 3383
rect 19337 3343 19395 3349
rect 19521 3383 19579 3389
rect 19521 3349 19533 3383
rect 19567 3380 19579 3383
rect 24136 3380 24164 3420
rect 26418 3408 26424 3460
rect 26476 3448 26482 3460
rect 28166 3448 28172 3460
rect 26476 3420 28028 3448
rect 28127 3420 28172 3448
rect 26476 3408 26482 3420
rect 19567 3352 24164 3380
rect 19567 3349 19579 3352
rect 19521 3343 19579 3349
rect 24486 3340 24492 3392
rect 24544 3380 24550 3392
rect 27890 3380 27896 3392
rect 24544 3352 27896 3380
rect 24544 3340 24550 3352
rect 27890 3340 27896 3352
rect 27948 3340 27954 3392
rect 28000 3380 28028 3420
rect 28166 3408 28172 3420
rect 28224 3408 28230 3460
rect 29270 3380 29276 3392
rect 28000 3352 29276 3380
rect 29270 3340 29276 3352
rect 29328 3340 29334 3392
rect 1104 3290 28888 3312
rect 1104 3238 5614 3290
rect 5666 3238 5678 3290
rect 5730 3238 5742 3290
rect 5794 3238 5806 3290
rect 5858 3238 14878 3290
rect 14930 3238 14942 3290
rect 14994 3238 15006 3290
rect 15058 3238 15070 3290
rect 15122 3238 24142 3290
rect 24194 3238 24206 3290
rect 24258 3238 24270 3290
rect 24322 3238 24334 3290
rect 24386 3238 28888 3290
rect 1104 3216 28888 3238
rect 2866 3176 2872 3188
rect 2827 3148 2872 3176
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 10873 3179 10931 3185
rect 5092 3148 10824 3176
rect 1857 3111 1915 3117
rect 1857 3077 1869 3111
rect 1903 3108 1915 3111
rect 5092 3108 5120 3148
rect 1903 3080 5120 3108
rect 6457 3111 6515 3117
rect 1903 3077 1915 3080
rect 1857 3071 1915 3077
rect 6457 3077 6469 3111
rect 6503 3108 6515 3111
rect 6638 3108 6644 3120
rect 6503 3080 6644 3108
rect 6503 3077 6515 3080
rect 6457 3071 6515 3077
rect 6638 3068 6644 3080
rect 6696 3068 6702 3120
rect 10796 3108 10824 3148
rect 10873 3145 10885 3179
rect 10919 3176 10931 3179
rect 11606 3176 11612 3188
rect 10919 3148 11612 3176
rect 10919 3145 10931 3148
rect 10873 3139 10931 3145
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 11790 3136 11796 3188
rect 11848 3176 11854 3188
rect 12805 3179 12863 3185
rect 12805 3176 12817 3179
rect 11848 3148 12817 3176
rect 11848 3136 11854 3148
rect 12805 3145 12817 3148
rect 12851 3145 12863 3179
rect 12805 3139 12863 3145
rect 13541 3179 13599 3185
rect 13541 3145 13553 3179
rect 13587 3176 13599 3179
rect 15562 3176 15568 3188
rect 13587 3148 15568 3176
rect 13587 3145 13599 3148
rect 13541 3139 13599 3145
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 16298 3136 16304 3188
rect 16356 3176 16362 3188
rect 16393 3179 16451 3185
rect 16393 3176 16405 3179
rect 16356 3148 16405 3176
rect 16356 3136 16362 3148
rect 16393 3145 16405 3148
rect 16439 3145 16451 3179
rect 17034 3176 17040 3188
rect 16995 3148 17040 3176
rect 16393 3139 16451 3145
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 27433 3179 27491 3185
rect 17276 3148 26234 3176
rect 17276 3136 17282 3148
rect 11146 3108 11152 3120
rect 10796 3080 11152 3108
rect 11146 3068 11152 3080
rect 11204 3068 11210 3120
rect 11517 3111 11575 3117
rect 11517 3077 11529 3111
rect 11563 3108 11575 3111
rect 12618 3108 12624 3120
rect 11563 3080 12624 3108
rect 11563 3077 11575 3080
rect 11517 3071 11575 3077
rect 12618 3068 12624 3080
rect 12676 3068 12682 3120
rect 12894 3068 12900 3120
rect 12952 3108 12958 3120
rect 15746 3108 15752 3120
rect 12952 3080 15752 3108
rect 12952 3068 12958 3080
rect 15746 3068 15752 3080
rect 15804 3068 15810 3120
rect 16206 3068 16212 3120
rect 16264 3108 16270 3120
rect 18969 3111 19027 3117
rect 18969 3108 18981 3111
rect 16264 3080 18981 3108
rect 16264 3068 16270 3080
rect 18969 3077 18981 3080
rect 19015 3108 19027 3111
rect 19150 3108 19156 3120
rect 19015 3080 19156 3108
rect 19015 3077 19027 3080
rect 18969 3071 19027 3077
rect 19150 3068 19156 3080
rect 19208 3068 19214 3120
rect 19886 3068 19892 3120
rect 19944 3108 19950 3120
rect 20073 3111 20131 3117
rect 20073 3108 20085 3111
rect 19944 3080 20085 3108
rect 19944 3068 19950 3080
rect 20073 3077 20085 3080
rect 20119 3077 20131 3111
rect 22370 3108 22376 3120
rect 22331 3080 22376 3108
rect 20073 3071 20131 3077
rect 22370 3068 22376 3080
rect 22428 3068 22434 3120
rect 22922 3108 22928 3120
rect 22883 3080 22928 3108
rect 22922 3068 22928 3080
rect 22980 3068 22986 3120
rect 23014 3068 23020 3120
rect 23072 3108 23078 3120
rect 25130 3108 25136 3120
rect 23072 3080 25136 3108
rect 23072 3068 23078 3080
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 2958 3040 2964 3052
rect 2639 3012 2964 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 4890 3000 4896 3052
rect 4948 3040 4954 3052
rect 5077 3043 5135 3049
rect 5077 3040 5089 3043
rect 4948 3012 5089 3040
rect 4948 3000 4954 3012
rect 5077 3009 5089 3012
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 7009 3043 7067 3049
rect 7009 3040 7021 3043
rect 6972 3012 7021 3040
rect 6972 3000 6978 3012
rect 7009 3009 7021 3012
rect 7055 3009 7067 3043
rect 12158 3040 12164 3052
rect 12119 3012 12164 3040
rect 7009 3003 7067 3009
rect 12158 3000 12164 3012
rect 12216 3000 12222 3052
rect 13354 3000 13360 3052
rect 13412 3040 13418 3052
rect 13725 3043 13783 3049
rect 13725 3040 13737 3043
rect 13412 3012 13737 3040
rect 13412 3000 13418 3012
rect 13725 3009 13737 3012
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 15194 3000 15200 3052
rect 15252 3040 15258 3052
rect 15381 3043 15439 3049
rect 15381 3040 15393 3043
rect 15252 3012 15393 3040
rect 15252 3000 15258 3012
rect 15381 3009 15393 3012
rect 15427 3009 15439 3043
rect 17678 3040 17684 3052
rect 17639 3012 17684 3040
rect 15381 3003 15439 3009
rect 17678 3000 17684 3012
rect 17736 3000 17742 3052
rect 20162 3040 20168 3052
rect 18248 3012 20168 3040
rect 1670 2972 1676 2984
rect 1631 2944 1676 2972
rect 1670 2932 1676 2944
rect 1728 2932 1734 2984
rect 2501 2975 2559 2981
rect 2501 2941 2513 2975
rect 2547 2972 2559 2975
rect 3142 2972 3148 2984
rect 2547 2944 3148 2972
rect 2547 2941 2559 2944
rect 2501 2935 2559 2941
rect 3142 2932 3148 2944
rect 3200 2932 3206 2984
rect 3510 2932 3516 2984
rect 3568 2972 3574 2984
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 3568 2944 4261 2972
rect 3568 2932 3574 2944
rect 4249 2941 4261 2944
rect 4295 2941 4307 2975
rect 4249 2935 4307 2941
rect 5344 2975 5402 2981
rect 5344 2941 5356 2975
rect 5390 2972 5402 2975
rect 6178 2972 6184 2984
rect 5390 2944 6184 2972
rect 5390 2941 5402 2944
rect 5344 2935 5402 2941
rect 6178 2932 6184 2944
rect 6236 2932 6242 2984
rect 7098 2932 7104 2984
rect 7156 2972 7162 2984
rect 7265 2975 7323 2981
rect 7265 2972 7277 2975
rect 7156 2944 7277 2972
rect 7156 2932 7162 2944
rect 7265 2941 7277 2944
rect 7311 2941 7323 2975
rect 7265 2935 7323 2941
rect 7558 2932 7564 2984
rect 7616 2972 7622 2984
rect 9493 2975 9551 2981
rect 9493 2972 9505 2975
rect 7616 2944 9505 2972
rect 7616 2932 7622 2944
rect 9493 2941 9505 2944
rect 9539 2941 9551 2975
rect 9493 2935 9551 2941
rect 9582 2932 9588 2984
rect 9640 2972 9646 2984
rect 9749 2975 9807 2981
rect 9749 2972 9761 2975
rect 9640 2944 9761 2972
rect 9640 2932 9646 2944
rect 9749 2941 9761 2944
rect 9795 2941 9807 2975
rect 9749 2935 9807 2941
rect 10042 2932 10048 2984
rect 10100 2972 10106 2984
rect 12713 2975 12771 2981
rect 10100 2944 12434 2972
rect 10100 2932 10106 2944
rect 4341 2907 4399 2913
rect 4341 2873 4353 2907
rect 4387 2904 4399 2907
rect 11885 2907 11943 2913
rect 11885 2904 11897 2907
rect 4387 2876 11897 2904
rect 4387 2873 4399 2876
rect 4341 2867 4399 2873
rect 11885 2873 11897 2876
rect 11931 2873 11943 2907
rect 12406 2904 12434 2944
rect 12713 2941 12725 2975
rect 12759 2972 12771 2975
rect 13541 2975 13599 2981
rect 13541 2972 13553 2975
rect 12759 2944 13553 2972
rect 12759 2941 12771 2944
rect 12713 2935 12771 2941
rect 13541 2941 13553 2944
rect 13587 2941 13599 2975
rect 13541 2935 13599 2941
rect 13633 2975 13691 2981
rect 13633 2941 13645 2975
rect 13679 2972 13691 2975
rect 16206 2972 16212 2984
rect 13679 2944 16212 2972
rect 13679 2941 13691 2944
rect 13633 2935 13691 2941
rect 16206 2932 16212 2944
rect 16264 2932 16270 2984
rect 16301 2975 16359 2981
rect 16301 2941 16313 2975
rect 16347 2972 16359 2975
rect 17310 2972 17316 2984
rect 16347 2944 17316 2972
rect 16347 2941 16359 2944
rect 16301 2935 16359 2941
rect 17310 2932 17316 2944
rect 17368 2932 17374 2984
rect 18248 2981 18276 3012
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 18233 2975 18291 2981
rect 18233 2941 18245 2975
rect 18279 2941 18291 2975
rect 18233 2935 18291 2941
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2972 18383 2975
rect 18414 2972 18420 2984
rect 18371 2944 18420 2972
rect 18371 2941 18383 2944
rect 18325 2935 18383 2941
rect 18414 2932 18420 2944
rect 18472 2932 18478 2984
rect 18877 2975 18935 2981
rect 18877 2941 18889 2975
rect 18923 2972 18935 2975
rect 19334 2972 19340 2984
rect 18923 2944 19340 2972
rect 18923 2941 18935 2944
rect 18877 2935 18935 2941
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 19978 2972 19984 2984
rect 19939 2944 19984 2972
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 20070 2932 20076 2984
rect 20128 2972 20134 2984
rect 20993 2975 21051 2981
rect 20993 2972 21005 2975
rect 20128 2944 21005 2972
rect 20128 2932 20134 2944
rect 20993 2941 21005 2944
rect 21039 2941 21051 2975
rect 20993 2935 21051 2941
rect 21082 2932 21088 2984
rect 21140 2972 21146 2984
rect 21249 2975 21307 2981
rect 21249 2972 21261 2975
rect 21140 2944 21261 2972
rect 21140 2932 21146 2944
rect 21249 2941 21261 2944
rect 21295 2941 21307 2975
rect 21249 2935 21307 2941
rect 23106 2932 23112 2984
rect 23164 2981 23170 2984
rect 23308 2981 23336 3080
rect 25130 3068 25136 3080
rect 25188 3068 25194 3120
rect 25317 3111 25375 3117
rect 25317 3077 25329 3111
rect 25363 3108 25375 3111
rect 25866 3108 25872 3120
rect 25363 3080 25872 3108
rect 25363 3077 25375 3080
rect 25317 3071 25375 3077
rect 25866 3068 25872 3080
rect 25924 3068 25930 3120
rect 25148 3040 25176 3068
rect 25148 3012 25708 3040
rect 23164 2975 23213 2981
rect 23164 2941 23167 2975
rect 23201 2941 23213 2975
rect 23164 2935 23213 2941
rect 23293 2975 23351 2981
rect 23293 2941 23305 2975
rect 23339 2941 23351 2975
rect 23293 2935 23351 2941
rect 23385 2975 23443 2981
rect 23385 2941 23397 2975
rect 23431 2972 23443 2975
rect 23569 2975 23627 2981
rect 23431 2944 23500 2972
rect 23431 2941 23443 2944
rect 23385 2935 23443 2941
rect 23164 2932 23170 2935
rect 15197 2907 15255 2913
rect 15197 2904 15209 2907
rect 12406 2876 15209 2904
rect 11885 2867 11943 2873
rect 15197 2873 15209 2876
rect 15243 2873 15255 2907
rect 15197 2867 15255 2873
rect 17126 2864 17132 2916
rect 17184 2904 17190 2916
rect 17405 2907 17463 2913
rect 17405 2904 17417 2907
rect 17184 2876 17417 2904
rect 17184 2864 17190 2876
rect 17405 2873 17417 2876
rect 17451 2873 17463 2907
rect 17405 2867 17463 2873
rect 17497 2907 17555 2913
rect 17497 2873 17509 2907
rect 17543 2904 17555 2907
rect 21910 2904 21916 2916
rect 17543 2876 21916 2904
rect 17543 2873 17555 2876
rect 17497 2867 17555 2873
rect 21910 2864 21916 2876
rect 21968 2864 21974 2916
rect 22002 2864 22008 2916
rect 22060 2904 22066 2916
rect 23014 2904 23020 2916
rect 22060 2876 23020 2904
rect 22060 2864 22066 2876
rect 23014 2864 23020 2876
rect 23072 2864 23078 2916
rect 6914 2796 6920 2848
rect 6972 2836 6978 2848
rect 7558 2836 7564 2848
rect 6972 2808 7564 2836
rect 6972 2796 6978 2808
rect 7558 2796 7564 2808
rect 7616 2796 7622 2848
rect 7742 2796 7748 2848
rect 7800 2836 7806 2848
rect 8389 2839 8447 2845
rect 8389 2836 8401 2839
rect 7800 2808 8401 2836
rect 7800 2796 7806 2808
rect 8389 2805 8401 2808
rect 8435 2805 8447 2839
rect 11974 2836 11980 2848
rect 11935 2808 11980 2836
rect 8389 2799 8447 2805
rect 11974 2796 11980 2808
rect 12032 2796 12038 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 14090 2836 14096 2848
rect 12492 2808 14096 2836
rect 12492 2796 12498 2808
rect 14090 2796 14096 2808
rect 14148 2796 14154 2848
rect 14829 2839 14887 2845
rect 14829 2805 14841 2839
rect 14875 2836 14887 2839
rect 15102 2836 15108 2848
rect 14875 2808 15108 2836
rect 14875 2805 14887 2808
rect 14829 2799 14887 2805
rect 15102 2796 15108 2808
rect 15160 2796 15166 2848
rect 15289 2839 15347 2845
rect 15289 2805 15301 2839
rect 15335 2836 15347 2839
rect 15378 2836 15384 2848
rect 15335 2808 15384 2836
rect 15335 2805 15347 2808
rect 15289 2799 15347 2805
rect 15378 2796 15384 2808
rect 15436 2836 15442 2848
rect 21358 2836 21364 2848
rect 15436 2808 21364 2836
rect 15436 2796 15442 2808
rect 21358 2796 21364 2808
rect 21416 2796 21422 2848
rect 21542 2796 21548 2848
rect 21600 2836 21606 2848
rect 23472 2836 23500 2944
rect 23569 2941 23581 2975
rect 23615 2972 23627 2975
rect 23658 2972 23664 2984
rect 23615 2944 23664 2972
rect 23615 2941 23627 2944
rect 23569 2935 23627 2941
rect 23658 2932 23664 2944
rect 23716 2932 23722 2984
rect 25680 2981 25708 3012
rect 25573 2975 25631 2981
rect 25573 2941 25585 2975
rect 25619 2941 25631 2975
rect 25573 2935 25631 2941
rect 25666 2975 25724 2981
rect 25666 2941 25678 2975
rect 25712 2941 25724 2975
rect 25666 2935 25724 2941
rect 23934 2864 23940 2916
rect 23992 2904 23998 2916
rect 24121 2907 24179 2913
rect 24121 2904 24133 2907
rect 23992 2876 24133 2904
rect 23992 2864 23998 2876
rect 24121 2873 24133 2876
rect 24167 2904 24179 2907
rect 24486 2904 24492 2916
rect 24167 2876 24492 2904
rect 24167 2873 24179 2876
rect 24121 2867 24179 2873
rect 24486 2864 24492 2876
rect 24544 2864 24550 2916
rect 21600 2808 23500 2836
rect 24213 2839 24271 2845
rect 21600 2796 21606 2808
rect 24213 2805 24225 2839
rect 24259 2836 24271 2839
rect 24762 2836 24768 2848
rect 24259 2808 24768 2836
rect 24259 2805 24271 2808
rect 24213 2799 24271 2805
rect 24762 2796 24768 2808
rect 24820 2796 24826 2848
rect 25599 2836 25627 2935
rect 25774 2932 25780 2984
rect 25832 2981 25838 2984
rect 25832 2972 25840 2981
rect 25832 2944 25877 2972
rect 25832 2935 25840 2944
rect 25832 2932 25838 2935
rect 25958 2932 25964 2984
rect 26016 2972 26022 2984
rect 26206 2972 26234 3148
rect 27433 3145 27445 3179
rect 27479 3176 27491 3179
rect 27522 3176 27528 3188
rect 27479 3148 27528 3176
rect 27479 3145 27491 3148
rect 27433 3139 27491 3145
rect 27522 3136 27528 3148
rect 27580 3136 27586 3188
rect 27246 3068 27252 3120
rect 27304 3108 27310 3120
rect 27304 3080 28028 3108
rect 27304 3068 27310 3080
rect 27890 3040 27896 3052
rect 27851 3012 27896 3040
rect 27890 3000 27896 3012
rect 27948 3000 27954 3052
rect 28000 3049 28028 3080
rect 27985 3043 28043 3049
rect 27985 3009 27997 3043
rect 28031 3009 28043 3043
rect 27985 3003 28043 3009
rect 27801 2975 27859 2981
rect 27801 2972 27813 2975
rect 26016 2944 26061 2972
rect 26206 2944 27813 2972
rect 26016 2932 26022 2944
rect 27801 2941 27813 2944
rect 27847 2941 27859 2975
rect 27801 2935 27859 2941
rect 26786 2904 26792 2916
rect 26747 2876 26792 2904
rect 26786 2864 26792 2876
rect 26844 2864 26850 2916
rect 26970 2904 26976 2916
rect 26931 2876 26976 2904
rect 26970 2864 26976 2876
rect 27028 2864 27034 2916
rect 27246 2836 27252 2848
rect 25599 2808 27252 2836
rect 27246 2796 27252 2808
rect 27304 2796 27310 2848
rect 27338 2796 27344 2848
rect 27396 2836 27402 2848
rect 27890 2836 27896 2848
rect 27396 2808 27896 2836
rect 27396 2796 27402 2808
rect 27890 2796 27896 2808
rect 27948 2796 27954 2848
rect 1104 2746 28888 2768
rect 1104 2694 10246 2746
rect 10298 2694 10310 2746
rect 10362 2694 10374 2746
rect 10426 2694 10438 2746
rect 10490 2694 19510 2746
rect 19562 2694 19574 2746
rect 19626 2694 19638 2746
rect 19690 2694 19702 2746
rect 19754 2694 28888 2746
rect 1104 2672 28888 2694
rect 4341 2635 4399 2641
rect 4341 2601 4353 2635
rect 4387 2632 4399 2635
rect 4522 2632 4528 2644
rect 4387 2604 4528 2632
rect 4387 2601 4399 2604
rect 4341 2595 4399 2601
rect 4522 2592 4528 2604
rect 4580 2592 4586 2644
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 5077 2635 5135 2641
rect 5077 2632 5089 2635
rect 5040 2604 5089 2632
rect 5040 2592 5046 2604
rect 5077 2601 5089 2604
rect 5123 2601 5135 2635
rect 8389 2635 8447 2641
rect 8389 2632 8401 2635
rect 5077 2595 5135 2601
rect 6886 2604 8401 2632
rect 6886 2564 6914 2604
rect 8389 2601 8401 2604
rect 8435 2601 8447 2635
rect 8389 2595 8447 2601
rect 9398 2592 9404 2644
rect 9456 2632 9462 2644
rect 9585 2635 9643 2641
rect 9585 2632 9597 2635
rect 9456 2604 9597 2632
rect 9456 2592 9462 2604
rect 9585 2601 9597 2604
rect 9631 2601 9643 2635
rect 9585 2595 9643 2601
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 10594 2632 10600 2644
rect 10275 2604 10600 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10594 2592 10600 2604
rect 10652 2592 10658 2644
rect 11241 2635 11299 2641
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 11974 2632 11980 2644
rect 11287 2604 11980 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12158 2592 12164 2644
rect 12216 2632 12222 2644
rect 12345 2635 12403 2641
rect 12345 2632 12357 2635
rect 12216 2604 12357 2632
rect 12216 2592 12222 2604
rect 12345 2601 12357 2604
rect 12391 2601 12403 2635
rect 12345 2595 12403 2601
rect 13538 2592 13544 2644
rect 13596 2632 13602 2644
rect 15013 2635 15071 2641
rect 15013 2632 15025 2635
rect 13596 2604 15025 2632
rect 13596 2592 13602 2604
rect 15013 2601 15025 2604
rect 15059 2601 15071 2635
rect 15562 2632 15568 2644
rect 15523 2604 15568 2632
rect 15013 2595 15071 2601
rect 15562 2592 15568 2604
rect 15620 2592 15626 2644
rect 16206 2632 16212 2644
rect 16167 2604 16212 2632
rect 16206 2592 16212 2604
rect 16264 2592 16270 2644
rect 17310 2592 17316 2644
rect 17368 2632 17374 2644
rect 18233 2635 18291 2641
rect 18233 2632 18245 2635
rect 17368 2604 18245 2632
rect 17368 2592 17374 2604
rect 18233 2601 18245 2604
rect 18279 2601 18291 2635
rect 18233 2595 18291 2601
rect 19978 2592 19984 2644
rect 20036 2632 20042 2644
rect 20257 2635 20315 2641
rect 20257 2632 20269 2635
rect 20036 2604 20269 2632
rect 20036 2592 20042 2604
rect 20257 2601 20269 2604
rect 20303 2601 20315 2635
rect 20257 2595 20315 2601
rect 20901 2635 20959 2641
rect 20901 2601 20913 2635
rect 20947 2601 20959 2635
rect 20901 2595 20959 2601
rect 4264 2536 6914 2564
rect 7929 2567 7987 2573
rect 658 2456 664 2508
rect 716 2496 722 2508
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 716 2468 1869 2496
rect 716 2456 722 2468
rect 1857 2465 1869 2468
rect 1903 2465 1915 2499
rect 2590 2496 2596 2508
rect 2551 2468 2596 2496
rect 1857 2459 1915 2465
rect 2590 2456 2596 2468
rect 2648 2456 2654 2508
rect 4264 2505 4292 2536
rect 7929 2533 7941 2567
rect 7975 2564 7987 2567
rect 12710 2564 12716 2576
rect 7975 2536 12716 2564
rect 7975 2533 7987 2536
rect 7929 2527 7987 2533
rect 12710 2524 12716 2536
rect 12768 2524 12774 2576
rect 14274 2524 14280 2576
rect 14332 2564 14338 2576
rect 20916 2564 20944 2595
rect 21358 2592 21364 2644
rect 21416 2632 21422 2644
rect 21416 2604 26464 2632
rect 21416 2592 21422 2604
rect 14332 2536 16436 2564
rect 20916 2536 21588 2564
rect 14332 2524 14338 2536
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2465 4307 2499
rect 4249 2459 4307 2465
rect 4893 2499 4951 2505
rect 4893 2465 4905 2499
rect 4939 2465 4951 2499
rect 4893 2459 4951 2465
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 6086 2496 6092 2508
rect 5767 2468 6092 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2777 2431 2835 2437
rect 2777 2428 2789 2431
rect 2004 2400 2789 2428
rect 2004 2388 2010 2400
rect 2777 2397 2789 2400
rect 2823 2397 2835 2431
rect 2777 2391 2835 2397
rect 3326 2388 3332 2440
rect 3384 2428 3390 2440
rect 4908 2428 4936 2459
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 7466 2456 7472 2508
rect 7524 2496 7530 2508
rect 7561 2499 7619 2505
rect 7561 2496 7573 2499
rect 7524 2468 7573 2496
rect 7524 2456 7530 2468
rect 7561 2465 7573 2468
rect 7607 2465 7619 2499
rect 8570 2496 8576 2508
rect 8531 2468 8576 2496
rect 7561 2459 7619 2465
rect 8570 2456 8576 2468
rect 8628 2456 8634 2508
rect 8754 2456 8760 2508
rect 8812 2496 8818 2508
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 8812 2468 9781 2496
rect 8812 2456 8818 2468
rect 9769 2465 9781 2468
rect 9815 2465 9827 2499
rect 9769 2459 9827 2465
rect 10134 2456 10140 2508
rect 10192 2496 10198 2508
rect 10413 2499 10471 2505
rect 10413 2496 10425 2499
rect 10192 2468 10425 2496
rect 10192 2456 10198 2468
rect 10413 2465 10425 2468
rect 10459 2465 10471 2499
rect 11146 2496 11152 2508
rect 11107 2468 11152 2496
rect 10413 2459 10471 2465
rect 11146 2456 11152 2468
rect 11204 2456 11210 2508
rect 12250 2496 12256 2508
rect 12211 2468 12256 2496
rect 12250 2456 12256 2468
rect 12308 2456 12314 2508
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 12584 2468 12909 2496
rect 12584 2456 12590 2468
rect 12897 2465 12909 2468
rect 12943 2465 12955 2499
rect 12897 2459 12955 2465
rect 13817 2499 13875 2505
rect 13817 2465 13829 2499
rect 13863 2496 13875 2499
rect 14642 2496 14648 2508
rect 13863 2468 14648 2496
rect 13863 2465 13875 2468
rect 13817 2459 13875 2465
rect 14642 2456 14648 2468
rect 14700 2456 14706 2508
rect 14921 2499 14979 2505
rect 14921 2465 14933 2499
rect 14967 2465 14979 2499
rect 15746 2496 15752 2508
rect 15707 2468 15752 2496
rect 14921 2459 14979 2465
rect 11882 2428 11888 2440
rect 3384 2400 4936 2428
rect 6886 2400 11888 2428
rect 3384 2388 3390 2400
rect 2041 2363 2099 2369
rect 2041 2329 2053 2363
rect 2087 2360 2099 2363
rect 5905 2363 5963 2369
rect 2087 2332 4476 2360
rect 2087 2329 2099 2332
rect 2041 2323 2099 2329
rect 4448 2292 4476 2332
rect 5905 2329 5917 2363
rect 5951 2360 5963 2363
rect 6886 2360 6914 2400
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 7926 2360 7932 2372
rect 5951 2332 6914 2360
rect 7392 2332 7932 2360
rect 5951 2329 5963 2332
rect 5905 2323 5963 2329
rect 7392 2292 7420 2332
rect 7926 2320 7932 2332
rect 7984 2320 7990 2372
rect 14936 2360 14964 2459
rect 15746 2456 15752 2468
rect 15804 2456 15810 2508
rect 16408 2505 16436 2536
rect 16393 2499 16451 2505
rect 16393 2465 16405 2499
rect 16439 2465 16451 2499
rect 17773 2499 17831 2505
rect 17773 2496 17785 2499
rect 16393 2459 16451 2465
rect 16500 2468 17785 2496
rect 15654 2388 15660 2440
rect 15712 2428 15718 2440
rect 16500 2428 16528 2468
rect 17773 2465 17785 2468
rect 17819 2465 17831 2499
rect 17773 2459 17831 2465
rect 18417 2499 18475 2505
rect 18417 2465 18429 2499
rect 18463 2465 18475 2499
rect 19334 2496 19340 2508
rect 19295 2468 19340 2496
rect 18417 2459 18475 2465
rect 15712 2400 16528 2428
rect 15712 2388 15718 2400
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 18432 2428 18460 2459
rect 19334 2456 19340 2468
rect 19392 2456 19398 2508
rect 20438 2496 20444 2508
rect 20399 2468 20444 2496
rect 20438 2456 20444 2468
rect 20496 2456 20502 2508
rect 21560 2505 21588 2536
rect 21634 2524 21640 2576
rect 21692 2564 21698 2576
rect 26436 2573 26464 2604
rect 23109 2567 23167 2573
rect 21692 2536 21737 2564
rect 21692 2524 21698 2536
rect 23109 2533 23121 2567
rect 23155 2564 23167 2567
rect 25685 2567 25743 2573
rect 25685 2564 25697 2567
rect 23155 2536 25697 2564
rect 23155 2533 23167 2536
rect 23109 2527 23167 2533
rect 25685 2533 25697 2536
rect 25731 2533 25743 2567
rect 25685 2527 25743 2533
rect 26421 2567 26479 2573
rect 26421 2533 26433 2567
rect 26467 2533 26479 2567
rect 26421 2527 26479 2533
rect 21093 2499 21151 2505
rect 21093 2465 21105 2499
rect 21139 2496 21151 2499
rect 21545 2499 21603 2505
rect 21139 2468 21496 2496
rect 21139 2465 21151 2468
rect 21093 2459 21151 2465
rect 21358 2428 21364 2440
rect 17000 2400 18460 2428
rect 19306 2400 21364 2428
rect 17000 2388 17006 2400
rect 17589 2363 17647 2369
rect 17589 2360 17601 2363
rect 14936 2332 17601 2360
rect 17589 2329 17601 2332
rect 17635 2329 17647 2363
rect 19306 2360 19334 2400
rect 21358 2388 21364 2400
rect 21416 2388 21422 2440
rect 21468 2428 21496 2468
rect 21545 2465 21557 2499
rect 21591 2465 21603 2499
rect 23014 2496 23020 2508
rect 22975 2468 23020 2496
rect 21545 2459 21603 2465
rect 23014 2456 23020 2468
rect 23072 2456 23078 2508
rect 23382 2456 23388 2508
rect 23440 2496 23446 2508
rect 23753 2499 23811 2505
rect 23753 2496 23765 2499
rect 23440 2468 23765 2496
rect 23440 2456 23446 2468
rect 23753 2465 23765 2468
rect 23799 2465 23811 2499
rect 24486 2496 24492 2508
rect 24447 2468 24492 2496
rect 23753 2459 23811 2465
rect 24486 2456 24492 2468
rect 24544 2456 24550 2508
rect 27154 2496 27160 2508
rect 27115 2468 27160 2496
rect 27154 2456 27160 2468
rect 27212 2456 27218 2508
rect 22462 2428 22468 2440
rect 21468 2400 22468 2428
rect 22462 2388 22468 2400
rect 22520 2388 22526 2440
rect 25222 2428 25228 2440
rect 23860 2400 25228 2428
rect 17589 2323 17647 2329
rect 17972 2332 19334 2360
rect 12986 2292 12992 2304
rect 4448 2264 7420 2292
rect 12947 2264 12992 2292
rect 12986 2252 12992 2264
rect 13044 2252 13050 2304
rect 13909 2295 13967 2301
rect 13909 2261 13921 2295
rect 13955 2292 13967 2295
rect 17972 2292 18000 2332
rect 13955 2264 18000 2292
rect 19153 2295 19211 2301
rect 13955 2261 13967 2264
rect 13909 2255 13967 2261
rect 19153 2261 19165 2295
rect 19199 2292 19211 2295
rect 23860 2292 23888 2400
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 23937 2363 23995 2369
rect 23937 2329 23949 2363
rect 23983 2360 23995 2363
rect 25038 2360 25044 2372
rect 23983 2332 25044 2360
rect 23983 2329 23995 2332
rect 23937 2323 23995 2329
rect 25038 2320 25044 2332
rect 25096 2320 25102 2372
rect 25866 2360 25872 2372
rect 25827 2332 25872 2360
rect 25866 2320 25872 2332
rect 25924 2320 25930 2372
rect 26050 2320 26056 2372
rect 26108 2360 26114 2372
rect 27341 2363 27399 2369
rect 27341 2360 27353 2363
rect 26108 2332 27353 2360
rect 26108 2320 26114 2332
rect 27341 2329 27353 2332
rect 27387 2329 27399 2363
rect 27341 2323 27399 2329
rect 19199 2264 23888 2292
rect 24581 2295 24639 2301
rect 19199 2261 19211 2264
rect 19153 2255 19211 2261
rect 24581 2261 24593 2295
rect 24627 2292 24639 2295
rect 25406 2292 25412 2304
rect 24627 2264 25412 2292
rect 24627 2261 24639 2264
rect 24581 2255 24639 2261
rect 25406 2252 25412 2264
rect 25464 2252 25470 2304
rect 26142 2252 26148 2304
rect 26200 2292 26206 2304
rect 26513 2295 26571 2301
rect 26513 2292 26525 2295
rect 26200 2264 26525 2292
rect 26200 2252 26206 2264
rect 26513 2261 26525 2264
rect 26559 2261 26571 2295
rect 26513 2255 26571 2261
rect 1104 2202 28888 2224
rect 1104 2150 5614 2202
rect 5666 2150 5678 2202
rect 5730 2150 5742 2202
rect 5794 2150 5806 2202
rect 5858 2150 14878 2202
rect 14930 2150 14942 2202
rect 14994 2150 15006 2202
rect 15058 2150 15070 2202
rect 15122 2150 24142 2202
rect 24194 2150 24206 2202
rect 24258 2150 24270 2202
rect 24322 2150 24334 2202
rect 24386 2150 28888 2202
rect 1104 2128 28888 2150
rect 2590 2048 2596 2100
rect 2648 2088 2654 2100
rect 2648 2060 12434 2088
rect 2648 2048 2654 2060
rect 3510 1980 3516 2032
rect 3568 2020 3574 2032
rect 6822 2020 6828 2032
rect 3568 1992 6828 2020
rect 3568 1980 3574 1992
rect 6822 1980 6828 1992
rect 6880 1980 6886 2032
rect 2774 1912 2780 1964
rect 2832 1952 2838 1964
rect 5902 1952 5908 1964
rect 2832 1924 5908 1952
rect 2832 1912 2838 1924
rect 5902 1912 5908 1924
rect 5960 1912 5966 1964
rect 12406 1952 12434 2060
rect 19334 2048 19340 2100
rect 19392 2088 19398 2100
rect 26510 2088 26516 2100
rect 19392 2060 26516 2088
rect 19392 2048 19398 2060
rect 26510 2048 26516 2060
rect 26568 2048 26574 2100
rect 12986 1980 12992 2032
rect 13044 2020 13050 2032
rect 27154 2020 27160 2032
rect 13044 1992 27160 2020
rect 13044 1980 13050 1992
rect 27154 1980 27160 1992
rect 27212 1980 27218 2032
rect 25590 1952 25596 1964
rect 12406 1924 25596 1952
rect 25590 1912 25596 1924
rect 25648 1912 25654 1964
rect 3418 1844 3424 1896
rect 3476 1884 3482 1896
rect 7650 1884 7656 1896
rect 3476 1856 7656 1884
rect 3476 1844 3482 1856
rect 7650 1844 7656 1856
rect 7708 1844 7714 1896
rect 20438 1232 20444 1284
rect 20496 1272 20502 1284
rect 23750 1272 23756 1284
rect 20496 1244 23756 1272
rect 20496 1232 20502 1244
rect 23750 1232 23756 1244
rect 23808 1232 23814 1284
rect 2958 1028 2964 1080
rect 3016 1068 3022 1080
rect 8570 1068 8576 1080
rect 3016 1040 8576 1068
rect 3016 1028 3022 1040
rect 8570 1028 8576 1040
rect 8628 1028 8634 1080
<< via1 >>
rect 3884 54000 3936 54052
rect 5908 54000 5960 54052
rect 24032 53864 24084 53916
rect 25044 53864 25096 53916
rect 20720 53728 20772 53780
rect 27068 53728 27120 53780
rect 19156 53660 19208 53712
rect 26700 53660 26752 53712
rect 20904 53592 20956 53644
rect 25688 53592 25740 53644
rect 23204 53524 23256 53576
rect 25504 53524 25556 53576
rect 22836 53456 22888 53508
rect 24860 53456 24912 53508
rect 21180 53388 21232 53440
rect 27252 53388 27304 53440
rect 5614 53286 5666 53338
rect 5678 53286 5730 53338
rect 5742 53286 5794 53338
rect 5806 53286 5858 53338
rect 14878 53286 14930 53338
rect 14942 53286 14994 53338
rect 15006 53286 15058 53338
rect 15070 53286 15122 53338
rect 24142 53286 24194 53338
rect 24206 53286 24258 53338
rect 24270 53286 24322 53338
rect 24334 53286 24386 53338
rect 4344 53184 4396 53236
rect 6092 53184 6144 53236
rect 7840 53184 7892 53236
rect 9588 53184 9640 53236
rect 11428 53184 11480 53236
rect 13176 53184 13228 53236
rect 18420 53184 18472 53236
rect 19156 53227 19208 53236
rect 19156 53193 19165 53227
rect 19165 53193 19199 53227
rect 19199 53193 19208 53227
rect 19156 53184 19208 53193
rect 20168 53184 20220 53236
rect 21180 53227 21232 53236
rect 21180 53193 21189 53227
rect 21189 53193 21223 53227
rect 21223 53193 21232 53227
rect 21180 53184 21232 53193
rect 23204 53227 23256 53236
rect 23204 53193 23213 53227
rect 23213 53193 23247 53227
rect 23247 53193 23256 53227
rect 23204 53184 23256 53193
rect 23756 53184 23808 53236
rect 2596 53116 2648 53168
rect 15200 53159 15252 53168
rect 15200 53125 15209 53159
rect 15209 53125 15243 53159
rect 15243 53125 15252 53159
rect 15200 53116 15252 53125
rect 16672 53159 16724 53168
rect 16672 53125 16681 53159
rect 16681 53125 16715 53159
rect 16715 53125 16724 53159
rect 16672 53116 16724 53125
rect 22008 53159 22060 53168
rect 22008 53125 22017 53159
rect 22017 53125 22051 53159
rect 22051 53125 22060 53159
rect 22008 53116 22060 53125
rect 2780 53048 2832 53100
rect 4068 53048 4120 53100
rect 5356 52980 5408 53032
rect 24032 53048 24084 53100
rect 23296 52980 23348 53032
rect 27896 53184 27948 53236
rect 27988 53116 28040 53168
rect 24860 53048 24912 53100
rect 27252 53048 27304 53100
rect 24584 52980 24636 53032
rect 25780 53023 25832 53032
rect 25780 52989 25789 53023
rect 25789 52989 25823 53023
rect 25823 52989 25832 53023
rect 25780 52980 25832 52989
rect 27068 53023 27120 53032
rect 27068 52989 27077 53023
rect 27077 52989 27111 53023
rect 27111 52989 27120 53023
rect 27068 52980 27120 52989
rect 3976 52912 4028 52964
rect 5816 52955 5868 52964
rect 2044 52844 2096 52896
rect 2872 52887 2924 52896
rect 2872 52853 2881 52887
rect 2881 52853 2915 52887
rect 2915 52853 2924 52887
rect 2872 52844 2924 52853
rect 5816 52921 5825 52955
rect 5825 52921 5859 52955
rect 5859 52921 5868 52955
rect 5816 52912 5868 52921
rect 7012 52955 7064 52964
rect 7012 52921 7021 52955
rect 7021 52921 7055 52955
rect 7055 52921 7064 52955
rect 7012 52912 7064 52921
rect 7840 52912 7892 52964
rect 9956 52912 10008 52964
rect 12072 52912 12124 52964
rect 13268 52955 13320 52964
rect 13268 52921 13277 52955
rect 13277 52921 13311 52955
rect 13311 52921 13320 52955
rect 13268 52912 13320 52921
rect 14372 52912 14424 52964
rect 16488 52955 16540 52964
rect 16488 52921 16497 52955
rect 16497 52921 16531 52955
rect 16531 52921 16540 52955
rect 16488 52912 16540 52921
rect 18512 52955 18564 52964
rect 18512 52921 18521 52955
rect 18521 52921 18555 52955
rect 18555 52921 18564 52955
rect 18512 52912 18564 52921
rect 20352 52955 20404 52964
rect 20352 52921 20361 52955
rect 20361 52921 20395 52955
rect 20395 52921 20404 52955
rect 20352 52912 20404 52921
rect 11520 52844 11572 52896
rect 21640 52912 21692 52964
rect 22100 52912 22152 52964
rect 23756 52912 23808 52964
rect 22008 52844 22060 52896
rect 22652 52844 22704 52896
rect 26240 52912 26292 52964
rect 26608 52912 26660 52964
rect 24676 52844 24728 52896
rect 24768 52844 24820 52896
rect 25504 52844 25556 52896
rect 26424 52887 26476 52896
rect 26424 52853 26433 52887
rect 26433 52853 26467 52887
rect 26467 52853 26476 52887
rect 26424 52844 26476 52853
rect 27160 52887 27212 52896
rect 27160 52853 27169 52887
rect 27169 52853 27203 52887
rect 27203 52853 27212 52887
rect 27160 52844 27212 52853
rect 10246 52742 10298 52794
rect 10310 52742 10362 52794
rect 10374 52742 10426 52794
rect 10438 52742 10490 52794
rect 19510 52742 19562 52794
rect 19574 52742 19626 52794
rect 19638 52742 19690 52794
rect 19702 52742 19754 52794
rect 22652 52683 22704 52692
rect 22652 52649 22661 52683
rect 22661 52649 22695 52683
rect 22695 52649 22704 52683
rect 22652 52640 22704 52649
rect 23296 52683 23348 52692
rect 23296 52649 23305 52683
rect 23305 52649 23339 52683
rect 23339 52649 23348 52683
rect 23296 52640 23348 52649
rect 26516 52640 26568 52692
rect 1860 52547 1912 52556
rect 1860 52513 1869 52547
rect 1869 52513 1903 52547
rect 1903 52513 1912 52547
rect 1860 52504 1912 52513
rect 2596 52547 2648 52556
rect 2596 52513 2605 52547
rect 2605 52513 2639 52547
rect 2639 52513 2648 52547
rect 2596 52504 2648 52513
rect 4068 52547 4120 52556
rect 4068 52513 4102 52547
rect 4102 52513 4120 52547
rect 4068 52504 4120 52513
rect 5172 52504 5224 52556
rect 7564 52504 7616 52556
rect 2780 52479 2832 52488
rect 2780 52445 2789 52479
rect 2789 52445 2823 52479
rect 2823 52445 2832 52479
rect 3792 52479 3844 52488
rect 2780 52436 2832 52445
rect 3792 52445 3801 52479
rect 3801 52445 3835 52479
rect 3835 52445 3844 52479
rect 3792 52436 3844 52445
rect 8024 52436 8076 52488
rect 848 52368 900 52420
rect 2872 52368 2924 52420
rect 9680 52368 9732 52420
rect 11612 52368 11664 52420
rect 14096 52504 14148 52556
rect 18236 52547 18288 52556
rect 18236 52513 18270 52547
rect 18270 52513 18288 52547
rect 20260 52547 20312 52556
rect 18236 52504 18288 52513
rect 20260 52513 20269 52547
rect 20269 52513 20303 52547
rect 20303 52513 20312 52547
rect 20260 52504 20312 52513
rect 20904 52547 20956 52556
rect 20904 52513 20913 52547
rect 20913 52513 20947 52547
rect 20947 52513 20956 52547
rect 20904 52504 20956 52513
rect 21364 52547 21416 52556
rect 21364 52513 21373 52547
rect 21373 52513 21407 52547
rect 21407 52513 21416 52547
rect 21364 52504 21416 52513
rect 22836 52547 22888 52556
rect 22836 52513 22845 52547
rect 22845 52513 22879 52547
rect 22879 52513 22888 52547
rect 22836 52504 22888 52513
rect 12716 52436 12768 52488
rect 12992 52436 13044 52488
rect 16120 52436 16172 52488
rect 21456 52479 21508 52488
rect 21456 52445 21465 52479
rect 21465 52445 21499 52479
rect 21499 52445 21508 52479
rect 21456 52436 21508 52445
rect 24860 52572 24912 52624
rect 24676 52504 24728 52556
rect 25044 52504 25096 52556
rect 24492 52436 24544 52488
rect 27528 52572 27580 52624
rect 27896 52615 27948 52624
rect 27896 52581 27905 52615
rect 27905 52581 27939 52615
rect 27939 52581 27948 52615
rect 27896 52572 27948 52581
rect 25412 52547 25464 52556
rect 25412 52513 25421 52547
rect 25421 52513 25455 52547
rect 25455 52513 25464 52547
rect 25412 52504 25464 52513
rect 25504 52504 25556 52556
rect 26240 52504 26292 52556
rect 26332 52436 26384 52488
rect 27620 52436 27672 52488
rect 1952 52343 2004 52352
rect 1952 52309 1961 52343
rect 1961 52309 1995 52343
rect 1995 52309 2004 52343
rect 1952 52300 2004 52309
rect 5172 52343 5224 52352
rect 5172 52309 5181 52343
rect 5181 52309 5215 52343
rect 5215 52309 5224 52343
rect 5172 52300 5224 52309
rect 6552 52300 6604 52352
rect 7748 52343 7800 52352
rect 7748 52309 7757 52343
rect 7757 52309 7791 52343
rect 7791 52309 7800 52343
rect 7748 52300 7800 52309
rect 8300 52343 8352 52352
rect 8300 52309 8309 52343
rect 8309 52309 8343 52343
rect 8343 52309 8352 52343
rect 8300 52300 8352 52309
rect 8392 52300 8444 52352
rect 19340 52343 19392 52352
rect 19340 52309 19349 52343
rect 19349 52309 19383 52343
rect 19383 52309 19392 52343
rect 19340 52300 19392 52309
rect 20720 52343 20772 52352
rect 20720 52309 20729 52343
rect 20729 52309 20763 52343
rect 20763 52309 20772 52343
rect 20720 52300 20772 52309
rect 26056 52343 26108 52352
rect 26056 52309 26065 52343
rect 26065 52309 26099 52343
rect 26099 52309 26108 52343
rect 26056 52300 26108 52309
rect 5614 52198 5666 52250
rect 5678 52198 5730 52250
rect 5742 52198 5794 52250
rect 5806 52198 5858 52250
rect 14878 52198 14930 52250
rect 14942 52198 14994 52250
rect 15006 52198 15058 52250
rect 15070 52198 15122 52250
rect 24142 52198 24194 52250
rect 24206 52198 24258 52250
rect 24270 52198 24322 52250
rect 24334 52198 24386 52250
rect 2596 52096 2648 52148
rect 3608 52028 3660 52080
rect 2780 52003 2832 52012
rect 2780 51969 2789 52003
rect 2789 51969 2823 52003
rect 2823 51969 2832 52003
rect 2780 51960 2832 51969
rect 6000 51935 6052 51944
rect 6000 51901 6009 51935
rect 6009 51901 6043 51935
rect 6043 51901 6052 51935
rect 6000 51892 6052 51901
rect 6368 51935 6420 51944
rect 6368 51901 6377 51935
rect 6377 51901 6411 51935
rect 6411 51901 6420 51935
rect 6368 51892 6420 51901
rect 2688 51824 2740 51876
rect 1492 51756 1544 51808
rect 7564 51824 7616 51876
rect 8116 51960 8168 52012
rect 8484 51960 8536 52012
rect 10600 52028 10652 52080
rect 7748 51892 7800 51944
rect 9772 51935 9824 51944
rect 7932 51824 7984 51876
rect 9772 51901 9781 51935
rect 9781 51901 9815 51935
rect 9815 51901 9824 51935
rect 9772 51892 9824 51901
rect 11244 51824 11296 51876
rect 22928 52028 22980 52080
rect 11612 52003 11664 52012
rect 11612 51969 11621 52003
rect 11621 51969 11655 52003
rect 11655 51969 11664 52003
rect 11612 51960 11664 51969
rect 12164 51892 12216 51944
rect 14648 51960 14700 52012
rect 15476 51960 15528 52012
rect 16120 52003 16172 52012
rect 16120 51969 16129 52003
rect 16129 51969 16163 52003
rect 16163 51969 16172 52003
rect 16120 51960 16172 51969
rect 13820 51824 13872 51876
rect 8208 51756 8260 51808
rect 9588 51756 9640 51808
rect 10784 51756 10836 51808
rect 13636 51756 13688 51808
rect 14740 51799 14792 51808
rect 14740 51765 14749 51799
rect 14749 51765 14783 51799
rect 14783 51765 14792 51799
rect 14740 51756 14792 51765
rect 15108 51799 15160 51808
rect 15108 51765 15117 51799
rect 15117 51765 15151 51799
rect 15151 51765 15160 51799
rect 15108 51756 15160 51765
rect 21824 51935 21876 51944
rect 21824 51901 21833 51935
rect 21833 51901 21867 51935
rect 21867 51901 21876 51935
rect 21824 51892 21876 51901
rect 23848 52028 23900 52080
rect 29000 52028 29052 52080
rect 16396 51867 16448 51876
rect 16396 51833 16430 51867
rect 16430 51833 16448 51867
rect 16396 51824 16448 51833
rect 17500 51799 17552 51808
rect 17500 51765 17509 51799
rect 17509 51765 17543 51799
rect 17543 51765 17552 51799
rect 17500 51756 17552 51765
rect 20444 51824 20496 51876
rect 22560 51824 22612 51876
rect 24492 51892 24544 51944
rect 26516 51935 26568 51944
rect 26516 51901 26525 51935
rect 26525 51901 26559 51935
rect 26559 51901 26568 51935
rect 26516 51892 26568 51901
rect 27252 51935 27304 51944
rect 27252 51901 27261 51935
rect 27261 51901 27295 51935
rect 27295 51901 27304 51935
rect 27252 51892 27304 51901
rect 27528 51892 27580 51944
rect 23940 51824 23992 51876
rect 26424 51824 26476 51876
rect 20812 51756 20864 51808
rect 21364 51799 21416 51808
rect 21364 51765 21373 51799
rect 21373 51765 21407 51799
rect 21407 51765 21416 51799
rect 21364 51756 21416 51765
rect 23388 51756 23440 51808
rect 25872 51799 25924 51808
rect 25872 51765 25881 51799
rect 25881 51765 25915 51799
rect 25915 51765 25924 51799
rect 25872 51756 25924 51765
rect 28080 51799 28132 51808
rect 28080 51765 28089 51799
rect 28089 51765 28123 51799
rect 28123 51765 28132 51799
rect 28080 51756 28132 51765
rect 10246 51654 10298 51706
rect 10310 51654 10362 51706
rect 10374 51654 10426 51706
rect 10438 51654 10490 51706
rect 19510 51654 19562 51706
rect 19574 51654 19626 51706
rect 19638 51654 19690 51706
rect 19702 51654 19754 51706
rect 3424 51595 3476 51604
rect 3424 51561 3433 51595
rect 3433 51561 3467 51595
rect 3467 51561 3476 51595
rect 3424 51552 3476 51561
rect 4068 51552 4120 51604
rect 5172 51552 5224 51604
rect 5908 51552 5960 51604
rect 6552 51552 6604 51604
rect 8116 51552 8168 51604
rect 10600 51552 10652 51604
rect 10784 51595 10836 51604
rect 10784 51561 10793 51595
rect 10793 51561 10827 51595
rect 10827 51561 10836 51595
rect 10784 51552 10836 51561
rect 12532 51552 12584 51604
rect 12348 51484 12400 51536
rect 1860 51459 1912 51468
rect 1860 51425 1869 51459
rect 1869 51425 1903 51459
rect 1903 51425 1912 51459
rect 1860 51416 1912 51425
rect 3332 51459 3384 51468
rect 3332 51425 3341 51459
rect 3341 51425 3375 51459
rect 3375 51425 3384 51459
rect 3332 51416 3384 51425
rect 6368 51416 6420 51468
rect 7656 51416 7708 51468
rect 7932 51416 7984 51468
rect 8208 51416 8260 51468
rect 8484 51416 8536 51468
rect 9864 51416 9916 51468
rect 10784 51416 10836 51468
rect 11888 51416 11940 51468
rect 15108 51552 15160 51604
rect 14740 51484 14792 51536
rect 13636 51459 13688 51468
rect 13636 51425 13645 51459
rect 13645 51425 13679 51459
rect 13679 51425 13688 51459
rect 13636 51416 13688 51425
rect 18236 51552 18288 51604
rect 20444 51595 20496 51604
rect 20444 51561 20453 51595
rect 20453 51561 20487 51595
rect 20487 51561 20496 51595
rect 20444 51552 20496 51561
rect 20812 51595 20864 51604
rect 20812 51561 20821 51595
rect 20821 51561 20855 51595
rect 20855 51561 20864 51595
rect 20812 51552 20864 51561
rect 22560 51595 22612 51604
rect 22560 51561 22569 51595
rect 22569 51561 22603 51595
rect 22603 51561 22612 51595
rect 22560 51552 22612 51561
rect 22928 51595 22980 51604
rect 22928 51561 22937 51595
rect 22937 51561 22971 51595
rect 22971 51561 22980 51595
rect 22928 51552 22980 51561
rect 23112 51552 23164 51604
rect 26056 51552 26108 51604
rect 15844 51484 15896 51536
rect 19340 51416 19392 51468
rect 22376 51416 22428 51468
rect 23940 51416 23992 51468
rect 24032 51416 24084 51468
rect 26700 51459 26752 51468
rect 26700 51425 26709 51459
rect 26709 51425 26743 51459
rect 26743 51425 26752 51459
rect 26700 51416 26752 51425
rect 27988 51459 28040 51468
rect 27988 51425 27997 51459
rect 27997 51425 28031 51459
rect 28031 51425 28040 51459
rect 27988 51416 28040 51425
rect 2780 51323 2832 51332
rect 2780 51289 2789 51323
rect 2789 51289 2823 51323
rect 2823 51289 2832 51323
rect 5172 51348 5224 51400
rect 10968 51391 11020 51400
rect 10968 51357 10977 51391
rect 10977 51357 11011 51391
rect 11011 51357 11020 51391
rect 10968 51348 11020 51357
rect 12164 51348 12216 51400
rect 12808 51348 12860 51400
rect 12992 51348 13044 51400
rect 13176 51348 13228 51400
rect 14096 51348 14148 51400
rect 18788 51391 18840 51400
rect 18788 51357 18797 51391
rect 18797 51357 18831 51391
rect 18831 51357 18840 51391
rect 18788 51348 18840 51357
rect 18880 51391 18932 51400
rect 18880 51357 18889 51391
rect 18889 51357 18923 51391
rect 18923 51357 18932 51391
rect 20904 51391 20956 51400
rect 18880 51348 18932 51357
rect 20904 51357 20913 51391
rect 20913 51357 20947 51391
rect 20947 51357 20956 51391
rect 20904 51348 20956 51357
rect 21364 51348 21416 51400
rect 23020 51391 23072 51400
rect 2780 51280 2832 51289
rect 12716 51280 12768 51332
rect 1400 51212 1452 51264
rect 5908 51212 5960 51264
rect 8576 51212 8628 51264
rect 9680 51255 9732 51264
rect 9680 51221 9689 51255
rect 9689 51221 9723 51255
rect 9723 51221 9732 51255
rect 9680 51212 9732 51221
rect 12440 51212 12492 51264
rect 13912 51212 13964 51264
rect 16304 51255 16356 51264
rect 16304 51221 16313 51255
rect 16313 51221 16347 51255
rect 16347 51221 16356 51255
rect 16304 51212 16356 51221
rect 19616 51255 19668 51264
rect 19616 51221 19625 51255
rect 19625 51221 19659 51255
rect 19659 51221 19668 51255
rect 19616 51212 19668 51221
rect 21824 51280 21876 51332
rect 23020 51357 23029 51391
rect 23029 51357 23063 51391
rect 23063 51357 23072 51391
rect 23020 51348 23072 51357
rect 22376 51212 22428 51264
rect 23940 51212 23992 51264
rect 25688 51212 25740 51264
rect 26792 51255 26844 51264
rect 26792 51221 26801 51255
rect 26801 51221 26835 51255
rect 26835 51221 26844 51255
rect 26792 51212 26844 51221
rect 5614 51110 5666 51162
rect 5678 51110 5730 51162
rect 5742 51110 5794 51162
rect 5806 51110 5858 51162
rect 14878 51110 14930 51162
rect 14942 51110 14994 51162
rect 15006 51110 15058 51162
rect 15070 51110 15122 51162
rect 24142 51110 24194 51162
rect 24206 51110 24258 51162
rect 24270 51110 24322 51162
rect 24334 51110 24386 51162
rect 3240 51008 3292 51060
rect 2964 50940 3016 50992
rect 23112 51008 23164 51060
rect 23204 51008 23256 51060
rect 2596 50779 2648 50788
rect 2596 50745 2605 50779
rect 2605 50745 2639 50779
rect 2639 50745 2648 50779
rect 2596 50736 2648 50745
rect 1952 50711 2004 50720
rect 1952 50677 1961 50711
rect 1961 50677 1995 50711
rect 1995 50677 2004 50711
rect 1952 50668 2004 50677
rect 5908 50940 5960 50992
rect 5816 50847 5868 50856
rect 5816 50813 5825 50847
rect 5825 50813 5859 50847
rect 5859 50813 5868 50847
rect 5816 50804 5868 50813
rect 11336 50940 11388 50992
rect 9496 50872 9548 50924
rect 10968 50872 11020 50924
rect 12532 50940 12584 50992
rect 12716 50872 12768 50924
rect 16396 50940 16448 50992
rect 17224 50940 17276 50992
rect 22468 50940 22520 50992
rect 6828 50804 6880 50856
rect 7104 50804 7156 50856
rect 7564 50804 7616 50856
rect 12440 50804 12492 50856
rect 12992 50847 13044 50856
rect 12992 50813 13001 50847
rect 13001 50813 13035 50847
rect 13035 50813 13044 50847
rect 12992 50804 13044 50813
rect 13084 50804 13136 50856
rect 13728 50804 13780 50856
rect 16304 50804 16356 50856
rect 17500 50804 17552 50856
rect 18420 50872 18472 50924
rect 18328 50804 18380 50856
rect 18880 50804 18932 50856
rect 19616 50804 19668 50856
rect 21456 50804 21508 50856
rect 22192 50804 22244 50856
rect 23572 50940 23624 50992
rect 23480 50872 23532 50924
rect 23940 51008 23992 51060
rect 25320 51008 25372 51060
rect 27344 51051 27396 51060
rect 27344 51017 27353 51051
rect 27353 51017 27387 51051
rect 27387 51017 27396 51051
rect 27344 51008 27396 51017
rect 26608 50872 26660 50924
rect 23388 50847 23440 50856
rect 23388 50813 23397 50847
rect 23397 50813 23431 50847
rect 23431 50813 23440 50847
rect 23388 50804 23440 50813
rect 25688 50804 25740 50856
rect 26056 50847 26108 50856
rect 26056 50813 26065 50847
rect 26065 50813 26099 50847
rect 26099 50813 26108 50847
rect 26056 50804 26108 50813
rect 26700 50847 26752 50856
rect 26700 50813 26709 50847
rect 26709 50813 26743 50847
rect 26743 50813 26752 50847
rect 26700 50804 26752 50813
rect 5540 50736 5592 50788
rect 6000 50736 6052 50788
rect 6460 50736 6512 50788
rect 8116 50779 8168 50788
rect 8116 50745 8125 50779
rect 8125 50745 8159 50779
rect 8159 50745 8168 50779
rect 8116 50736 8168 50745
rect 22284 50736 22336 50788
rect 26332 50736 26384 50788
rect 27436 50736 27488 50788
rect 8300 50711 8352 50720
rect 8300 50677 8309 50711
rect 8309 50677 8343 50711
rect 8343 50677 8352 50711
rect 8300 50668 8352 50677
rect 9220 50668 9272 50720
rect 11796 50711 11848 50720
rect 11796 50677 11805 50711
rect 11805 50677 11839 50711
rect 11839 50677 11848 50711
rect 11796 50668 11848 50677
rect 14188 50668 14240 50720
rect 14280 50668 14332 50720
rect 15292 50711 15344 50720
rect 15292 50677 15301 50711
rect 15301 50677 15335 50711
rect 15335 50677 15344 50711
rect 15292 50668 15344 50677
rect 16856 50668 16908 50720
rect 18236 50668 18288 50720
rect 19984 50711 20036 50720
rect 19984 50677 19993 50711
rect 19993 50677 20027 50711
rect 20027 50677 20036 50711
rect 19984 50668 20036 50677
rect 20076 50668 20128 50720
rect 21272 50668 21324 50720
rect 21824 50668 21876 50720
rect 22928 50668 22980 50720
rect 23112 50668 23164 50720
rect 24124 50668 24176 50720
rect 25872 50711 25924 50720
rect 25872 50677 25881 50711
rect 25881 50677 25915 50711
rect 25915 50677 25924 50711
rect 25872 50668 25924 50677
rect 27160 50668 27212 50720
rect 28080 50711 28132 50720
rect 28080 50677 28089 50711
rect 28089 50677 28123 50711
rect 28123 50677 28132 50711
rect 28080 50668 28132 50677
rect 10246 50566 10298 50618
rect 10310 50566 10362 50618
rect 10374 50566 10426 50618
rect 10438 50566 10490 50618
rect 19510 50566 19562 50618
rect 19574 50566 19626 50618
rect 19638 50566 19690 50618
rect 19702 50566 19754 50618
rect 3148 50464 3200 50516
rect 8116 50464 8168 50516
rect 9772 50464 9824 50516
rect 11796 50464 11848 50516
rect 14188 50507 14240 50516
rect 14188 50473 14197 50507
rect 14197 50473 14231 50507
rect 14231 50473 14240 50507
rect 14188 50464 14240 50473
rect 14280 50507 14332 50516
rect 14280 50473 14289 50507
rect 14289 50473 14323 50507
rect 14323 50473 14332 50507
rect 18236 50507 18288 50516
rect 14280 50464 14332 50473
rect 18236 50473 18245 50507
rect 18245 50473 18279 50507
rect 18279 50473 18288 50507
rect 18236 50464 18288 50473
rect 21272 50507 21324 50516
rect 17224 50396 17276 50448
rect 2504 50328 2556 50380
rect 5540 50371 5592 50380
rect 5540 50337 5549 50371
rect 5549 50337 5583 50371
rect 5583 50337 5592 50371
rect 5540 50328 5592 50337
rect 6092 50328 6144 50380
rect 6368 50328 6420 50380
rect 7104 50371 7156 50380
rect 7104 50337 7113 50371
rect 7113 50337 7147 50371
rect 7147 50337 7156 50371
rect 7104 50328 7156 50337
rect 7564 50371 7616 50380
rect 7564 50337 7573 50371
rect 7573 50337 7607 50371
rect 7607 50337 7616 50371
rect 7564 50328 7616 50337
rect 8024 50371 8076 50380
rect 8024 50337 8033 50371
rect 8033 50337 8067 50371
rect 8067 50337 8076 50371
rect 8024 50328 8076 50337
rect 8300 50328 8352 50380
rect 9220 50371 9272 50380
rect 9220 50337 9229 50371
rect 9229 50337 9263 50371
rect 9263 50337 9272 50371
rect 9220 50328 9272 50337
rect 9496 50371 9548 50380
rect 9496 50337 9505 50371
rect 9505 50337 9539 50371
rect 9539 50337 9548 50371
rect 9496 50328 9548 50337
rect 9864 50328 9916 50380
rect 16396 50371 16448 50380
rect 2780 50235 2832 50244
rect 2780 50201 2789 50235
rect 2789 50201 2823 50235
rect 2823 50201 2832 50235
rect 7656 50303 7708 50312
rect 7656 50269 7665 50303
rect 7665 50269 7699 50303
rect 7699 50269 7708 50303
rect 7656 50260 7708 50269
rect 11980 50260 12032 50312
rect 12624 50260 12676 50312
rect 16396 50337 16405 50371
rect 16405 50337 16439 50371
rect 16439 50337 16448 50371
rect 16396 50328 16448 50337
rect 16856 50260 16908 50312
rect 19248 50328 19300 50380
rect 19984 50396 20036 50448
rect 21272 50473 21281 50507
rect 21281 50473 21315 50507
rect 21315 50473 21324 50507
rect 21272 50464 21324 50473
rect 22192 50464 22244 50516
rect 23204 50464 23256 50516
rect 21916 50396 21968 50448
rect 18420 50303 18472 50312
rect 18420 50269 18429 50303
rect 18429 50269 18463 50303
rect 18463 50269 18472 50303
rect 18420 50260 18472 50269
rect 18512 50260 18564 50312
rect 2780 50192 2832 50201
rect 1400 50124 1452 50176
rect 11060 50124 11112 50176
rect 13636 50124 13688 50176
rect 16304 50167 16356 50176
rect 16304 50133 16313 50167
rect 16313 50133 16347 50167
rect 16347 50133 16356 50167
rect 16304 50124 16356 50133
rect 17684 50124 17736 50176
rect 18236 50124 18288 50176
rect 22560 50328 22612 50380
rect 23848 50396 23900 50448
rect 24032 50464 24084 50516
rect 27436 50464 27488 50516
rect 24676 50396 24728 50448
rect 25872 50396 25924 50448
rect 20260 50260 20312 50312
rect 21180 50303 21232 50312
rect 21180 50269 21189 50303
rect 21189 50269 21223 50303
rect 21223 50269 21232 50303
rect 21180 50260 21232 50269
rect 22284 50192 22336 50244
rect 23572 50328 23624 50380
rect 24124 50328 24176 50380
rect 24952 50371 25004 50380
rect 24952 50337 24961 50371
rect 24961 50337 24995 50371
rect 24995 50337 25004 50371
rect 24952 50328 25004 50337
rect 25596 50371 25648 50380
rect 25596 50337 25605 50371
rect 25605 50337 25639 50371
rect 25639 50337 25648 50371
rect 25596 50328 25648 50337
rect 26240 50371 26292 50380
rect 26240 50337 26249 50371
rect 26249 50337 26283 50371
rect 26283 50337 26292 50371
rect 26240 50328 26292 50337
rect 26976 50328 27028 50380
rect 24768 50260 24820 50312
rect 20168 50124 20220 50176
rect 20996 50124 21048 50176
rect 22744 50124 22796 50176
rect 23020 50124 23072 50176
rect 25136 50192 25188 50244
rect 27896 50192 27948 50244
rect 25872 50124 25924 50176
rect 27988 50124 28040 50176
rect 5614 50022 5666 50074
rect 5678 50022 5730 50074
rect 5742 50022 5794 50074
rect 5806 50022 5858 50074
rect 14878 50022 14930 50074
rect 14942 50022 14994 50074
rect 15006 50022 15058 50074
rect 15070 50022 15122 50074
rect 24142 50022 24194 50074
rect 24206 50022 24258 50074
rect 24270 50022 24322 50074
rect 24334 50022 24386 50074
rect 11980 49963 12032 49972
rect 11980 49929 11989 49963
rect 11989 49929 12023 49963
rect 12023 49929 12032 49963
rect 11980 49920 12032 49929
rect 18512 49963 18564 49972
rect 18512 49929 18521 49963
rect 18521 49929 18555 49963
rect 18555 49929 18564 49963
rect 18512 49920 18564 49929
rect 20076 49963 20128 49972
rect 20076 49929 20085 49963
rect 20085 49929 20119 49963
rect 20119 49929 20128 49963
rect 20076 49920 20128 49929
rect 21180 49963 21232 49972
rect 21180 49929 21189 49963
rect 21189 49929 21223 49963
rect 21223 49929 21232 49963
rect 21180 49920 21232 49929
rect 21824 49963 21876 49972
rect 21824 49929 21833 49963
rect 21833 49929 21867 49963
rect 21867 49929 21876 49963
rect 21824 49920 21876 49929
rect 21916 49920 21968 49972
rect 16396 49852 16448 49904
rect 2964 49784 3016 49836
rect 2688 49716 2740 49768
rect 2872 49716 2924 49768
rect 6000 49716 6052 49768
rect 11336 49784 11388 49836
rect 8208 49716 8260 49768
rect 11888 49759 11940 49768
rect 11888 49725 11897 49759
rect 11897 49725 11931 49759
rect 11931 49725 11940 49759
rect 11888 49716 11940 49725
rect 12716 49716 12768 49768
rect 15476 49784 15528 49836
rect 17684 49827 17736 49836
rect 17684 49793 17693 49827
rect 17693 49793 17727 49827
rect 17727 49793 17736 49827
rect 17684 49784 17736 49793
rect 18236 49784 18288 49836
rect 13084 49716 13136 49768
rect 13636 49759 13688 49768
rect 13636 49725 13645 49759
rect 13645 49725 13679 49759
rect 13679 49725 13688 49759
rect 13636 49716 13688 49725
rect 15384 49759 15436 49768
rect 15384 49725 15393 49759
rect 15393 49725 15427 49759
rect 15427 49725 15436 49759
rect 15384 49716 15436 49725
rect 16948 49716 17000 49768
rect 20904 49784 20956 49836
rect 2504 49580 2556 49632
rect 15200 49648 15252 49700
rect 16304 49648 16356 49700
rect 18788 49716 18840 49768
rect 19340 49716 19392 49768
rect 20996 49716 21048 49768
rect 25136 49852 25188 49904
rect 23020 49784 23072 49836
rect 26424 49784 26476 49836
rect 22652 49716 22704 49768
rect 22928 49716 22980 49768
rect 22836 49648 22888 49700
rect 23848 49716 23900 49768
rect 24032 49716 24084 49768
rect 12900 49623 12952 49632
rect 12900 49589 12909 49623
rect 12909 49589 12943 49623
rect 12943 49589 12952 49623
rect 12900 49580 12952 49589
rect 13912 49580 13964 49632
rect 17500 49580 17552 49632
rect 22744 49623 22796 49632
rect 22744 49589 22753 49623
rect 22753 49589 22787 49623
rect 22787 49589 22796 49623
rect 22744 49580 22796 49589
rect 24032 49623 24084 49632
rect 24032 49589 24041 49623
rect 24041 49589 24075 49623
rect 24075 49589 24084 49623
rect 24032 49580 24084 49589
rect 25412 49716 25464 49768
rect 25780 49759 25832 49768
rect 25780 49725 25789 49759
rect 25789 49725 25823 49759
rect 25823 49725 25832 49759
rect 25780 49716 25832 49725
rect 25872 49716 25924 49768
rect 25872 49580 25924 49632
rect 10246 49478 10298 49530
rect 10310 49478 10362 49530
rect 10374 49478 10426 49530
rect 10438 49478 10490 49530
rect 19510 49478 19562 49530
rect 19574 49478 19626 49530
rect 19638 49478 19690 49530
rect 19702 49478 19754 49530
rect 5908 49419 5960 49428
rect 5908 49385 5917 49419
rect 5917 49385 5951 49419
rect 5951 49385 5960 49419
rect 5908 49376 5960 49385
rect 6000 49376 6052 49428
rect 2688 49308 2740 49360
rect 18420 49308 18472 49360
rect 19340 49308 19392 49360
rect 1860 49283 1912 49292
rect 1860 49249 1869 49283
rect 1869 49249 1903 49283
rect 1903 49249 1912 49283
rect 1860 49240 1912 49249
rect 4712 49240 4764 49292
rect 2688 49172 2740 49224
rect 3792 49172 3844 49224
rect 6184 49240 6236 49292
rect 2780 49147 2832 49156
rect 2780 49113 2789 49147
rect 2789 49113 2823 49147
rect 2823 49113 2832 49147
rect 2780 49104 2832 49113
rect 1952 49079 2004 49088
rect 1952 49045 1961 49079
rect 1961 49045 1995 49079
rect 1995 49045 2004 49079
rect 1952 49036 2004 49045
rect 6092 49172 6144 49224
rect 6644 49172 6696 49224
rect 7748 49240 7800 49292
rect 7932 49283 7984 49292
rect 7932 49249 7966 49283
rect 7966 49249 7984 49283
rect 7932 49240 7984 49249
rect 9864 49240 9916 49292
rect 9588 49172 9640 49224
rect 11060 49240 11112 49292
rect 10692 49172 10744 49224
rect 11888 49240 11940 49292
rect 12256 49283 12308 49292
rect 12256 49249 12265 49283
rect 12265 49249 12299 49283
rect 12299 49249 12308 49283
rect 12256 49240 12308 49249
rect 13176 49240 13228 49292
rect 13544 49283 13596 49292
rect 13544 49249 13553 49283
rect 13553 49249 13587 49283
rect 13587 49249 13596 49283
rect 13544 49240 13596 49249
rect 13912 49240 13964 49292
rect 14740 49283 14792 49292
rect 12348 49215 12400 49224
rect 12348 49181 12357 49215
rect 12357 49181 12391 49215
rect 12391 49181 12400 49215
rect 12348 49172 12400 49181
rect 12808 49172 12860 49224
rect 12900 49172 12952 49224
rect 14740 49249 14749 49283
rect 14749 49249 14783 49283
rect 14783 49249 14792 49283
rect 14740 49240 14792 49249
rect 16948 49240 17000 49292
rect 20444 49308 20496 49360
rect 22744 49376 22796 49428
rect 23112 49419 23164 49428
rect 23112 49385 23121 49419
rect 23121 49385 23155 49419
rect 23155 49385 23164 49419
rect 23112 49376 23164 49385
rect 25780 49376 25832 49428
rect 27896 49351 27948 49360
rect 27896 49317 27905 49351
rect 27905 49317 27939 49351
rect 27939 49317 27948 49351
rect 27896 49308 27948 49317
rect 20260 49283 20312 49292
rect 20260 49249 20269 49283
rect 20269 49249 20303 49283
rect 20303 49249 20312 49283
rect 20260 49240 20312 49249
rect 23848 49240 23900 49292
rect 21364 49215 21416 49224
rect 21364 49181 21373 49215
rect 21373 49181 21407 49215
rect 21407 49181 21416 49215
rect 21364 49172 21416 49181
rect 22560 49172 22612 49224
rect 22928 49172 22980 49224
rect 23940 49172 23992 49224
rect 24676 49283 24728 49292
rect 24676 49249 24685 49283
rect 24685 49249 24719 49283
rect 24719 49249 24728 49283
rect 24860 49283 24912 49292
rect 24676 49240 24728 49249
rect 24860 49249 24869 49283
rect 24869 49249 24903 49283
rect 24903 49249 24912 49283
rect 24860 49240 24912 49249
rect 25780 49283 25832 49292
rect 25780 49249 25789 49283
rect 25789 49249 25823 49283
rect 25823 49249 25832 49283
rect 25780 49240 25832 49249
rect 26884 49283 26936 49292
rect 26884 49249 26893 49283
rect 26893 49249 26927 49283
rect 26927 49249 26936 49283
rect 26884 49240 26936 49249
rect 25596 49172 25648 49224
rect 25872 49215 25924 49224
rect 25872 49181 25881 49215
rect 25881 49181 25915 49215
rect 25915 49181 25924 49215
rect 25872 49172 25924 49181
rect 26148 49172 26200 49224
rect 13912 49104 13964 49156
rect 28080 49104 28132 49156
rect 5264 49079 5316 49088
rect 5264 49045 5273 49079
rect 5273 49045 5307 49079
rect 5307 49045 5316 49079
rect 5264 49036 5316 49045
rect 9036 49079 9088 49088
rect 9036 49045 9045 49079
rect 9045 49045 9079 49079
rect 9079 49045 9088 49079
rect 9036 49036 9088 49045
rect 10048 49036 10100 49088
rect 10968 49079 11020 49088
rect 10968 49045 10977 49079
rect 10977 49045 11011 49079
rect 11011 49045 11020 49079
rect 10968 49036 11020 49045
rect 13360 49079 13412 49088
rect 13360 49045 13369 49079
rect 13369 49045 13403 49079
rect 13403 49045 13412 49079
rect 13360 49036 13412 49045
rect 13544 49036 13596 49088
rect 14648 49079 14700 49088
rect 14648 49045 14657 49079
rect 14657 49045 14691 49079
rect 14691 49045 14700 49079
rect 16120 49079 16172 49088
rect 14648 49036 14700 49045
rect 16120 49045 16129 49079
rect 16129 49045 16163 49079
rect 16163 49045 16172 49079
rect 16120 49036 16172 49045
rect 16396 49036 16448 49088
rect 23204 49036 23256 49088
rect 25504 49036 25556 49088
rect 27896 49036 27948 49088
rect 5614 48934 5666 48986
rect 5678 48934 5730 48986
rect 5742 48934 5794 48986
rect 5806 48934 5858 48986
rect 14878 48934 14930 48986
rect 14942 48934 14994 48986
rect 15006 48934 15058 48986
rect 15070 48934 15122 48986
rect 24142 48934 24194 48986
rect 24206 48934 24258 48986
rect 24270 48934 24322 48986
rect 24334 48934 24386 48986
rect 5172 48832 5224 48884
rect 5448 48832 5500 48884
rect 7932 48832 7984 48884
rect 15384 48832 15436 48884
rect 25780 48832 25832 48884
rect 28080 48875 28132 48884
rect 28080 48841 28089 48875
rect 28089 48841 28123 48875
rect 28123 48841 28132 48875
rect 28080 48832 28132 48841
rect 4160 48764 4212 48816
rect 6276 48807 6328 48816
rect 6276 48773 6285 48807
rect 6285 48773 6319 48807
rect 6319 48773 6328 48807
rect 6276 48764 6328 48773
rect 8024 48764 8076 48816
rect 5172 48696 5224 48748
rect 5448 48696 5500 48748
rect 2872 48628 2924 48680
rect 3792 48628 3844 48680
rect 5264 48628 5316 48680
rect 8300 48628 8352 48680
rect 10600 48764 10652 48816
rect 13360 48764 13412 48816
rect 15200 48764 15252 48816
rect 2596 48560 2648 48612
rect 4436 48560 4488 48612
rect 6552 48603 6604 48612
rect 6552 48569 6561 48603
rect 6561 48569 6595 48603
rect 6595 48569 6604 48603
rect 6552 48560 6604 48569
rect 6920 48560 6972 48612
rect 9036 48560 9088 48612
rect 4252 48535 4304 48544
rect 4252 48501 4261 48535
rect 4261 48501 4295 48535
rect 4295 48501 4304 48535
rect 4252 48492 4304 48501
rect 4620 48535 4672 48544
rect 4620 48501 4629 48535
rect 4629 48501 4663 48535
rect 4663 48501 4672 48535
rect 4620 48492 4672 48501
rect 6736 48535 6788 48544
rect 6736 48501 6745 48535
rect 6745 48501 6779 48535
rect 6779 48501 6788 48535
rect 6736 48492 6788 48501
rect 9588 48492 9640 48544
rect 11152 48696 11204 48748
rect 12256 48696 12308 48748
rect 12348 48696 12400 48748
rect 14648 48696 14700 48748
rect 15292 48696 15344 48748
rect 16120 48696 16172 48748
rect 21180 48696 21232 48748
rect 24032 48696 24084 48748
rect 24768 48764 24820 48816
rect 10140 48628 10192 48680
rect 10692 48628 10744 48680
rect 11060 48628 11112 48680
rect 11060 48492 11112 48544
rect 12900 48671 12952 48680
rect 12900 48637 12909 48671
rect 12909 48637 12943 48671
rect 12943 48637 12952 48671
rect 12900 48628 12952 48637
rect 13176 48628 13228 48680
rect 13912 48628 13964 48680
rect 14556 48628 14608 48680
rect 16856 48628 16908 48680
rect 17500 48671 17552 48680
rect 17500 48637 17509 48671
rect 17509 48637 17543 48671
rect 17543 48637 17552 48671
rect 17500 48628 17552 48637
rect 21364 48671 21416 48680
rect 21364 48637 21373 48671
rect 21373 48637 21407 48671
rect 21407 48637 21416 48671
rect 21364 48628 21416 48637
rect 22836 48628 22888 48680
rect 23204 48671 23256 48680
rect 23204 48637 23213 48671
rect 23213 48637 23247 48671
rect 23247 48637 23256 48671
rect 23204 48628 23256 48637
rect 24676 48628 24728 48680
rect 25320 48628 25372 48680
rect 25504 48671 25556 48680
rect 25504 48637 25513 48671
rect 25513 48637 25547 48671
rect 25547 48637 25556 48671
rect 25504 48628 25556 48637
rect 26700 48671 26752 48680
rect 22192 48560 22244 48612
rect 22744 48560 22796 48612
rect 23940 48560 23992 48612
rect 24032 48560 24084 48612
rect 26700 48637 26709 48671
rect 26709 48637 26743 48671
rect 26743 48637 26752 48671
rect 26700 48628 26752 48637
rect 27160 48628 27212 48680
rect 27988 48671 28040 48680
rect 27988 48637 27997 48671
rect 27997 48637 28031 48671
rect 28031 48637 28040 48671
rect 27988 48628 28040 48637
rect 17684 48535 17736 48544
rect 17684 48501 17693 48535
rect 17693 48501 17727 48535
rect 17727 48501 17736 48535
rect 17684 48492 17736 48501
rect 24584 48492 24636 48544
rect 24768 48492 24820 48544
rect 25320 48492 25372 48544
rect 26148 48492 26200 48544
rect 26516 48535 26568 48544
rect 26516 48501 26525 48535
rect 26525 48501 26559 48535
rect 26559 48501 26568 48535
rect 26516 48492 26568 48501
rect 10246 48390 10298 48442
rect 10310 48390 10362 48442
rect 10374 48390 10426 48442
rect 10438 48390 10490 48442
rect 19510 48390 19562 48442
rect 19574 48390 19626 48442
rect 19638 48390 19690 48442
rect 19702 48390 19754 48442
rect 4620 48288 4672 48340
rect 4712 48288 4764 48340
rect 5264 48288 5316 48340
rect 7104 48331 7156 48340
rect 7104 48297 7113 48331
rect 7113 48297 7147 48331
rect 7147 48297 7156 48331
rect 7104 48288 7156 48297
rect 10140 48288 10192 48340
rect 11060 48331 11112 48340
rect 11060 48297 11069 48331
rect 11069 48297 11103 48331
rect 11103 48297 11112 48331
rect 11060 48288 11112 48297
rect 4252 48220 4304 48272
rect 8208 48220 8260 48272
rect 7104 48195 7156 48204
rect 1216 48084 1268 48136
rect 2964 48127 3016 48136
rect 2964 48093 2973 48127
rect 2973 48093 3007 48127
rect 3007 48093 3016 48127
rect 2964 48084 3016 48093
rect 5448 48127 5500 48136
rect 2872 48016 2924 48068
rect 5448 48093 5457 48127
rect 5457 48093 5491 48127
rect 5491 48093 5500 48127
rect 5448 48084 5500 48093
rect 7104 48161 7113 48195
rect 7113 48161 7147 48195
rect 7147 48161 7156 48195
rect 7104 48152 7156 48161
rect 7196 48152 7248 48204
rect 8300 48152 8352 48204
rect 9588 48152 9640 48204
rect 9864 48195 9916 48204
rect 9864 48161 9873 48195
rect 9873 48161 9907 48195
rect 9907 48161 9916 48195
rect 9864 48152 9916 48161
rect 8576 48127 8628 48136
rect 8576 48093 8585 48127
rect 8585 48093 8619 48127
rect 8619 48093 8628 48127
rect 10048 48127 10100 48136
rect 8576 48084 8628 48093
rect 10048 48093 10057 48127
rect 10057 48093 10091 48127
rect 10091 48093 10100 48127
rect 10048 48084 10100 48093
rect 10968 48220 11020 48272
rect 11152 48195 11204 48204
rect 11152 48161 11161 48195
rect 11161 48161 11195 48195
rect 11195 48161 11204 48195
rect 11152 48152 11204 48161
rect 16856 48220 16908 48272
rect 17408 48152 17460 48204
rect 17684 48220 17736 48272
rect 18144 48195 18196 48204
rect 18144 48161 18153 48195
rect 18153 48161 18187 48195
rect 18187 48161 18196 48195
rect 18144 48152 18196 48161
rect 18880 48152 18932 48204
rect 5908 48016 5960 48068
rect 6736 48016 6788 48068
rect 18052 48084 18104 48136
rect 18512 48084 18564 48136
rect 2688 47948 2740 48000
rect 10876 47991 10928 48000
rect 10876 47957 10885 47991
rect 10885 47957 10919 47991
rect 10919 47957 10928 47991
rect 10876 47948 10928 47957
rect 20260 48288 20312 48340
rect 24584 48288 24636 48340
rect 23940 48220 23992 48272
rect 20444 48152 20496 48204
rect 20628 48152 20680 48204
rect 19984 48084 20036 48136
rect 21088 48152 21140 48204
rect 21364 48152 21416 48204
rect 23204 48195 23256 48204
rect 23204 48161 23213 48195
rect 23213 48161 23247 48195
rect 23247 48161 23256 48195
rect 23204 48152 23256 48161
rect 24032 48152 24084 48204
rect 24492 48152 24544 48204
rect 27896 48220 27948 48272
rect 25596 48195 25648 48204
rect 25596 48161 25605 48195
rect 25605 48161 25639 48195
rect 25639 48161 25648 48195
rect 25596 48152 25648 48161
rect 26240 48195 26292 48204
rect 26240 48161 26249 48195
rect 26249 48161 26283 48195
rect 26283 48161 26292 48195
rect 26240 48152 26292 48161
rect 26976 48152 27028 48204
rect 21180 48084 21232 48136
rect 22836 48084 22888 48136
rect 21364 48016 21416 48068
rect 24676 48084 24728 48136
rect 18788 47948 18840 48000
rect 19064 47991 19116 48000
rect 19064 47957 19073 47991
rect 19073 47957 19107 47991
rect 19107 47957 19116 47991
rect 19064 47948 19116 47957
rect 19248 47948 19300 48000
rect 20260 47948 20312 48000
rect 20444 47948 20496 48000
rect 21272 47948 21324 48000
rect 23848 47948 23900 48000
rect 23940 47948 23992 48000
rect 25964 47948 26016 48000
rect 26056 47991 26108 48000
rect 26056 47957 26065 47991
rect 26065 47957 26099 47991
rect 26099 47957 26108 47991
rect 26056 47948 26108 47957
rect 27896 47948 27948 48000
rect 5614 47846 5666 47898
rect 5678 47846 5730 47898
rect 5742 47846 5794 47898
rect 5806 47846 5858 47898
rect 14878 47846 14930 47898
rect 14942 47846 14994 47898
rect 15006 47846 15058 47898
rect 15070 47846 15122 47898
rect 24142 47846 24194 47898
rect 24206 47846 24258 47898
rect 24270 47846 24322 47898
rect 24334 47846 24386 47898
rect 2596 47787 2648 47796
rect 2596 47753 2605 47787
rect 2605 47753 2639 47787
rect 2639 47753 2648 47787
rect 2596 47744 2648 47753
rect 1860 47676 1912 47728
rect 23940 47744 23992 47796
rect 24492 47744 24544 47796
rect 7288 47676 7340 47728
rect 19984 47676 20036 47728
rect 20168 47676 20220 47728
rect 5172 47608 5224 47660
rect 9036 47608 9088 47660
rect 4620 47540 4672 47592
rect 5816 47583 5868 47592
rect 5816 47549 5825 47583
rect 5825 47549 5859 47583
rect 5859 47549 5868 47583
rect 5816 47540 5868 47549
rect 6460 47583 6512 47592
rect 2596 47472 2648 47524
rect 4160 47472 4212 47524
rect 4896 47472 4948 47524
rect 5724 47472 5776 47524
rect 6460 47549 6469 47583
rect 6469 47549 6503 47583
rect 6503 47549 6512 47583
rect 6460 47540 6512 47549
rect 6644 47540 6696 47592
rect 6828 47540 6880 47592
rect 6276 47472 6328 47524
rect 8944 47540 8996 47592
rect 9864 47540 9916 47592
rect 15200 47608 15252 47660
rect 15476 47608 15528 47660
rect 17684 47608 17736 47660
rect 18052 47583 18104 47592
rect 8392 47515 8444 47524
rect 8392 47481 8401 47515
rect 8401 47481 8435 47515
rect 8435 47481 8444 47515
rect 8392 47472 8444 47481
rect 8576 47472 8628 47524
rect 9588 47472 9640 47524
rect 18052 47549 18061 47583
rect 18061 47549 18095 47583
rect 18095 47549 18104 47583
rect 18052 47540 18104 47549
rect 18144 47540 18196 47592
rect 19800 47608 19852 47660
rect 21272 47651 21324 47660
rect 21272 47617 21281 47651
rect 21281 47617 21315 47651
rect 21315 47617 21324 47651
rect 21272 47608 21324 47617
rect 20076 47540 20128 47592
rect 20904 47540 20956 47592
rect 20996 47540 21048 47592
rect 16212 47472 16264 47524
rect 18788 47472 18840 47524
rect 23848 47540 23900 47592
rect 25412 47540 25464 47592
rect 25872 47583 25924 47592
rect 25872 47549 25881 47583
rect 25881 47549 25915 47583
rect 25915 47549 25924 47583
rect 25872 47540 25924 47549
rect 25964 47540 26016 47592
rect 1952 47447 2004 47456
rect 1952 47413 1961 47447
rect 1961 47413 1995 47447
rect 1995 47413 2004 47447
rect 1952 47404 2004 47413
rect 3056 47447 3108 47456
rect 3056 47413 3065 47447
rect 3065 47413 3099 47447
rect 3099 47413 3108 47447
rect 3056 47404 3108 47413
rect 4620 47447 4672 47456
rect 4620 47413 4629 47447
rect 4629 47413 4663 47447
rect 4663 47413 4672 47447
rect 4620 47404 4672 47413
rect 7104 47404 7156 47456
rect 8668 47404 8720 47456
rect 9864 47447 9916 47456
rect 9864 47413 9873 47447
rect 9873 47413 9907 47447
rect 9907 47413 9916 47447
rect 9864 47404 9916 47413
rect 10140 47404 10192 47456
rect 11060 47447 11112 47456
rect 11060 47413 11069 47447
rect 11069 47413 11103 47447
rect 11103 47413 11112 47447
rect 11060 47404 11112 47413
rect 17040 47447 17092 47456
rect 17040 47413 17049 47447
rect 17049 47413 17083 47447
rect 17083 47413 17092 47447
rect 17040 47404 17092 47413
rect 21272 47404 21324 47456
rect 21732 47447 21784 47456
rect 21732 47413 21741 47447
rect 21741 47413 21775 47447
rect 21775 47413 21784 47447
rect 21732 47404 21784 47413
rect 25964 47404 26016 47456
rect 10246 47302 10298 47354
rect 10310 47302 10362 47354
rect 10374 47302 10426 47354
rect 10438 47302 10490 47354
rect 19510 47302 19562 47354
rect 19574 47302 19626 47354
rect 19638 47302 19690 47354
rect 19702 47302 19754 47354
rect 3792 47200 3844 47252
rect 7196 47200 7248 47252
rect 2964 47132 3016 47184
rect 9588 47175 9640 47184
rect 9588 47141 9597 47175
rect 9597 47141 9631 47175
rect 9631 47141 9640 47175
rect 9588 47132 9640 47141
rect 9864 47132 9916 47184
rect 10600 47175 10652 47184
rect 2504 47064 2556 47116
rect 2688 47064 2740 47116
rect 3332 47107 3384 47116
rect 3332 47073 3341 47107
rect 3341 47073 3375 47107
rect 3375 47073 3384 47107
rect 3332 47064 3384 47073
rect 5724 47107 5776 47116
rect 2780 46971 2832 46980
rect 2780 46937 2789 46971
rect 2789 46937 2823 46971
rect 2823 46937 2832 46971
rect 5724 47073 5733 47107
rect 5733 47073 5767 47107
rect 5767 47073 5776 47107
rect 5724 47064 5776 47073
rect 7104 47107 7156 47116
rect 7104 47073 7113 47107
rect 7113 47073 7147 47107
rect 7147 47073 7156 47107
rect 7104 47064 7156 47073
rect 7288 47107 7340 47116
rect 7288 47073 7297 47107
rect 7297 47073 7331 47107
rect 7331 47073 7340 47107
rect 7288 47064 7340 47073
rect 8944 47064 8996 47116
rect 9404 47107 9456 47116
rect 9404 47073 9413 47107
rect 9413 47073 9447 47107
rect 9447 47073 9456 47107
rect 9404 47064 9456 47073
rect 10140 47064 10192 47116
rect 10600 47141 10609 47175
rect 10609 47141 10643 47175
rect 10643 47141 10652 47175
rect 10600 47132 10652 47141
rect 10508 47064 10560 47116
rect 12440 47064 12492 47116
rect 12624 47107 12676 47116
rect 12624 47073 12633 47107
rect 12633 47073 12667 47107
rect 12667 47073 12676 47107
rect 12624 47064 12676 47073
rect 5908 46996 5960 47048
rect 6828 46996 6880 47048
rect 7564 47039 7616 47048
rect 7564 47005 7573 47039
rect 7573 47005 7607 47039
rect 7607 47005 7616 47039
rect 7564 46996 7616 47005
rect 10968 46996 11020 47048
rect 12532 46996 12584 47048
rect 12808 47039 12860 47048
rect 12808 47005 12817 47039
rect 12817 47005 12851 47039
rect 12851 47005 12860 47039
rect 12808 46996 12860 47005
rect 14096 47064 14148 47116
rect 14648 47107 14700 47116
rect 14648 47073 14682 47107
rect 14682 47073 14700 47107
rect 14648 47064 14700 47073
rect 18052 47064 18104 47116
rect 14188 46996 14240 47048
rect 2780 46928 2832 46937
rect 3424 46903 3476 46912
rect 3424 46869 3433 46903
rect 3433 46869 3467 46903
rect 3467 46869 3476 46903
rect 3424 46860 3476 46869
rect 3516 46860 3568 46912
rect 9772 46928 9824 46980
rect 11152 46928 11204 46980
rect 14096 46928 14148 46980
rect 17684 46928 17736 46980
rect 18144 46971 18196 46980
rect 18144 46937 18153 46971
rect 18153 46937 18187 46971
rect 18187 46937 18196 46971
rect 18144 46928 18196 46937
rect 18512 47200 18564 47252
rect 19800 47243 19852 47252
rect 19800 47209 19809 47243
rect 19809 47209 19843 47243
rect 19843 47209 19852 47243
rect 19800 47200 19852 47209
rect 20168 47200 20220 47252
rect 23664 47200 23716 47252
rect 24032 47200 24084 47252
rect 25872 47200 25924 47252
rect 18328 47107 18380 47116
rect 18328 47073 18337 47107
rect 18337 47073 18371 47107
rect 18371 47073 18380 47107
rect 18328 47064 18380 47073
rect 19892 47064 19944 47116
rect 21732 47132 21784 47184
rect 26516 47132 26568 47184
rect 27896 47175 27948 47184
rect 27896 47141 27905 47175
rect 27905 47141 27939 47175
rect 27939 47141 27948 47175
rect 27896 47132 27948 47141
rect 20076 47107 20128 47116
rect 20076 47073 20085 47107
rect 20085 47073 20119 47107
rect 20119 47073 20128 47107
rect 20260 47107 20312 47116
rect 20076 47064 20128 47073
rect 20260 47073 20269 47107
rect 20269 47073 20303 47107
rect 20303 47073 20312 47107
rect 20260 47064 20312 47073
rect 20444 47064 20496 47116
rect 20996 47107 21048 47116
rect 20996 47073 21005 47107
rect 21005 47073 21039 47107
rect 21039 47073 21048 47107
rect 20996 47064 21048 47073
rect 21088 47107 21140 47116
rect 21088 47073 21097 47107
rect 21097 47073 21131 47107
rect 21131 47073 21140 47107
rect 21272 47107 21324 47116
rect 21088 47064 21140 47073
rect 21272 47073 21281 47107
rect 21281 47073 21315 47107
rect 21315 47073 21324 47107
rect 21272 47064 21324 47073
rect 22560 47064 22612 47116
rect 24308 47064 24360 47116
rect 20904 46996 20956 47048
rect 21180 47039 21232 47048
rect 21180 47005 21189 47039
rect 21189 47005 21223 47039
rect 21223 47005 21232 47039
rect 21180 46996 21232 47005
rect 25044 46996 25096 47048
rect 25964 46996 26016 47048
rect 26148 46996 26200 47048
rect 21364 46928 21416 46980
rect 8208 46860 8260 46912
rect 8484 46860 8536 46912
rect 13728 46903 13780 46912
rect 13728 46869 13737 46903
rect 13737 46869 13771 46903
rect 13771 46869 13780 46903
rect 13728 46860 13780 46869
rect 15752 46903 15804 46912
rect 15752 46869 15761 46903
rect 15761 46869 15795 46903
rect 15795 46869 15804 46903
rect 15752 46860 15804 46869
rect 20260 46860 20312 46912
rect 20628 46860 20680 46912
rect 23388 46860 23440 46912
rect 5614 46758 5666 46810
rect 5678 46758 5730 46810
rect 5742 46758 5794 46810
rect 5806 46758 5858 46810
rect 14878 46758 14930 46810
rect 14942 46758 14994 46810
rect 15006 46758 15058 46810
rect 15070 46758 15122 46810
rect 24142 46758 24194 46810
rect 24206 46758 24258 46810
rect 24270 46758 24322 46810
rect 24334 46758 24386 46810
rect 6552 46656 6604 46708
rect 9404 46656 9456 46708
rect 9588 46699 9640 46708
rect 9588 46665 9597 46699
rect 9597 46665 9631 46699
rect 9631 46665 9640 46699
rect 9588 46656 9640 46665
rect 3332 46588 3384 46640
rect 13268 46588 13320 46640
rect 14648 46588 14700 46640
rect 16212 46631 16264 46640
rect 16212 46597 16221 46631
rect 16221 46597 16255 46631
rect 16255 46597 16264 46631
rect 16212 46588 16264 46597
rect 20996 46588 21048 46640
rect 23204 46588 23256 46640
rect 2596 46520 2648 46572
rect 1216 46452 1268 46504
rect 3976 46452 4028 46504
rect 4436 46495 4488 46504
rect 4436 46461 4445 46495
rect 4445 46461 4479 46495
rect 4479 46461 4488 46495
rect 4436 46452 4488 46461
rect 4896 46495 4948 46504
rect 4896 46461 4905 46495
rect 4905 46461 4939 46495
rect 4939 46461 4948 46495
rect 4896 46452 4948 46461
rect 5908 46452 5960 46504
rect 6276 46452 6328 46504
rect 1584 46384 1636 46436
rect 8300 46520 8352 46572
rect 10508 46520 10560 46572
rect 10784 46520 10836 46572
rect 13728 46520 13780 46572
rect 14832 46520 14884 46572
rect 18328 46520 18380 46572
rect 23020 46520 23072 46572
rect 8484 46452 8536 46504
rect 8668 46452 8720 46504
rect 11060 46452 11112 46504
rect 13544 46452 13596 46504
rect 11796 46384 11848 46436
rect 12532 46384 12584 46436
rect 15752 46384 15804 46436
rect 17040 46452 17092 46504
rect 19892 46452 19944 46504
rect 20168 46495 20220 46504
rect 20168 46461 20177 46495
rect 20177 46461 20211 46495
rect 20211 46461 20220 46495
rect 20168 46452 20220 46461
rect 20904 46452 20956 46504
rect 23848 46452 23900 46504
rect 25964 46495 26016 46504
rect 25964 46461 25973 46495
rect 25973 46461 26007 46495
rect 26007 46461 26016 46495
rect 25964 46452 26016 46461
rect 26424 46495 26476 46504
rect 26424 46461 26433 46495
rect 26433 46461 26467 46495
rect 26467 46461 26476 46495
rect 26424 46452 26476 46461
rect 26056 46384 26108 46436
rect 3148 46316 3200 46368
rect 4344 46359 4396 46368
rect 4344 46325 4353 46359
rect 4353 46325 4387 46359
rect 4387 46325 4396 46359
rect 4344 46316 4396 46325
rect 4988 46359 5040 46368
rect 4988 46325 4997 46359
rect 4997 46325 5031 46359
rect 5031 46325 5040 46359
rect 4988 46316 5040 46325
rect 6276 46316 6328 46368
rect 8668 46316 8720 46368
rect 10048 46359 10100 46368
rect 10048 46325 10057 46359
rect 10057 46325 10091 46359
rect 10091 46325 10100 46359
rect 10048 46316 10100 46325
rect 11428 46316 11480 46368
rect 11612 46359 11664 46368
rect 11612 46325 11621 46359
rect 11621 46325 11655 46359
rect 11655 46325 11664 46359
rect 11612 46316 11664 46325
rect 11704 46359 11756 46368
rect 11704 46325 11713 46359
rect 11713 46325 11747 46359
rect 11747 46325 11756 46359
rect 13636 46359 13688 46368
rect 11704 46316 11756 46325
rect 13636 46325 13645 46359
rect 13645 46325 13679 46359
rect 13679 46325 13688 46359
rect 13636 46316 13688 46325
rect 14188 46316 14240 46368
rect 17316 46316 17368 46368
rect 17500 46359 17552 46368
rect 17500 46325 17509 46359
rect 17509 46325 17543 46359
rect 17543 46325 17552 46359
rect 17500 46316 17552 46325
rect 23112 46359 23164 46368
rect 23112 46325 23121 46359
rect 23121 46325 23155 46359
rect 23155 46325 23164 46359
rect 23112 46316 23164 46325
rect 23204 46359 23256 46368
rect 23204 46325 23213 46359
rect 23213 46325 23247 46359
rect 23247 46325 23256 46359
rect 23204 46316 23256 46325
rect 24492 46316 24544 46368
rect 25872 46316 25924 46368
rect 10246 46214 10298 46266
rect 10310 46214 10362 46266
rect 10374 46214 10426 46266
rect 10438 46214 10490 46266
rect 19510 46214 19562 46266
rect 19574 46214 19626 46266
rect 19638 46214 19690 46266
rect 19702 46214 19754 46266
rect 4620 46112 4672 46164
rect 6092 46112 6144 46164
rect 10048 46155 10100 46164
rect 10048 46121 10057 46155
rect 10057 46121 10091 46155
rect 10091 46121 10100 46155
rect 10048 46112 10100 46121
rect 11612 46112 11664 46164
rect 11796 46112 11848 46164
rect 4252 46044 4304 46096
rect 8208 46044 8260 46096
rect 13544 46044 13596 46096
rect 1768 45976 1820 46028
rect 3148 45976 3200 46028
rect 3332 45976 3384 46028
rect 3516 45951 3568 45960
rect 3516 45917 3525 45951
rect 3525 45917 3559 45951
rect 3559 45917 3568 45951
rect 3516 45908 3568 45917
rect 3608 45951 3660 45960
rect 3608 45917 3617 45951
rect 3617 45917 3651 45951
rect 3651 45917 3660 45951
rect 3608 45908 3660 45917
rect 4804 45908 4856 45960
rect 2780 45840 2832 45892
rect 4160 45840 4212 45892
rect 10600 45976 10652 46028
rect 13728 46044 13780 46096
rect 19984 46087 20036 46096
rect 19984 46053 19993 46087
rect 19993 46053 20027 46087
rect 20027 46053 20036 46087
rect 19984 46044 20036 46053
rect 23204 46112 23256 46164
rect 23388 46155 23440 46164
rect 23388 46121 23397 46155
rect 23397 46121 23431 46155
rect 23431 46121 23440 46155
rect 23388 46112 23440 46121
rect 24584 46112 24636 46164
rect 10876 45951 10928 45960
rect 10876 45917 10885 45951
rect 10885 45917 10919 45951
rect 10919 45917 10928 45951
rect 10876 45908 10928 45917
rect 11704 45840 11756 45892
rect 14188 45976 14240 46028
rect 13544 45908 13596 45960
rect 3148 45772 3200 45824
rect 4528 45815 4580 45824
rect 4528 45781 4537 45815
rect 4537 45781 4571 45815
rect 4571 45781 4580 45815
rect 4528 45772 4580 45781
rect 12348 45815 12400 45824
rect 12348 45781 12357 45815
rect 12357 45781 12391 45815
rect 12391 45781 12400 45815
rect 12348 45772 12400 45781
rect 13176 45772 13228 45824
rect 13268 45772 13320 45824
rect 15752 45976 15804 46028
rect 17132 45976 17184 46028
rect 17408 45976 17460 46028
rect 18144 46019 18196 46028
rect 18144 45985 18153 46019
rect 18153 45985 18187 46019
rect 18187 45985 18196 46019
rect 18144 45976 18196 45985
rect 19892 45976 19944 46028
rect 23480 45951 23532 45960
rect 23480 45917 23489 45951
rect 23489 45917 23523 45951
rect 23523 45917 23532 45951
rect 23480 45908 23532 45917
rect 24032 45976 24084 46028
rect 24584 46019 24636 46028
rect 24584 45985 24593 46019
rect 24593 45985 24627 46019
rect 24627 45985 24636 46019
rect 24584 45976 24636 45985
rect 24860 45976 24912 46028
rect 25596 46019 25648 46028
rect 25596 45985 25605 46019
rect 25605 45985 25639 46019
rect 25639 45985 25648 46019
rect 25596 45976 25648 45985
rect 26240 46019 26292 46028
rect 26240 45985 26249 46019
rect 26249 45985 26283 46019
rect 26283 45985 26292 46019
rect 26240 45976 26292 45985
rect 26976 45976 27028 46028
rect 22192 45840 22244 45892
rect 27620 45840 27672 45892
rect 15752 45815 15804 45824
rect 15752 45781 15761 45815
rect 15761 45781 15795 45815
rect 15795 45781 15804 45815
rect 15752 45772 15804 45781
rect 18236 45815 18288 45824
rect 18236 45781 18245 45815
rect 18245 45781 18279 45815
rect 18279 45781 18288 45815
rect 18236 45772 18288 45781
rect 27896 45772 27948 45824
rect 5614 45670 5666 45722
rect 5678 45670 5730 45722
rect 5742 45670 5794 45722
rect 5806 45670 5858 45722
rect 14878 45670 14930 45722
rect 14942 45670 14994 45722
rect 15006 45670 15058 45722
rect 15070 45670 15122 45722
rect 24142 45670 24194 45722
rect 24206 45670 24258 45722
rect 24270 45670 24322 45722
rect 24334 45670 24386 45722
rect 1584 45611 1636 45620
rect 1584 45577 1593 45611
rect 1593 45577 1627 45611
rect 1627 45577 1636 45611
rect 1584 45568 1636 45577
rect 2504 45500 2556 45552
rect 2136 45432 2188 45484
rect 2320 45432 2372 45484
rect 3332 45568 3384 45620
rect 7564 45568 7616 45620
rect 13636 45568 13688 45620
rect 3516 45500 3568 45552
rect 4620 45500 4672 45552
rect 10784 45500 10836 45552
rect 12348 45500 12400 45552
rect 21456 45568 21508 45620
rect 4804 45475 4856 45484
rect 4804 45441 4813 45475
rect 4813 45441 4847 45475
rect 4847 45441 4856 45475
rect 4804 45432 4856 45441
rect 6920 45432 6972 45484
rect 7472 45432 7524 45484
rect 11152 45475 11204 45484
rect 11152 45441 11161 45475
rect 11161 45441 11195 45475
rect 11195 45441 11204 45475
rect 11152 45432 11204 45441
rect 11428 45475 11480 45484
rect 11428 45441 11437 45475
rect 11437 45441 11471 45475
rect 11471 45441 11480 45475
rect 11428 45432 11480 45441
rect 3240 45364 3292 45416
rect 4988 45364 5040 45416
rect 9312 45364 9364 45416
rect 13544 45364 13596 45416
rect 17132 45500 17184 45552
rect 18052 45500 18104 45552
rect 22560 45543 22612 45552
rect 22560 45509 22569 45543
rect 22569 45509 22603 45543
rect 22603 45509 22612 45543
rect 22560 45500 22612 45509
rect 24584 45500 24636 45552
rect 25688 45500 25740 45552
rect 14280 45432 14332 45484
rect 13728 45407 13780 45416
rect 13728 45373 13737 45407
rect 13737 45373 13771 45407
rect 13771 45373 13780 45407
rect 13728 45364 13780 45373
rect 15752 45364 15804 45416
rect 16028 45364 16080 45416
rect 18144 45407 18196 45416
rect 2228 45228 2280 45280
rect 3608 45296 3660 45348
rect 7656 45296 7708 45348
rect 8024 45296 8076 45348
rect 14096 45296 14148 45348
rect 16120 45296 16172 45348
rect 18144 45373 18153 45407
rect 18153 45373 18187 45407
rect 18187 45373 18196 45407
rect 18144 45364 18196 45373
rect 18420 45407 18472 45416
rect 18420 45373 18429 45407
rect 18429 45373 18463 45407
rect 18463 45373 18472 45407
rect 18420 45364 18472 45373
rect 21180 45407 21232 45416
rect 21180 45373 21189 45407
rect 21189 45373 21223 45407
rect 21223 45373 21232 45407
rect 21180 45364 21232 45373
rect 21456 45339 21508 45348
rect 21456 45305 21490 45339
rect 21490 45305 21508 45339
rect 21456 45296 21508 45305
rect 22560 45364 22612 45416
rect 23020 45296 23072 45348
rect 24492 45432 24544 45484
rect 24124 45364 24176 45416
rect 25596 45364 25648 45416
rect 27068 45407 27120 45416
rect 27068 45373 27077 45407
rect 27077 45373 27111 45407
rect 27111 45373 27120 45407
rect 27068 45364 27120 45373
rect 27620 45407 27672 45416
rect 27620 45373 27629 45407
rect 27629 45373 27663 45407
rect 27663 45373 27672 45407
rect 27620 45364 27672 45373
rect 3332 45228 3384 45280
rect 3976 45228 4028 45280
rect 4712 45271 4764 45280
rect 4712 45237 4721 45271
rect 4721 45237 4755 45271
rect 4755 45237 4764 45271
rect 4712 45228 4764 45237
rect 6000 45228 6052 45280
rect 6184 45271 6236 45280
rect 6184 45237 6193 45271
rect 6193 45237 6227 45271
rect 6227 45237 6236 45271
rect 6184 45228 6236 45237
rect 6460 45228 6512 45280
rect 7748 45228 7800 45280
rect 9496 45228 9548 45280
rect 11796 45228 11848 45280
rect 12624 45228 12676 45280
rect 14280 45228 14332 45280
rect 15568 45228 15620 45280
rect 15660 45228 15712 45280
rect 18144 45228 18196 45280
rect 21548 45228 21600 45280
rect 23940 45296 23992 45348
rect 23388 45228 23440 45280
rect 23848 45228 23900 45280
rect 24308 45228 24360 45280
rect 26884 45271 26936 45280
rect 26884 45237 26893 45271
rect 26893 45237 26927 45271
rect 26927 45237 26936 45271
rect 26884 45228 26936 45237
rect 10246 45126 10298 45178
rect 10310 45126 10362 45178
rect 10374 45126 10426 45178
rect 10438 45126 10490 45178
rect 19510 45126 19562 45178
rect 19574 45126 19626 45178
rect 19638 45126 19690 45178
rect 19702 45126 19754 45178
rect 4160 45024 4212 45076
rect 4344 45067 4396 45076
rect 4344 45033 4353 45067
rect 4353 45033 4387 45067
rect 4387 45033 4396 45067
rect 4344 45024 4396 45033
rect 4528 45024 4580 45076
rect 2136 44956 2188 45008
rect 17500 44956 17552 45008
rect 18328 44956 18380 45008
rect 19064 44956 19116 45008
rect 20076 44956 20128 45008
rect 23112 45024 23164 45076
rect 24124 45024 24176 45076
rect 23940 44956 23992 45008
rect 24032 44999 24084 45008
rect 24032 44965 24041 44999
rect 24041 44965 24075 44999
rect 24075 44965 24084 44999
rect 24032 44956 24084 44965
rect 24308 44956 24360 45008
rect 2596 44888 2648 44940
rect 5080 44888 5132 44940
rect 5724 44931 5776 44940
rect 5724 44897 5733 44931
rect 5733 44897 5767 44931
rect 5767 44897 5776 44931
rect 5724 44888 5776 44897
rect 6000 44888 6052 44940
rect 6828 44931 6880 44940
rect 6828 44897 6837 44931
rect 6837 44897 6871 44931
rect 6871 44897 6880 44931
rect 6828 44888 6880 44897
rect 7564 44931 7616 44940
rect 3240 44820 3292 44872
rect 3516 44820 3568 44872
rect 3608 44820 3660 44872
rect 6368 44820 6420 44872
rect 7564 44897 7573 44931
rect 7573 44897 7607 44931
rect 7607 44897 7616 44931
rect 7564 44888 7616 44897
rect 7932 44931 7984 44940
rect 7932 44897 7941 44931
rect 7941 44897 7975 44931
rect 7975 44897 7984 44931
rect 7932 44888 7984 44897
rect 8024 44888 8076 44940
rect 9496 44931 9548 44940
rect 9496 44897 9505 44931
rect 9505 44897 9539 44931
rect 9539 44897 9548 44931
rect 9496 44888 9548 44897
rect 9680 44931 9732 44940
rect 9680 44897 9689 44931
rect 9689 44897 9723 44931
rect 9723 44897 9732 44931
rect 9680 44888 9732 44897
rect 12348 44888 12400 44940
rect 15568 44888 15620 44940
rect 17592 44888 17644 44940
rect 18144 44931 18196 44940
rect 18144 44897 18153 44931
rect 18153 44897 18187 44931
rect 18187 44897 18196 44931
rect 18144 44888 18196 44897
rect 18236 44888 18288 44940
rect 18972 44931 19024 44940
rect 18972 44897 18981 44931
rect 18981 44897 19015 44931
rect 19015 44897 19024 44931
rect 18972 44888 19024 44897
rect 22560 44888 22612 44940
rect 8760 44863 8812 44872
rect 8760 44829 8769 44863
rect 8769 44829 8803 44863
rect 8803 44829 8812 44863
rect 8760 44820 8812 44829
rect 12900 44863 12952 44872
rect 12900 44829 12909 44863
rect 12909 44829 12943 44863
rect 12943 44829 12952 44863
rect 12900 44820 12952 44829
rect 13544 44820 13596 44872
rect 14096 44863 14148 44872
rect 4804 44752 4856 44804
rect 6644 44752 6696 44804
rect 10784 44752 10836 44804
rect 14096 44829 14105 44863
rect 14105 44829 14139 44863
rect 14139 44829 14148 44863
rect 14096 44820 14148 44829
rect 14556 44820 14608 44872
rect 22744 44888 22796 44940
rect 23296 44931 23348 44940
rect 23296 44897 23305 44931
rect 23305 44897 23339 44931
rect 23339 44897 23348 44931
rect 23296 44888 23348 44897
rect 27896 44999 27948 45008
rect 27896 44965 27905 44999
rect 27905 44965 27939 44999
rect 27939 44965 27948 44999
rect 27896 44956 27948 44965
rect 25320 44931 25372 44940
rect 14464 44752 14516 44804
rect 15660 44795 15712 44804
rect 15660 44761 15669 44795
rect 15669 44761 15703 44795
rect 15703 44761 15712 44795
rect 15660 44752 15712 44761
rect 18788 44752 18840 44804
rect 1952 44727 2004 44736
rect 1952 44693 1961 44727
rect 1961 44693 1995 44727
rect 1995 44693 2004 44727
rect 1952 44684 2004 44693
rect 2412 44684 2464 44736
rect 3608 44684 3660 44736
rect 6736 44684 6788 44736
rect 7104 44684 7156 44736
rect 8392 44684 8444 44736
rect 9312 44684 9364 44736
rect 9772 44684 9824 44736
rect 19156 44727 19208 44736
rect 19156 44693 19165 44727
rect 19165 44693 19199 44727
rect 19199 44693 19208 44727
rect 19156 44684 19208 44693
rect 23388 44820 23440 44872
rect 25320 44897 25329 44931
rect 25329 44897 25363 44931
rect 25363 44897 25372 44931
rect 25320 44888 25372 44897
rect 26148 44888 26200 44940
rect 27160 44888 27212 44940
rect 22192 44752 22244 44804
rect 23940 44752 23992 44804
rect 21640 44684 21692 44736
rect 24768 44684 24820 44736
rect 24952 44684 25004 44736
rect 25136 44727 25188 44736
rect 25136 44693 25145 44727
rect 25145 44693 25179 44727
rect 25179 44693 25188 44727
rect 25136 44684 25188 44693
rect 26056 44727 26108 44736
rect 26056 44693 26065 44727
rect 26065 44693 26099 44727
rect 26099 44693 26108 44727
rect 26056 44684 26108 44693
rect 26700 44727 26752 44736
rect 26700 44693 26709 44727
rect 26709 44693 26743 44727
rect 26743 44693 26752 44727
rect 26700 44684 26752 44693
rect 5614 44582 5666 44634
rect 5678 44582 5730 44634
rect 5742 44582 5794 44634
rect 5806 44582 5858 44634
rect 14878 44582 14930 44634
rect 14942 44582 14994 44634
rect 15006 44582 15058 44634
rect 15070 44582 15122 44634
rect 24142 44582 24194 44634
rect 24206 44582 24258 44634
rect 24270 44582 24322 44634
rect 24334 44582 24386 44634
rect 3056 44480 3108 44532
rect 4988 44480 5040 44532
rect 6460 44523 6512 44532
rect 6460 44489 6469 44523
rect 6469 44489 6503 44523
rect 6503 44489 6512 44523
rect 6460 44480 6512 44489
rect 1860 44412 1912 44464
rect 2688 44412 2740 44464
rect 23940 44480 23992 44532
rect 25320 44480 25372 44532
rect 9680 44412 9732 44464
rect 11152 44455 11204 44464
rect 11152 44421 11161 44455
rect 11161 44421 11195 44455
rect 11195 44421 11204 44455
rect 11152 44412 11204 44421
rect 16120 44455 16172 44464
rect 16120 44421 16129 44455
rect 16129 44421 16163 44455
rect 16163 44421 16172 44455
rect 16120 44412 16172 44421
rect 18236 44455 18288 44464
rect 18236 44421 18245 44455
rect 18245 44421 18279 44455
rect 18279 44421 18288 44455
rect 18236 44412 18288 44421
rect 18696 44412 18748 44464
rect 4344 44344 4396 44396
rect 5448 44387 5500 44396
rect 5448 44353 5457 44387
rect 5457 44353 5491 44387
rect 5491 44353 5500 44387
rect 5448 44344 5500 44353
rect 7104 44387 7156 44396
rect 7104 44353 7113 44387
rect 7113 44353 7147 44387
rect 7147 44353 7156 44387
rect 7104 44344 7156 44353
rect 2228 44276 2280 44328
rect 3056 44319 3108 44328
rect 3056 44285 3065 44319
rect 3065 44285 3099 44319
rect 3099 44285 3108 44319
rect 3056 44276 3108 44285
rect 6736 44276 6788 44328
rect 9772 44387 9824 44396
rect 7564 44276 7616 44328
rect 9404 44276 9456 44328
rect 2412 44251 2464 44260
rect 2412 44217 2421 44251
rect 2421 44217 2455 44251
rect 2455 44217 2464 44251
rect 2412 44208 2464 44217
rect 5908 44208 5960 44260
rect 7748 44251 7800 44260
rect 7748 44217 7757 44251
rect 7757 44217 7791 44251
rect 7791 44217 7800 44251
rect 7748 44208 7800 44217
rect 8208 44208 8260 44260
rect 9772 44353 9781 44387
rect 9781 44353 9815 44387
rect 9815 44353 9824 44387
rect 9772 44344 9824 44353
rect 12900 44344 12952 44396
rect 13728 44344 13780 44396
rect 15476 44344 15528 44396
rect 16396 44344 16448 44396
rect 18144 44344 18196 44396
rect 20076 44412 20128 44464
rect 21180 44412 21232 44464
rect 23480 44455 23532 44464
rect 23480 44421 23489 44455
rect 23489 44421 23523 44455
rect 23523 44421 23532 44455
rect 23480 44412 23532 44421
rect 10048 44276 10100 44328
rect 10692 44276 10744 44328
rect 13268 44319 13320 44328
rect 13268 44285 13277 44319
rect 13277 44285 13311 44319
rect 13311 44285 13320 44319
rect 13268 44276 13320 44285
rect 14096 44276 14148 44328
rect 17132 44319 17184 44328
rect 17132 44285 17141 44319
rect 17141 44285 17175 44319
rect 17175 44285 17184 44319
rect 17132 44276 17184 44285
rect 17592 44276 17644 44328
rect 19800 44276 19852 44328
rect 20720 44276 20772 44328
rect 21272 44319 21324 44328
rect 21272 44285 21281 44319
rect 21281 44285 21315 44319
rect 21315 44285 21324 44319
rect 21272 44276 21324 44285
rect 21824 44276 21876 44328
rect 23572 44344 23624 44396
rect 23848 44344 23900 44396
rect 25412 44412 25464 44464
rect 24492 44344 24544 44396
rect 24860 44344 24912 44396
rect 17316 44208 17368 44260
rect 19340 44208 19392 44260
rect 25412 44276 25464 44328
rect 25596 44276 25648 44328
rect 26884 44276 26936 44328
rect 23572 44208 23624 44260
rect 4804 44183 4856 44192
rect 4804 44149 4813 44183
rect 4813 44149 4847 44183
rect 4847 44149 4856 44183
rect 4804 44140 4856 44149
rect 6368 44140 6420 44192
rect 8024 44140 8076 44192
rect 9772 44183 9824 44192
rect 9772 44149 9781 44183
rect 9781 44149 9815 44183
rect 9815 44149 9824 44183
rect 9772 44140 9824 44149
rect 12808 44140 12860 44192
rect 13268 44140 13320 44192
rect 18972 44183 19024 44192
rect 18972 44149 18981 44183
rect 18981 44149 19015 44183
rect 19015 44149 19024 44183
rect 18972 44140 19024 44149
rect 19800 44140 19852 44192
rect 21272 44140 21324 44192
rect 21548 44140 21600 44192
rect 23940 44140 23992 44192
rect 24860 44208 24912 44260
rect 28080 44183 28132 44192
rect 28080 44149 28089 44183
rect 28089 44149 28123 44183
rect 28123 44149 28132 44183
rect 28080 44140 28132 44149
rect 10246 44038 10298 44090
rect 10310 44038 10362 44090
rect 10374 44038 10426 44090
rect 10438 44038 10490 44090
rect 19510 44038 19562 44090
rect 19574 44038 19626 44090
rect 19638 44038 19690 44090
rect 19702 44038 19754 44090
rect 3424 43979 3476 43988
rect 3424 43945 3433 43979
rect 3433 43945 3467 43979
rect 3467 43945 3476 43979
rect 3424 43936 3476 43945
rect 5908 43936 5960 43988
rect 6644 43936 6696 43988
rect 2688 43800 2740 43852
rect 2780 43707 2832 43716
rect 2780 43673 2789 43707
rect 2789 43673 2823 43707
rect 2823 43673 2832 43707
rect 2780 43664 2832 43673
rect 1400 43596 1452 43648
rect 4804 43868 4856 43920
rect 6828 43868 6880 43920
rect 7932 43936 7984 43988
rect 8208 43936 8260 43988
rect 3976 43732 4028 43784
rect 6368 43732 6420 43784
rect 7748 43732 7800 43784
rect 9772 43868 9824 43920
rect 10048 43936 10100 43988
rect 13544 43868 13596 43920
rect 14740 43868 14792 43920
rect 18420 43868 18472 43920
rect 21364 43868 21416 43920
rect 21456 43868 21508 43920
rect 23848 43868 23900 43920
rect 10692 43800 10744 43852
rect 12624 43800 12676 43852
rect 14648 43800 14700 43852
rect 17592 43843 17644 43852
rect 17592 43809 17601 43843
rect 17601 43809 17635 43843
rect 17635 43809 17644 43843
rect 17592 43800 17644 43809
rect 18788 43843 18840 43852
rect 18788 43809 18797 43843
rect 18797 43809 18831 43843
rect 18831 43809 18840 43843
rect 18788 43800 18840 43809
rect 19064 43800 19116 43852
rect 19156 43800 19208 43852
rect 9220 43732 9272 43784
rect 18880 43775 18932 43784
rect 18880 43741 18889 43775
rect 18889 43741 18923 43775
rect 18923 43741 18932 43775
rect 18880 43732 18932 43741
rect 19340 43775 19392 43784
rect 19340 43741 19349 43775
rect 19349 43741 19383 43775
rect 19383 43741 19392 43775
rect 19340 43732 19392 43741
rect 20996 43775 21048 43784
rect 20996 43741 21005 43775
rect 21005 43741 21039 43775
rect 21039 43741 21048 43775
rect 20996 43732 21048 43741
rect 21548 43732 21600 43784
rect 21824 43732 21876 43784
rect 23388 43800 23440 43852
rect 24860 43936 24912 43988
rect 25504 43936 25556 43988
rect 25688 43936 25740 43988
rect 24952 43868 25004 43920
rect 25320 43911 25372 43920
rect 25320 43877 25329 43911
rect 25329 43877 25363 43911
rect 25363 43877 25372 43911
rect 25320 43868 25372 43877
rect 26056 43868 26108 43920
rect 23480 43732 23532 43784
rect 25136 43732 25188 43784
rect 25964 43800 26016 43852
rect 26148 43843 26200 43852
rect 26148 43809 26157 43843
rect 26157 43809 26191 43843
rect 26191 43809 26200 43843
rect 26148 43800 26200 43809
rect 26240 43800 26292 43852
rect 28080 43732 28132 43784
rect 9036 43596 9088 43648
rect 10600 43664 10652 43716
rect 10784 43596 10836 43648
rect 18328 43664 18380 43716
rect 20260 43596 20312 43648
rect 22376 43596 22428 43648
rect 23848 43596 23900 43648
rect 27252 43664 27304 43716
rect 28080 43639 28132 43648
rect 28080 43605 28089 43639
rect 28089 43605 28123 43639
rect 28123 43605 28132 43639
rect 28080 43596 28132 43605
rect 5614 43494 5666 43546
rect 5678 43494 5730 43546
rect 5742 43494 5794 43546
rect 5806 43494 5858 43546
rect 14878 43494 14930 43546
rect 14942 43494 14994 43546
rect 15006 43494 15058 43546
rect 15070 43494 15122 43546
rect 24142 43494 24194 43546
rect 24206 43494 24258 43546
rect 24270 43494 24322 43546
rect 24334 43494 24386 43546
rect 1308 43392 1360 43444
rect 4436 43392 4488 43444
rect 4620 43392 4672 43444
rect 6184 43392 6236 43444
rect 10692 43392 10744 43444
rect 10784 43392 10836 43444
rect 21364 43435 21416 43444
rect 1768 43324 1820 43376
rect 10600 43324 10652 43376
rect 12900 43324 12952 43376
rect 13084 43324 13136 43376
rect 21364 43401 21373 43435
rect 21373 43401 21407 43435
rect 21407 43401 21416 43435
rect 21364 43392 21416 43401
rect 23020 43392 23072 43444
rect 25320 43435 25372 43444
rect 25320 43401 25329 43435
rect 25329 43401 25363 43435
rect 25363 43401 25372 43435
rect 25320 43392 25372 43401
rect 27988 43324 28040 43376
rect 4160 43188 4212 43240
rect 4620 43188 4672 43240
rect 4896 43231 4948 43240
rect 4896 43197 4905 43231
rect 4905 43197 4939 43231
rect 4939 43197 4948 43231
rect 4896 43188 4948 43197
rect 2504 43120 2556 43172
rect 3332 43120 3384 43172
rect 4436 43120 4488 43172
rect 6184 43188 6236 43240
rect 6552 43188 6604 43240
rect 9496 43231 9548 43240
rect 9496 43197 9505 43231
rect 9505 43197 9539 43231
rect 9539 43197 9548 43231
rect 9496 43188 9548 43197
rect 10692 43188 10744 43240
rect 6276 43120 6328 43172
rect 11152 43163 11204 43172
rect 11152 43129 11186 43163
rect 11186 43129 11204 43163
rect 15108 43188 15160 43240
rect 18696 43188 18748 43240
rect 18788 43231 18840 43240
rect 18788 43197 18797 43231
rect 18797 43197 18831 43231
rect 18831 43197 18840 43231
rect 18788 43188 18840 43197
rect 11152 43120 11204 43129
rect 15292 43163 15344 43172
rect 15292 43129 15326 43163
rect 15326 43129 15344 43163
rect 15292 43120 15344 43129
rect 2964 43052 3016 43104
rect 9312 43052 9364 43104
rect 11060 43052 11112 43104
rect 11612 43052 11664 43104
rect 12348 43052 12400 43104
rect 15200 43052 15252 43104
rect 15384 43052 15436 43104
rect 16396 43095 16448 43104
rect 16396 43061 16405 43095
rect 16405 43061 16439 43095
rect 16439 43061 16448 43095
rect 16396 43052 16448 43061
rect 18972 43163 19024 43172
rect 18420 43052 18472 43104
rect 18972 43129 18981 43163
rect 18981 43129 19015 43163
rect 19015 43129 19024 43163
rect 18972 43120 19024 43129
rect 22284 43256 22336 43308
rect 20076 43188 20128 43240
rect 20260 43231 20312 43240
rect 20260 43197 20294 43231
rect 20294 43197 20312 43231
rect 20260 43188 20312 43197
rect 23020 43231 23072 43240
rect 23020 43197 23029 43231
rect 23029 43197 23063 43231
rect 23063 43197 23072 43231
rect 23020 43188 23072 43197
rect 24860 43188 24912 43240
rect 25136 43188 25188 43240
rect 26056 43231 26108 43240
rect 26056 43197 26065 43231
rect 26065 43197 26099 43231
rect 26099 43197 26108 43231
rect 26056 43188 26108 43197
rect 26792 43188 26844 43240
rect 18880 43052 18932 43104
rect 21456 43052 21508 43104
rect 21824 43095 21876 43104
rect 21824 43061 21833 43095
rect 21833 43061 21867 43095
rect 21867 43061 21876 43095
rect 21824 43052 21876 43061
rect 22284 43095 22336 43104
rect 22284 43061 22293 43095
rect 22293 43061 22327 43095
rect 22327 43061 22336 43095
rect 22284 43052 22336 43061
rect 26240 43120 26292 43172
rect 27252 43163 27304 43172
rect 27252 43129 27261 43163
rect 27261 43129 27295 43163
rect 27295 43129 27304 43163
rect 27252 43120 27304 43129
rect 10246 42950 10298 43002
rect 10310 42950 10362 43002
rect 10374 42950 10426 43002
rect 10438 42950 10490 43002
rect 19510 42950 19562 43002
rect 19574 42950 19626 43002
rect 19638 42950 19690 43002
rect 19702 42950 19754 43002
rect 2596 42848 2648 42900
rect 28080 42848 28132 42900
rect 1584 42780 1636 42832
rect 4896 42780 4948 42832
rect 11152 42823 11204 42832
rect 11152 42789 11161 42823
rect 11161 42789 11195 42823
rect 11195 42789 11204 42823
rect 11152 42780 11204 42789
rect 11244 42780 11296 42832
rect 12532 42823 12584 42832
rect 12532 42789 12541 42823
rect 12541 42789 12575 42823
rect 12575 42789 12584 42823
rect 12532 42780 12584 42789
rect 18972 42780 19024 42832
rect 21824 42780 21876 42832
rect 23388 42780 23440 42832
rect 25136 42823 25188 42832
rect 25136 42789 25145 42823
rect 25145 42789 25179 42823
rect 25179 42789 25188 42823
rect 25136 42780 25188 42789
rect 2412 42712 2464 42764
rect 2596 42755 2648 42764
rect 2596 42721 2605 42755
rect 2605 42721 2639 42755
rect 2639 42721 2648 42755
rect 2596 42712 2648 42721
rect 3608 42687 3660 42696
rect 3608 42653 3617 42687
rect 3617 42653 3651 42687
rect 3651 42653 3660 42687
rect 3608 42644 3660 42653
rect 4160 42644 4212 42696
rect 4436 42644 4488 42696
rect 4988 42712 5040 42764
rect 7748 42712 7800 42764
rect 9496 42712 9548 42764
rect 10784 42755 10836 42764
rect 10784 42721 10793 42755
rect 10793 42721 10827 42755
rect 10827 42721 10836 42755
rect 10784 42712 10836 42721
rect 12348 42712 12400 42764
rect 9404 42644 9456 42696
rect 14280 42712 14332 42764
rect 18420 42755 18472 42764
rect 18420 42721 18429 42755
rect 18429 42721 18463 42755
rect 18463 42721 18472 42755
rect 18420 42712 18472 42721
rect 13636 42644 13688 42696
rect 13728 42687 13780 42696
rect 13728 42653 13737 42687
rect 13737 42653 13771 42687
rect 13771 42653 13780 42687
rect 14004 42687 14056 42696
rect 13728 42644 13780 42653
rect 14004 42653 14013 42687
rect 14013 42653 14047 42687
rect 14047 42653 14056 42687
rect 14004 42644 14056 42653
rect 14188 42644 14240 42696
rect 2780 42619 2832 42628
rect 2780 42585 2789 42619
rect 2789 42585 2823 42619
rect 2823 42585 2832 42619
rect 2780 42576 2832 42585
rect 4896 42576 4948 42628
rect 5448 42576 5500 42628
rect 7380 42576 7432 42628
rect 11612 42576 11664 42628
rect 12256 42576 12308 42628
rect 22284 42712 22336 42764
rect 23848 42755 23900 42764
rect 23848 42721 23857 42755
rect 23857 42721 23891 42755
rect 23891 42721 23900 42755
rect 23848 42712 23900 42721
rect 24032 42755 24084 42764
rect 24032 42721 24041 42755
rect 24041 42721 24075 42755
rect 24075 42721 24084 42755
rect 24032 42712 24084 42721
rect 26700 42755 26752 42764
rect 26700 42721 26709 42755
rect 26709 42721 26743 42755
rect 26743 42721 26752 42755
rect 26700 42712 26752 42721
rect 27988 42755 28040 42764
rect 27988 42721 27997 42755
rect 27997 42721 28031 42755
rect 28031 42721 28040 42755
rect 27988 42712 28040 42721
rect 22192 42644 22244 42696
rect 23204 42687 23256 42696
rect 23204 42653 23213 42687
rect 23213 42653 23247 42687
rect 23247 42653 23256 42687
rect 23204 42644 23256 42653
rect 24492 42644 24544 42696
rect 25504 42576 25556 42628
rect 1952 42551 2004 42560
rect 1952 42517 1961 42551
rect 1961 42517 1995 42551
rect 1995 42517 2004 42551
rect 1952 42508 2004 42517
rect 3884 42508 3936 42560
rect 4252 42508 4304 42560
rect 8852 42508 8904 42560
rect 11060 42508 11112 42560
rect 13176 42508 13228 42560
rect 19800 42551 19852 42560
rect 19800 42517 19809 42551
rect 19809 42517 19843 42551
rect 19843 42517 19852 42551
rect 19800 42508 19852 42517
rect 23296 42508 23348 42560
rect 26148 42508 26200 42560
rect 26608 42508 26660 42560
rect 28080 42551 28132 42560
rect 28080 42517 28089 42551
rect 28089 42517 28123 42551
rect 28123 42517 28132 42551
rect 28080 42508 28132 42517
rect 5614 42406 5666 42458
rect 5678 42406 5730 42458
rect 5742 42406 5794 42458
rect 5806 42406 5858 42458
rect 14878 42406 14930 42458
rect 14942 42406 14994 42458
rect 15006 42406 15058 42458
rect 15070 42406 15122 42458
rect 24142 42406 24194 42458
rect 24206 42406 24258 42458
rect 24270 42406 24322 42458
rect 24334 42406 24386 42458
rect 2596 42304 2648 42356
rect 22192 42347 22244 42356
rect 2872 42236 2924 42288
rect 13636 42279 13688 42288
rect 4344 42211 4396 42220
rect 4344 42177 4353 42211
rect 4353 42177 4387 42211
rect 4387 42177 4396 42211
rect 4344 42168 4396 42177
rect 1216 42100 1268 42152
rect 3976 42100 4028 42152
rect 4252 42143 4304 42152
rect 4252 42109 4261 42143
rect 4261 42109 4295 42143
rect 4295 42109 4304 42143
rect 4252 42100 4304 42109
rect 4528 42100 4580 42152
rect 13636 42245 13645 42279
rect 13645 42245 13679 42279
rect 13679 42245 13688 42279
rect 13636 42236 13688 42245
rect 15292 42279 15344 42288
rect 15292 42245 15301 42279
rect 15301 42245 15335 42279
rect 15335 42245 15344 42279
rect 15292 42236 15344 42245
rect 7656 42168 7708 42220
rect 9404 42100 9456 42152
rect 9680 42168 9732 42220
rect 12256 42211 12308 42220
rect 12256 42177 12265 42211
rect 12265 42177 12299 42211
rect 12299 42177 12308 42211
rect 12256 42168 12308 42177
rect 16672 42211 16724 42220
rect 10140 42100 10192 42152
rect 12348 42100 12400 42152
rect 16672 42177 16681 42211
rect 16681 42177 16715 42211
rect 16715 42177 16724 42211
rect 16672 42168 16724 42177
rect 19340 42236 19392 42288
rect 19708 42236 19760 42288
rect 22192 42313 22201 42347
rect 22201 42313 22235 42347
rect 22235 42313 22244 42347
rect 22192 42304 22244 42313
rect 24032 42304 24084 42356
rect 28080 42304 28132 42356
rect 25412 42236 25464 42288
rect 18788 42168 18840 42220
rect 22376 42168 22428 42220
rect 23020 42168 23072 42220
rect 1492 42032 1544 42084
rect 2688 42032 2740 42084
rect 4988 42007 5040 42016
rect 4988 41973 4997 42007
rect 4997 41973 5031 42007
rect 5031 41973 5040 42007
rect 4988 41964 5040 41973
rect 9772 42007 9824 42016
rect 9772 41973 9781 42007
rect 9781 41973 9815 42007
rect 9815 41973 9824 42007
rect 9772 41964 9824 41973
rect 12440 42032 12492 42084
rect 14280 42032 14332 42084
rect 14556 42032 14608 42084
rect 16396 42007 16448 42016
rect 16396 41973 16405 42007
rect 16405 41973 16439 42007
rect 16439 41973 16448 42007
rect 16396 41964 16448 41973
rect 16580 41964 16632 42016
rect 17500 42032 17552 42084
rect 17868 42075 17920 42084
rect 17868 42041 17877 42075
rect 17877 42041 17911 42075
rect 17911 42041 17920 42075
rect 17868 42032 17920 42041
rect 22192 42100 22244 42152
rect 22744 42100 22796 42152
rect 23296 42143 23348 42152
rect 23296 42109 23305 42143
rect 23305 42109 23339 42143
rect 23339 42109 23348 42143
rect 23296 42100 23348 42109
rect 23848 42168 23900 42220
rect 25596 42168 25648 42220
rect 25412 42143 25464 42152
rect 18420 42032 18472 42084
rect 25412 42109 25421 42143
rect 25421 42109 25455 42143
rect 25455 42109 25464 42143
rect 25412 42100 25464 42109
rect 26608 42100 26660 42152
rect 27436 42100 27488 42152
rect 26332 42075 26384 42084
rect 26332 42041 26366 42075
rect 26366 42041 26384 42075
rect 26332 42032 26384 42041
rect 25596 41964 25648 42016
rect 27896 41964 27948 42016
rect 10246 41862 10298 41914
rect 10310 41862 10362 41914
rect 10374 41862 10426 41914
rect 10438 41862 10490 41914
rect 19510 41862 19562 41914
rect 19574 41862 19626 41914
rect 19638 41862 19690 41914
rect 19702 41862 19754 41914
rect 1492 41803 1544 41812
rect 1492 41769 1501 41803
rect 1501 41769 1535 41803
rect 1535 41769 1544 41803
rect 1492 41760 1544 41769
rect 2872 41760 2924 41812
rect 4252 41760 4304 41812
rect 5356 41760 5408 41812
rect 7656 41803 7708 41812
rect 7656 41769 7665 41803
rect 7665 41769 7699 41803
rect 7699 41769 7708 41803
rect 7656 41760 7708 41769
rect 8760 41803 8812 41812
rect 8760 41769 8769 41803
rect 8769 41769 8803 41803
rect 8803 41769 8812 41803
rect 8760 41760 8812 41769
rect 9680 41760 9732 41812
rect 10140 41760 10192 41812
rect 17500 41803 17552 41812
rect 2504 41692 2556 41744
rect 13176 41735 13228 41744
rect 13176 41701 13185 41735
rect 13185 41701 13219 41735
rect 13219 41701 13228 41735
rect 13176 41692 13228 41701
rect 17500 41769 17509 41803
rect 17509 41769 17543 41803
rect 17543 41769 17552 41803
rect 17500 41760 17552 41769
rect 19340 41760 19392 41812
rect 19800 41760 19852 41812
rect 26332 41803 26384 41812
rect 26332 41769 26341 41803
rect 26341 41769 26375 41803
rect 26375 41769 26384 41803
rect 26332 41760 26384 41769
rect 3056 41624 3108 41676
rect 3700 41667 3752 41676
rect 3700 41633 3709 41667
rect 3709 41633 3743 41667
rect 3743 41633 3752 41667
rect 3700 41624 3752 41633
rect 8116 41624 8168 41676
rect 8484 41624 8536 41676
rect 8852 41667 8904 41676
rect 8852 41633 8861 41667
rect 8861 41633 8895 41667
rect 8895 41633 8904 41667
rect 8852 41624 8904 41633
rect 9312 41667 9364 41676
rect 9312 41633 9321 41667
rect 9321 41633 9355 41667
rect 9355 41633 9364 41667
rect 9312 41624 9364 41633
rect 9588 41667 9640 41676
rect 9588 41633 9597 41667
rect 9597 41633 9631 41667
rect 9631 41633 9640 41667
rect 9588 41624 9640 41633
rect 2320 41556 2372 41608
rect 3148 41556 3200 41608
rect 3792 41556 3844 41608
rect 4620 41599 4672 41608
rect 4620 41565 4629 41599
rect 4629 41565 4663 41599
rect 4663 41565 4672 41599
rect 4620 41556 4672 41565
rect 3516 41488 3568 41540
rect 6184 41556 6236 41608
rect 7104 41556 7156 41608
rect 8300 41556 8352 41608
rect 9864 41624 9916 41676
rect 10140 41624 10192 41676
rect 12532 41624 12584 41676
rect 13636 41624 13688 41676
rect 4896 41531 4948 41540
rect 4896 41497 4905 41531
rect 4905 41497 4939 41531
rect 4939 41497 4948 41531
rect 4896 41488 4948 41497
rect 9864 41488 9916 41540
rect 13544 41556 13596 41608
rect 16120 41624 16172 41676
rect 16672 41624 16724 41676
rect 21456 41667 21508 41676
rect 21456 41633 21465 41667
rect 21465 41633 21499 41667
rect 21499 41633 21508 41667
rect 21456 41624 21508 41633
rect 23664 41624 23716 41676
rect 24124 41624 24176 41676
rect 24492 41667 24544 41676
rect 24492 41633 24501 41667
rect 24501 41633 24535 41667
rect 24535 41633 24544 41667
rect 24492 41624 24544 41633
rect 18052 41556 18104 41608
rect 19340 41556 19392 41608
rect 25228 41599 25280 41608
rect 25228 41565 25237 41599
rect 25237 41565 25271 41599
rect 25271 41565 25280 41599
rect 25228 41556 25280 41565
rect 26148 41599 26200 41608
rect 26148 41565 26157 41599
rect 26157 41565 26191 41599
rect 26191 41565 26200 41599
rect 26148 41556 26200 41565
rect 16396 41488 16448 41540
rect 23940 41488 23992 41540
rect 25964 41488 26016 41540
rect 27068 41624 27120 41676
rect 4252 41420 4304 41472
rect 5908 41420 5960 41472
rect 7196 41463 7248 41472
rect 7196 41429 7205 41463
rect 7205 41429 7239 41463
rect 7239 41429 7248 41463
rect 7196 41420 7248 41429
rect 9496 41420 9548 41472
rect 14648 41420 14700 41472
rect 18880 41420 18932 41472
rect 21088 41420 21140 41472
rect 5614 41318 5666 41370
rect 5678 41318 5730 41370
rect 5742 41318 5794 41370
rect 5806 41318 5858 41370
rect 14878 41318 14930 41370
rect 14942 41318 14994 41370
rect 15006 41318 15058 41370
rect 15070 41318 15122 41370
rect 24142 41318 24194 41370
rect 24206 41318 24258 41370
rect 24270 41318 24322 41370
rect 24334 41318 24386 41370
rect 2412 41216 2464 41268
rect 8116 41259 8168 41268
rect 1492 41148 1544 41200
rect 3976 41080 4028 41132
rect 4252 41055 4304 41064
rect 4252 41021 4261 41055
rect 4261 41021 4295 41055
rect 4295 41021 4304 41055
rect 4252 41012 4304 41021
rect 5540 41012 5592 41064
rect 6644 41148 6696 41200
rect 8116 41225 8125 41259
rect 8125 41225 8159 41259
rect 8159 41225 8168 41259
rect 8116 41216 8168 41225
rect 27068 41216 27120 41268
rect 7380 41123 7432 41132
rect 7380 41089 7389 41123
rect 7389 41089 7423 41123
rect 7423 41089 7432 41123
rect 7380 41080 7432 41089
rect 9220 41080 9272 41132
rect 9772 41055 9824 41064
rect 9772 41021 9806 41055
rect 9806 41021 9824 41055
rect 9772 41012 9824 41021
rect 12808 41012 12860 41064
rect 13452 41148 13504 41200
rect 25412 41148 25464 41200
rect 13636 41080 13688 41132
rect 15200 41080 15252 41132
rect 16120 41080 16172 41132
rect 16488 41080 16540 41132
rect 2136 40987 2188 40996
rect 2136 40953 2145 40987
rect 2145 40953 2179 40987
rect 2179 40953 2188 40987
rect 2136 40944 2188 40953
rect 2228 40944 2280 40996
rect 3056 40987 3108 40996
rect 3056 40953 3065 40987
rect 3065 40953 3099 40987
rect 3099 40953 3108 40987
rect 3056 40944 3108 40953
rect 6644 40944 6696 40996
rect 7840 40944 7892 40996
rect 2504 40876 2556 40928
rect 3148 40919 3200 40928
rect 3148 40885 3157 40919
rect 3157 40885 3191 40919
rect 3191 40885 3200 40919
rect 3148 40876 3200 40885
rect 4344 40919 4396 40928
rect 4344 40885 4353 40919
rect 4353 40885 4387 40919
rect 4387 40885 4396 40919
rect 4344 40876 4396 40885
rect 7104 40876 7156 40928
rect 9864 40876 9916 40928
rect 12716 40944 12768 40996
rect 14648 41012 14700 41064
rect 15384 41012 15436 41064
rect 20996 41080 21048 41132
rect 23296 41123 23348 41132
rect 23296 41089 23305 41123
rect 23305 41089 23339 41123
rect 23339 41089 23348 41123
rect 23296 41080 23348 41089
rect 23664 41080 23716 41132
rect 13268 40987 13320 40996
rect 13268 40953 13277 40987
rect 13277 40953 13311 40987
rect 13311 40953 13320 40987
rect 13268 40944 13320 40953
rect 16764 40944 16816 40996
rect 17040 40919 17092 40928
rect 17040 40885 17049 40919
rect 17049 40885 17083 40919
rect 17083 40885 17092 40919
rect 17040 40876 17092 40885
rect 22192 41055 22244 41064
rect 22192 41021 22201 41055
rect 22201 41021 22235 41055
rect 22235 41021 22244 41055
rect 22192 41012 22244 41021
rect 23020 41012 23072 41064
rect 23848 41055 23900 41064
rect 23848 41021 23857 41055
rect 23857 41021 23891 41055
rect 23891 41021 23900 41055
rect 23848 41012 23900 41021
rect 24952 41012 25004 41064
rect 25320 41012 25372 41064
rect 25504 41055 25556 41064
rect 25504 41021 25513 41055
rect 25513 41021 25547 41055
rect 25547 41021 25556 41055
rect 25504 41012 25556 41021
rect 26148 41055 26200 41064
rect 26148 41021 26157 41055
rect 26157 41021 26191 41055
rect 26191 41021 26200 41055
rect 26148 41012 26200 41021
rect 26792 41055 26844 41064
rect 26792 41021 26801 41055
rect 26801 41021 26835 41055
rect 26835 41021 26844 41055
rect 26792 41012 26844 41021
rect 27528 41012 27580 41064
rect 23664 40944 23716 40996
rect 20536 40919 20588 40928
rect 20536 40885 20545 40919
rect 20545 40885 20579 40919
rect 20579 40885 20588 40919
rect 20536 40876 20588 40885
rect 21456 40876 21508 40928
rect 22192 40919 22244 40928
rect 22192 40885 22201 40919
rect 22201 40885 22235 40919
rect 22235 40885 22244 40919
rect 22192 40876 22244 40885
rect 26608 40919 26660 40928
rect 26608 40885 26617 40919
rect 26617 40885 26651 40919
rect 26651 40885 26660 40919
rect 26608 40876 26660 40885
rect 27252 40876 27304 40928
rect 10246 40774 10298 40826
rect 10310 40774 10362 40826
rect 10374 40774 10426 40826
rect 10438 40774 10490 40826
rect 19510 40774 19562 40826
rect 19574 40774 19626 40826
rect 19638 40774 19690 40826
rect 19702 40774 19754 40826
rect 2504 40715 2556 40724
rect 2504 40681 2513 40715
rect 2513 40681 2547 40715
rect 2547 40681 2556 40715
rect 2504 40672 2556 40681
rect 2136 40604 2188 40656
rect 7196 40672 7248 40724
rect 2688 40536 2740 40588
rect 3700 40579 3752 40588
rect 3700 40545 3709 40579
rect 3709 40545 3743 40579
rect 3743 40545 3752 40579
rect 3700 40536 3752 40545
rect 4896 40604 4948 40656
rect 7656 40672 7708 40724
rect 10968 40672 11020 40724
rect 13820 40672 13872 40724
rect 21456 40672 21508 40724
rect 4988 40536 5040 40588
rect 5356 40536 5408 40588
rect 6184 40536 6236 40588
rect 7196 40579 7248 40588
rect 7196 40545 7205 40579
rect 7205 40545 7239 40579
rect 7239 40545 7248 40579
rect 7196 40536 7248 40545
rect 12716 40579 12768 40588
rect 12716 40545 12725 40579
rect 12725 40545 12759 40579
rect 12759 40545 12768 40579
rect 12716 40536 12768 40545
rect 13084 40579 13136 40588
rect 3332 40468 3384 40520
rect 3608 40468 3660 40520
rect 4896 40468 4948 40520
rect 5264 40468 5316 40520
rect 9956 40468 10008 40520
rect 11888 40468 11940 40520
rect 12440 40468 12492 40520
rect 4252 40400 4304 40452
rect 4620 40400 4672 40452
rect 4988 40443 5040 40452
rect 4988 40409 4997 40443
rect 4997 40409 5031 40443
rect 5031 40409 5040 40443
rect 4988 40400 5040 40409
rect 7012 40400 7064 40452
rect 9772 40400 9824 40452
rect 12716 40400 12768 40452
rect 13084 40545 13093 40579
rect 13093 40545 13127 40579
rect 13127 40545 13136 40579
rect 13084 40536 13136 40545
rect 13728 40536 13780 40588
rect 14740 40536 14792 40588
rect 19432 40604 19484 40656
rect 20536 40604 20588 40656
rect 24032 40604 24084 40656
rect 26608 40604 26660 40656
rect 18052 40579 18104 40588
rect 18052 40545 18061 40579
rect 18061 40545 18095 40579
rect 18095 40545 18104 40579
rect 18052 40536 18104 40545
rect 18880 40579 18932 40588
rect 18880 40545 18889 40579
rect 18889 40545 18923 40579
rect 18923 40545 18932 40579
rect 18880 40536 18932 40545
rect 18972 40536 19024 40588
rect 20076 40536 20128 40588
rect 23664 40536 23716 40588
rect 23848 40579 23900 40588
rect 23848 40545 23857 40579
rect 23857 40545 23891 40579
rect 23891 40545 23900 40579
rect 23848 40536 23900 40545
rect 24860 40536 24912 40588
rect 14280 40511 14332 40520
rect 14280 40477 14289 40511
rect 14289 40477 14323 40511
rect 14323 40477 14332 40511
rect 14280 40468 14332 40477
rect 19524 40511 19576 40520
rect 19524 40477 19533 40511
rect 19533 40477 19567 40511
rect 19567 40477 19576 40511
rect 19524 40468 19576 40477
rect 24492 40468 24544 40520
rect 26148 40511 26200 40520
rect 26148 40477 26157 40511
rect 26157 40477 26191 40511
rect 26191 40477 26200 40511
rect 26148 40468 26200 40477
rect 1952 40375 2004 40384
rect 1952 40341 1961 40375
rect 1961 40341 1995 40375
rect 1995 40341 2004 40375
rect 1952 40332 2004 40341
rect 3792 40375 3844 40384
rect 3792 40341 3801 40375
rect 3801 40341 3835 40375
rect 3835 40341 3844 40375
rect 3792 40332 3844 40341
rect 4160 40375 4212 40384
rect 4160 40341 4169 40375
rect 4169 40341 4203 40375
rect 4203 40341 4212 40375
rect 4160 40332 4212 40341
rect 5448 40332 5500 40384
rect 6920 40375 6972 40384
rect 6920 40341 6929 40375
rect 6929 40341 6963 40375
rect 6963 40341 6972 40375
rect 6920 40332 6972 40341
rect 9496 40332 9548 40384
rect 10692 40332 10744 40384
rect 12348 40332 12400 40384
rect 12808 40332 12860 40384
rect 13176 40332 13228 40384
rect 16672 40332 16724 40384
rect 25964 40332 26016 40384
rect 27988 40375 28040 40384
rect 27988 40341 27997 40375
rect 27997 40341 28031 40375
rect 28031 40341 28040 40375
rect 27988 40332 28040 40341
rect 5614 40230 5666 40282
rect 5678 40230 5730 40282
rect 5742 40230 5794 40282
rect 5806 40230 5858 40282
rect 14878 40230 14930 40282
rect 14942 40230 14994 40282
rect 15006 40230 15058 40282
rect 15070 40230 15122 40282
rect 24142 40230 24194 40282
rect 24206 40230 24258 40282
rect 24270 40230 24322 40282
rect 24334 40230 24386 40282
rect 3056 40128 3108 40180
rect 27988 40128 28040 40180
rect 13452 40060 13504 40112
rect 15108 40060 15160 40112
rect 17040 40060 17092 40112
rect 5448 39992 5500 40044
rect 7196 39992 7248 40044
rect 9588 39992 9640 40044
rect 9864 39992 9916 40044
rect 14004 39992 14056 40044
rect 4344 39924 4396 39976
rect 5080 39967 5132 39976
rect 5080 39933 5089 39967
rect 5089 39933 5123 39967
rect 5123 39933 5132 39967
rect 5080 39924 5132 39933
rect 6368 39967 6420 39976
rect 2412 39856 2464 39908
rect 2596 39899 2648 39908
rect 2596 39865 2605 39899
rect 2605 39865 2639 39899
rect 2639 39865 2648 39899
rect 2596 39856 2648 39865
rect 2780 39899 2832 39908
rect 2780 39865 2789 39899
rect 2789 39865 2823 39899
rect 2823 39865 2832 39899
rect 2780 39856 2832 39865
rect 4528 39856 4580 39908
rect 6368 39933 6377 39967
rect 6377 39933 6411 39967
rect 6411 39933 6420 39967
rect 6368 39924 6420 39933
rect 6552 39967 6604 39976
rect 6552 39933 6561 39967
rect 6561 39933 6595 39967
rect 6595 39933 6604 39967
rect 6552 39924 6604 39933
rect 7748 39924 7800 39976
rect 8484 39924 8536 39976
rect 8668 39924 8720 39976
rect 1400 39788 1452 39840
rect 6552 39788 6604 39840
rect 8116 39788 8168 39840
rect 10784 39924 10836 39976
rect 12532 39924 12584 39976
rect 13268 39924 13320 39976
rect 11980 39856 12032 39908
rect 13636 39967 13688 39976
rect 13636 39933 13645 39967
rect 13645 39933 13679 39967
rect 13679 39933 13688 39967
rect 13636 39924 13688 39933
rect 13912 39924 13964 39976
rect 13728 39856 13780 39908
rect 16764 39992 16816 40044
rect 18052 39992 18104 40044
rect 22468 40060 22520 40112
rect 22192 40035 22244 40044
rect 22192 40001 22201 40035
rect 22201 40001 22235 40035
rect 22235 40001 22244 40035
rect 22192 39992 22244 40001
rect 15384 39967 15436 39976
rect 15384 39933 15393 39967
rect 15393 39933 15427 39967
rect 15427 39933 15436 39967
rect 15384 39924 15436 39933
rect 16120 39924 16172 39976
rect 16488 39967 16540 39976
rect 16488 39933 16497 39967
rect 16497 39933 16531 39967
rect 16531 39933 16540 39967
rect 16488 39924 16540 39933
rect 15476 39856 15528 39908
rect 11060 39788 11112 39840
rect 12072 39831 12124 39840
rect 12072 39797 12081 39831
rect 12081 39797 12115 39831
rect 12115 39797 12124 39831
rect 12072 39788 12124 39797
rect 14372 39788 14424 39840
rect 14832 39788 14884 39840
rect 15200 39788 15252 39840
rect 15292 39788 15344 39840
rect 16672 39967 16724 39976
rect 16672 39933 16681 39967
rect 16681 39933 16715 39967
rect 16715 39933 16724 39967
rect 16672 39924 16724 39933
rect 16948 39924 17000 39976
rect 18420 39967 18472 39976
rect 18420 39933 18429 39967
rect 18429 39933 18463 39967
rect 18463 39933 18472 39967
rect 18420 39924 18472 39933
rect 21088 39967 21140 39976
rect 21088 39933 21097 39967
rect 21097 39933 21131 39967
rect 21131 39933 21140 39967
rect 21088 39924 21140 39933
rect 16764 39856 16816 39908
rect 18052 39856 18104 39908
rect 18604 39899 18656 39908
rect 18604 39865 18613 39899
rect 18613 39865 18647 39899
rect 18647 39865 18656 39899
rect 18604 39856 18656 39865
rect 18420 39788 18472 39840
rect 19524 39856 19576 39908
rect 20168 39856 20220 39908
rect 23204 39924 23256 39976
rect 23848 39992 23900 40044
rect 25228 39992 25280 40044
rect 25320 39992 25372 40044
rect 23664 39924 23716 39976
rect 24216 39924 24268 39976
rect 25412 39967 25464 39976
rect 25412 39933 25421 39967
rect 25421 39933 25455 39967
rect 25455 39933 25464 39967
rect 25412 39924 25464 39933
rect 25964 39924 26016 39976
rect 27896 39967 27948 39976
rect 27896 39933 27905 39967
rect 27905 39933 27939 39967
rect 27939 39933 27948 39967
rect 27896 39924 27948 39933
rect 24492 39856 24544 39908
rect 22652 39788 22704 39840
rect 23572 39788 23624 39840
rect 24400 39788 24452 39840
rect 25228 39831 25280 39840
rect 25228 39797 25237 39831
rect 25237 39797 25271 39831
rect 25271 39797 25280 39831
rect 25228 39788 25280 39797
rect 27344 39788 27396 39840
rect 10246 39686 10298 39738
rect 10310 39686 10362 39738
rect 10374 39686 10426 39738
rect 10438 39686 10490 39738
rect 19510 39686 19562 39738
rect 19574 39686 19626 39738
rect 19638 39686 19690 39738
rect 19702 39686 19754 39738
rect 3608 39584 3660 39636
rect 4160 39516 4212 39568
rect 11704 39584 11756 39636
rect 11980 39584 12032 39636
rect 12716 39584 12768 39636
rect 14280 39584 14332 39636
rect 10232 39516 10284 39568
rect 2228 39448 2280 39500
rect 2504 39448 2556 39500
rect 3884 39491 3936 39500
rect 3884 39457 3893 39491
rect 3893 39457 3927 39491
rect 3927 39457 3936 39491
rect 3884 39448 3936 39457
rect 3976 39491 4028 39500
rect 3976 39457 3985 39491
rect 3985 39457 4019 39491
rect 4019 39457 4028 39491
rect 3976 39448 4028 39457
rect 6920 39448 6972 39500
rect 2688 39380 2740 39432
rect 2872 39312 2924 39364
rect 2964 39244 3016 39296
rect 3792 39380 3844 39432
rect 6368 39380 6420 39432
rect 7104 39380 7156 39432
rect 8484 39448 8536 39500
rect 8668 39491 8720 39500
rect 8668 39457 8677 39491
rect 8677 39457 8711 39491
rect 8711 39457 8720 39491
rect 8668 39448 8720 39457
rect 9220 39448 9272 39500
rect 9864 39491 9916 39500
rect 9864 39457 9873 39491
rect 9873 39457 9907 39491
rect 9907 39457 9916 39491
rect 9864 39448 9916 39457
rect 10324 39491 10376 39500
rect 10324 39457 10333 39491
rect 10333 39457 10367 39491
rect 10367 39457 10376 39491
rect 10324 39448 10376 39457
rect 10508 39491 10560 39500
rect 10508 39457 10515 39491
rect 10515 39457 10560 39491
rect 10508 39448 10560 39457
rect 8576 39380 8628 39432
rect 5264 39312 5316 39364
rect 7748 39244 7800 39296
rect 8116 39312 8168 39364
rect 10232 39380 10284 39432
rect 10876 39448 10928 39500
rect 11060 39448 11112 39500
rect 11244 39448 11296 39500
rect 11428 39448 11480 39500
rect 12072 39448 12124 39500
rect 12440 39491 12492 39500
rect 12440 39457 12449 39491
rect 12449 39457 12483 39491
rect 12483 39457 12492 39491
rect 12440 39448 12492 39457
rect 12808 39448 12860 39500
rect 13820 39448 13872 39500
rect 14004 39448 14056 39500
rect 15384 39584 15436 39636
rect 20720 39584 20772 39636
rect 22652 39627 22704 39636
rect 22652 39593 22661 39627
rect 22661 39593 22695 39627
rect 22695 39593 22704 39627
rect 22652 39584 22704 39593
rect 14740 39516 14792 39568
rect 14556 39491 14608 39500
rect 13728 39380 13780 39432
rect 9312 39312 9364 39364
rect 12532 39312 12584 39364
rect 9680 39244 9732 39296
rect 9864 39244 9916 39296
rect 13636 39244 13688 39296
rect 14556 39457 14565 39491
rect 14565 39457 14599 39491
rect 14599 39457 14608 39491
rect 14556 39448 14608 39457
rect 14832 39448 14884 39500
rect 15108 39491 15160 39500
rect 15108 39457 15118 39491
rect 15118 39457 15152 39491
rect 15152 39457 15160 39491
rect 15292 39491 15344 39500
rect 15108 39448 15160 39457
rect 15292 39457 15301 39491
rect 15301 39457 15335 39491
rect 15335 39457 15344 39491
rect 15292 39448 15344 39457
rect 15384 39491 15436 39500
rect 15384 39457 15393 39491
rect 15393 39457 15427 39491
rect 15427 39457 15436 39491
rect 15384 39448 15436 39457
rect 15844 39516 15896 39568
rect 27344 39584 27396 39636
rect 25228 39516 25280 39568
rect 14648 39380 14700 39432
rect 18604 39448 18656 39500
rect 23664 39448 23716 39500
rect 24216 39448 24268 39500
rect 26884 39491 26936 39500
rect 26884 39457 26893 39491
rect 26893 39457 26927 39491
rect 26927 39457 26936 39491
rect 26884 39448 26936 39457
rect 17224 39380 17276 39432
rect 24400 39423 24452 39432
rect 24400 39389 24409 39423
rect 24409 39389 24443 39423
rect 24443 39389 24452 39423
rect 24400 39380 24452 39389
rect 24860 39423 24912 39432
rect 24860 39389 24869 39423
rect 24869 39389 24903 39423
rect 24903 39389 24912 39423
rect 24860 39380 24912 39389
rect 15476 39312 15528 39364
rect 15660 39287 15712 39296
rect 15660 39253 15669 39287
rect 15669 39253 15703 39287
rect 15703 39253 15712 39287
rect 15660 39244 15712 39253
rect 15844 39244 15896 39296
rect 28172 39312 28224 39364
rect 20076 39287 20128 39296
rect 20076 39253 20085 39287
rect 20085 39253 20119 39287
rect 20119 39253 20128 39287
rect 20076 39244 20128 39253
rect 23664 39244 23716 39296
rect 24492 39244 24544 39296
rect 27896 39244 27948 39296
rect 28080 39287 28132 39296
rect 28080 39253 28089 39287
rect 28089 39253 28123 39287
rect 28123 39253 28132 39287
rect 28080 39244 28132 39253
rect 5614 39142 5666 39194
rect 5678 39142 5730 39194
rect 5742 39142 5794 39194
rect 5806 39142 5858 39194
rect 14878 39142 14930 39194
rect 14942 39142 14994 39194
rect 15006 39142 15058 39194
rect 15070 39142 15122 39194
rect 24142 39142 24194 39194
rect 24206 39142 24258 39194
rect 24270 39142 24322 39194
rect 24334 39142 24386 39194
rect 2044 39040 2096 39092
rect 2688 39040 2740 39092
rect 3976 39040 4028 39092
rect 6184 39040 6236 39092
rect 8300 39040 8352 39092
rect 8484 39083 8536 39092
rect 8484 39049 8493 39083
rect 8493 39049 8527 39083
rect 8527 39049 8536 39083
rect 8484 39040 8536 39049
rect 1860 39015 1912 39024
rect 1860 38981 1869 39015
rect 1869 38981 1903 39015
rect 1903 38981 1912 39015
rect 1860 38972 1912 38981
rect 2596 38972 2648 39024
rect 1584 38904 1636 38956
rect 2044 38904 2096 38956
rect 3240 38879 3292 38888
rect 3240 38845 3249 38879
rect 3249 38845 3283 38879
rect 3283 38845 3292 38879
rect 3240 38836 3292 38845
rect 3884 38836 3936 38888
rect 3056 38768 3108 38820
rect 4528 38879 4580 38888
rect 4528 38845 4537 38879
rect 4537 38845 4571 38879
rect 4571 38845 4580 38879
rect 4528 38836 4580 38845
rect 5264 38836 5316 38888
rect 6920 38836 6972 38888
rect 7748 38879 7800 38888
rect 7748 38845 7757 38879
rect 7757 38845 7791 38879
rect 7791 38845 7800 38879
rect 7748 38836 7800 38845
rect 8116 38904 8168 38956
rect 9680 38904 9732 38956
rect 11428 38972 11480 39024
rect 11612 39015 11664 39024
rect 11612 38981 11621 39015
rect 11621 38981 11655 39015
rect 11655 38981 11664 39015
rect 11612 38972 11664 38981
rect 12164 39040 12216 39092
rect 15660 39040 15712 39092
rect 22284 39040 22336 39092
rect 16672 38972 16724 39024
rect 18972 39015 19024 39024
rect 18972 38981 18981 39015
rect 18981 38981 19015 39015
rect 19015 38981 19024 39015
rect 18972 38972 19024 38981
rect 7104 38768 7156 38820
rect 9864 38879 9916 38888
rect 9864 38845 9873 38879
rect 9873 38845 9907 38879
rect 9907 38845 9916 38879
rect 9864 38836 9916 38845
rect 10232 38836 10284 38888
rect 9588 38768 9640 38820
rect 11244 38904 11296 38956
rect 10508 38768 10560 38820
rect 11520 38836 11572 38888
rect 12072 38836 12124 38888
rect 14648 38836 14700 38888
rect 16580 38836 16632 38888
rect 16764 38879 16816 38888
rect 16764 38845 16773 38879
rect 16773 38845 16807 38879
rect 16807 38845 16816 38879
rect 16764 38836 16816 38845
rect 17040 38879 17092 38888
rect 17040 38845 17049 38879
rect 17049 38845 17083 38879
rect 17083 38845 17092 38879
rect 17040 38836 17092 38845
rect 3884 38700 3936 38752
rect 4344 38700 4396 38752
rect 4804 38700 4856 38752
rect 11704 38768 11756 38820
rect 17224 38836 17276 38888
rect 28080 39040 28132 39092
rect 22468 38904 22520 38956
rect 27804 38972 27856 39024
rect 28172 39015 28224 39024
rect 28172 38981 28181 39015
rect 28181 38981 28215 39015
rect 28215 38981 28224 39015
rect 28172 38972 28224 38981
rect 22652 38836 22704 38888
rect 17408 38768 17460 38820
rect 11612 38700 11664 38752
rect 11980 38700 12032 38752
rect 12532 38700 12584 38752
rect 14740 38743 14792 38752
rect 14740 38709 14749 38743
rect 14749 38709 14783 38743
rect 14783 38709 14792 38743
rect 14740 38700 14792 38709
rect 16396 38743 16448 38752
rect 16396 38709 16405 38743
rect 16405 38709 16439 38743
rect 16439 38709 16448 38743
rect 16396 38700 16448 38709
rect 20168 38700 20220 38752
rect 26056 38879 26108 38888
rect 26056 38845 26065 38879
rect 26065 38845 26099 38879
rect 26099 38845 26108 38879
rect 26056 38836 26108 38845
rect 26792 38836 26844 38888
rect 27252 38879 27304 38888
rect 27252 38845 27261 38879
rect 27261 38845 27295 38879
rect 27295 38845 27304 38879
rect 27252 38836 27304 38845
rect 22744 38743 22796 38752
rect 22744 38709 22753 38743
rect 22753 38709 22787 38743
rect 22787 38709 22796 38743
rect 22744 38700 22796 38709
rect 25504 38700 25556 38752
rect 25872 38700 25924 38752
rect 10246 38598 10298 38650
rect 10310 38598 10362 38650
rect 10374 38598 10426 38650
rect 10438 38598 10490 38650
rect 19510 38598 19562 38650
rect 19574 38598 19626 38650
rect 19638 38598 19690 38650
rect 19702 38598 19754 38650
rect 1860 38428 1912 38480
rect 20076 38539 20128 38548
rect 20076 38505 20085 38539
rect 20085 38505 20119 38539
rect 20119 38505 20128 38539
rect 20076 38496 20128 38505
rect 3056 38428 3108 38480
rect 2596 38360 2648 38412
rect 1584 38224 1636 38276
rect 2228 38156 2280 38208
rect 2780 38199 2832 38208
rect 2780 38165 2789 38199
rect 2789 38165 2823 38199
rect 2823 38165 2832 38199
rect 4160 38428 4212 38480
rect 4528 38471 4580 38480
rect 4528 38437 4537 38471
rect 4537 38437 4571 38471
rect 4571 38437 4580 38471
rect 4528 38428 4580 38437
rect 5080 38428 5132 38480
rect 9496 38428 9548 38480
rect 9680 38428 9732 38480
rect 11520 38428 11572 38480
rect 4620 38360 4672 38412
rect 3884 38292 3936 38344
rect 5908 38360 5960 38412
rect 8852 38360 8904 38412
rect 9036 38335 9088 38344
rect 9036 38301 9045 38335
rect 9045 38301 9079 38335
rect 9079 38301 9088 38335
rect 9036 38292 9088 38301
rect 9220 38335 9272 38344
rect 9220 38301 9229 38335
rect 9229 38301 9263 38335
rect 9263 38301 9272 38335
rect 9220 38292 9272 38301
rect 9404 38292 9456 38344
rect 10508 38403 10560 38412
rect 10508 38369 10518 38403
rect 10518 38369 10552 38403
rect 10552 38369 10560 38403
rect 10784 38403 10836 38412
rect 10508 38360 10560 38369
rect 10784 38369 10793 38403
rect 10793 38369 10827 38403
rect 10827 38369 10836 38403
rect 10784 38360 10836 38369
rect 10876 38403 10928 38412
rect 10876 38369 10890 38403
rect 10890 38369 10924 38403
rect 10924 38369 10928 38403
rect 10876 38360 10928 38369
rect 9864 38224 9916 38276
rect 11428 38292 11480 38344
rect 13268 38360 13320 38412
rect 15292 38360 15344 38412
rect 16396 38428 16448 38480
rect 28080 38496 28132 38548
rect 11980 38292 12032 38344
rect 17224 38292 17276 38344
rect 18420 38292 18472 38344
rect 27252 38428 27304 38480
rect 27896 38471 27948 38480
rect 27896 38437 27905 38471
rect 27905 38437 27939 38471
rect 27939 38437 27948 38471
rect 27896 38428 27948 38437
rect 20904 38360 20956 38412
rect 20352 38292 20404 38344
rect 21272 38360 21324 38412
rect 25044 38360 25096 38412
rect 26148 38360 26200 38412
rect 26884 38403 26936 38412
rect 26884 38369 26893 38403
rect 26893 38369 26927 38403
rect 26927 38369 26936 38403
rect 26884 38360 26936 38369
rect 18788 38224 18840 38276
rect 22192 38292 22244 38344
rect 21364 38224 21416 38276
rect 22652 38224 22704 38276
rect 2780 38156 2832 38165
rect 4160 38156 4212 38208
rect 4528 38156 4580 38208
rect 5356 38156 5408 38208
rect 6184 38156 6236 38208
rect 11336 38156 11388 38208
rect 12072 38156 12124 38208
rect 13544 38156 13596 38208
rect 14372 38156 14424 38208
rect 15200 38199 15252 38208
rect 15200 38165 15209 38199
rect 15209 38165 15243 38199
rect 15243 38165 15252 38199
rect 15200 38156 15252 38165
rect 17960 38156 18012 38208
rect 20444 38156 20496 38208
rect 21088 38156 21140 38208
rect 23112 38156 23164 38208
rect 23204 38156 23256 38208
rect 24860 38156 24912 38208
rect 25320 38156 25372 38208
rect 25872 38156 25924 38208
rect 26056 38199 26108 38208
rect 26056 38165 26065 38199
rect 26065 38165 26099 38199
rect 26099 38165 26108 38199
rect 26056 38156 26108 38165
rect 26700 38199 26752 38208
rect 26700 38165 26709 38199
rect 26709 38165 26743 38199
rect 26743 38165 26752 38199
rect 26700 38156 26752 38165
rect 27988 38199 28040 38208
rect 27988 38165 27997 38199
rect 27997 38165 28031 38199
rect 28031 38165 28040 38199
rect 27988 38156 28040 38165
rect 5614 38054 5666 38106
rect 5678 38054 5730 38106
rect 5742 38054 5794 38106
rect 5806 38054 5858 38106
rect 14878 38054 14930 38106
rect 14942 38054 14994 38106
rect 15006 38054 15058 38106
rect 15070 38054 15122 38106
rect 24142 38054 24194 38106
rect 24206 38054 24258 38106
rect 24270 38054 24322 38106
rect 24334 38054 24386 38106
rect 2872 37952 2924 38004
rect 3240 37952 3292 38004
rect 22192 37995 22244 38004
rect 1400 37816 1452 37868
rect 1584 37816 1636 37868
rect 13360 37884 13412 37936
rect 16672 37884 16724 37936
rect 20076 37884 20128 37936
rect 20352 37884 20404 37936
rect 22192 37961 22201 37995
rect 22201 37961 22235 37995
rect 22235 37961 22244 37995
rect 22192 37952 22244 37961
rect 27252 37995 27304 38004
rect 27252 37961 27261 37995
rect 27261 37961 27295 37995
rect 27295 37961 27304 37995
rect 27252 37952 27304 37961
rect 27988 37884 28040 37936
rect 4160 37816 4212 37868
rect 11612 37816 11664 37868
rect 2228 37748 2280 37800
rect 1584 37723 1636 37732
rect 1584 37689 1593 37723
rect 1593 37689 1627 37723
rect 1627 37689 1636 37723
rect 1584 37680 1636 37689
rect 2596 37748 2648 37800
rect 3148 37791 3200 37800
rect 3148 37757 3157 37791
rect 3157 37757 3191 37791
rect 3191 37757 3200 37791
rect 4252 37791 4304 37800
rect 3148 37748 3200 37757
rect 4252 37757 4261 37791
rect 4261 37757 4295 37791
rect 4295 37757 4304 37791
rect 4252 37748 4304 37757
rect 3056 37680 3108 37732
rect 1676 37655 1728 37664
rect 1676 37621 1685 37655
rect 1685 37621 1719 37655
rect 1719 37621 1728 37655
rect 1676 37612 1728 37621
rect 2504 37612 2556 37664
rect 2872 37612 2924 37664
rect 3424 37612 3476 37664
rect 5908 37748 5960 37800
rect 11152 37748 11204 37800
rect 11980 37791 12032 37800
rect 11980 37757 11989 37791
rect 11989 37757 12023 37791
rect 12023 37757 12032 37791
rect 11980 37748 12032 37757
rect 5356 37723 5408 37732
rect 5356 37689 5390 37723
rect 5390 37689 5408 37723
rect 5356 37680 5408 37689
rect 9956 37680 10008 37732
rect 10232 37680 10284 37732
rect 10968 37680 11020 37732
rect 12072 37680 12124 37732
rect 13360 37748 13412 37800
rect 13728 37748 13780 37800
rect 14004 37748 14056 37800
rect 14740 37748 14792 37800
rect 15384 37748 15436 37800
rect 15660 37791 15712 37800
rect 15660 37757 15667 37791
rect 15667 37757 15712 37791
rect 15660 37748 15712 37757
rect 16028 37816 16080 37868
rect 18604 37816 18656 37868
rect 20812 37859 20864 37868
rect 20812 37825 20821 37859
rect 20821 37825 20855 37859
rect 20855 37825 20864 37859
rect 20812 37816 20864 37825
rect 22744 37816 22796 37868
rect 25872 37859 25924 37868
rect 25872 37825 25881 37859
rect 25881 37825 25915 37859
rect 25915 37825 25924 37859
rect 25872 37816 25924 37825
rect 25964 37859 26016 37868
rect 25964 37825 25973 37859
rect 25973 37825 26007 37859
rect 26007 37825 26016 37859
rect 25964 37816 26016 37825
rect 15936 37791 15988 37800
rect 15936 37757 15950 37791
rect 15950 37757 15984 37791
rect 15984 37757 15988 37791
rect 15936 37748 15988 37757
rect 14832 37723 14884 37732
rect 14832 37689 14841 37723
rect 14841 37689 14875 37723
rect 14875 37689 14884 37723
rect 14832 37680 14884 37689
rect 16580 37748 16632 37800
rect 20076 37791 20128 37800
rect 20076 37757 20085 37791
rect 20085 37757 20119 37791
rect 20119 37757 20128 37791
rect 20076 37748 20128 37757
rect 20168 37748 20220 37800
rect 21088 37791 21140 37800
rect 21088 37757 21122 37791
rect 21122 37757 21140 37791
rect 21088 37748 21140 37757
rect 23112 37791 23164 37800
rect 23112 37757 23121 37791
rect 23121 37757 23155 37791
rect 23155 37757 23164 37791
rect 23112 37748 23164 37757
rect 24032 37748 24084 37800
rect 26056 37748 26108 37800
rect 27804 37748 27856 37800
rect 16488 37680 16540 37732
rect 25320 37680 25372 37732
rect 6828 37612 6880 37664
rect 11520 37655 11572 37664
rect 11520 37621 11529 37655
rect 11529 37621 11563 37655
rect 11563 37621 11572 37655
rect 11520 37612 11572 37621
rect 11980 37612 12032 37664
rect 12348 37612 12400 37664
rect 13452 37612 13504 37664
rect 13820 37612 13872 37664
rect 15476 37612 15528 37664
rect 15568 37612 15620 37664
rect 15936 37612 15988 37664
rect 20352 37612 20404 37664
rect 25412 37655 25464 37664
rect 25412 37621 25421 37655
rect 25421 37621 25455 37655
rect 25455 37621 25464 37655
rect 25412 37612 25464 37621
rect 27344 37612 27396 37664
rect 10246 37510 10298 37562
rect 10310 37510 10362 37562
rect 10374 37510 10426 37562
rect 10438 37510 10490 37562
rect 19510 37510 19562 37562
rect 19574 37510 19626 37562
rect 19638 37510 19690 37562
rect 19702 37510 19754 37562
rect 2412 37408 2464 37460
rect 13452 37408 13504 37460
rect 13820 37408 13872 37460
rect 27344 37408 27396 37460
rect 28080 37451 28132 37460
rect 28080 37417 28089 37451
rect 28089 37417 28123 37451
rect 28123 37417 28132 37451
rect 28080 37408 28132 37417
rect 2872 37340 2924 37392
rect 5356 37383 5408 37392
rect 2412 37272 2464 37324
rect 2596 37315 2648 37324
rect 2596 37281 2605 37315
rect 2605 37281 2639 37315
rect 2639 37281 2648 37315
rect 2596 37272 2648 37281
rect 3516 37315 3568 37324
rect 3516 37281 3525 37315
rect 3525 37281 3559 37315
rect 3559 37281 3568 37315
rect 3516 37272 3568 37281
rect 4528 37272 4580 37324
rect 4804 37315 4856 37324
rect 3608 37247 3660 37256
rect 3608 37213 3617 37247
rect 3617 37213 3651 37247
rect 3651 37213 3660 37247
rect 3608 37204 3660 37213
rect 4804 37281 4813 37315
rect 4813 37281 4847 37315
rect 4847 37281 4856 37315
rect 4804 37272 4856 37281
rect 4896 37204 4948 37256
rect 5356 37349 5365 37383
rect 5365 37349 5399 37383
rect 5399 37349 5408 37383
rect 5356 37340 5408 37349
rect 8760 37340 8812 37392
rect 5264 37315 5316 37324
rect 5264 37281 5273 37315
rect 5273 37281 5307 37315
rect 5307 37281 5316 37315
rect 5264 37272 5316 37281
rect 2780 37179 2832 37188
rect 2780 37145 2789 37179
rect 2789 37145 2823 37179
rect 2823 37145 2832 37179
rect 2780 37136 2832 37145
rect 3976 37136 4028 37188
rect 4436 37136 4488 37188
rect 8852 37272 8904 37324
rect 9864 37315 9916 37324
rect 9864 37281 9873 37315
rect 9873 37281 9907 37315
rect 9907 37281 9916 37315
rect 9864 37272 9916 37281
rect 10876 37340 10928 37392
rect 12072 37383 12124 37392
rect 12072 37349 12081 37383
rect 12081 37349 12115 37383
rect 12115 37349 12124 37383
rect 12072 37340 12124 37349
rect 12164 37340 12216 37392
rect 11520 37272 11572 37324
rect 12256 37272 12308 37324
rect 12716 37315 12768 37324
rect 12164 37204 12216 37256
rect 12716 37281 12725 37315
rect 12725 37281 12759 37315
rect 12759 37281 12768 37315
rect 12716 37272 12768 37281
rect 13268 37340 13320 37392
rect 13728 37340 13780 37392
rect 14004 37340 14056 37392
rect 13452 37315 13504 37324
rect 13452 37281 13461 37315
rect 13461 37281 13495 37315
rect 13495 37281 13504 37315
rect 13452 37272 13504 37281
rect 13820 37281 13829 37286
rect 13829 37281 13863 37286
rect 13863 37281 13872 37286
rect 13820 37234 13872 37281
rect 14832 37340 14884 37392
rect 15568 37340 15620 37392
rect 15660 37340 15712 37392
rect 20352 37383 20404 37392
rect 14740 37315 14792 37324
rect 14740 37281 14749 37315
rect 14749 37281 14783 37315
rect 14783 37281 14792 37315
rect 14740 37272 14792 37281
rect 15292 37272 15344 37324
rect 17960 37272 18012 37324
rect 20352 37349 20361 37383
rect 20361 37349 20395 37383
rect 20395 37349 20404 37383
rect 20352 37340 20404 37349
rect 20444 37383 20496 37392
rect 20444 37349 20453 37383
rect 20453 37349 20487 37383
rect 20487 37349 20496 37383
rect 20444 37340 20496 37349
rect 20904 37340 20956 37392
rect 21272 37383 21324 37392
rect 21272 37349 21281 37383
rect 21281 37349 21315 37383
rect 21315 37349 21324 37383
rect 21272 37340 21324 37349
rect 21364 37340 21416 37392
rect 25044 37383 25096 37392
rect 21088 37272 21140 37324
rect 22744 37272 22796 37324
rect 25044 37349 25053 37383
rect 25053 37349 25087 37383
rect 25087 37349 25096 37383
rect 25044 37340 25096 37349
rect 26700 37340 26752 37392
rect 15660 37204 15712 37256
rect 17224 37204 17276 37256
rect 18052 37247 18104 37256
rect 18052 37213 18061 37247
rect 18061 37213 18095 37247
rect 18095 37213 18104 37247
rect 18052 37204 18104 37213
rect 20352 37204 20404 37256
rect 25320 37272 25372 37324
rect 25412 37272 25464 37324
rect 25780 37247 25832 37256
rect 11152 37136 11204 37188
rect 11520 37136 11572 37188
rect 14372 37136 14424 37188
rect 7288 37068 7340 37120
rect 15200 37136 15252 37188
rect 17868 37136 17920 37188
rect 14740 37068 14792 37120
rect 19340 37068 19392 37120
rect 20904 37068 20956 37120
rect 20996 37068 21048 37120
rect 25780 37213 25789 37247
rect 25789 37213 25823 37247
rect 25823 37213 25832 37247
rect 25780 37204 25832 37213
rect 26976 37272 27028 37324
rect 26608 37204 26660 37256
rect 23020 37068 23072 37120
rect 23204 37068 23256 37120
rect 24032 37068 24084 37120
rect 5614 36966 5666 37018
rect 5678 36966 5730 37018
rect 5742 36966 5794 37018
rect 5806 36966 5858 37018
rect 14878 36966 14930 37018
rect 14942 36966 14994 37018
rect 15006 36966 15058 37018
rect 15070 36966 15122 37018
rect 24142 36966 24194 37018
rect 24206 36966 24258 37018
rect 24270 36966 24322 37018
rect 24334 36966 24386 37018
rect 2596 36796 2648 36848
rect 3608 36796 3660 36848
rect 9036 36796 9088 36848
rect 10968 36796 11020 36848
rect 13728 36796 13780 36848
rect 16764 36796 16816 36848
rect 17500 36796 17552 36848
rect 25780 36864 25832 36916
rect 27896 36796 27948 36848
rect 2688 36728 2740 36780
rect 4160 36660 4212 36712
rect 4620 36660 4672 36712
rect 1860 36635 1912 36644
rect 1860 36601 1869 36635
rect 1869 36601 1903 36635
rect 1903 36601 1912 36635
rect 1860 36592 1912 36601
rect 2596 36635 2648 36644
rect 2596 36601 2605 36635
rect 2605 36601 2639 36635
rect 2639 36601 2648 36635
rect 2596 36592 2648 36601
rect 2780 36635 2832 36644
rect 2780 36601 2789 36635
rect 2789 36601 2823 36635
rect 2823 36601 2832 36635
rect 2780 36592 2832 36601
rect 4712 36592 4764 36644
rect 1952 36567 2004 36576
rect 1952 36533 1961 36567
rect 1961 36533 1995 36567
rect 1995 36533 2004 36567
rect 1952 36524 2004 36533
rect 5908 36660 5960 36712
rect 6368 36660 6420 36712
rect 9680 36703 9732 36712
rect 9680 36669 9689 36703
rect 9689 36669 9723 36703
rect 9723 36669 9732 36703
rect 9680 36660 9732 36669
rect 11980 36703 12032 36712
rect 11980 36669 11989 36703
rect 11989 36669 12023 36703
rect 12023 36669 12032 36703
rect 11980 36660 12032 36669
rect 12440 36728 12492 36780
rect 15476 36728 15528 36780
rect 16028 36728 16080 36780
rect 17224 36728 17276 36780
rect 18972 36728 19024 36780
rect 25504 36728 25556 36780
rect 12164 36703 12216 36712
rect 12164 36669 12173 36703
rect 12173 36669 12207 36703
rect 12207 36669 12216 36703
rect 12164 36660 12216 36669
rect 13268 36660 13320 36712
rect 14096 36592 14148 36644
rect 14372 36592 14424 36644
rect 15200 36592 15252 36644
rect 7288 36524 7340 36576
rect 9496 36567 9548 36576
rect 9496 36533 9505 36567
rect 9505 36533 9539 36567
rect 9539 36533 9548 36567
rect 9496 36524 9548 36533
rect 10876 36524 10928 36576
rect 13360 36524 13412 36576
rect 15660 36703 15712 36712
rect 15660 36669 15669 36703
rect 15669 36669 15703 36703
rect 15703 36669 15712 36703
rect 15936 36703 15988 36712
rect 15660 36660 15712 36669
rect 15936 36669 15945 36703
rect 15945 36669 15979 36703
rect 15979 36669 15988 36703
rect 15936 36660 15988 36669
rect 16212 36660 16264 36712
rect 16396 36660 16448 36712
rect 20720 36703 20772 36712
rect 16580 36524 16632 36576
rect 20720 36669 20729 36703
rect 20729 36669 20763 36703
rect 20763 36669 20772 36703
rect 20720 36660 20772 36669
rect 21272 36660 21324 36712
rect 25412 36703 25464 36712
rect 25412 36669 25421 36703
rect 25421 36669 25455 36703
rect 25455 36669 25464 36703
rect 25412 36660 25464 36669
rect 25780 36660 25832 36712
rect 26792 36703 26844 36712
rect 26792 36669 26801 36703
rect 26801 36669 26835 36703
rect 26835 36669 26844 36703
rect 26792 36660 26844 36669
rect 27436 36703 27488 36712
rect 27436 36669 27445 36703
rect 27445 36669 27479 36703
rect 27479 36669 27488 36703
rect 27436 36660 27488 36669
rect 25504 36592 25556 36644
rect 18052 36524 18104 36576
rect 18604 36524 18656 36576
rect 18696 36524 18748 36576
rect 20536 36567 20588 36576
rect 20536 36533 20545 36567
rect 20545 36533 20579 36567
rect 20579 36533 20588 36567
rect 20536 36524 20588 36533
rect 21916 36524 21968 36576
rect 25228 36567 25280 36576
rect 25228 36533 25237 36567
rect 25237 36533 25271 36567
rect 25271 36533 25280 36567
rect 25228 36524 25280 36533
rect 25780 36524 25832 36576
rect 26056 36524 26108 36576
rect 27804 36524 27856 36576
rect 10246 36422 10298 36474
rect 10310 36422 10362 36474
rect 10374 36422 10426 36474
rect 10438 36422 10490 36474
rect 19510 36422 19562 36474
rect 19574 36422 19626 36474
rect 19638 36422 19690 36474
rect 19702 36422 19754 36474
rect 4252 36320 4304 36372
rect 5264 36320 5316 36372
rect 6092 36320 6144 36372
rect 9496 36320 9548 36372
rect 11612 36320 11664 36372
rect 14556 36320 14608 36372
rect 15936 36320 15988 36372
rect 22744 36363 22796 36372
rect 1400 36184 1452 36236
rect 1676 36227 1728 36236
rect 1676 36193 1685 36227
rect 1685 36193 1719 36227
rect 1719 36193 1728 36227
rect 1676 36184 1728 36193
rect 1768 36159 1820 36168
rect 1768 36125 1777 36159
rect 1777 36125 1811 36159
rect 1811 36125 1820 36159
rect 1768 36116 1820 36125
rect 2228 36116 2280 36168
rect 1584 36048 1636 36100
rect 18512 36252 18564 36304
rect 18880 36252 18932 36304
rect 3056 36184 3108 36236
rect 3148 36227 3200 36236
rect 3148 36193 3157 36227
rect 3157 36193 3191 36227
rect 3191 36193 3200 36227
rect 3148 36184 3200 36193
rect 4436 36184 4488 36236
rect 4344 36116 4396 36168
rect 6828 36184 6880 36236
rect 7196 36227 7248 36236
rect 7196 36193 7230 36227
rect 7230 36193 7248 36227
rect 9128 36227 9180 36236
rect 7196 36184 7248 36193
rect 9128 36193 9137 36227
rect 9137 36193 9171 36227
rect 9171 36193 9180 36227
rect 9128 36184 9180 36193
rect 10416 36184 10468 36236
rect 10876 36227 10928 36236
rect 10876 36193 10885 36227
rect 10885 36193 10919 36227
rect 10919 36193 10928 36227
rect 10876 36184 10928 36193
rect 11152 36227 11204 36236
rect 6368 36116 6420 36168
rect 9864 36116 9916 36168
rect 11152 36193 11161 36227
rect 11161 36193 11195 36227
rect 11195 36193 11204 36227
rect 11152 36184 11204 36193
rect 11612 36184 11664 36236
rect 14004 36184 14056 36236
rect 15476 36227 15528 36236
rect 8760 36091 8812 36100
rect 8760 36057 8769 36091
rect 8769 36057 8803 36091
rect 8803 36057 8812 36091
rect 8760 36048 8812 36057
rect 3884 36023 3936 36032
rect 3884 35989 3893 36023
rect 3893 35989 3927 36023
rect 3927 35989 3936 36023
rect 3884 35980 3936 35989
rect 9680 35980 9732 36032
rect 9956 35980 10008 36032
rect 10508 36023 10560 36032
rect 10508 35989 10517 36023
rect 10517 35989 10551 36023
rect 10551 35989 10560 36023
rect 10508 35980 10560 35989
rect 10876 36048 10928 36100
rect 13728 36116 13780 36168
rect 11980 36048 12032 36100
rect 13636 36048 13688 36100
rect 15476 36193 15485 36227
rect 15485 36193 15519 36227
rect 15519 36193 15528 36227
rect 15476 36184 15528 36193
rect 15844 36227 15896 36236
rect 14556 36116 14608 36168
rect 15108 36116 15160 36168
rect 15844 36193 15853 36227
rect 15853 36193 15887 36227
rect 15887 36193 15896 36227
rect 15844 36184 15896 36193
rect 17224 36184 17276 36236
rect 18052 36227 18104 36236
rect 16488 36116 16540 36168
rect 16856 36116 16908 36168
rect 17316 36116 17368 36168
rect 17408 36159 17460 36168
rect 17408 36125 17417 36159
rect 17417 36125 17451 36159
rect 17451 36125 17460 36159
rect 17408 36116 17460 36125
rect 17500 36048 17552 36100
rect 18052 36193 18061 36227
rect 18061 36193 18095 36227
rect 18095 36193 18104 36227
rect 18052 36184 18104 36193
rect 18604 36184 18656 36236
rect 18972 36227 19024 36236
rect 18972 36193 19006 36227
rect 19006 36193 19024 36227
rect 18972 36184 19024 36193
rect 17868 36048 17920 36100
rect 22744 36329 22753 36363
rect 22753 36329 22787 36363
rect 22787 36329 22796 36363
rect 22744 36320 22796 36329
rect 25504 36320 25556 36372
rect 25228 36252 25280 36304
rect 23112 36227 23164 36236
rect 23112 36193 23121 36227
rect 23121 36193 23155 36227
rect 23155 36193 23164 36227
rect 23112 36184 23164 36193
rect 23204 36227 23256 36236
rect 23204 36193 23213 36227
rect 23213 36193 23247 36227
rect 23247 36193 23256 36227
rect 23388 36227 23440 36236
rect 23204 36184 23256 36193
rect 23388 36193 23397 36227
rect 23397 36193 23431 36227
rect 23431 36193 23440 36227
rect 23388 36184 23440 36193
rect 25872 36184 25924 36236
rect 26148 36184 26200 36236
rect 26884 36227 26936 36236
rect 26884 36193 26893 36227
rect 26893 36193 26927 36227
rect 26927 36193 26936 36227
rect 26884 36184 26936 36193
rect 23664 36116 23716 36168
rect 24032 36116 24084 36168
rect 11520 35980 11572 36032
rect 12164 35980 12216 36032
rect 16212 35980 16264 36032
rect 16304 35980 16356 36032
rect 18144 35980 18196 36032
rect 18236 35980 18288 36032
rect 18972 35980 19024 36032
rect 19892 35980 19944 36032
rect 20076 36023 20128 36032
rect 20076 35989 20085 36023
rect 20085 35989 20119 36023
rect 20119 35989 20128 36023
rect 20076 35980 20128 35989
rect 21180 35980 21232 36032
rect 22652 35980 22704 36032
rect 22744 35980 22796 36032
rect 23388 35980 23440 36032
rect 26056 36023 26108 36032
rect 26056 35989 26065 36023
rect 26065 35989 26099 36023
rect 26099 35989 26108 36023
rect 26056 35980 26108 35989
rect 27988 35980 28040 36032
rect 5614 35878 5666 35930
rect 5678 35878 5730 35930
rect 5742 35878 5794 35930
rect 5806 35878 5858 35930
rect 14878 35878 14930 35930
rect 14942 35878 14994 35930
rect 15006 35878 15058 35930
rect 15070 35878 15122 35930
rect 24142 35878 24194 35930
rect 24206 35878 24258 35930
rect 24270 35878 24322 35930
rect 24334 35878 24386 35930
rect 2412 35776 2464 35828
rect 1768 35708 1820 35760
rect 3148 35708 3200 35760
rect 3332 35708 3384 35760
rect 3516 35708 3568 35760
rect 6644 35708 6696 35760
rect 2044 35572 2096 35624
rect 3884 35640 3936 35692
rect 7196 35776 7248 35828
rect 9956 35776 10008 35828
rect 10416 35776 10468 35828
rect 11060 35819 11112 35828
rect 11060 35785 11069 35819
rect 11069 35785 11103 35819
rect 11103 35785 11112 35819
rect 11060 35776 11112 35785
rect 12808 35776 12860 35828
rect 13820 35776 13872 35828
rect 3608 35572 3660 35624
rect 7288 35572 7340 35624
rect 9404 35572 9456 35624
rect 10508 35640 10560 35692
rect 11612 35640 11664 35692
rect 11704 35615 11756 35624
rect 1492 35504 1544 35556
rect 1860 35504 1912 35556
rect 6920 35504 6972 35556
rect 8024 35504 8076 35556
rect 9128 35504 9180 35556
rect 11704 35581 11713 35615
rect 11713 35581 11747 35615
rect 11747 35581 11756 35615
rect 11704 35572 11756 35581
rect 13544 35708 13596 35760
rect 15568 35708 15620 35760
rect 16120 35708 16172 35760
rect 18236 35751 18288 35760
rect 18236 35717 18245 35751
rect 18245 35717 18279 35751
rect 18279 35717 18288 35751
rect 18236 35708 18288 35717
rect 18788 35708 18840 35760
rect 19432 35708 19484 35760
rect 22652 35708 22704 35760
rect 23020 35751 23072 35760
rect 23020 35717 23029 35751
rect 23029 35717 23063 35751
rect 23063 35717 23072 35751
rect 23020 35708 23072 35717
rect 23204 35708 23256 35760
rect 14188 35640 14240 35692
rect 16672 35640 16724 35692
rect 17500 35640 17552 35692
rect 2872 35479 2924 35488
rect 2872 35445 2881 35479
rect 2881 35445 2915 35479
rect 2915 35445 2924 35479
rect 2872 35436 2924 35445
rect 3240 35479 3292 35488
rect 3240 35445 3249 35479
rect 3249 35445 3283 35479
rect 3283 35445 3292 35479
rect 3240 35436 3292 35445
rect 4344 35436 4396 35488
rect 9864 35436 9916 35488
rect 11612 35436 11664 35488
rect 11704 35436 11756 35488
rect 12348 35436 12400 35488
rect 13544 35572 13596 35624
rect 14556 35572 14608 35624
rect 15200 35572 15252 35624
rect 16120 35572 16172 35624
rect 16488 35572 16540 35624
rect 18512 35615 18564 35624
rect 18512 35581 18521 35615
rect 18521 35581 18555 35615
rect 18555 35581 18564 35615
rect 18512 35572 18564 35581
rect 20536 35640 20588 35692
rect 13636 35504 13688 35556
rect 14004 35504 14056 35556
rect 17868 35504 17920 35556
rect 18236 35504 18288 35556
rect 19156 35572 19208 35624
rect 20812 35572 20864 35624
rect 23112 35640 23164 35692
rect 23848 35572 23900 35624
rect 24400 35640 24452 35692
rect 24860 35640 24912 35692
rect 24584 35572 24636 35624
rect 26056 35572 26108 35624
rect 27896 35572 27948 35624
rect 20076 35504 20128 35556
rect 20720 35504 20772 35556
rect 13728 35436 13780 35488
rect 14556 35436 14608 35488
rect 16028 35479 16080 35488
rect 16028 35445 16037 35479
rect 16037 35445 16071 35479
rect 16071 35445 16080 35479
rect 16028 35436 16080 35445
rect 16212 35436 16264 35488
rect 26608 35479 26660 35488
rect 26608 35445 26617 35479
rect 26617 35445 26651 35479
rect 26651 35445 26660 35479
rect 26608 35436 26660 35445
rect 10246 35334 10298 35386
rect 10310 35334 10362 35386
rect 10374 35334 10426 35386
rect 10438 35334 10490 35386
rect 19510 35334 19562 35386
rect 19574 35334 19626 35386
rect 19638 35334 19690 35386
rect 19702 35334 19754 35386
rect 3240 35232 3292 35284
rect 3608 35275 3660 35284
rect 3608 35241 3617 35275
rect 3617 35241 3651 35275
rect 3651 35241 3660 35275
rect 3608 35232 3660 35241
rect 11152 35232 11204 35284
rect 13084 35232 13136 35284
rect 13912 35232 13964 35284
rect 14556 35232 14608 35284
rect 10324 35164 10376 35216
rect 3240 35139 3292 35148
rect 3240 35105 3249 35139
rect 3249 35105 3283 35139
rect 3283 35105 3292 35139
rect 3240 35096 3292 35105
rect 3148 35028 3200 35080
rect 3424 35139 3476 35148
rect 3424 35105 3433 35139
rect 3433 35105 3467 35139
rect 3467 35105 3476 35139
rect 3424 35096 3476 35105
rect 4528 35096 4580 35148
rect 4988 35096 5040 35148
rect 9496 35096 9548 35148
rect 9864 35096 9916 35148
rect 10508 35096 10560 35148
rect 10968 35164 11020 35216
rect 15568 35232 15620 35284
rect 16120 35275 16172 35284
rect 16120 35241 16129 35275
rect 16129 35241 16163 35275
rect 16163 35241 16172 35275
rect 16120 35232 16172 35241
rect 17960 35232 18012 35284
rect 18512 35232 18564 35284
rect 19892 35232 19944 35284
rect 1676 34935 1728 34944
rect 1676 34901 1685 34935
rect 1685 34901 1719 34935
rect 1719 34901 1728 34935
rect 1676 34892 1728 34901
rect 2228 34935 2280 34944
rect 2228 34901 2237 34935
rect 2237 34901 2271 34935
rect 2271 34901 2280 34935
rect 2228 34892 2280 34901
rect 2412 34892 2464 34944
rect 10416 35028 10468 35080
rect 10876 35139 10928 35148
rect 10876 35105 10885 35139
rect 10885 35105 10919 35139
rect 10919 35105 10928 35139
rect 11060 35139 11112 35148
rect 10876 35096 10928 35105
rect 11060 35105 11069 35139
rect 11069 35105 11103 35139
rect 11103 35105 11112 35139
rect 11060 35096 11112 35105
rect 12348 35096 12400 35148
rect 12532 35139 12584 35148
rect 12532 35105 12541 35139
rect 12541 35105 12575 35139
rect 12575 35105 12584 35139
rect 12532 35096 12584 35105
rect 12808 35096 12860 35148
rect 13452 35139 13504 35148
rect 13452 35105 13461 35139
rect 13461 35105 13495 35139
rect 13495 35105 13504 35139
rect 13452 35096 13504 35105
rect 14004 35096 14056 35148
rect 14832 35096 14884 35148
rect 15292 35139 15344 35148
rect 15292 35105 15301 35139
rect 15301 35105 15335 35139
rect 15335 35105 15344 35139
rect 17500 35164 17552 35216
rect 15292 35096 15344 35105
rect 17408 35096 17460 35148
rect 18236 35096 18288 35148
rect 18604 35096 18656 35148
rect 18696 35096 18748 35148
rect 19708 35096 19760 35148
rect 20076 35139 20128 35148
rect 20076 35105 20085 35139
rect 20085 35105 20119 35139
rect 20119 35105 20128 35139
rect 20076 35096 20128 35105
rect 20444 35096 20496 35148
rect 20720 35164 20772 35216
rect 21180 35139 21232 35148
rect 11336 35028 11388 35080
rect 12072 35028 12124 35080
rect 20996 35028 21048 35080
rect 21180 35105 21203 35139
rect 21203 35105 21232 35139
rect 21180 35096 21232 35105
rect 23112 35232 23164 35284
rect 24584 35232 24636 35284
rect 24860 35232 24912 35284
rect 25780 35232 25832 35284
rect 21548 35139 21600 35148
rect 21548 35105 21557 35139
rect 21557 35105 21591 35139
rect 21591 35105 21600 35139
rect 21548 35096 21600 35105
rect 22468 35096 22520 35148
rect 23204 35139 23256 35148
rect 23204 35105 23237 35139
rect 23237 35105 23256 35139
rect 23204 35096 23256 35105
rect 23388 35096 23440 35148
rect 27988 35207 28040 35216
rect 27988 35173 27997 35207
rect 27997 35173 28031 35207
rect 28031 35173 28040 35207
rect 27988 35164 28040 35173
rect 24216 35139 24268 35148
rect 24216 35105 24225 35139
rect 24225 35105 24259 35139
rect 24259 35105 24268 35139
rect 24216 35096 24268 35105
rect 24400 35139 24452 35148
rect 24400 35105 24409 35139
rect 24409 35105 24443 35139
rect 24443 35105 24452 35139
rect 24584 35139 24636 35148
rect 24400 35096 24452 35105
rect 24584 35105 24593 35139
rect 24593 35105 24627 35139
rect 24627 35105 24636 35139
rect 24584 35096 24636 35105
rect 24768 35096 24820 35148
rect 6920 34960 6972 35012
rect 5908 34892 5960 34944
rect 7748 34935 7800 34944
rect 7748 34901 7757 34935
rect 7757 34901 7791 34935
rect 7791 34901 7800 34935
rect 7748 34892 7800 34901
rect 10416 34935 10468 34944
rect 10416 34901 10425 34935
rect 10425 34901 10459 34935
rect 10459 34901 10468 34935
rect 10416 34892 10468 34901
rect 12808 34892 12860 34944
rect 13544 34892 13596 34944
rect 16028 34892 16080 34944
rect 17224 34892 17276 34944
rect 17500 34892 17552 34944
rect 19616 34935 19668 34944
rect 19616 34901 19625 34935
rect 19625 34901 19659 34935
rect 19659 34901 19668 34935
rect 19616 34892 19668 34901
rect 19984 34960 20036 35012
rect 22376 34960 22428 35012
rect 23020 34960 23072 35012
rect 24216 34960 24268 35012
rect 24860 34960 24912 35012
rect 5614 34790 5666 34842
rect 5678 34790 5730 34842
rect 5742 34790 5794 34842
rect 5806 34790 5858 34842
rect 14878 34790 14930 34842
rect 14942 34790 14994 34842
rect 15006 34790 15058 34842
rect 15070 34790 15122 34842
rect 24142 34790 24194 34842
rect 24206 34790 24258 34842
rect 24270 34790 24322 34842
rect 24334 34790 24386 34842
rect 2412 34688 2464 34740
rect 4988 34731 5040 34740
rect 4988 34697 4997 34731
rect 4997 34697 5031 34731
rect 5031 34697 5040 34731
rect 4988 34688 5040 34697
rect 2596 34620 2648 34672
rect 16120 34688 16172 34740
rect 16948 34688 17000 34740
rect 18052 34688 18104 34740
rect 18604 34688 18656 34740
rect 19708 34688 19760 34740
rect 20352 34688 20404 34740
rect 22744 34688 22796 34740
rect 24584 34688 24636 34740
rect 25964 34688 26016 34740
rect 27344 34731 27396 34740
rect 27344 34697 27353 34731
rect 27353 34697 27387 34731
rect 27387 34697 27396 34731
rect 27344 34688 27396 34697
rect 9404 34620 9456 34672
rect 3976 34552 4028 34604
rect 2044 34527 2096 34536
rect 2044 34493 2053 34527
rect 2053 34493 2087 34527
rect 2087 34493 2096 34527
rect 2044 34484 2096 34493
rect 2780 34527 2832 34536
rect 2780 34493 2789 34527
rect 2789 34493 2823 34527
rect 2823 34493 2832 34527
rect 4528 34527 4580 34536
rect 2780 34484 2832 34493
rect 4528 34493 4537 34527
rect 4537 34493 4571 34527
rect 4571 34493 4580 34527
rect 4528 34484 4580 34493
rect 4712 34484 4764 34536
rect 5540 34552 5592 34604
rect 6368 34552 6420 34604
rect 6644 34552 6696 34604
rect 2596 34459 2648 34468
rect 2596 34425 2605 34459
rect 2605 34425 2639 34459
rect 2639 34425 2648 34459
rect 2596 34416 2648 34425
rect 4436 34416 4488 34468
rect 4988 34459 5040 34468
rect 4988 34425 4997 34459
rect 4997 34425 5031 34459
rect 5031 34425 5040 34459
rect 4988 34416 5040 34425
rect 9404 34484 9456 34536
rect 10508 34620 10560 34672
rect 11152 34620 11204 34672
rect 12716 34620 12768 34672
rect 13360 34620 13412 34672
rect 19616 34620 19668 34672
rect 10416 34552 10468 34604
rect 11520 34484 11572 34536
rect 12348 34552 12400 34604
rect 13728 34552 13780 34604
rect 14004 34552 14056 34604
rect 15200 34552 15252 34604
rect 10968 34416 11020 34468
rect 12808 34484 12860 34536
rect 13544 34484 13596 34536
rect 13084 34416 13136 34468
rect 16028 34527 16080 34536
rect 16028 34493 16037 34527
rect 16037 34493 16071 34527
rect 16071 34493 16080 34527
rect 17224 34552 17276 34604
rect 16028 34484 16080 34493
rect 4896 34348 4948 34400
rect 5264 34348 5316 34400
rect 10876 34391 10928 34400
rect 10876 34357 10885 34391
rect 10885 34357 10919 34391
rect 10919 34357 10928 34391
rect 10876 34348 10928 34357
rect 11888 34348 11940 34400
rect 13820 34348 13872 34400
rect 16488 34416 16540 34468
rect 17684 34484 17736 34536
rect 18236 34552 18288 34604
rect 19892 34552 19944 34604
rect 19156 34484 19208 34536
rect 22468 34527 22520 34536
rect 22468 34493 22477 34527
rect 22477 34493 22511 34527
rect 22511 34493 22520 34527
rect 22468 34484 22520 34493
rect 23388 34552 23440 34604
rect 23848 34552 23900 34604
rect 25228 34552 25280 34604
rect 26608 34552 26660 34604
rect 16028 34348 16080 34400
rect 16212 34348 16264 34400
rect 17868 34348 17920 34400
rect 17960 34348 18012 34400
rect 22192 34416 22244 34468
rect 20352 34348 20404 34400
rect 22468 34348 22520 34400
rect 25412 34527 25464 34536
rect 25412 34493 25421 34527
rect 25421 34493 25455 34527
rect 25455 34493 25464 34527
rect 25412 34484 25464 34493
rect 26056 34527 26108 34536
rect 26056 34493 26065 34527
rect 26065 34493 26099 34527
rect 26099 34493 26108 34527
rect 26056 34484 26108 34493
rect 26700 34527 26752 34536
rect 26700 34493 26709 34527
rect 26709 34493 26743 34527
rect 26743 34493 26752 34527
rect 26700 34484 26752 34493
rect 23572 34348 23624 34400
rect 27804 34416 27856 34468
rect 26516 34391 26568 34400
rect 26516 34357 26525 34391
rect 26525 34357 26559 34391
rect 26559 34357 26568 34391
rect 26516 34348 26568 34357
rect 10246 34246 10298 34298
rect 10310 34246 10362 34298
rect 10374 34246 10426 34298
rect 10438 34246 10490 34298
rect 19510 34246 19562 34298
rect 19574 34246 19626 34298
rect 19638 34246 19690 34298
rect 19702 34246 19754 34298
rect 3884 34187 3936 34196
rect 3884 34153 3893 34187
rect 3893 34153 3927 34187
rect 3927 34153 3936 34187
rect 3884 34144 3936 34153
rect 4896 34144 4948 34196
rect 4988 34144 5040 34196
rect 11060 34187 11112 34196
rect 11060 34153 11069 34187
rect 11069 34153 11103 34187
rect 11103 34153 11112 34187
rect 11060 34144 11112 34153
rect 2044 34051 2096 34060
rect 2044 34017 2053 34051
rect 2053 34017 2087 34051
rect 2087 34017 2096 34051
rect 2044 34008 2096 34017
rect 2412 34008 2464 34060
rect 4436 34008 4488 34060
rect 5172 34051 5224 34060
rect 5172 34017 5181 34051
rect 5181 34017 5215 34051
rect 5215 34017 5224 34051
rect 5172 34008 5224 34017
rect 5264 34008 5316 34060
rect 7656 34051 7708 34060
rect 7656 34017 7690 34051
rect 7690 34017 7708 34051
rect 7656 34008 7708 34017
rect 3056 33872 3108 33924
rect 6368 33872 6420 33924
rect 10968 34051 11020 34060
rect 10968 34017 10977 34051
rect 10977 34017 11011 34051
rect 11011 34017 11020 34051
rect 10968 34008 11020 34017
rect 11152 34051 11204 34060
rect 11152 34017 11161 34051
rect 11161 34017 11195 34051
rect 11195 34017 11204 34051
rect 13452 34076 13504 34128
rect 14188 34076 14240 34128
rect 11152 34008 11204 34017
rect 13084 34008 13136 34060
rect 14004 34051 14056 34060
rect 14004 34017 14013 34051
rect 14013 34017 14047 34051
rect 14047 34017 14056 34051
rect 14004 34008 14056 34017
rect 14280 34008 14332 34060
rect 15844 34076 15896 34128
rect 17040 34076 17092 34128
rect 18052 34119 18104 34128
rect 18052 34085 18061 34119
rect 18061 34085 18095 34119
rect 18095 34085 18104 34119
rect 18052 34076 18104 34085
rect 18696 34076 18748 34128
rect 12808 33940 12860 33992
rect 13452 33940 13504 33992
rect 13912 33940 13964 33992
rect 15660 34008 15712 34060
rect 16028 34051 16080 34060
rect 16028 34017 16037 34051
rect 16037 34017 16071 34051
rect 16071 34017 16080 34051
rect 16028 34008 16080 34017
rect 15568 33940 15620 33992
rect 16212 34051 16264 34060
rect 16212 34017 16221 34051
rect 16221 34017 16255 34051
rect 16255 34017 16264 34051
rect 16212 34008 16264 34017
rect 16488 34008 16540 34060
rect 17684 34051 17736 34060
rect 17684 34017 17693 34051
rect 17693 34017 17727 34051
rect 17727 34017 17736 34051
rect 17684 34008 17736 34017
rect 17316 33940 17368 33992
rect 17868 34051 17920 34060
rect 17868 34017 17877 34051
rect 17877 34017 17911 34051
rect 17911 34017 17920 34051
rect 17868 34008 17920 34017
rect 18788 34008 18840 34060
rect 20444 34076 20496 34128
rect 21548 34076 21600 34128
rect 25780 34144 25832 34196
rect 19156 34008 19208 34060
rect 20996 34051 21048 34060
rect 20996 34017 21005 34051
rect 21005 34017 21039 34051
rect 21039 34017 21048 34051
rect 20996 34008 21048 34017
rect 21088 34051 21140 34060
rect 21088 34017 21097 34051
rect 21097 34017 21131 34051
rect 21131 34017 21140 34051
rect 21088 34008 21140 34017
rect 23388 34008 23440 34060
rect 24860 34051 24912 34060
rect 24860 34017 24869 34051
rect 24869 34017 24903 34051
rect 24903 34017 24912 34051
rect 24860 34008 24912 34017
rect 25504 34051 25556 34060
rect 25504 34017 25513 34051
rect 25513 34017 25547 34051
rect 25547 34017 25556 34051
rect 25504 34008 25556 34017
rect 26148 34051 26200 34060
rect 26148 34017 26157 34051
rect 26157 34017 26191 34051
rect 26191 34017 26200 34051
rect 26148 34008 26200 34017
rect 26516 34076 26568 34128
rect 22468 33940 22520 33992
rect 23112 33940 23164 33992
rect 23296 33940 23348 33992
rect 24492 33940 24544 33992
rect 24676 33940 24728 33992
rect 4160 33804 4212 33856
rect 27252 33872 27304 33924
rect 7748 33804 7800 33856
rect 9496 33804 9548 33856
rect 13544 33804 13596 33856
rect 15476 33804 15528 33856
rect 15844 33804 15896 33856
rect 17960 33804 18012 33856
rect 18420 33804 18472 33856
rect 22008 33804 22060 33856
rect 24492 33804 24544 33856
rect 26516 33804 26568 33856
rect 26792 33847 26844 33856
rect 26792 33813 26801 33847
rect 26801 33813 26835 33847
rect 26835 33813 26844 33847
rect 26792 33804 26844 33813
rect 5614 33702 5666 33754
rect 5678 33702 5730 33754
rect 5742 33702 5794 33754
rect 5806 33702 5858 33754
rect 14878 33702 14930 33754
rect 14942 33702 14994 33754
rect 15006 33702 15058 33754
rect 15070 33702 15122 33754
rect 24142 33702 24194 33754
rect 24206 33702 24258 33754
rect 24270 33702 24322 33754
rect 24334 33702 24386 33754
rect 1400 33600 1452 33652
rect 3148 33600 3200 33652
rect 7656 33600 7708 33652
rect 4804 33532 4856 33584
rect 5264 33532 5316 33584
rect 26792 33600 26844 33652
rect 27252 33643 27304 33652
rect 27252 33609 27261 33643
rect 27261 33609 27295 33643
rect 27295 33609 27304 33643
rect 27252 33600 27304 33609
rect 27988 33643 28040 33652
rect 27988 33609 27997 33643
rect 27997 33609 28031 33643
rect 28031 33609 28040 33643
rect 27988 33600 28040 33609
rect 2504 33396 2556 33448
rect 2688 33439 2740 33448
rect 2688 33405 2697 33439
rect 2697 33405 2731 33439
rect 2731 33405 2740 33439
rect 2688 33396 2740 33405
rect 3148 33439 3200 33448
rect 3148 33405 3157 33439
rect 3157 33405 3191 33439
rect 3191 33405 3200 33439
rect 3148 33396 3200 33405
rect 3424 33396 3476 33448
rect 5172 33396 5224 33448
rect 5908 33396 5960 33448
rect 6644 33396 6696 33448
rect 23848 33532 23900 33584
rect 24400 33532 24452 33584
rect 24676 33532 24728 33584
rect 25780 33532 25832 33584
rect 9128 33464 9180 33516
rect 12808 33507 12860 33516
rect 12808 33473 12817 33507
rect 12817 33473 12851 33507
rect 12851 33473 12860 33507
rect 12808 33464 12860 33473
rect 14188 33464 14240 33516
rect 14556 33464 14608 33516
rect 14832 33464 14884 33516
rect 9956 33396 10008 33448
rect 10876 33396 10928 33448
rect 9496 33328 9548 33380
rect 3608 33260 3660 33312
rect 5172 33260 5224 33312
rect 5448 33260 5500 33312
rect 8116 33260 8168 33312
rect 11060 33260 11112 33312
rect 11336 33260 11388 33312
rect 13084 33396 13136 33448
rect 13360 33439 13412 33448
rect 13360 33405 13369 33439
rect 13369 33405 13403 33439
rect 13403 33405 13412 33439
rect 13360 33396 13412 33405
rect 12808 33328 12860 33380
rect 13912 33396 13964 33448
rect 15016 33439 15068 33448
rect 15016 33405 15025 33439
rect 15025 33405 15059 33439
rect 15059 33405 15068 33439
rect 15016 33396 15068 33405
rect 20720 33464 20772 33516
rect 14004 33260 14056 33312
rect 15292 33260 15344 33312
rect 16948 33396 17000 33448
rect 21180 33396 21232 33448
rect 21548 33396 21600 33448
rect 23664 33439 23716 33448
rect 23664 33405 23673 33439
rect 23673 33405 23707 33439
rect 23707 33405 23716 33439
rect 23664 33396 23716 33405
rect 24492 33464 24544 33516
rect 26332 33464 26384 33516
rect 24308 33396 24360 33448
rect 18420 33328 18472 33380
rect 20444 33328 20496 33380
rect 23848 33371 23900 33380
rect 23848 33337 23857 33371
rect 23857 33337 23891 33371
rect 23891 33337 23900 33371
rect 23848 33328 23900 33337
rect 23940 33371 23992 33380
rect 23940 33337 23949 33371
rect 23949 33337 23983 33371
rect 23983 33337 23992 33371
rect 23940 33328 23992 33337
rect 16212 33303 16264 33312
rect 16212 33269 16221 33303
rect 16221 33269 16255 33303
rect 16255 33269 16264 33303
rect 16212 33260 16264 33269
rect 16488 33260 16540 33312
rect 18788 33260 18840 33312
rect 22008 33303 22060 33312
rect 22008 33269 22017 33303
rect 22017 33269 22051 33303
rect 22051 33269 22060 33303
rect 22008 33260 22060 33269
rect 24032 33260 24084 33312
rect 26056 33439 26108 33448
rect 26056 33405 26065 33439
rect 26065 33405 26099 33439
rect 26099 33405 26108 33439
rect 26056 33396 26108 33405
rect 26240 33396 26292 33448
rect 26424 33328 26476 33380
rect 26240 33260 26292 33312
rect 10246 33158 10298 33210
rect 10310 33158 10362 33210
rect 10374 33158 10426 33210
rect 10438 33158 10490 33210
rect 19510 33158 19562 33210
rect 19574 33158 19626 33210
rect 19638 33158 19690 33210
rect 19702 33158 19754 33210
rect 2596 32988 2648 33040
rect 4252 32988 4304 33040
rect 4436 32988 4488 33040
rect 13084 33031 13136 33040
rect 13084 32997 13093 33031
rect 13093 32997 13127 33031
rect 13127 32997 13136 33031
rect 13084 32988 13136 32997
rect 14004 32988 14056 33040
rect 15016 32988 15068 33040
rect 18420 32988 18472 33040
rect 18696 32988 18748 33040
rect 19984 32988 20036 33040
rect 24768 32988 24820 33040
rect 1492 32963 1544 32972
rect 1492 32929 1501 32963
rect 1501 32929 1535 32963
rect 1535 32929 1544 32963
rect 1492 32920 1544 32929
rect 1768 32920 1820 32972
rect 2044 32920 2096 32972
rect 4988 32920 5040 32972
rect 8668 32963 8720 32972
rect 8668 32929 8677 32963
rect 8677 32929 8711 32963
rect 8711 32929 8720 32963
rect 8668 32920 8720 32929
rect 9496 32963 9548 32972
rect 9496 32929 9505 32963
rect 9505 32929 9539 32963
rect 9539 32929 9548 32963
rect 9496 32920 9548 32929
rect 3424 32852 3476 32904
rect 4252 32895 4304 32904
rect 2688 32827 2740 32836
rect 2688 32793 2697 32827
rect 2697 32793 2731 32827
rect 2731 32793 2740 32827
rect 2688 32784 2740 32793
rect 3884 32784 3936 32836
rect 4252 32861 4261 32895
rect 4261 32861 4295 32895
rect 4295 32861 4304 32895
rect 4252 32852 4304 32861
rect 8760 32895 8812 32904
rect 8760 32861 8769 32895
rect 8769 32861 8803 32895
rect 8803 32861 8812 32895
rect 8760 32852 8812 32861
rect 8484 32784 8536 32836
rect 9864 32852 9916 32904
rect 11152 32920 11204 32972
rect 12164 32963 12216 32972
rect 12164 32929 12173 32963
rect 12173 32929 12207 32963
rect 12207 32929 12216 32963
rect 12164 32920 12216 32929
rect 12072 32852 12124 32904
rect 12348 32963 12400 32972
rect 12348 32929 12357 32963
rect 12357 32929 12391 32963
rect 12391 32929 12400 32963
rect 12348 32920 12400 32929
rect 12808 32920 12860 32972
rect 12716 32784 12768 32836
rect 13360 32920 13412 32972
rect 13820 32920 13872 32972
rect 14188 32784 14240 32836
rect 14556 32963 14608 32972
rect 14556 32929 14565 32963
rect 14565 32929 14599 32963
rect 14599 32929 14608 32963
rect 14740 32963 14792 32972
rect 14556 32920 14608 32929
rect 14740 32929 14749 32963
rect 14749 32929 14783 32963
rect 14783 32929 14792 32963
rect 14740 32920 14792 32929
rect 18512 32920 18564 32972
rect 16120 32852 16172 32904
rect 16488 32852 16540 32904
rect 19156 32784 19208 32836
rect 3792 32759 3844 32768
rect 3792 32725 3801 32759
rect 3801 32725 3835 32759
rect 3835 32725 3844 32759
rect 3792 32716 3844 32725
rect 7840 32716 7892 32768
rect 9864 32716 9916 32768
rect 11336 32716 11388 32768
rect 11980 32716 12032 32768
rect 12164 32716 12216 32768
rect 13268 32716 13320 32768
rect 17868 32716 17920 32768
rect 18696 32716 18748 32768
rect 18972 32716 19024 32768
rect 19892 32920 19944 32972
rect 22100 32920 22152 32972
rect 24492 32920 24544 32972
rect 24860 32920 24912 32972
rect 20260 32895 20312 32904
rect 20260 32861 20269 32895
rect 20269 32861 20303 32895
rect 20303 32861 20312 32895
rect 20260 32852 20312 32861
rect 20536 32895 20588 32904
rect 20536 32861 20545 32895
rect 20545 32861 20579 32895
rect 20579 32861 20588 32895
rect 20536 32852 20588 32861
rect 20812 32852 20864 32904
rect 22376 32852 22428 32904
rect 22836 32895 22888 32904
rect 22836 32861 22845 32895
rect 22845 32861 22879 32895
rect 22879 32861 22888 32895
rect 22836 32852 22888 32861
rect 23848 32852 23900 32904
rect 21088 32784 21140 32836
rect 20720 32716 20772 32768
rect 23020 32716 23072 32768
rect 23940 32759 23992 32768
rect 23940 32725 23949 32759
rect 23949 32725 23983 32759
rect 23983 32725 23992 32759
rect 23940 32716 23992 32725
rect 24308 32784 24360 32836
rect 24768 32784 24820 32836
rect 24860 32784 24912 32836
rect 25136 32784 25188 32836
rect 27252 32920 27304 32972
rect 26240 32895 26292 32904
rect 26240 32861 26249 32895
rect 26249 32861 26283 32895
rect 26283 32861 26292 32895
rect 26240 32852 26292 32861
rect 26332 32895 26384 32904
rect 26332 32861 26341 32895
rect 26341 32861 26375 32895
rect 26375 32861 26384 32895
rect 26332 32852 26384 32861
rect 25780 32716 25832 32768
rect 5614 32614 5666 32666
rect 5678 32614 5730 32666
rect 5742 32614 5794 32666
rect 5806 32614 5858 32666
rect 14878 32614 14930 32666
rect 14942 32614 14994 32666
rect 15006 32614 15058 32666
rect 15070 32614 15122 32666
rect 24142 32614 24194 32666
rect 24206 32614 24258 32666
rect 24270 32614 24322 32666
rect 24334 32614 24386 32666
rect 4620 32512 4672 32564
rect 2412 32444 2464 32496
rect 6276 32444 6328 32496
rect 7104 32444 7156 32496
rect 8116 32512 8168 32564
rect 4436 32376 4488 32428
rect 4620 32376 4672 32428
rect 5632 32376 5684 32428
rect 2228 32308 2280 32360
rect 2596 32308 2648 32360
rect 2780 32308 2832 32360
rect 2964 32308 3016 32360
rect 2136 32240 2188 32292
rect 6092 32308 6144 32360
rect 6184 32308 6236 32360
rect 6368 32308 6420 32360
rect 9680 32376 9732 32428
rect 9956 32376 10008 32428
rect 10784 32376 10836 32428
rect 8300 32351 8352 32360
rect 8300 32317 8309 32351
rect 8309 32317 8343 32351
rect 8343 32317 8352 32351
rect 8300 32308 8352 32317
rect 9864 32351 9916 32360
rect 9864 32317 9873 32351
rect 9873 32317 9907 32351
rect 9907 32317 9916 32351
rect 9864 32308 9916 32317
rect 11336 32351 11388 32360
rect 5540 32240 5592 32292
rect 4896 32172 4948 32224
rect 6368 32215 6420 32224
rect 6368 32181 6377 32215
rect 6377 32181 6411 32215
rect 6411 32181 6420 32215
rect 7104 32240 7156 32292
rect 9404 32240 9456 32292
rect 11336 32317 11345 32351
rect 11345 32317 11379 32351
rect 11379 32317 11388 32351
rect 11336 32308 11388 32317
rect 11888 32308 11940 32360
rect 12440 32351 12492 32360
rect 12440 32317 12449 32351
rect 12449 32317 12483 32351
rect 12483 32317 12492 32351
rect 12808 32376 12860 32428
rect 13268 32376 13320 32428
rect 13544 32444 13596 32496
rect 13912 32444 13964 32496
rect 15936 32444 15988 32496
rect 16488 32444 16540 32496
rect 18604 32512 18656 32564
rect 18788 32512 18840 32564
rect 20536 32512 20588 32564
rect 20812 32555 20864 32564
rect 20812 32521 20821 32555
rect 20821 32521 20855 32555
rect 20855 32521 20864 32555
rect 20812 32512 20864 32521
rect 21732 32512 21784 32564
rect 22376 32512 22428 32564
rect 22652 32512 22704 32564
rect 23020 32555 23072 32564
rect 23020 32521 23029 32555
rect 23029 32521 23063 32555
rect 23063 32521 23072 32555
rect 23020 32512 23072 32521
rect 23756 32512 23808 32564
rect 26056 32512 26108 32564
rect 15108 32376 15160 32428
rect 12440 32308 12492 32317
rect 15292 32308 15344 32360
rect 16028 32308 16080 32360
rect 17500 32376 17552 32428
rect 18512 32376 18564 32428
rect 18972 32419 19024 32428
rect 18972 32385 18981 32419
rect 18981 32385 19015 32419
rect 19015 32385 19024 32419
rect 18972 32376 19024 32385
rect 19156 32444 19208 32496
rect 17776 32351 17828 32360
rect 6368 32172 6420 32181
rect 8760 32172 8812 32224
rect 9588 32172 9640 32224
rect 9864 32172 9916 32224
rect 9956 32215 10008 32224
rect 9956 32181 9965 32215
rect 9965 32181 9999 32215
rect 9999 32181 10008 32215
rect 10692 32215 10744 32224
rect 9956 32172 10008 32181
rect 10692 32181 10701 32215
rect 10701 32181 10735 32215
rect 10735 32181 10744 32215
rect 10692 32172 10744 32181
rect 13452 32240 13504 32292
rect 14924 32240 14976 32292
rect 17776 32317 17785 32351
rect 17785 32317 17819 32351
rect 17819 32317 17828 32351
rect 17776 32308 17828 32317
rect 18788 32351 18840 32360
rect 18788 32317 18797 32351
rect 18797 32317 18831 32351
rect 18831 32317 18840 32351
rect 18788 32308 18840 32317
rect 15936 32172 15988 32224
rect 16580 32172 16632 32224
rect 17040 32172 17092 32224
rect 17684 32283 17736 32292
rect 17684 32249 17693 32283
rect 17693 32249 17727 32283
rect 17727 32249 17736 32283
rect 17684 32240 17736 32249
rect 18052 32240 18104 32292
rect 17868 32172 17920 32224
rect 19156 32240 19208 32292
rect 20352 32376 20404 32428
rect 20536 32376 20588 32428
rect 22008 32376 22060 32428
rect 24124 32444 24176 32496
rect 26332 32444 26384 32496
rect 20444 32351 20496 32360
rect 20444 32317 20453 32351
rect 20453 32317 20487 32351
rect 20487 32317 20496 32351
rect 20444 32308 20496 32317
rect 20720 32308 20772 32360
rect 21088 32308 21140 32360
rect 22100 32308 22152 32360
rect 20536 32283 20588 32292
rect 20536 32249 20545 32283
rect 20545 32249 20579 32283
rect 20579 32249 20588 32283
rect 20536 32240 20588 32249
rect 23296 32240 23348 32292
rect 23664 32308 23716 32360
rect 24400 32376 24452 32428
rect 25228 32351 25280 32360
rect 23848 32172 23900 32224
rect 24032 32240 24084 32292
rect 25228 32317 25237 32351
rect 25237 32317 25271 32351
rect 25271 32317 25280 32351
rect 25228 32308 25280 32317
rect 25780 32308 25832 32360
rect 24860 32240 24912 32292
rect 25872 32240 25924 32292
rect 27436 32240 27488 32292
rect 26240 32172 26292 32224
rect 27620 32172 27672 32224
rect 10246 32070 10298 32122
rect 10310 32070 10362 32122
rect 10374 32070 10426 32122
rect 10438 32070 10490 32122
rect 19510 32070 19562 32122
rect 19574 32070 19626 32122
rect 19638 32070 19690 32122
rect 19702 32070 19754 32122
rect 2044 32011 2096 32020
rect 2044 31977 2053 32011
rect 2053 31977 2087 32011
rect 2087 31977 2096 32011
rect 2044 31968 2096 31977
rect 2780 31968 2832 32020
rect 3148 31968 3200 32020
rect 3608 31968 3660 32020
rect 4896 32011 4948 32020
rect 4896 31977 4905 32011
rect 4905 31977 4939 32011
rect 4939 31977 4948 32011
rect 4896 31968 4948 31977
rect 5264 32011 5316 32020
rect 5264 31977 5273 32011
rect 5273 31977 5307 32011
rect 5307 31977 5316 32011
rect 5264 31968 5316 31977
rect 5540 31968 5592 32020
rect 6276 31968 6328 32020
rect 8668 31968 8720 32020
rect 12440 31968 12492 32020
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 2596 31900 2648 31952
rect 3792 31900 3844 31952
rect 2504 31875 2556 31884
rect 2504 31841 2513 31875
rect 2513 31841 2547 31875
rect 2547 31841 2556 31875
rect 2504 31832 2556 31841
rect 3056 31832 3108 31884
rect 6736 31832 6788 31884
rect 5448 31764 5500 31816
rect 5632 31764 5684 31816
rect 7288 31900 7340 31952
rect 7840 31943 7892 31952
rect 7840 31909 7849 31943
rect 7849 31909 7883 31943
rect 7883 31909 7892 31943
rect 7840 31900 7892 31909
rect 8116 31900 8168 31952
rect 7012 31832 7064 31884
rect 8300 31832 8352 31884
rect 8760 31875 8812 31884
rect 8760 31841 8769 31875
rect 8769 31841 8803 31875
rect 8803 31841 8812 31875
rect 8760 31832 8812 31841
rect 10048 31900 10100 31952
rect 10324 31900 10376 31952
rect 13268 31968 13320 32020
rect 14556 32011 14608 32020
rect 14556 31977 14565 32011
rect 14565 31977 14599 32011
rect 14599 31977 14608 32011
rect 14556 31968 14608 31977
rect 18144 31968 18196 32020
rect 18512 31968 18564 32020
rect 21088 31968 21140 32020
rect 21180 31968 21232 32020
rect 13728 31900 13780 31952
rect 14924 31900 14976 31952
rect 9220 31832 9272 31884
rect 9772 31832 9824 31884
rect 11152 31832 11204 31884
rect 13544 31875 13596 31884
rect 13544 31841 13553 31875
rect 13553 31841 13587 31875
rect 13587 31841 13596 31875
rect 13544 31832 13596 31841
rect 13820 31832 13872 31884
rect 15292 31900 15344 31952
rect 15476 31900 15528 31952
rect 11336 31764 11388 31816
rect 12256 31764 12308 31816
rect 8576 31696 8628 31748
rect 12808 31696 12860 31748
rect 4988 31628 5040 31680
rect 7104 31628 7156 31680
rect 8300 31671 8352 31680
rect 8300 31637 8309 31671
rect 8309 31637 8343 31671
rect 8343 31637 8352 31671
rect 8300 31628 8352 31637
rect 10324 31628 10376 31680
rect 11152 31628 11204 31680
rect 12716 31628 12768 31680
rect 13912 31764 13964 31816
rect 15108 31875 15160 31884
rect 15108 31841 15117 31875
rect 15117 31841 15151 31875
rect 15151 31841 15160 31875
rect 15108 31832 15160 31841
rect 14556 31628 14608 31680
rect 15936 31875 15988 31884
rect 15936 31841 15945 31875
rect 15945 31841 15979 31875
rect 15979 31841 15988 31875
rect 15936 31832 15988 31841
rect 16304 31900 16356 31952
rect 18788 31900 18840 31952
rect 22560 31900 22612 31952
rect 16488 31832 16540 31884
rect 17408 31832 17460 31884
rect 16580 31764 16632 31816
rect 17040 31764 17092 31816
rect 17500 31696 17552 31748
rect 17776 31832 17828 31884
rect 18512 31875 18564 31884
rect 18512 31841 18521 31875
rect 18521 31841 18555 31875
rect 18555 31841 18564 31875
rect 18512 31832 18564 31841
rect 18604 31807 18656 31816
rect 18604 31773 18613 31807
rect 18613 31773 18647 31807
rect 18647 31773 18656 31807
rect 18604 31764 18656 31773
rect 19156 31832 19208 31884
rect 20444 31832 20496 31884
rect 21180 31832 21232 31884
rect 21364 31875 21416 31884
rect 21364 31841 21373 31875
rect 21373 31841 21407 31875
rect 21407 31841 21416 31875
rect 21364 31832 21416 31841
rect 22192 31832 22244 31884
rect 22744 31832 22796 31884
rect 23112 31968 23164 32020
rect 24032 31968 24084 32020
rect 24768 31968 24820 32020
rect 26608 31968 26660 32020
rect 15568 31671 15620 31680
rect 15568 31637 15577 31671
rect 15577 31637 15611 31671
rect 15611 31637 15620 31671
rect 15568 31628 15620 31637
rect 17868 31671 17920 31680
rect 17868 31637 17877 31671
rect 17877 31637 17911 31671
rect 17911 31637 17920 31671
rect 17868 31628 17920 31637
rect 18604 31628 18656 31680
rect 18972 31764 19024 31816
rect 21088 31764 21140 31816
rect 23572 31832 23624 31884
rect 23756 31832 23808 31884
rect 23296 31764 23348 31816
rect 24400 31832 24452 31884
rect 25228 31832 25280 31884
rect 26148 31875 26200 31884
rect 26148 31841 26157 31875
rect 26157 31841 26191 31875
rect 26191 31841 26200 31875
rect 26148 31832 26200 31841
rect 26516 31832 26568 31884
rect 22468 31696 22520 31748
rect 23940 31696 23992 31748
rect 18880 31628 18932 31680
rect 21272 31628 21324 31680
rect 21640 31671 21692 31680
rect 21640 31637 21649 31671
rect 21649 31637 21683 31671
rect 21683 31637 21692 31671
rect 21640 31628 21692 31637
rect 21732 31628 21784 31680
rect 22100 31628 22152 31680
rect 22652 31628 22704 31680
rect 22928 31628 22980 31680
rect 23388 31628 23440 31680
rect 23848 31628 23900 31680
rect 27988 31671 28040 31680
rect 27988 31637 27997 31671
rect 27997 31637 28031 31671
rect 28031 31637 28040 31671
rect 27988 31628 28040 31637
rect 5614 31526 5666 31578
rect 5678 31526 5730 31578
rect 5742 31526 5794 31578
rect 5806 31526 5858 31578
rect 14878 31526 14930 31578
rect 14942 31526 14994 31578
rect 15006 31526 15058 31578
rect 15070 31526 15122 31578
rect 24142 31526 24194 31578
rect 24206 31526 24258 31578
rect 24270 31526 24322 31578
rect 24334 31526 24386 31578
rect 1400 31424 1452 31476
rect 4252 31424 4304 31476
rect 6368 31467 6420 31476
rect 6368 31433 6377 31467
rect 6377 31433 6411 31467
rect 6411 31433 6420 31467
rect 6368 31424 6420 31433
rect 2504 31399 2556 31408
rect 2504 31365 2513 31399
rect 2513 31365 2547 31399
rect 2547 31365 2556 31399
rect 2504 31356 2556 31365
rect 4988 31356 5040 31408
rect 8576 31424 8628 31476
rect 8668 31424 8720 31476
rect 7288 31399 7340 31408
rect 7288 31365 7297 31399
rect 7297 31365 7331 31399
rect 7331 31365 7340 31399
rect 7288 31356 7340 31365
rect 10876 31356 10928 31408
rect 12440 31356 12492 31408
rect 14556 31356 14608 31408
rect 16580 31356 16632 31408
rect 2688 31220 2740 31272
rect 7196 31288 7248 31340
rect 4160 31220 4212 31272
rect 4528 31220 4580 31272
rect 5908 31220 5960 31272
rect 6368 31220 6420 31272
rect 10692 31288 10744 31340
rect 11520 31220 11572 31272
rect 11888 31263 11940 31272
rect 11888 31229 11897 31263
rect 11897 31229 11931 31263
rect 11931 31229 11940 31263
rect 11888 31220 11940 31229
rect 14188 31288 14240 31340
rect 2136 31195 2188 31204
rect 2136 31161 2145 31195
rect 2145 31161 2179 31195
rect 2179 31161 2188 31195
rect 2136 31152 2188 31161
rect 7012 31152 7064 31204
rect 7288 31152 7340 31204
rect 11980 31195 12032 31204
rect 1400 31084 1452 31136
rect 3240 31127 3292 31136
rect 3240 31093 3249 31127
rect 3249 31093 3283 31127
rect 3283 31093 3292 31127
rect 3240 31084 3292 31093
rect 3332 31084 3384 31136
rect 7932 31127 7984 31136
rect 7932 31093 7941 31127
rect 7941 31093 7975 31127
rect 7975 31093 7984 31127
rect 7932 31084 7984 31093
rect 11980 31161 11989 31195
rect 11989 31161 12023 31195
rect 12023 31161 12032 31195
rect 11980 31152 12032 31161
rect 12716 31220 12768 31272
rect 13176 31220 13228 31272
rect 15476 31220 15528 31272
rect 16028 31220 16080 31272
rect 17408 31220 17460 31272
rect 18512 31288 18564 31340
rect 21732 31356 21784 31408
rect 22836 31424 22888 31476
rect 24124 31356 24176 31408
rect 24768 31356 24820 31408
rect 18328 31220 18380 31272
rect 18972 31220 19024 31272
rect 20260 31263 20312 31272
rect 20260 31229 20269 31263
rect 20269 31229 20303 31263
rect 20303 31229 20312 31263
rect 20260 31220 20312 31229
rect 20536 31220 20588 31272
rect 21640 31288 21692 31340
rect 22468 31263 22520 31272
rect 22468 31229 22477 31263
rect 22477 31229 22511 31263
rect 22511 31229 22520 31263
rect 22468 31220 22520 31229
rect 15844 31152 15896 31204
rect 21916 31152 21968 31204
rect 22652 31263 22704 31272
rect 22652 31229 22661 31263
rect 22661 31229 22695 31263
rect 22695 31229 22704 31263
rect 22652 31220 22704 31229
rect 23940 31263 23992 31272
rect 23940 31229 23949 31263
rect 23949 31229 23983 31263
rect 23983 31229 23992 31263
rect 23940 31220 23992 31229
rect 24124 31263 24176 31272
rect 24124 31229 24133 31263
rect 24133 31229 24167 31263
rect 24167 31229 24176 31263
rect 24124 31220 24176 31229
rect 25228 31263 25280 31272
rect 10876 31084 10928 31136
rect 12164 31084 12216 31136
rect 12440 31084 12492 31136
rect 12716 31084 12768 31136
rect 13820 31084 13872 31136
rect 14188 31084 14240 31136
rect 18512 31084 18564 31136
rect 18972 31127 19024 31136
rect 18972 31093 18981 31127
rect 18981 31093 19015 31127
rect 19015 31093 19024 31127
rect 18972 31084 19024 31093
rect 21364 31084 21416 31136
rect 24032 31084 24084 31136
rect 25228 31229 25237 31263
rect 25237 31229 25271 31263
rect 25271 31229 25280 31263
rect 25228 31220 25280 31229
rect 25780 31220 25832 31272
rect 26332 31152 26384 31204
rect 25872 31084 25924 31136
rect 10246 30982 10298 31034
rect 10310 30982 10362 31034
rect 10374 30982 10426 31034
rect 10438 30982 10490 31034
rect 19510 30982 19562 31034
rect 19574 30982 19626 31034
rect 19638 30982 19690 31034
rect 19702 30982 19754 31034
rect 3792 30880 3844 30932
rect 27988 30880 28040 30932
rect 1860 30787 1912 30796
rect 1860 30753 1869 30787
rect 1869 30753 1903 30787
rect 1903 30753 1912 30787
rect 1860 30744 1912 30753
rect 2596 30787 2648 30796
rect 2596 30753 2605 30787
rect 2605 30753 2639 30787
rect 2639 30753 2648 30787
rect 2596 30744 2648 30753
rect 3516 30744 3568 30796
rect 8668 30812 8720 30864
rect 10048 30812 10100 30864
rect 11060 30812 11112 30864
rect 11336 30812 11388 30864
rect 7564 30787 7616 30796
rect 7564 30753 7573 30787
rect 7573 30753 7607 30787
rect 7607 30753 7616 30787
rect 7564 30744 7616 30753
rect 7932 30787 7984 30796
rect 7932 30753 7941 30787
rect 7941 30753 7975 30787
rect 7975 30753 7984 30787
rect 7932 30744 7984 30753
rect 1952 30676 2004 30728
rect 3240 30676 3292 30728
rect 4068 30676 4120 30728
rect 7472 30676 7524 30728
rect 8300 30744 8352 30796
rect 12256 30744 12308 30796
rect 12440 30787 12492 30796
rect 12440 30753 12449 30787
rect 12449 30753 12483 30787
rect 12483 30753 12492 30787
rect 12440 30744 12492 30753
rect 13912 30787 13964 30796
rect 12716 30676 12768 30728
rect 2780 30651 2832 30660
rect 2780 30617 2789 30651
rect 2789 30617 2823 30651
rect 2823 30617 2832 30651
rect 2780 30608 2832 30617
rect 8944 30608 8996 30660
rect 9956 30608 10008 30660
rect 10692 30608 10744 30660
rect 11336 30608 11388 30660
rect 11520 30608 11572 30660
rect 1952 30583 2004 30592
rect 1952 30549 1961 30583
rect 1961 30549 1995 30583
rect 1995 30549 2004 30583
rect 1952 30540 2004 30549
rect 3884 30540 3936 30592
rect 11888 30540 11940 30592
rect 12440 30583 12492 30592
rect 12440 30549 12449 30583
rect 12449 30549 12483 30583
rect 12483 30549 12492 30583
rect 13912 30753 13921 30787
rect 13921 30753 13955 30787
rect 13955 30753 13964 30787
rect 13912 30744 13964 30753
rect 14280 30787 14332 30796
rect 14280 30753 14289 30787
rect 14289 30753 14323 30787
rect 14323 30753 14332 30787
rect 14280 30744 14332 30753
rect 15108 30744 15160 30796
rect 16212 30812 16264 30864
rect 18512 30855 18564 30864
rect 18512 30821 18521 30855
rect 18521 30821 18555 30855
rect 18555 30821 18564 30855
rect 18512 30812 18564 30821
rect 20260 30812 20312 30864
rect 15476 30744 15528 30796
rect 16120 30787 16172 30796
rect 16120 30753 16129 30787
rect 16129 30753 16163 30787
rect 16163 30753 16172 30787
rect 16120 30744 16172 30753
rect 17408 30744 17460 30796
rect 17868 30744 17920 30796
rect 19432 30787 19484 30796
rect 19432 30753 19441 30787
rect 19441 30753 19475 30787
rect 19475 30753 19484 30787
rect 19432 30744 19484 30753
rect 16672 30676 16724 30728
rect 17408 30608 17460 30660
rect 12440 30540 12492 30549
rect 13820 30540 13872 30592
rect 16028 30540 16080 30592
rect 16580 30540 16632 30592
rect 19708 30744 19760 30796
rect 20444 30744 20496 30796
rect 21364 30812 21416 30864
rect 20996 30787 21048 30796
rect 20996 30753 21005 30787
rect 21005 30753 21039 30787
rect 21039 30753 21048 30787
rect 20996 30744 21048 30753
rect 21180 30744 21232 30796
rect 23020 30744 23072 30796
rect 17776 30608 17828 30660
rect 20076 30676 20128 30728
rect 21916 30676 21968 30728
rect 20812 30608 20864 30660
rect 20904 30608 20956 30660
rect 22652 30608 22704 30660
rect 23388 30744 23440 30796
rect 26608 30812 26660 30864
rect 25412 30744 25464 30796
rect 25780 30744 25832 30796
rect 27528 30744 27580 30796
rect 25228 30676 25280 30728
rect 18696 30540 18748 30592
rect 19432 30540 19484 30592
rect 20536 30540 20588 30592
rect 20996 30540 21048 30592
rect 21272 30540 21324 30592
rect 25228 30540 25280 30592
rect 27988 30583 28040 30592
rect 27988 30549 27997 30583
rect 27997 30549 28031 30583
rect 28031 30549 28040 30583
rect 27988 30540 28040 30549
rect 5614 30438 5666 30490
rect 5678 30438 5730 30490
rect 5742 30438 5794 30490
rect 5806 30438 5858 30490
rect 14878 30438 14930 30490
rect 14942 30438 14994 30490
rect 15006 30438 15058 30490
rect 15070 30438 15122 30490
rect 24142 30438 24194 30490
rect 24206 30438 24258 30490
rect 24270 30438 24322 30490
rect 24334 30438 24386 30490
rect 4988 30336 5040 30388
rect 5264 30336 5316 30388
rect 6644 30336 6696 30388
rect 6920 30336 6972 30388
rect 12348 30336 12400 30388
rect 13728 30336 13780 30388
rect 17408 30336 17460 30388
rect 1860 30268 1912 30320
rect 6092 30311 6144 30320
rect 2872 30200 2924 30252
rect 6092 30277 6101 30311
rect 6101 30277 6135 30311
rect 6135 30277 6144 30311
rect 6092 30268 6144 30277
rect 6736 30311 6788 30320
rect 6736 30277 6745 30311
rect 6745 30277 6779 30311
rect 6779 30277 6788 30311
rect 6736 30268 6788 30277
rect 1860 30107 1912 30116
rect 1860 30073 1869 30107
rect 1869 30073 1903 30107
rect 1903 30073 1912 30107
rect 1860 30064 1912 30073
rect 4344 30132 4396 30184
rect 4804 30175 4856 30184
rect 4804 30141 4813 30175
rect 4813 30141 4847 30175
rect 4847 30141 4856 30175
rect 4804 30132 4856 30141
rect 4896 30175 4948 30184
rect 4896 30141 4905 30175
rect 4905 30141 4939 30175
rect 4939 30141 4948 30175
rect 4896 30132 4948 30141
rect 4068 30064 4120 30116
rect 4712 30064 4764 30116
rect 5908 30132 5960 30184
rect 6092 30132 6144 30184
rect 6644 30175 6696 30184
rect 6644 30141 6653 30175
rect 6653 30141 6687 30175
rect 6687 30141 6696 30175
rect 6644 30132 6696 30141
rect 9588 30175 9640 30184
rect 9588 30141 9597 30175
rect 9597 30141 9631 30175
rect 9631 30141 9640 30175
rect 9588 30132 9640 30141
rect 11980 30175 12032 30184
rect 11980 30141 11989 30175
rect 11989 30141 12023 30175
rect 12023 30141 12032 30175
rect 11980 30132 12032 30141
rect 12440 30132 12492 30184
rect 12808 30175 12860 30184
rect 12808 30141 12817 30175
rect 12817 30141 12851 30175
rect 12851 30141 12860 30175
rect 12808 30132 12860 30141
rect 6184 30064 6236 30116
rect 2412 29996 2464 30048
rect 3332 30039 3384 30048
rect 3332 30005 3341 30039
rect 3341 30005 3375 30039
rect 3375 30005 3384 30039
rect 3332 29996 3384 30005
rect 3976 29996 4028 30048
rect 9680 30039 9732 30048
rect 9680 30005 9689 30039
rect 9689 30005 9723 30039
rect 9723 30005 9732 30039
rect 9680 29996 9732 30005
rect 16580 30311 16632 30320
rect 13728 30200 13780 30252
rect 16580 30277 16589 30311
rect 16589 30277 16623 30311
rect 16623 30277 16632 30311
rect 16580 30268 16632 30277
rect 15108 30200 15160 30252
rect 16948 30200 17000 30252
rect 19708 30268 19760 30320
rect 20812 30268 20864 30320
rect 13452 30175 13504 30184
rect 13452 30141 13461 30175
rect 13461 30141 13495 30175
rect 13495 30141 13504 30175
rect 13452 30132 13504 30141
rect 13820 30132 13872 30184
rect 14556 30132 14608 30184
rect 13912 30064 13964 30116
rect 16120 30132 16172 30184
rect 20444 30200 20496 30252
rect 22100 30336 22152 30388
rect 23020 30336 23072 30388
rect 24032 30379 24084 30388
rect 23296 30268 23348 30320
rect 24032 30345 24041 30379
rect 24041 30345 24075 30379
rect 24075 30345 24084 30379
rect 24032 30336 24084 30345
rect 15844 30107 15896 30116
rect 15844 30073 15853 30107
rect 15853 30073 15887 30107
rect 15887 30073 15896 30107
rect 15844 30064 15896 30073
rect 16672 30064 16724 30116
rect 18788 30175 18840 30184
rect 18788 30141 18797 30175
rect 18797 30141 18831 30175
rect 18831 30141 18840 30175
rect 18788 30132 18840 30141
rect 18972 30064 19024 30116
rect 20352 30107 20404 30116
rect 20352 30073 20361 30107
rect 20361 30073 20395 30107
rect 20395 30073 20404 30107
rect 20352 30064 20404 30073
rect 20812 30175 20864 30184
rect 20812 30141 20821 30175
rect 20821 30141 20855 30175
rect 20855 30141 20864 30175
rect 20996 30175 21048 30184
rect 20812 30132 20864 30141
rect 20996 30141 21005 30175
rect 21005 30141 21039 30175
rect 21039 30141 21048 30175
rect 20996 30132 21048 30141
rect 21732 30175 21784 30184
rect 21732 30141 21741 30175
rect 21741 30141 21775 30175
rect 21775 30141 21784 30175
rect 21732 30132 21784 30141
rect 22928 30132 22980 30184
rect 25228 30268 25280 30320
rect 25688 30175 25740 30184
rect 17040 29996 17092 30048
rect 23204 30064 23256 30116
rect 25688 30141 25697 30175
rect 25697 30141 25731 30175
rect 25731 30141 25740 30175
rect 25688 30132 25740 30141
rect 26148 30132 26200 30184
rect 21456 29996 21508 30048
rect 22468 29996 22520 30048
rect 25596 29996 25648 30048
rect 27068 29996 27120 30048
rect 10246 29894 10298 29946
rect 10310 29894 10362 29946
rect 10374 29894 10426 29946
rect 10438 29894 10490 29946
rect 19510 29894 19562 29946
rect 19574 29894 19626 29946
rect 19638 29894 19690 29946
rect 19702 29894 19754 29946
rect 2596 29792 2648 29844
rect 13820 29792 13872 29844
rect 13912 29792 13964 29844
rect 14188 29792 14240 29844
rect 3332 29724 3384 29776
rect 2780 29656 2832 29708
rect 2228 29631 2280 29640
rect 2228 29597 2237 29631
rect 2237 29597 2271 29631
rect 2271 29597 2280 29631
rect 2228 29588 2280 29597
rect 2320 29631 2372 29640
rect 2320 29597 2329 29631
rect 2329 29597 2363 29631
rect 2363 29597 2372 29631
rect 5448 29656 5500 29708
rect 5908 29656 5960 29708
rect 2320 29588 2372 29597
rect 1400 29520 1452 29572
rect 3056 29520 3108 29572
rect 4988 29588 5040 29640
rect 5724 29631 5776 29640
rect 5724 29597 5733 29631
rect 5733 29597 5767 29631
rect 5767 29597 5776 29631
rect 5724 29588 5776 29597
rect 5540 29520 5592 29572
rect 1676 29452 1728 29504
rect 4528 29495 4580 29504
rect 4528 29461 4537 29495
rect 4537 29461 4571 29495
rect 4571 29461 4580 29495
rect 4528 29452 4580 29461
rect 9128 29724 9180 29776
rect 6644 29656 6696 29708
rect 9956 29724 10008 29776
rect 12164 29724 12216 29776
rect 7748 29588 7800 29640
rect 12716 29656 12768 29708
rect 14280 29699 14332 29708
rect 6276 29520 6328 29572
rect 9588 29563 9640 29572
rect 9588 29529 9597 29563
rect 9597 29529 9631 29563
rect 9631 29529 9640 29563
rect 9588 29520 9640 29529
rect 9956 29520 10008 29572
rect 14280 29665 14289 29699
rect 14289 29665 14323 29699
rect 14323 29665 14332 29699
rect 14280 29656 14332 29665
rect 14556 29656 14608 29708
rect 15292 29792 15344 29844
rect 15384 29792 15436 29844
rect 20076 29792 20128 29844
rect 20812 29792 20864 29844
rect 26332 29792 26384 29844
rect 15568 29724 15620 29776
rect 27068 29724 27120 29776
rect 27988 29767 28040 29776
rect 27988 29733 27997 29767
rect 27997 29733 28031 29767
rect 28031 29733 28040 29767
rect 27988 29724 28040 29733
rect 16120 29699 16172 29708
rect 6828 29452 6880 29504
rect 8392 29452 8444 29504
rect 16120 29665 16129 29699
rect 16129 29665 16163 29699
rect 16163 29665 16172 29699
rect 16120 29656 16172 29665
rect 16948 29656 17000 29708
rect 17224 29656 17276 29708
rect 26056 29656 26108 29708
rect 26700 29699 26752 29708
rect 26700 29665 26709 29699
rect 26709 29665 26743 29699
rect 26743 29665 26752 29699
rect 26700 29656 26752 29665
rect 17040 29588 17092 29640
rect 15292 29520 15344 29572
rect 15568 29520 15620 29572
rect 26240 29520 26292 29572
rect 26884 29563 26936 29572
rect 26884 29529 26893 29563
rect 26893 29529 26927 29563
rect 26927 29529 26936 29563
rect 26884 29520 26936 29529
rect 12440 29452 12492 29504
rect 13452 29452 13504 29504
rect 15476 29452 15528 29504
rect 20444 29452 20496 29504
rect 5614 29350 5666 29402
rect 5678 29350 5730 29402
rect 5742 29350 5794 29402
rect 5806 29350 5858 29402
rect 14878 29350 14930 29402
rect 14942 29350 14994 29402
rect 15006 29350 15058 29402
rect 15070 29350 15122 29402
rect 24142 29350 24194 29402
rect 24206 29350 24258 29402
rect 24270 29350 24322 29402
rect 24334 29350 24386 29402
rect 25596 29248 25648 29300
rect 27436 29248 27488 29300
rect 4896 29180 4948 29232
rect 6828 29223 6880 29232
rect 6828 29189 6837 29223
rect 6837 29189 6871 29223
rect 6871 29189 6880 29223
rect 6828 29180 6880 29189
rect 7564 29180 7616 29232
rect 1400 29155 1452 29164
rect 1400 29121 1409 29155
rect 1409 29121 1443 29155
rect 1443 29121 1452 29155
rect 1400 29112 1452 29121
rect 2688 29112 2740 29164
rect 4988 29112 5040 29164
rect 5448 29155 5500 29164
rect 5448 29121 5457 29155
rect 5457 29121 5491 29155
rect 5491 29121 5500 29155
rect 5448 29112 5500 29121
rect 10508 29180 10560 29232
rect 11704 29180 11756 29232
rect 22376 29180 22428 29232
rect 22928 29180 22980 29232
rect 26516 29180 26568 29232
rect 9128 29112 9180 29164
rect 9404 29112 9456 29164
rect 11060 29112 11112 29164
rect 1676 29087 1728 29096
rect 1676 29053 1710 29087
rect 1710 29053 1728 29087
rect 1676 29044 1728 29053
rect 2780 29044 2832 29096
rect 4344 29044 4396 29096
rect 5356 29044 5408 29096
rect 7748 29044 7800 29096
rect 7932 29087 7984 29096
rect 7932 29053 7941 29087
rect 7941 29053 7975 29087
rect 7975 29053 7984 29087
rect 7932 29044 7984 29053
rect 8392 29044 8444 29096
rect 4252 28976 4304 29028
rect 4712 29019 4764 29028
rect 4712 28985 4721 29019
rect 4721 28985 4755 29019
rect 4755 28985 4764 29019
rect 4712 28976 4764 28985
rect 5816 28976 5868 29028
rect 10784 29087 10836 29096
rect 10784 29053 10793 29087
rect 10793 29053 10827 29087
rect 10827 29053 10836 29087
rect 10784 29044 10836 29053
rect 12256 29112 12308 29164
rect 25688 29155 25740 29164
rect 11704 29044 11756 29096
rect 11888 29087 11940 29096
rect 11888 29053 11897 29087
rect 11897 29053 11931 29087
rect 11931 29053 11940 29087
rect 11888 29044 11940 29053
rect 13452 29044 13504 29096
rect 14556 29044 14608 29096
rect 25688 29121 25697 29155
rect 25697 29121 25731 29155
rect 25731 29121 25740 29155
rect 25688 29112 25740 29121
rect 15844 29044 15896 29096
rect 26516 29044 26568 29096
rect 27620 29087 27672 29096
rect 27620 29053 27629 29087
rect 27629 29053 27663 29087
rect 27663 29053 27672 29087
rect 27620 29044 27672 29053
rect 27712 29044 27764 29096
rect 28264 29044 28316 29096
rect 3976 28908 4028 28960
rect 10232 28976 10284 29028
rect 9864 28951 9916 28960
rect 9864 28917 9873 28951
rect 9873 28917 9907 28951
rect 9907 28917 9916 28951
rect 9864 28908 9916 28917
rect 11336 28908 11388 28960
rect 14280 28908 14332 28960
rect 25596 28976 25648 29028
rect 26424 29019 26476 29028
rect 26424 28985 26433 29019
rect 26433 28985 26467 29019
rect 26467 28985 26476 29019
rect 26424 28976 26476 28985
rect 27160 29019 27212 29028
rect 27160 28985 27169 29019
rect 27169 28985 27203 29019
rect 27203 28985 27212 29019
rect 27160 28976 27212 28985
rect 16120 28908 16172 28960
rect 20168 28908 20220 28960
rect 24860 28908 24912 28960
rect 25136 28908 25188 28960
rect 26700 28908 26752 28960
rect 27896 28908 27948 28960
rect 10246 28806 10298 28858
rect 10310 28806 10362 28858
rect 10374 28806 10426 28858
rect 10438 28806 10490 28858
rect 19510 28806 19562 28858
rect 19574 28806 19626 28858
rect 19638 28806 19690 28858
rect 19702 28806 19754 28858
rect 2228 28704 2280 28756
rect 1860 28679 1912 28688
rect 1860 28645 1869 28679
rect 1869 28645 1903 28679
rect 1903 28645 1912 28679
rect 1860 28636 1912 28645
rect 4344 28704 4396 28756
rect 4804 28704 4856 28756
rect 5816 28747 5868 28756
rect 5816 28713 5825 28747
rect 5825 28713 5859 28747
rect 5859 28713 5868 28747
rect 5816 28704 5868 28713
rect 7932 28747 7984 28756
rect 2136 28568 2188 28620
rect 4528 28636 4580 28688
rect 5264 28636 5316 28688
rect 4988 28611 5040 28620
rect 4988 28577 4997 28611
rect 4997 28577 5031 28611
rect 5031 28577 5040 28611
rect 4988 28568 5040 28577
rect 7104 28611 7156 28620
rect 5172 28500 5224 28552
rect 5448 28500 5500 28552
rect 6184 28500 6236 28552
rect 7104 28577 7113 28611
rect 7113 28577 7147 28611
rect 7147 28577 7156 28611
rect 7104 28568 7156 28577
rect 7564 28636 7616 28688
rect 7932 28713 7941 28747
rect 7941 28713 7975 28747
rect 7975 28713 7984 28747
rect 7932 28704 7984 28713
rect 9680 28704 9732 28756
rect 9864 28704 9916 28756
rect 11060 28704 11112 28756
rect 10692 28679 10744 28688
rect 7472 28568 7524 28620
rect 8300 28611 8352 28620
rect 8300 28577 8309 28611
rect 8309 28577 8343 28611
rect 8343 28577 8352 28611
rect 8300 28568 8352 28577
rect 10692 28645 10701 28679
rect 10701 28645 10735 28679
rect 10735 28645 10744 28679
rect 10692 28636 10744 28645
rect 21272 28704 21324 28756
rect 25136 28704 25188 28756
rect 26700 28704 26752 28756
rect 12808 28636 12860 28688
rect 14096 28636 14148 28688
rect 11336 28568 11388 28620
rect 14188 28611 14240 28620
rect 7380 28500 7432 28552
rect 8576 28543 8628 28552
rect 8576 28509 8585 28543
rect 8585 28509 8619 28543
rect 8619 28509 8628 28543
rect 8576 28500 8628 28509
rect 9772 28543 9824 28552
rect 2044 28475 2096 28484
rect 2044 28441 2053 28475
rect 2053 28441 2087 28475
rect 2087 28441 2096 28475
rect 2044 28432 2096 28441
rect 3148 28364 3200 28416
rect 4068 28432 4120 28484
rect 4528 28432 4580 28484
rect 6644 28432 6696 28484
rect 9772 28509 9781 28543
rect 9781 28509 9815 28543
rect 9815 28509 9824 28543
rect 9772 28500 9824 28509
rect 11060 28500 11112 28552
rect 14188 28577 14197 28611
rect 14197 28577 14231 28611
rect 14231 28577 14240 28611
rect 14188 28568 14240 28577
rect 6368 28364 6420 28416
rect 7104 28364 7156 28416
rect 9864 28432 9916 28484
rect 10784 28432 10836 28484
rect 12808 28364 12860 28416
rect 14280 28500 14332 28552
rect 15476 28543 15528 28552
rect 15476 28509 15485 28543
rect 15485 28509 15519 28543
rect 15519 28509 15528 28543
rect 15476 28500 15528 28509
rect 16028 28568 16080 28620
rect 16396 28568 16448 28620
rect 18972 28611 19024 28620
rect 18972 28577 18981 28611
rect 18981 28577 19015 28611
rect 19015 28577 19024 28611
rect 18972 28568 19024 28577
rect 20260 28611 20312 28620
rect 20260 28577 20294 28611
rect 20294 28577 20312 28611
rect 20260 28568 20312 28577
rect 16212 28500 16264 28552
rect 19340 28500 19392 28552
rect 24860 28500 24912 28552
rect 25136 28568 25188 28620
rect 25228 28500 25280 28552
rect 26148 28568 26200 28620
rect 27988 28611 28040 28620
rect 27988 28577 27997 28611
rect 27997 28577 28031 28611
rect 28031 28577 28040 28611
rect 27988 28568 28040 28577
rect 13728 28432 13780 28484
rect 19248 28432 19300 28484
rect 15936 28364 15988 28416
rect 21364 28407 21416 28416
rect 21364 28373 21373 28407
rect 21373 28373 21407 28407
rect 21407 28373 21416 28407
rect 21364 28364 21416 28373
rect 22928 28364 22980 28416
rect 24860 28407 24912 28416
rect 24860 28373 24869 28407
rect 24869 28373 24903 28407
rect 24903 28373 24912 28407
rect 24860 28364 24912 28373
rect 28264 28432 28316 28484
rect 26056 28364 26108 28416
rect 5614 28262 5666 28314
rect 5678 28262 5730 28314
rect 5742 28262 5794 28314
rect 5806 28262 5858 28314
rect 14878 28262 14930 28314
rect 14942 28262 14994 28314
rect 15006 28262 15058 28314
rect 15070 28262 15122 28314
rect 24142 28262 24194 28314
rect 24206 28262 24258 28314
rect 24270 28262 24322 28314
rect 24334 28262 24386 28314
rect 2504 28160 2556 28212
rect 4896 28160 4948 28212
rect 5448 28160 5500 28212
rect 6184 28203 6236 28212
rect 6184 28169 6193 28203
rect 6193 28169 6227 28203
rect 6227 28169 6236 28203
rect 6184 28160 6236 28169
rect 1768 28135 1820 28144
rect 1768 28101 1777 28135
rect 1777 28101 1811 28135
rect 1811 28101 1820 28135
rect 1768 28092 1820 28101
rect 6828 28160 6880 28212
rect 7380 28160 7432 28212
rect 7932 28203 7984 28212
rect 7932 28169 7941 28203
rect 7941 28169 7975 28203
rect 7975 28169 7984 28203
rect 7932 28160 7984 28169
rect 11336 28160 11388 28212
rect 12808 28160 12860 28212
rect 3148 28067 3200 28076
rect 3148 28033 3157 28067
rect 3157 28033 3191 28067
rect 3191 28033 3200 28067
rect 3148 28024 3200 28033
rect 3792 28024 3844 28076
rect 1952 27999 2004 28008
rect 1952 27965 1961 27999
rect 1961 27965 1995 27999
rect 1995 27965 2004 27999
rect 1952 27956 2004 27965
rect 4252 27999 4304 28008
rect 4252 27965 4261 27999
rect 4261 27965 4295 27999
rect 4295 27965 4304 27999
rect 4252 27956 4304 27965
rect 6736 27956 6788 28008
rect 3240 27931 3292 27940
rect 3240 27897 3249 27931
rect 3249 27897 3283 27931
rect 3283 27897 3292 27931
rect 3240 27888 3292 27897
rect 3148 27863 3200 27872
rect 3148 27829 3157 27863
rect 3157 27829 3191 27863
rect 3191 27829 3200 27863
rect 3148 27820 3200 27829
rect 4344 27863 4396 27872
rect 4344 27829 4353 27863
rect 4353 27829 4387 27863
rect 4387 27829 4396 27863
rect 4344 27820 4396 27829
rect 11428 28092 11480 28144
rect 14648 28092 14700 28144
rect 14924 28092 14976 28144
rect 7380 28024 7432 28076
rect 7104 27999 7156 28008
rect 7104 27965 7113 27999
rect 7113 27965 7147 27999
rect 7147 27965 7156 27999
rect 7104 27956 7156 27965
rect 7196 27999 7248 28008
rect 7196 27965 7205 27999
rect 7205 27965 7239 27999
rect 7239 27965 7248 27999
rect 7656 27999 7708 28008
rect 7196 27956 7248 27965
rect 7656 27965 7665 27999
rect 7665 27965 7699 27999
rect 7699 27965 7708 27999
rect 7656 27956 7708 27965
rect 8760 27956 8812 28008
rect 9496 27999 9548 28008
rect 9496 27965 9505 27999
rect 9505 27965 9539 27999
rect 9539 27965 9548 27999
rect 9496 27956 9548 27965
rect 11060 28024 11112 28076
rect 11336 28024 11388 28076
rect 12348 28024 12400 28076
rect 12532 28024 12584 28076
rect 14096 28024 14148 28076
rect 16212 28024 16264 28076
rect 11428 27956 11480 28008
rect 11612 27956 11664 28008
rect 11980 27999 12032 28008
rect 11980 27965 11989 27999
rect 11989 27965 12023 27999
rect 12023 27965 12032 27999
rect 11980 27956 12032 27965
rect 13268 27956 13320 28008
rect 15200 27956 15252 28008
rect 15568 27999 15620 28008
rect 15568 27965 15577 27999
rect 15577 27965 15611 27999
rect 15611 27965 15620 27999
rect 15568 27956 15620 27965
rect 20168 28160 20220 28212
rect 25136 28160 25188 28212
rect 27988 28203 28040 28212
rect 27988 28169 27997 28203
rect 27997 28169 28031 28203
rect 28031 28169 28040 28203
rect 27988 28160 28040 28169
rect 17224 28024 17276 28076
rect 17500 28092 17552 28144
rect 19984 28024 20036 28076
rect 17868 27999 17920 28008
rect 17868 27965 17877 27999
rect 17877 27965 17911 27999
rect 17911 27965 17920 27999
rect 17868 27956 17920 27965
rect 9220 27888 9272 27940
rect 6920 27820 6972 27872
rect 7748 27820 7800 27872
rect 8208 27820 8260 27872
rect 11612 27863 11664 27872
rect 11612 27829 11621 27863
rect 11621 27829 11655 27863
rect 11655 27829 11664 27863
rect 11612 27820 11664 27829
rect 12532 27820 12584 27872
rect 13452 27820 13504 27872
rect 13820 27820 13872 27872
rect 17684 27888 17736 27940
rect 18512 27820 18564 27872
rect 18880 27863 18932 27872
rect 18880 27829 18889 27863
rect 18889 27829 18923 27863
rect 18923 27829 18932 27863
rect 18880 27820 18932 27829
rect 20076 27956 20128 28008
rect 21364 27956 21416 28008
rect 25228 28024 25280 28076
rect 24032 27956 24084 28008
rect 24124 27999 24176 28008
rect 24124 27965 24133 27999
rect 24133 27965 24167 27999
rect 24167 27965 24176 27999
rect 24124 27956 24176 27965
rect 24860 27956 24912 28008
rect 25688 27956 25740 28008
rect 20168 27931 20220 27940
rect 20168 27897 20177 27931
rect 20177 27897 20211 27931
rect 20211 27897 20220 27931
rect 20168 27888 20220 27897
rect 20444 27931 20496 27940
rect 20444 27897 20453 27931
rect 20453 27897 20487 27931
rect 20487 27897 20496 27931
rect 20444 27888 20496 27897
rect 20536 27931 20588 27940
rect 20536 27897 20545 27931
rect 20545 27897 20579 27931
rect 20579 27897 20588 27931
rect 21272 27931 21324 27940
rect 20536 27888 20588 27897
rect 21272 27897 21281 27931
rect 21281 27897 21315 27931
rect 21315 27897 21324 27931
rect 21272 27888 21324 27897
rect 21088 27820 21140 27872
rect 21640 27820 21692 27872
rect 21732 27820 21784 27872
rect 23388 27820 23440 27872
rect 23572 27820 23624 27872
rect 25596 27863 25648 27872
rect 25596 27829 25605 27863
rect 25605 27829 25639 27863
rect 25639 27829 25648 27863
rect 25596 27820 25648 27829
rect 25964 27931 26016 27940
rect 25964 27897 25973 27931
rect 25973 27897 26007 27931
rect 26007 27897 26016 27931
rect 26700 27956 26752 28008
rect 27988 28024 28040 28076
rect 27528 27956 27580 28008
rect 25964 27888 26016 27897
rect 27252 27888 27304 27940
rect 27804 27931 27856 27940
rect 26056 27820 26108 27872
rect 26240 27820 26292 27872
rect 27804 27897 27813 27931
rect 27813 27897 27847 27931
rect 27847 27897 27856 27931
rect 27804 27888 27856 27897
rect 27620 27863 27672 27872
rect 27620 27829 27629 27863
rect 27629 27829 27663 27863
rect 27663 27829 27672 27863
rect 27620 27820 27672 27829
rect 10246 27718 10298 27770
rect 10310 27718 10362 27770
rect 10374 27718 10426 27770
rect 10438 27718 10490 27770
rect 19510 27718 19562 27770
rect 19574 27718 19626 27770
rect 19638 27718 19690 27770
rect 19702 27718 19754 27770
rect 2044 27616 2096 27668
rect 3148 27616 3200 27668
rect 7196 27659 7248 27668
rect 7196 27625 7205 27659
rect 7205 27625 7239 27659
rect 7239 27625 7248 27659
rect 7196 27616 7248 27625
rect 7656 27616 7708 27668
rect 8300 27616 8352 27668
rect 1768 27548 1820 27600
rect 4344 27548 4396 27600
rect 6920 27591 6972 27600
rect 6920 27557 6929 27591
rect 6929 27557 6963 27591
rect 6963 27557 6972 27591
rect 6920 27548 6972 27557
rect 7012 27548 7064 27600
rect 8484 27591 8536 27600
rect 1676 27480 1728 27532
rect 2044 27480 2096 27532
rect 2412 27480 2464 27532
rect 7196 27523 7248 27532
rect 7196 27489 7205 27523
rect 7205 27489 7239 27523
rect 7239 27489 7248 27523
rect 7196 27480 7248 27489
rect 8208 27480 8260 27532
rect 8484 27557 8493 27591
rect 8493 27557 8527 27591
rect 8527 27557 8536 27591
rect 8484 27548 8536 27557
rect 8668 27480 8720 27532
rect 10876 27548 10928 27600
rect 17868 27616 17920 27668
rect 11704 27480 11756 27532
rect 2688 27412 2740 27464
rect 3884 27455 3936 27464
rect 3884 27421 3893 27455
rect 3893 27421 3927 27455
rect 3927 27421 3936 27455
rect 3884 27412 3936 27421
rect 3516 27344 3568 27396
rect 6828 27412 6880 27464
rect 12348 27412 12400 27464
rect 12808 27480 12860 27532
rect 13176 27480 13228 27532
rect 13820 27548 13872 27600
rect 14924 27548 14976 27600
rect 16396 27548 16448 27600
rect 13452 27523 13504 27532
rect 13452 27489 13473 27523
rect 13473 27489 13504 27523
rect 13452 27480 13504 27489
rect 17408 27480 17460 27532
rect 17500 27480 17552 27532
rect 18880 27548 18932 27600
rect 20076 27616 20128 27668
rect 20260 27616 20312 27668
rect 21732 27616 21784 27668
rect 22560 27548 22612 27600
rect 22928 27548 22980 27600
rect 23940 27616 23992 27668
rect 24676 27616 24728 27668
rect 23572 27548 23624 27600
rect 24032 27548 24084 27600
rect 25964 27616 26016 27668
rect 26148 27616 26200 27668
rect 27528 27616 27580 27668
rect 14556 27412 14608 27464
rect 15108 27412 15160 27464
rect 18788 27480 18840 27532
rect 19248 27480 19300 27532
rect 18604 27412 18656 27464
rect 20352 27412 20404 27464
rect 21088 27480 21140 27532
rect 23296 27480 23348 27532
rect 22468 27412 22520 27464
rect 5080 27344 5132 27396
rect 6368 27344 6420 27396
rect 21456 27344 21508 27396
rect 24860 27344 24912 27396
rect 4160 27276 4212 27328
rect 5908 27276 5960 27328
rect 6736 27276 6788 27328
rect 7380 27276 7432 27328
rect 9680 27276 9732 27328
rect 9956 27276 10008 27328
rect 16120 27276 16172 27328
rect 17868 27276 17920 27328
rect 19524 27276 19576 27328
rect 20536 27319 20588 27328
rect 20536 27285 20545 27319
rect 20545 27285 20579 27319
rect 20579 27285 20588 27319
rect 20536 27276 20588 27285
rect 25320 27276 25372 27328
rect 26332 27548 26384 27600
rect 26700 27591 26752 27600
rect 26700 27557 26709 27591
rect 26709 27557 26743 27591
rect 26743 27557 26752 27591
rect 26700 27548 26752 27557
rect 27252 27548 27304 27600
rect 26240 27480 26292 27532
rect 25780 27344 25832 27396
rect 26424 27344 26476 27396
rect 26240 27276 26292 27328
rect 26792 27319 26844 27328
rect 26792 27285 26801 27319
rect 26801 27285 26835 27319
rect 26835 27285 26844 27319
rect 26792 27276 26844 27285
rect 27620 27276 27672 27328
rect 28172 27319 28224 27328
rect 28172 27285 28181 27319
rect 28181 27285 28215 27319
rect 28215 27285 28224 27319
rect 28172 27276 28224 27285
rect 5614 27174 5666 27226
rect 5678 27174 5730 27226
rect 5742 27174 5794 27226
rect 5806 27174 5858 27226
rect 14878 27174 14930 27226
rect 14942 27174 14994 27226
rect 15006 27174 15058 27226
rect 15070 27174 15122 27226
rect 24142 27174 24194 27226
rect 24206 27174 24258 27226
rect 24270 27174 24322 27226
rect 24334 27174 24386 27226
rect 4160 27072 4212 27124
rect 7288 27072 7340 27124
rect 1676 27004 1728 27056
rect 1952 26911 2004 26920
rect 1952 26877 1961 26911
rect 1961 26877 1995 26911
rect 1995 26877 2004 26911
rect 1952 26868 2004 26877
rect 2780 26868 2832 26920
rect 3056 26911 3108 26920
rect 3056 26877 3065 26911
rect 3065 26877 3099 26911
rect 3099 26877 3108 26911
rect 3056 26868 3108 26877
rect 6368 27004 6420 27056
rect 11060 27072 11112 27124
rect 11612 27072 11664 27124
rect 13544 27072 13596 27124
rect 13728 27072 13780 27124
rect 17500 27115 17552 27124
rect 17500 27081 17509 27115
rect 17509 27081 17543 27115
rect 17543 27081 17552 27115
rect 17500 27072 17552 27081
rect 20536 27072 20588 27124
rect 23940 27072 23992 27124
rect 25780 27072 25832 27124
rect 27712 27072 27764 27124
rect 9956 27004 10008 27056
rect 10600 27004 10652 27056
rect 12164 27004 12216 27056
rect 6276 26936 6328 26988
rect 11612 26936 11664 26988
rect 11888 26936 11940 26988
rect 3976 26732 4028 26784
rect 4896 26800 4948 26852
rect 5080 26843 5132 26852
rect 5080 26809 5089 26843
rect 5089 26809 5123 26843
rect 5123 26809 5132 26843
rect 5080 26800 5132 26809
rect 10784 26868 10836 26920
rect 12532 26936 12584 26988
rect 6644 26732 6696 26784
rect 10876 26732 10928 26784
rect 11888 26800 11940 26852
rect 12532 26800 12584 26852
rect 18972 27004 19024 27056
rect 23572 27047 23624 27056
rect 23572 27013 23581 27047
rect 23581 27013 23615 27047
rect 23615 27013 23624 27047
rect 23572 27004 23624 27013
rect 13820 26979 13872 26988
rect 13820 26945 13829 26979
rect 13829 26945 13863 26979
rect 13863 26945 13872 26979
rect 13820 26936 13872 26945
rect 17224 26936 17276 26988
rect 17500 26936 17552 26988
rect 22468 26936 22520 26988
rect 12808 26911 12860 26920
rect 12808 26877 12817 26911
rect 12817 26877 12851 26911
rect 12851 26877 12860 26911
rect 12808 26868 12860 26877
rect 13544 26911 13596 26920
rect 12716 26732 12768 26784
rect 13544 26877 13553 26911
rect 13553 26877 13587 26911
rect 13587 26877 13596 26911
rect 13544 26868 13596 26877
rect 15844 26868 15896 26920
rect 16120 26868 16172 26920
rect 17684 26868 17736 26920
rect 17868 26868 17920 26920
rect 18788 26911 18840 26920
rect 13084 26800 13136 26852
rect 14740 26843 14792 26852
rect 14740 26809 14749 26843
rect 14749 26809 14783 26843
rect 14783 26809 14792 26843
rect 14740 26800 14792 26809
rect 14832 26800 14884 26852
rect 15936 26800 15988 26852
rect 18788 26877 18797 26911
rect 18797 26877 18831 26911
rect 18831 26877 18840 26911
rect 18788 26868 18840 26877
rect 18880 26868 18932 26920
rect 19524 26868 19576 26920
rect 26332 27004 26384 27056
rect 28356 27004 28408 27056
rect 24860 26936 24912 26988
rect 25412 26936 25464 26988
rect 25320 26911 25372 26920
rect 13728 26732 13780 26784
rect 14280 26732 14332 26784
rect 17040 26732 17092 26784
rect 20168 26732 20220 26784
rect 21916 26732 21968 26784
rect 22652 26843 22704 26852
rect 22652 26809 22661 26843
rect 22661 26809 22695 26843
rect 22695 26809 22704 26843
rect 23020 26843 23072 26852
rect 22652 26800 22704 26809
rect 23020 26809 23029 26843
rect 23029 26809 23063 26843
rect 23063 26809 23072 26843
rect 23020 26800 23072 26809
rect 25320 26877 25329 26911
rect 25329 26877 25363 26911
rect 25363 26877 25372 26911
rect 25320 26868 25372 26877
rect 28172 26936 28224 26988
rect 27804 26868 27856 26920
rect 24032 26800 24084 26852
rect 26424 26800 26476 26852
rect 26608 26843 26660 26852
rect 26608 26809 26617 26843
rect 26617 26809 26651 26843
rect 26651 26809 26660 26843
rect 26608 26800 26660 26809
rect 24952 26732 25004 26784
rect 25320 26732 25372 26784
rect 26700 26775 26752 26784
rect 26700 26741 26709 26775
rect 26709 26741 26743 26775
rect 26743 26741 26752 26775
rect 26700 26732 26752 26741
rect 10246 26630 10298 26682
rect 10310 26630 10362 26682
rect 10374 26630 10426 26682
rect 10438 26630 10490 26682
rect 19510 26630 19562 26682
rect 19574 26630 19626 26682
rect 19638 26630 19690 26682
rect 19702 26630 19754 26682
rect 1768 26571 1820 26580
rect 1768 26537 1777 26571
rect 1777 26537 1811 26571
rect 1811 26537 1820 26571
rect 1768 26528 1820 26537
rect 2412 26528 2464 26580
rect 2964 26528 3016 26580
rect 4620 26528 4672 26580
rect 5908 26528 5960 26580
rect 6828 26528 6880 26580
rect 9864 26571 9916 26580
rect 9864 26537 9873 26571
rect 9873 26537 9907 26571
rect 9907 26537 9916 26571
rect 9864 26528 9916 26537
rect 11704 26528 11756 26580
rect 12348 26528 12400 26580
rect 12716 26528 12768 26580
rect 13268 26528 13320 26580
rect 13820 26528 13872 26580
rect 15476 26528 15528 26580
rect 18788 26528 18840 26580
rect 20260 26528 20312 26580
rect 26608 26528 26660 26580
rect 10968 26503 11020 26512
rect 1952 26435 2004 26444
rect 1952 26401 1961 26435
rect 1961 26401 1995 26435
rect 1995 26401 2004 26435
rect 1952 26392 2004 26401
rect 2504 26392 2556 26444
rect 2228 26256 2280 26308
rect 3056 26435 3108 26444
rect 3056 26401 3065 26435
rect 3065 26401 3099 26435
rect 3099 26401 3108 26435
rect 3056 26392 3108 26401
rect 4160 26392 4212 26444
rect 8024 26435 8076 26444
rect 8024 26401 8033 26435
rect 8033 26401 8067 26435
rect 8067 26401 8076 26435
rect 8024 26392 8076 26401
rect 9036 26435 9088 26444
rect 9036 26401 9045 26435
rect 9045 26401 9079 26435
rect 9079 26401 9088 26435
rect 9036 26392 9088 26401
rect 4620 26367 4672 26376
rect 4620 26333 4629 26367
rect 4629 26333 4663 26367
rect 4663 26333 4672 26367
rect 4620 26324 4672 26333
rect 4896 26324 4948 26376
rect 8116 26367 8168 26376
rect 8116 26333 8125 26367
rect 8125 26333 8159 26367
rect 8159 26333 8168 26367
rect 8116 26324 8168 26333
rect 5172 26256 5224 26308
rect 6092 26256 6144 26308
rect 10968 26469 10977 26503
rect 10977 26469 11011 26503
rect 11011 26469 11020 26503
rect 10968 26460 11020 26469
rect 10140 26392 10192 26444
rect 10784 26435 10836 26444
rect 10784 26401 10793 26435
rect 10793 26401 10827 26435
rect 10827 26401 10836 26435
rect 10784 26392 10836 26401
rect 12256 26460 12308 26512
rect 14004 26460 14056 26512
rect 14832 26460 14884 26512
rect 17408 26460 17460 26512
rect 12532 26392 12584 26444
rect 13268 26392 13320 26444
rect 13544 26392 13596 26444
rect 14556 26392 14608 26444
rect 14648 26392 14700 26444
rect 10416 26324 10468 26376
rect 11152 26324 11204 26376
rect 15476 26392 15528 26444
rect 15936 26324 15988 26376
rect 18328 26392 18380 26444
rect 18604 26435 18656 26444
rect 18604 26401 18613 26435
rect 18613 26401 18647 26435
rect 18647 26401 18656 26435
rect 18604 26392 18656 26401
rect 23020 26460 23072 26512
rect 26148 26460 26200 26512
rect 27988 26503 28040 26512
rect 27988 26469 27997 26503
rect 27997 26469 28031 26503
rect 28031 26469 28040 26503
rect 27988 26460 28040 26469
rect 18788 26324 18840 26376
rect 9680 26256 9732 26308
rect 22284 26256 22336 26308
rect 22652 26256 22704 26308
rect 23296 26256 23348 26308
rect 26056 26392 26108 26444
rect 26240 26324 26292 26376
rect 25412 26299 25464 26308
rect 9588 26188 9640 26240
rect 13360 26188 13412 26240
rect 13544 26188 13596 26240
rect 13728 26188 13780 26240
rect 14096 26188 14148 26240
rect 14280 26188 14332 26240
rect 25412 26265 25421 26299
rect 25421 26265 25455 26299
rect 25455 26265 25464 26299
rect 25412 26256 25464 26265
rect 25688 26256 25740 26308
rect 26148 26299 26200 26308
rect 26148 26265 26157 26299
rect 26157 26265 26191 26299
rect 26191 26265 26200 26299
rect 26148 26256 26200 26265
rect 28172 26299 28224 26308
rect 28172 26265 28181 26299
rect 28181 26265 28215 26299
rect 28215 26265 28224 26299
rect 28172 26256 28224 26265
rect 5614 26086 5666 26138
rect 5678 26086 5730 26138
rect 5742 26086 5794 26138
rect 5806 26086 5858 26138
rect 14878 26086 14930 26138
rect 14942 26086 14994 26138
rect 15006 26086 15058 26138
rect 15070 26086 15122 26138
rect 24142 26086 24194 26138
rect 24206 26086 24258 26138
rect 24270 26086 24322 26138
rect 24334 26086 24386 26138
rect 1768 25848 1820 25900
rect 2044 25848 2096 25900
rect 6460 25984 6512 26036
rect 7196 25984 7248 26036
rect 7472 26027 7524 26036
rect 7472 25993 7481 26027
rect 7481 25993 7515 26027
rect 7515 25993 7524 26027
rect 7472 25984 7524 25993
rect 10968 25984 11020 26036
rect 12348 25984 12400 26036
rect 12624 25984 12676 26036
rect 12716 25984 12768 26036
rect 13360 25984 13412 26036
rect 16120 25984 16172 26036
rect 17408 25984 17460 26036
rect 20168 25984 20220 26036
rect 23848 25984 23900 26036
rect 25688 25984 25740 26036
rect 27804 25984 27856 26036
rect 11336 25916 11388 25968
rect 6184 25848 6236 25900
rect 10876 25848 10928 25900
rect 12256 25916 12308 25968
rect 14924 25916 14976 25968
rect 16212 25916 16264 25968
rect 17500 25916 17552 25968
rect 15476 25848 15528 25900
rect 19340 25916 19392 25968
rect 24676 25916 24728 25968
rect 18788 25848 18840 25900
rect 18972 25891 19024 25900
rect 18972 25857 18981 25891
rect 18981 25857 19015 25891
rect 19015 25857 19024 25891
rect 18972 25848 19024 25857
rect 23848 25848 23900 25900
rect 24952 25848 25004 25900
rect 1860 25823 1912 25832
rect 1860 25789 1869 25823
rect 1869 25789 1903 25823
rect 1903 25789 1912 25823
rect 1860 25780 1912 25789
rect 4252 25780 4304 25832
rect 5172 25780 5224 25832
rect 6920 25823 6972 25832
rect 6920 25789 6929 25823
rect 6929 25789 6963 25823
rect 6963 25789 6972 25823
rect 6920 25780 6972 25789
rect 7380 25823 7432 25832
rect 7380 25789 7389 25823
rect 7389 25789 7423 25823
rect 7423 25789 7432 25823
rect 7380 25780 7432 25789
rect 7748 25823 7800 25832
rect 7748 25789 7757 25823
rect 7757 25789 7791 25823
rect 7791 25789 7800 25823
rect 7748 25780 7800 25789
rect 8300 25823 8352 25832
rect 8300 25789 8309 25823
rect 8309 25789 8343 25823
rect 8343 25789 8352 25823
rect 8300 25780 8352 25789
rect 9496 25823 9548 25832
rect 9496 25789 9505 25823
rect 9505 25789 9539 25823
rect 9539 25789 9548 25823
rect 9496 25780 9548 25789
rect 9588 25780 9640 25832
rect 11704 25780 11756 25832
rect 14556 25780 14608 25832
rect 16580 25823 16632 25832
rect 16580 25789 16589 25823
rect 16589 25789 16623 25823
rect 16623 25789 16632 25823
rect 16580 25780 16632 25789
rect 18604 25823 18656 25832
rect 18604 25789 18613 25823
rect 18613 25789 18647 25823
rect 18647 25789 18656 25823
rect 18604 25780 18656 25789
rect 19340 25780 19392 25832
rect 24032 25780 24084 25832
rect 24492 25780 24544 25832
rect 26700 25780 26752 25832
rect 2044 25755 2096 25764
rect 2044 25721 2053 25755
rect 2053 25721 2087 25755
rect 2087 25721 2096 25755
rect 2044 25712 2096 25721
rect 6644 25755 6696 25764
rect 6644 25721 6653 25755
rect 6653 25721 6687 25755
rect 6687 25721 6696 25755
rect 6644 25712 6696 25721
rect 7564 25712 7616 25764
rect 13084 25712 13136 25764
rect 13268 25712 13320 25764
rect 13820 25712 13872 25764
rect 2320 25644 2372 25696
rect 4804 25644 4856 25696
rect 10876 25687 10928 25696
rect 10876 25653 10885 25687
rect 10885 25653 10919 25687
rect 10919 25653 10928 25687
rect 10876 25644 10928 25653
rect 11704 25644 11756 25696
rect 11980 25644 12032 25696
rect 12716 25644 12768 25696
rect 16120 25712 16172 25764
rect 21272 25712 21324 25764
rect 18052 25644 18104 25696
rect 22560 25687 22612 25696
rect 22560 25653 22569 25687
rect 22569 25653 22603 25687
rect 22603 25653 22612 25687
rect 22560 25644 22612 25653
rect 23020 25644 23072 25696
rect 26056 25712 26108 25764
rect 27988 25780 28040 25832
rect 27436 25712 27488 25764
rect 28080 25644 28132 25696
rect 10246 25542 10298 25594
rect 10310 25542 10362 25594
rect 10374 25542 10426 25594
rect 10438 25542 10490 25594
rect 19510 25542 19562 25594
rect 19574 25542 19626 25594
rect 19638 25542 19690 25594
rect 19702 25542 19754 25594
rect 4804 25483 4856 25492
rect 4804 25449 4813 25483
rect 4813 25449 4847 25483
rect 4847 25449 4856 25483
rect 4804 25440 4856 25449
rect 5356 25440 5408 25492
rect 5448 25440 5500 25492
rect 8024 25440 8076 25492
rect 8116 25440 8168 25492
rect 9036 25440 9088 25492
rect 10784 25440 10836 25492
rect 12532 25440 12584 25492
rect 13820 25440 13872 25492
rect 1768 25415 1820 25424
rect 1768 25381 1777 25415
rect 1777 25381 1811 25415
rect 1811 25381 1820 25415
rect 1768 25372 1820 25381
rect 2136 25372 2188 25424
rect 7380 25372 7432 25424
rect 2504 25347 2556 25356
rect 2504 25313 2513 25347
rect 2513 25313 2547 25347
rect 2547 25313 2556 25347
rect 2504 25304 2556 25313
rect 2596 25304 2648 25356
rect 4252 25304 4304 25356
rect 5448 25304 5500 25356
rect 7564 25304 7616 25356
rect 7840 25304 7892 25356
rect 10140 25372 10192 25424
rect 10876 25372 10928 25424
rect 14188 25440 14240 25492
rect 15568 25440 15620 25492
rect 9220 25347 9272 25356
rect 3424 25279 3476 25288
rect 3424 25245 3433 25279
rect 3433 25245 3467 25279
rect 3467 25245 3476 25279
rect 3424 25236 3476 25245
rect 8300 25236 8352 25288
rect 9220 25313 9229 25347
rect 9229 25313 9263 25347
rect 9263 25313 9272 25347
rect 9220 25304 9272 25313
rect 9404 25347 9456 25356
rect 9404 25313 9413 25347
rect 9413 25313 9447 25347
rect 9447 25313 9456 25347
rect 9404 25304 9456 25313
rect 10600 25347 10652 25356
rect 10600 25313 10609 25347
rect 10609 25313 10643 25347
rect 10643 25313 10652 25347
rect 10600 25304 10652 25313
rect 13268 25304 13320 25356
rect 11060 25236 11112 25288
rect 14280 25372 14332 25424
rect 18972 25440 19024 25492
rect 21824 25372 21876 25424
rect 1584 25168 1636 25220
rect 6368 25168 6420 25220
rect 12624 25168 12676 25220
rect 13176 25168 13228 25220
rect 14280 25168 14332 25220
rect 14924 25304 14976 25356
rect 15200 25236 15252 25288
rect 15476 25236 15528 25288
rect 15844 25347 15896 25356
rect 15844 25313 15853 25347
rect 15853 25313 15887 25347
rect 15887 25313 15896 25347
rect 16028 25347 16080 25356
rect 15844 25304 15896 25313
rect 16028 25313 16037 25347
rect 16037 25313 16071 25347
rect 16071 25313 16080 25347
rect 16028 25304 16080 25313
rect 17316 25304 17368 25356
rect 26700 25440 26752 25492
rect 27528 25440 27580 25492
rect 23020 25372 23072 25424
rect 25872 25415 25924 25424
rect 25872 25381 25881 25415
rect 25881 25381 25915 25415
rect 25915 25381 25924 25415
rect 26240 25415 26292 25424
rect 25872 25372 25924 25381
rect 26240 25381 26249 25415
rect 26249 25381 26283 25415
rect 26283 25381 26292 25415
rect 26240 25372 26292 25381
rect 22284 25304 22336 25356
rect 17040 25236 17092 25288
rect 15292 25168 15344 25220
rect 15568 25168 15620 25220
rect 4528 25100 4580 25152
rect 5264 25100 5316 25152
rect 6276 25100 6328 25152
rect 13728 25143 13780 25152
rect 13728 25109 13737 25143
rect 13737 25109 13771 25143
rect 13771 25109 13780 25143
rect 13728 25100 13780 25109
rect 14096 25100 14148 25152
rect 15200 25100 15252 25152
rect 15384 25100 15436 25152
rect 19248 25236 19300 25288
rect 19340 25236 19392 25288
rect 22744 25304 22796 25356
rect 24492 25347 24544 25356
rect 24492 25313 24501 25347
rect 24501 25313 24535 25347
rect 24535 25313 24544 25347
rect 24492 25304 24544 25313
rect 25688 25304 25740 25356
rect 23388 25236 23440 25288
rect 19064 25168 19116 25220
rect 22100 25168 22152 25220
rect 24952 25236 25004 25288
rect 25136 25236 25188 25288
rect 25504 25236 25556 25288
rect 20904 25143 20956 25152
rect 20904 25109 20913 25143
rect 20913 25109 20947 25143
rect 20947 25109 20956 25143
rect 20904 25100 20956 25109
rect 22928 25143 22980 25152
rect 22928 25109 22937 25143
rect 22937 25109 22971 25143
rect 22971 25109 22980 25143
rect 22928 25100 22980 25109
rect 23020 25143 23072 25152
rect 23020 25109 23029 25143
rect 23029 25109 23063 25143
rect 23063 25109 23072 25143
rect 23020 25100 23072 25109
rect 24768 25100 24820 25152
rect 25136 25100 25188 25152
rect 27528 25100 27580 25152
rect 5614 24998 5666 25050
rect 5678 24998 5730 25050
rect 5742 24998 5794 25050
rect 5806 24998 5858 25050
rect 14878 24998 14930 25050
rect 14942 24998 14994 25050
rect 15006 24998 15058 25050
rect 15070 24998 15122 25050
rect 24142 24998 24194 25050
rect 24206 24998 24258 25050
rect 24270 24998 24322 25050
rect 24334 24998 24386 25050
rect 10600 24896 10652 24948
rect 10876 24896 10928 24948
rect 14280 24896 14332 24948
rect 16028 24896 16080 24948
rect 16580 24896 16632 24948
rect 23388 24896 23440 24948
rect 25136 24896 25188 24948
rect 26240 24896 26292 24948
rect 27436 24939 27488 24948
rect 27436 24905 27445 24939
rect 27445 24905 27479 24939
rect 27479 24905 27488 24939
rect 27436 24896 27488 24905
rect 2228 24692 2280 24744
rect 2504 24692 2556 24744
rect 5264 24760 5316 24812
rect 6092 24828 6144 24880
rect 11336 24828 11388 24880
rect 2688 24692 2740 24744
rect 4896 24692 4948 24744
rect 5080 24735 5132 24744
rect 5080 24701 5089 24735
rect 5089 24701 5123 24735
rect 5123 24701 5132 24735
rect 5080 24692 5132 24701
rect 1584 24667 1636 24676
rect 1584 24633 1593 24667
rect 1593 24633 1627 24667
rect 1627 24633 1636 24667
rect 1584 24624 1636 24633
rect 1768 24624 1820 24676
rect 2044 24624 2096 24676
rect 5816 24692 5868 24744
rect 1492 24556 1544 24608
rect 2504 24556 2556 24608
rect 2688 24599 2740 24608
rect 2688 24565 2697 24599
rect 2697 24565 2731 24599
rect 2731 24565 2740 24599
rect 2688 24556 2740 24565
rect 3700 24556 3752 24608
rect 5540 24624 5592 24676
rect 6460 24760 6512 24812
rect 9220 24760 9272 24812
rect 9956 24760 10008 24812
rect 10784 24803 10836 24812
rect 10784 24769 10793 24803
rect 10793 24769 10827 24803
rect 10827 24769 10836 24803
rect 10784 24760 10836 24769
rect 10508 24692 10560 24744
rect 12716 24828 12768 24880
rect 12256 24760 12308 24812
rect 5816 24599 5868 24608
rect 5816 24565 5825 24599
rect 5825 24565 5859 24599
rect 5859 24565 5868 24599
rect 5816 24556 5868 24565
rect 7656 24624 7708 24676
rect 12716 24692 12768 24744
rect 13360 24828 13412 24880
rect 12256 24624 12308 24676
rect 15108 24692 15160 24744
rect 16120 24760 16172 24812
rect 15384 24735 15436 24744
rect 15384 24701 15393 24735
rect 15393 24701 15427 24735
rect 15427 24701 15436 24735
rect 15384 24692 15436 24701
rect 15660 24692 15712 24744
rect 16212 24692 16264 24744
rect 17500 24828 17552 24880
rect 22284 24871 22336 24880
rect 22284 24837 22293 24871
rect 22293 24837 22327 24871
rect 22327 24837 22336 24871
rect 22284 24828 22336 24837
rect 27896 24828 27948 24880
rect 17040 24760 17092 24812
rect 19984 24760 20036 24812
rect 21824 24760 21876 24812
rect 6092 24556 6144 24608
rect 11336 24556 11388 24608
rect 11520 24556 11572 24608
rect 15844 24624 15896 24676
rect 16672 24624 16724 24676
rect 17316 24692 17368 24744
rect 20444 24735 20496 24744
rect 20168 24667 20220 24676
rect 20168 24633 20177 24667
rect 20177 24633 20211 24667
rect 20211 24633 20220 24667
rect 20168 24624 20220 24633
rect 20444 24701 20453 24735
rect 20453 24701 20487 24735
rect 20487 24701 20496 24735
rect 20444 24692 20496 24701
rect 20904 24735 20956 24744
rect 20904 24701 20913 24735
rect 20913 24701 20947 24735
rect 20947 24701 20956 24735
rect 20904 24692 20956 24701
rect 21916 24692 21968 24744
rect 25964 24692 26016 24744
rect 27804 24735 27856 24744
rect 27804 24701 27813 24735
rect 27813 24701 27847 24735
rect 27847 24701 27856 24735
rect 27804 24692 27856 24701
rect 28080 24692 28132 24744
rect 20536 24667 20588 24676
rect 20536 24633 20545 24667
rect 20545 24633 20579 24667
rect 20579 24633 20588 24667
rect 20536 24624 20588 24633
rect 21732 24624 21784 24676
rect 22284 24624 22336 24676
rect 22652 24624 22704 24676
rect 22928 24624 22980 24676
rect 24768 24624 24820 24676
rect 20720 24556 20772 24608
rect 21456 24599 21508 24608
rect 21456 24565 21465 24599
rect 21465 24565 21499 24599
rect 21499 24565 21508 24599
rect 21456 24556 21508 24565
rect 10246 24454 10298 24506
rect 10310 24454 10362 24506
rect 10374 24454 10426 24506
rect 10438 24454 10490 24506
rect 19510 24454 19562 24506
rect 19574 24454 19626 24506
rect 19638 24454 19690 24506
rect 19702 24454 19754 24506
rect 5816 24352 5868 24404
rect 7380 24352 7432 24404
rect 13268 24395 13320 24404
rect 13268 24361 13277 24395
rect 13277 24361 13311 24395
rect 13311 24361 13320 24395
rect 13268 24352 13320 24361
rect 2504 24284 2556 24336
rect 6460 24284 6512 24336
rect 6644 24284 6696 24336
rect 14096 24352 14148 24404
rect 14188 24352 14240 24404
rect 15476 24352 15528 24404
rect 15844 24352 15896 24404
rect 16672 24352 16724 24404
rect 23020 24352 23072 24404
rect 1952 24259 2004 24268
rect 1952 24225 1961 24259
rect 1961 24225 1995 24259
rect 1995 24225 2004 24259
rect 1952 24216 2004 24225
rect 3148 24259 3200 24268
rect 3148 24225 3182 24259
rect 3182 24225 3200 24259
rect 6828 24259 6880 24268
rect 3148 24216 3200 24225
rect 6828 24225 6837 24259
rect 6837 24225 6871 24259
rect 6871 24225 6880 24259
rect 6828 24216 6880 24225
rect 11704 24216 11756 24268
rect 12072 24216 12124 24268
rect 13544 24284 13596 24336
rect 12716 24259 12768 24268
rect 2872 24191 2924 24200
rect 2872 24157 2881 24191
rect 2881 24157 2915 24191
rect 2915 24157 2924 24191
rect 2872 24148 2924 24157
rect 4804 24148 4856 24200
rect 5264 24148 5316 24200
rect 7012 24148 7064 24200
rect 12716 24225 12725 24259
rect 12725 24225 12759 24259
rect 12759 24225 12768 24259
rect 12716 24216 12768 24225
rect 13176 24259 13228 24268
rect 13176 24225 13185 24259
rect 13185 24225 13219 24259
rect 13219 24225 13228 24259
rect 13176 24216 13228 24225
rect 13360 24259 13412 24268
rect 13360 24225 13369 24259
rect 13369 24225 13403 24259
rect 13403 24225 13412 24259
rect 13360 24216 13412 24225
rect 13728 24216 13780 24268
rect 15108 24216 15160 24268
rect 16580 24284 16632 24336
rect 19984 24284 20036 24336
rect 20444 24284 20496 24336
rect 16120 24259 16172 24268
rect 16120 24225 16129 24259
rect 16129 24225 16163 24259
rect 16163 24225 16172 24259
rect 16120 24216 16172 24225
rect 13544 24148 13596 24200
rect 14188 24148 14240 24200
rect 15292 24148 15344 24200
rect 15844 24148 15896 24200
rect 16396 24148 16448 24200
rect 16672 24148 16724 24200
rect 17040 24148 17092 24200
rect 4896 24080 4948 24132
rect 11060 24080 11112 24132
rect 12716 24080 12768 24132
rect 13360 24080 13412 24132
rect 4252 24055 4304 24064
rect 4252 24021 4261 24055
rect 4261 24021 4295 24055
rect 4295 24021 4304 24055
rect 4252 24012 4304 24021
rect 6000 24012 6052 24064
rect 11704 24012 11756 24064
rect 12348 24012 12400 24064
rect 13268 24012 13320 24064
rect 19064 24216 19116 24268
rect 21180 24216 21232 24268
rect 21640 24259 21692 24268
rect 21640 24225 21649 24259
rect 21649 24225 21683 24259
rect 21683 24225 21692 24259
rect 21640 24216 21692 24225
rect 22560 24259 22612 24268
rect 22560 24225 22569 24259
rect 22569 24225 22603 24259
rect 22603 24225 22612 24259
rect 22560 24216 22612 24225
rect 22652 24216 22704 24268
rect 18328 24191 18380 24200
rect 18328 24157 18337 24191
rect 18337 24157 18371 24191
rect 18371 24157 18380 24191
rect 18328 24148 18380 24157
rect 21364 24148 21416 24200
rect 21824 24148 21876 24200
rect 21916 24148 21968 24200
rect 26148 24327 26200 24336
rect 26148 24293 26157 24327
rect 26157 24293 26191 24327
rect 26191 24293 26200 24327
rect 26148 24284 26200 24293
rect 26332 24284 26384 24336
rect 22100 24080 22152 24132
rect 23572 24080 23624 24132
rect 24492 24191 24544 24200
rect 24492 24157 24501 24191
rect 24501 24157 24535 24191
rect 24535 24157 24544 24191
rect 24492 24148 24544 24157
rect 24768 24080 24820 24132
rect 28172 24123 28224 24132
rect 28172 24089 28181 24123
rect 28181 24089 28215 24123
rect 28215 24089 28224 24123
rect 28172 24080 28224 24089
rect 18236 24012 18288 24064
rect 22652 24055 22704 24064
rect 22652 24021 22661 24055
rect 22661 24021 22695 24055
rect 22695 24021 22704 24055
rect 22652 24012 22704 24021
rect 26792 24055 26844 24064
rect 26792 24021 26801 24055
rect 26801 24021 26835 24055
rect 26835 24021 26844 24055
rect 26792 24012 26844 24021
rect 5614 23910 5666 23962
rect 5678 23910 5730 23962
rect 5742 23910 5794 23962
rect 5806 23910 5858 23962
rect 14878 23910 14930 23962
rect 14942 23910 14994 23962
rect 15006 23910 15058 23962
rect 15070 23910 15122 23962
rect 24142 23910 24194 23962
rect 24206 23910 24258 23962
rect 24270 23910 24322 23962
rect 24334 23910 24386 23962
rect 2504 23851 2556 23860
rect 2504 23817 2513 23851
rect 2513 23817 2547 23851
rect 2547 23817 2556 23851
rect 2504 23808 2556 23817
rect 6092 23808 6144 23860
rect 6644 23808 6696 23860
rect 4528 23740 4580 23792
rect 4896 23740 4948 23792
rect 5908 23740 5960 23792
rect 1860 23672 1912 23724
rect 2780 23604 2832 23656
rect 3332 23647 3384 23656
rect 3332 23613 3341 23647
rect 3341 23613 3375 23647
rect 3375 23613 3384 23647
rect 3332 23604 3384 23613
rect 4528 23604 4580 23656
rect 1584 23536 1636 23588
rect 2136 23536 2188 23588
rect 6092 23579 6144 23588
rect 6092 23545 6101 23579
rect 6101 23545 6135 23579
rect 6135 23545 6144 23579
rect 6092 23536 6144 23545
rect 4804 23468 4856 23520
rect 6736 23740 6788 23792
rect 18328 23808 18380 23860
rect 21272 23851 21324 23860
rect 21272 23817 21281 23851
rect 21281 23817 21315 23851
rect 21315 23817 21324 23851
rect 21272 23808 21324 23817
rect 27988 23851 28040 23860
rect 27988 23817 27997 23851
rect 27997 23817 28031 23851
rect 28031 23817 28040 23851
rect 27988 23808 28040 23817
rect 20720 23740 20772 23792
rect 8484 23672 8536 23724
rect 11704 23715 11756 23724
rect 11704 23681 11713 23715
rect 11713 23681 11747 23715
rect 11747 23681 11756 23715
rect 11704 23672 11756 23681
rect 12072 23672 12124 23724
rect 8576 23536 8628 23588
rect 9128 23536 9180 23588
rect 8392 23511 8444 23520
rect 8392 23477 8401 23511
rect 8401 23477 8435 23511
rect 8435 23477 8444 23511
rect 8392 23468 8444 23477
rect 14188 23672 14240 23724
rect 16028 23672 16080 23724
rect 14280 23604 14332 23656
rect 14740 23604 14792 23656
rect 16580 23604 16632 23656
rect 17224 23604 17276 23656
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 16396 23536 16448 23588
rect 16672 23536 16724 23588
rect 18328 23604 18380 23656
rect 21272 23672 21324 23724
rect 21732 23672 21784 23724
rect 26332 23672 26384 23724
rect 20996 23604 21048 23656
rect 21180 23647 21232 23656
rect 21180 23613 21189 23647
rect 21189 23613 21223 23647
rect 21223 23613 21232 23647
rect 21180 23604 21232 23613
rect 22652 23604 22704 23656
rect 26516 23604 26568 23656
rect 27620 23672 27672 23724
rect 26884 23647 26936 23656
rect 26884 23613 26893 23647
rect 26893 23613 26927 23647
rect 26927 23613 26936 23647
rect 26884 23604 26936 23613
rect 27160 23604 27212 23656
rect 20076 23536 20128 23588
rect 26240 23536 26292 23588
rect 12072 23468 12124 23520
rect 13360 23468 13412 23520
rect 13544 23468 13596 23520
rect 16948 23468 17000 23520
rect 17224 23468 17276 23520
rect 18052 23468 18104 23520
rect 19984 23468 20036 23520
rect 10246 23366 10298 23418
rect 10310 23366 10362 23418
rect 10374 23366 10426 23418
rect 10438 23366 10490 23418
rect 19510 23366 19562 23418
rect 19574 23366 19626 23418
rect 19638 23366 19690 23418
rect 19702 23366 19754 23418
rect 2688 23264 2740 23316
rect 3148 23264 3200 23316
rect 4252 23264 4304 23316
rect 4712 23264 4764 23316
rect 6828 23264 6880 23316
rect 8392 23264 8444 23316
rect 12256 23264 12308 23316
rect 14096 23264 14148 23316
rect 1768 23196 1820 23248
rect 17224 23264 17276 23316
rect 1400 23128 1452 23180
rect 2780 23128 2832 23180
rect 4160 23128 4212 23180
rect 14556 23196 14608 23248
rect 6736 23128 6788 23180
rect 8116 23171 8168 23180
rect 8116 23137 8150 23171
rect 8150 23137 8168 23171
rect 8116 23128 8168 23137
rect 9588 23128 9640 23180
rect 10600 23128 10652 23180
rect 10876 23171 10928 23180
rect 10876 23137 10885 23171
rect 10885 23137 10919 23171
rect 10919 23137 10928 23171
rect 10876 23128 10928 23137
rect 4344 23060 4396 23112
rect 12624 23128 12676 23180
rect 14740 23128 14792 23180
rect 16396 23196 16448 23248
rect 18328 23196 18380 23248
rect 28080 23264 28132 23316
rect 17040 23128 17092 23180
rect 17316 23128 17368 23180
rect 17408 23128 17460 23180
rect 25596 23128 25648 23180
rect 26516 23171 26568 23180
rect 26516 23137 26525 23171
rect 26525 23137 26559 23171
rect 26559 23137 26568 23171
rect 26516 23128 26568 23137
rect 6092 22992 6144 23044
rect 6644 22992 6696 23044
rect 2872 22924 2924 22976
rect 8944 22992 8996 23044
rect 9496 22992 9548 23044
rect 9772 22992 9824 23044
rect 26424 23060 26476 23112
rect 26700 23060 26752 23112
rect 27252 23060 27304 23112
rect 15476 22992 15528 23044
rect 15568 22992 15620 23044
rect 16580 22992 16632 23044
rect 25136 23035 25188 23044
rect 25136 23001 25145 23035
rect 25145 23001 25179 23035
rect 25179 23001 25188 23035
rect 25136 22992 25188 23001
rect 25872 23035 25924 23044
rect 25872 23001 25881 23035
rect 25881 23001 25915 23035
rect 25915 23001 25924 23035
rect 25872 22992 25924 23001
rect 28172 23035 28224 23044
rect 28172 23001 28181 23035
rect 28181 23001 28215 23035
rect 28215 23001 28224 23035
rect 28172 22992 28224 23001
rect 9220 22967 9272 22976
rect 9220 22933 9229 22967
rect 9229 22933 9263 22967
rect 9263 22933 9272 22967
rect 9220 22924 9272 22933
rect 10140 22924 10192 22976
rect 12532 22924 12584 22976
rect 27804 22924 27856 22976
rect 5614 22822 5666 22874
rect 5678 22822 5730 22874
rect 5742 22822 5794 22874
rect 5806 22822 5858 22874
rect 14878 22822 14930 22874
rect 14942 22822 14994 22874
rect 15006 22822 15058 22874
rect 15070 22822 15122 22874
rect 24142 22822 24194 22874
rect 24206 22822 24258 22874
rect 24270 22822 24322 22874
rect 24334 22822 24386 22874
rect 2044 22720 2096 22772
rect 2596 22720 2648 22772
rect 8484 22763 8536 22772
rect 8484 22729 8493 22763
rect 8493 22729 8527 22763
rect 8527 22729 8536 22763
rect 8484 22720 8536 22729
rect 9588 22763 9640 22772
rect 9588 22729 9597 22763
rect 9597 22729 9631 22763
rect 9631 22729 9640 22763
rect 9588 22720 9640 22729
rect 4068 22652 4120 22704
rect 10876 22652 10928 22704
rect 5540 22584 5592 22636
rect 6276 22584 6328 22636
rect 6460 22584 6512 22636
rect 6736 22627 6788 22636
rect 6736 22593 6745 22627
rect 6745 22593 6779 22627
rect 6779 22593 6788 22627
rect 6736 22584 6788 22593
rect 8668 22584 8720 22636
rect 10600 22584 10652 22636
rect 23112 22720 23164 22772
rect 24492 22720 24544 22772
rect 24768 22720 24820 22772
rect 25964 22720 26016 22772
rect 2872 22516 2924 22568
rect 4252 22559 4304 22568
rect 4252 22525 4261 22559
rect 4261 22525 4295 22559
rect 4295 22525 4304 22559
rect 4252 22516 4304 22525
rect 6644 22559 6696 22568
rect 6644 22525 6653 22559
rect 6653 22525 6687 22559
rect 6687 22525 6696 22559
rect 6644 22516 6696 22525
rect 8392 22559 8444 22568
rect 8392 22525 8401 22559
rect 8401 22525 8435 22559
rect 8435 22525 8444 22559
rect 8392 22516 8444 22525
rect 8576 22559 8628 22568
rect 8576 22525 8585 22559
rect 8585 22525 8619 22559
rect 8619 22525 8628 22559
rect 8576 22516 8628 22525
rect 10876 22559 10928 22568
rect 2044 22448 2096 22500
rect 8484 22448 8536 22500
rect 9220 22448 9272 22500
rect 10876 22525 10885 22559
rect 10885 22525 10919 22559
rect 10919 22525 10928 22559
rect 10876 22516 10928 22525
rect 11152 22559 11204 22568
rect 2780 22423 2832 22432
rect 2780 22389 2789 22423
rect 2789 22389 2823 22423
rect 2823 22389 2832 22423
rect 4344 22423 4396 22432
rect 2780 22380 2832 22389
rect 4344 22389 4353 22423
rect 4353 22389 4387 22423
rect 4387 22389 4396 22423
rect 4344 22380 4396 22389
rect 7472 22423 7524 22432
rect 7472 22389 7481 22423
rect 7481 22389 7515 22423
rect 7515 22389 7524 22423
rect 7472 22380 7524 22389
rect 11152 22525 11161 22559
rect 11161 22525 11195 22559
rect 11195 22525 11204 22559
rect 11152 22516 11204 22525
rect 12532 22627 12584 22636
rect 12532 22593 12541 22627
rect 12541 22593 12575 22627
rect 12575 22593 12584 22627
rect 12532 22584 12584 22593
rect 11520 22448 11572 22500
rect 13820 22584 13872 22636
rect 15568 22559 15620 22568
rect 15568 22525 15577 22559
rect 15577 22525 15611 22559
rect 15611 22525 15620 22559
rect 15568 22516 15620 22525
rect 16028 22652 16080 22704
rect 17684 22652 17736 22704
rect 18052 22652 18104 22704
rect 19064 22652 19116 22704
rect 22192 22652 22244 22704
rect 22744 22695 22796 22704
rect 22744 22661 22753 22695
rect 22753 22661 22787 22695
rect 22787 22661 22796 22695
rect 22744 22652 22796 22661
rect 23848 22652 23900 22704
rect 17316 22584 17368 22636
rect 22928 22584 22980 22636
rect 16672 22559 16724 22568
rect 14740 22448 14792 22500
rect 16304 22380 16356 22432
rect 16672 22525 16681 22559
rect 16681 22525 16715 22559
rect 16715 22525 16724 22559
rect 16672 22516 16724 22525
rect 20444 22516 20496 22568
rect 21640 22559 21692 22568
rect 21640 22525 21649 22559
rect 21649 22525 21683 22559
rect 21683 22525 21692 22559
rect 21640 22516 21692 22525
rect 23848 22559 23900 22568
rect 23848 22525 23857 22559
rect 23857 22525 23891 22559
rect 23891 22525 23900 22559
rect 23848 22516 23900 22525
rect 23940 22516 23992 22568
rect 24216 22559 24268 22568
rect 24216 22525 24225 22559
rect 24225 22525 24259 22559
rect 24259 22525 24268 22559
rect 24216 22516 24268 22525
rect 24952 22516 25004 22568
rect 25964 22584 26016 22636
rect 21364 22491 21416 22500
rect 21364 22457 21373 22491
rect 21373 22457 21407 22491
rect 21407 22457 21416 22491
rect 21364 22448 21416 22457
rect 21456 22448 21508 22500
rect 24676 22448 24728 22500
rect 25504 22516 25556 22568
rect 26240 22584 26292 22636
rect 28080 22720 28132 22772
rect 18052 22380 18104 22432
rect 20720 22380 20772 22432
rect 27436 22448 27488 22500
rect 21732 22423 21784 22432
rect 21732 22389 21741 22423
rect 21741 22389 21775 22423
rect 21775 22389 21784 22423
rect 21732 22380 21784 22389
rect 23940 22423 23992 22432
rect 23940 22389 23949 22423
rect 23949 22389 23983 22423
rect 23983 22389 23992 22423
rect 23940 22380 23992 22389
rect 24952 22380 25004 22432
rect 25504 22380 25556 22432
rect 10246 22278 10298 22330
rect 10310 22278 10362 22330
rect 10374 22278 10426 22330
rect 10438 22278 10490 22330
rect 19510 22278 19562 22330
rect 19574 22278 19626 22330
rect 19638 22278 19690 22330
rect 19702 22278 19754 22330
rect 2044 22219 2096 22228
rect 2044 22185 2053 22219
rect 2053 22185 2087 22219
rect 2087 22185 2096 22219
rect 2044 22176 2096 22185
rect 2780 22176 2832 22228
rect 2136 22108 2188 22160
rect 4068 22108 4120 22160
rect 4712 22151 4764 22160
rect 4712 22117 4721 22151
rect 4721 22117 4755 22151
rect 4755 22117 4764 22151
rect 4712 22108 4764 22117
rect 5080 22176 5132 22228
rect 5632 22176 5684 22228
rect 8116 22219 8168 22228
rect 8116 22185 8125 22219
rect 8125 22185 8159 22219
rect 8159 22185 8168 22219
rect 8116 22176 8168 22185
rect 8576 22219 8628 22228
rect 8576 22185 8585 22219
rect 8585 22185 8619 22219
rect 8619 22185 8628 22219
rect 8576 22176 8628 22185
rect 9772 22176 9824 22228
rect 10600 22176 10652 22228
rect 10876 22219 10928 22228
rect 10876 22185 10885 22219
rect 10885 22185 10919 22219
rect 10919 22185 10928 22219
rect 10876 22176 10928 22185
rect 11428 22176 11480 22228
rect 14648 22219 14700 22228
rect 1584 22083 1636 22092
rect 1584 22049 1593 22083
rect 1593 22049 1627 22083
rect 1627 22049 1636 22083
rect 1584 22040 1636 22049
rect 2320 22040 2372 22092
rect 2228 21972 2280 22024
rect 2780 22040 2832 22092
rect 5172 22083 5224 22092
rect 5172 22049 5181 22083
rect 5181 22049 5215 22083
rect 5215 22049 5224 22083
rect 5172 22040 5224 22049
rect 5908 22108 5960 22160
rect 6644 22108 6696 22160
rect 8484 22151 8536 22160
rect 8484 22117 8493 22151
rect 8493 22117 8527 22151
rect 8527 22117 8536 22151
rect 8484 22108 8536 22117
rect 5540 21972 5592 22024
rect 7104 22083 7156 22092
rect 7104 22049 7113 22083
rect 7113 22049 7147 22083
rect 7147 22049 7156 22083
rect 9680 22108 9732 22160
rect 10968 22108 11020 22160
rect 7104 22040 7156 22049
rect 8668 21972 8720 22024
rect 9404 21972 9456 22024
rect 5632 21904 5684 21956
rect 6000 21904 6052 21956
rect 6276 21904 6328 21956
rect 10232 22040 10284 22092
rect 11060 21972 11112 22024
rect 11612 22040 11664 22092
rect 12072 22040 12124 22092
rect 12256 22083 12308 22092
rect 12256 22049 12265 22083
rect 12265 22049 12299 22083
rect 12299 22049 12308 22083
rect 12256 22040 12308 22049
rect 14648 22185 14657 22219
rect 14657 22185 14691 22219
rect 14691 22185 14700 22219
rect 14648 22176 14700 22185
rect 16672 22176 16724 22228
rect 17224 22176 17276 22228
rect 24032 22219 24084 22228
rect 24032 22185 24041 22219
rect 24041 22185 24075 22219
rect 24075 22185 24084 22219
rect 24032 22176 24084 22185
rect 24216 22176 24268 22228
rect 15476 22108 15528 22160
rect 14188 22040 14240 22092
rect 16117 22083 16169 22092
rect 16117 22049 16144 22083
rect 16144 22049 16169 22083
rect 13544 22015 13596 22024
rect 13544 21981 13553 22015
rect 13553 21981 13587 22015
rect 13587 21981 13596 22015
rect 13544 21972 13596 21981
rect 1492 21836 1544 21888
rect 2412 21836 2464 21888
rect 3700 21836 3752 21888
rect 11060 21836 11112 21888
rect 11612 21836 11664 21888
rect 12164 21836 12216 21888
rect 12348 21836 12400 21888
rect 12716 21836 12768 21888
rect 15200 21836 15252 21888
rect 15568 21836 15620 21888
rect 16117 22040 16169 22049
rect 16304 21904 16356 21956
rect 17868 22040 17920 22092
rect 18052 22040 18104 22092
rect 19064 22040 19116 22092
rect 20720 22083 20772 22092
rect 20720 22049 20729 22083
rect 20729 22049 20763 22083
rect 20763 22049 20772 22083
rect 20720 22040 20772 22049
rect 20812 22040 20864 22092
rect 21732 22108 21784 22160
rect 22468 22108 22520 22160
rect 21640 22083 21692 22092
rect 20996 21972 21048 22024
rect 21640 22049 21649 22083
rect 21649 22049 21683 22083
rect 21683 22049 21692 22083
rect 21640 22040 21692 22049
rect 22744 22151 22796 22160
rect 22744 22117 22753 22151
rect 22753 22117 22787 22151
rect 22787 22117 22796 22151
rect 23112 22151 23164 22160
rect 22744 22108 22796 22117
rect 23112 22117 23121 22151
rect 23121 22117 23155 22151
rect 23155 22117 23164 22151
rect 23112 22108 23164 22117
rect 23296 22108 23348 22160
rect 23572 22108 23624 22160
rect 25596 22176 25648 22228
rect 26608 22176 26660 22228
rect 26700 22176 26752 22228
rect 26240 22108 26292 22160
rect 26424 22151 26476 22160
rect 26424 22117 26433 22151
rect 26433 22117 26467 22151
rect 26467 22117 26476 22151
rect 26424 22108 26476 22117
rect 24860 22040 24912 22092
rect 25688 22083 25740 22092
rect 25688 22049 25697 22083
rect 25697 22049 25731 22083
rect 25731 22049 25740 22083
rect 25688 22040 25740 22049
rect 26884 22040 26936 22092
rect 21916 21972 21968 22024
rect 22560 21972 22612 22024
rect 24952 21972 25004 22024
rect 27160 21972 27212 22024
rect 16672 21904 16724 21956
rect 17684 21904 17736 21956
rect 26516 21904 26568 21956
rect 20904 21836 20956 21888
rect 5614 21734 5666 21786
rect 5678 21734 5730 21786
rect 5742 21734 5794 21786
rect 5806 21734 5858 21786
rect 14878 21734 14930 21786
rect 14942 21734 14994 21786
rect 15006 21734 15058 21786
rect 15070 21734 15122 21786
rect 24142 21734 24194 21786
rect 24206 21734 24258 21786
rect 24270 21734 24322 21786
rect 24334 21734 24386 21786
rect 4988 21632 5040 21684
rect 6828 21632 6880 21684
rect 7104 21632 7156 21684
rect 10232 21675 10284 21684
rect 10232 21641 10241 21675
rect 10241 21641 10275 21675
rect 10275 21641 10284 21675
rect 10232 21632 10284 21641
rect 11060 21632 11112 21684
rect 12164 21632 12216 21684
rect 12532 21675 12584 21684
rect 12532 21641 12541 21675
rect 12541 21641 12575 21675
rect 12575 21641 12584 21675
rect 12532 21632 12584 21641
rect 13544 21632 13596 21684
rect 13636 21632 13688 21684
rect 14280 21632 14332 21684
rect 15292 21632 15344 21684
rect 15936 21632 15988 21684
rect 19064 21675 19116 21684
rect 19064 21641 19073 21675
rect 19073 21641 19107 21675
rect 19107 21641 19116 21675
rect 19064 21632 19116 21641
rect 19800 21632 19852 21684
rect 20168 21632 20220 21684
rect 21732 21632 21784 21684
rect 23572 21632 23624 21684
rect 26608 21675 26660 21684
rect 26608 21641 26617 21675
rect 26617 21641 26651 21675
rect 26651 21641 26660 21675
rect 26608 21632 26660 21641
rect 27436 21675 27488 21684
rect 27436 21641 27445 21675
rect 27445 21641 27479 21675
rect 27479 21641 27488 21675
rect 27436 21632 27488 21641
rect 1400 21496 1452 21548
rect 1676 21428 1728 21480
rect 6368 21564 6420 21616
rect 4252 21496 4304 21548
rect 5816 21496 5868 21548
rect 6276 21428 6328 21480
rect 1768 21360 1820 21412
rect 2044 21360 2096 21412
rect 2136 21360 2188 21412
rect 3332 21360 3384 21412
rect 4804 21360 4856 21412
rect 6644 21496 6696 21548
rect 9864 21564 9916 21616
rect 10600 21564 10652 21616
rect 10784 21496 10836 21548
rect 11060 21496 11112 21548
rect 11520 21496 11572 21548
rect 6460 21428 6512 21480
rect 8668 21428 8720 21480
rect 11244 21428 11296 21480
rect 12072 21428 12124 21480
rect 12256 21471 12308 21480
rect 12256 21437 12265 21471
rect 12265 21437 12299 21471
rect 12299 21437 12308 21471
rect 12256 21428 12308 21437
rect 13728 21564 13780 21616
rect 13820 21564 13872 21616
rect 14648 21496 14700 21548
rect 13360 21471 13412 21480
rect 13360 21437 13369 21471
rect 13369 21437 13403 21471
rect 13403 21437 13412 21471
rect 13360 21428 13412 21437
rect 17040 21564 17092 21616
rect 16120 21496 16172 21548
rect 16580 21496 16632 21548
rect 19248 21496 19300 21548
rect 19340 21496 19392 21548
rect 20076 21564 20128 21616
rect 27988 21539 28040 21548
rect 15936 21471 15988 21480
rect 2688 21335 2740 21344
rect 2688 21301 2697 21335
rect 2697 21301 2731 21335
rect 2731 21301 2740 21335
rect 2688 21292 2740 21301
rect 4160 21292 4212 21344
rect 11796 21292 11848 21344
rect 12900 21292 12952 21344
rect 13728 21360 13780 21412
rect 15200 21360 15252 21412
rect 15476 21360 15528 21412
rect 15936 21437 15945 21471
rect 15945 21437 15979 21471
rect 15979 21437 15988 21471
rect 15936 21428 15988 21437
rect 20996 21428 21048 21480
rect 22376 21471 22428 21480
rect 22376 21437 22385 21471
rect 22385 21437 22419 21471
rect 22419 21437 22428 21471
rect 22376 21428 22428 21437
rect 27988 21505 27997 21539
rect 27997 21505 28031 21539
rect 28031 21505 28040 21539
rect 27988 21496 28040 21505
rect 24860 21428 24912 21480
rect 25504 21471 25556 21480
rect 25504 21437 25538 21471
rect 25538 21437 25556 21471
rect 27804 21471 27856 21480
rect 20076 21360 20128 21412
rect 20536 21403 20588 21412
rect 20536 21369 20545 21403
rect 20545 21369 20579 21403
rect 20579 21369 20588 21403
rect 20904 21403 20956 21412
rect 20536 21360 20588 21369
rect 20904 21369 20913 21403
rect 20913 21369 20947 21403
rect 20947 21369 20956 21403
rect 20904 21360 20956 21369
rect 22284 21360 22336 21412
rect 22560 21360 22612 21412
rect 23296 21360 23348 21412
rect 25504 21428 25556 21437
rect 27804 21437 27813 21471
rect 27813 21437 27847 21471
rect 27847 21437 27856 21471
rect 27804 21428 27856 21437
rect 28080 21428 28132 21480
rect 26056 21360 26108 21412
rect 14096 21292 14148 21344
rect 16396 21292 16448 21344
rect 18236 21292 18288 21344
rect 19064 21292 19116 21344
rect 20260 21292 20312 21344
rect 22744 21292 22796 21344
rect 10246 21190 10298 21242
rect 10310 21190 10362 21242
rect 10374 21190 10426 21242
rect 10438 21190 10490 21242
rect 19510 21190 19562 21242
rect 19574 21190 19626 21242
rect 19638 21190 19690 21242
rect 19702 21190 19754 21242
rect 3700 21131 3752 21140
rect 3700 21097 3709 21131
rect 3709 21097 3743 21131
rect 3743 21097 3752 21131
rect 3700 21088 3752 21097
rect 5356 21088 5408 21140
rect 6920 21088 6972 21140
rect 9680 21088 9732 21140
rect 10784 21088 10836 21140
rect 5908 21020 5960 21072
rect 12256 21088 12308 21140
rect 1676 20995 1728 21004
rect 1676 20961 1685 20995
rect 1685 20961 1719 20995
rect 1719 20961 1728 20995
rect 1676 20952 1728 20961
rect 3240 20952 3292 21004
rect 3516 20952 3568 21004
rect 6828 20995 6880 21004
rect 2964 20816 3016 20868
rect 6828 20961 6837 20995
rect 6837 20961 6871 20995
rect 6871 20961 6880 20995
rect 6828 20952 6880 20961
rect 7104 20995 7156 21004
rect 7104 20961 7113 20995
rect 7113 20961 7147 20995
rect 7147 20961 7156 20995
rect 7104 20952 7156 20961
rect 7288 20995 7340 21004
rect 7288 20961 7297 20995
rect 7297 20961 7331 20995
rect 7331 20961 7340 20995
rect 7288 20952 7340 20961
rect 9680 20995 9732 21004
rect 3884 20927 3936 20936
rect 3884 20893 3893 20927
rect 3893 20893 3927 20927
rect 3927 20893 3936 20927
rect 3884 20884 3936 20893
rect 4804 20816 4856 20868
rect 9680 20961 9689 20995
rect 9689 20961 9723 20995
rect 9723 20961 9732 20995
rect 9680 20952 9732 20961
rect 11152 21020 11204 21072
rect 11520 21020 11572 21072
rect 12072 21020 12124 21072
rect 9956 20927 10008 20936
rect 9956 20893 9965 20927
rect 9965 20893 9999 20927
rect 9999 20893 10008 20927
rect 9956 20884 10008 20893
rect 10968 20995 11020 21004
rect 10968 20961 10977 20995
rect 10977 20961 11011 20995
rect 11011 20961 11020 20995
rect 10968 20952 11020 20961
rect 12164 20952 12216 21004
rect 12716 20995 12768 21004
rect 10968 20816 11020 20868
rect 12716 20961 12725 20995
rect 12725 20961 12759 20995
rect 12759 20961 12768 20995
rect 12716 20952 12768 20961
rect 15936 21088 15988 21140
rect 18236 21131 18288 21140
rect 18236 21097 18245 21131
rect 18245 21097 18279 21131
rect 18279 21097 18288 21131
rect 18236 21088 18288 21097
rect 19800 21088 19852 21140
rect 20536 21088 20588 21140
rect 20720 21088 20772 21140
rect 21180 21088 21232 21140
rect 22560 21131 22612 21140
rect 22560 21097 22569 21131
rect 22569 21097 22603 21131
rect 22603 21097 22612 21131
rect 22560 21088 22612 21097
rect 22928 21088 22980 21140
rect 23572 21088 23624 21140
rect 24032 21088 24084 21140
rect 24492 21131 24544 21140
rect 24492 21097 24501 21131
rect 24501 21097 24535 21131
rect 24535 21097 24544 21131
rect 24492 21088 24544 21097
rect 24860 21088 24912 21140
rect 14740 21020 14792 21072
rect 17960 21063 18012 21072
rect 12900 20884 12952 20936
rect 13728 20995 13780 21004
rect 13728 20961 13737 20995
rect 13737 20961 13771 20995
rect 13771 20961 13780 20995
rect 13728 20952 13780 20961
rect 14280 20952 14332 21004
rect 17960 21029 17969 21063
rect 17969 21029 18003 21063
rect 18003 21029 18012 21063
rect 17960 21020 18012 21029
rect 18052 21020 18104 21072
rect 18788 21020 18840 21072
rect 19064 21020 19116 21072
rect 20996 21020 21048 21072
rect 21732 21020 21784 21072
rect 15476 20952 15528 21004
rect 15568 20952 15620 21004
rect 18236 20995 18288 21004
rect 18236 20961 18245 20995
rect 18245 20961 18279 20995
rect 18279 20961 18288 20995
rect 18236 20952 18288 20961
rect 20904 20952 20956 21004
rect 22928 20995 22980 21004
rect 22928 20961 22937 20995
rect 22937 20961 22971 20995
rect 22971 20961 22980 20995
rect 22928 20952 22980 20961
rect 2136 20748 2188 20800
rect 8484 20748 8536 20800
rect 8944 20748 8996 20800
rect 9772 20791 9824 20800
rect 9772 20757 9781 20791
rect 9781 20757 9815 20791
rect 9815 20757 9824 20791
rect 9772 20748 9824 20757
rect 10048 20748 10100 20800
rect 12256 20748 12308 20800
rect 12532 20816 12584 20868
rect 12716 20816 12768 20868
rect 14556 20816 14608 20868
rect 15568 20816 15620 20868
rect 18788 20884 18840 20936
rect 20812 20927 20864 20936
rect 20812 20893 20821 20927
rect 20821 20893 20855 20927
rect 20855 20893 20864 20927
rect 20812 20884 20864 20893
rect 22100 20884 22152 20936
rect 23020 20884 23072 20936
rect 16120 20816 16172 20868
rect 23848 21020 23900 21072
rect 25964 21020 26016 21072
rect 23940 20952 23992 21004
rect 25412 20995 25464 21004
rect 23572 20884 23624 20936
rect 25412 20961 25421 20995
rect 25421 20961 25455 20995
rect 25455 20961 25464 20995
rect 25412 20952 25464 20961
rect 26884 20995 26936 21004
rect 26884 20961 26893 20995
rect 26893 20961 26927 20995
rect 26927 20961 26936 20995
rect 26884 20952 26936 20961
rect 12900 20748 12952 20800
rect 13912 20791 13964 20800
rect 13912 20757 13921 20791
rect 13921 20757 13955 20791
rect 13955 20757 13964 20791
rect 13912 20748 13964 20757
rect 14096 20748 14148 20800
rect 20260 20748 20312 20800
rect 24768 20816 24820 20868
rect 22468 20748 22520 20800
rect 28080 20791 28132 20800
rect 28080 20757 28089 20791
rect 28089 20757 28123 20791
rect 28123 20757 28132 20791
rect 28080 20748 28132 20757
rect 5614 20646 5666 20698
rect 5678 20646 5730 20698
rect 5742 20646 5794 20698
rect 5806 20646 5858 20698
rect 14878 20646 14930 20698
rect 14942 20646 14994 20698
rect 15006 20646 15058 20698
rect 15070 20646 15122 20698
rect 24142 20646 24194 20698
rect 24206 20646 24258 20698
rect 24270 20646 24322 20698
rect 24334 20646 24386 20698
rect 2688 20544 2740 20596
rect 2964 20587 3016 20596
rect 2964 20553 2973 20587
rect 2973 20553 3007 20587
rect 3007 20553 3016 20587
rect 2964 20544 3016 20553
rect 4620 20544 4672 20596
rect 11612 20544 11664 20596
rect 14188 20544 14240 20596
rect 20444 20544 20496 20596
rect 12532 20476 12584 20528
rect 13360 20476 13412 20528
rect 13912 20476 13964 20528
rect 1952 20383 2004 20392
rect 1952 20349 1961 20383
rect 1961 20349 1995 20383
rect 1995 20349 2004 20383
rect 1952 20340 2004 20349
rect 2964 20408 3016 20460
rect 3792 20408 3844 20460
rect 7656 20451 7708 20460
rect 7656 20417 7665 20451
rect 7665 20417 7699 20451
rect 7699 20417 7708 20451
rect 7656 20408 7708 20417
rect 9864 20408 9916 20460
rect 16028 20476 16080 20528
rect 22928 20544 22980 20596
rect 24492 20544 24544 20596
rect 26148 20544 26200 20596
rect 27528 20544 27580 20596
rect 2228 20272 2280 20324
rect 5080 20340 5132 20392
rect 6092 20383 6144 20392
rect 6092 20349 6101 20383
rect 6101 20349 6135 20383
rect 6135 20349 6144 20383
rect 6092 20340 6144 20349
rect 6368 20383 6420 20392
rect 6368 20349 6377 20383
rect 6377 20349 6411 20383
rect 6411 20349 6420 20383
rect 6368 20340 6420 20349
rect 7472 20340 7524 20392
rect 8484 20340 8536 20392
rect 10048 20340 10100 20392
rect 12348 20340 12400 20392
rect 12716 20340 12768 20392
rect 12900 20340 12952 20392
rect 13360 20340 13412 20392
rect 15016 20383 15068 20392
rect 15016 20349 15025 20383
rect 15025 20349 15059 20383
rect 15059 20349 15068 20383
rect 15016 20340 15068 20349
rect 15200 20383 15252 20392
rect 15200 20349 15209 20383
rect 15209 20349 15243 20383
rect 15243 20349 15252 20383
rect 15752 20408 15804 20460
rect 21364 20408 21416 20460
rect 15200 20340 15252 20349
rect 16028 20340 16080 20392
rect 16672 20383 16724 20392
rect 16672 20349 16681 20383
rect 16681 20349 16715 20383
rect 16715 20349 16724 20383
rect 16672 20340 16724 20349
rect 19064 20340 19116 20392
rect 20996 20383 21048 20392
rect 20996 20349 21005 20383
rect 21005 20349 21039 20383
rect 21039 20349 21048 20383
rect 20996 20340 21048 20349
rect 21640 20383 21692 20392
rect 21640 20349 21649 20383
rect 21649 20349 21683 20383
rect 21683 20349 21692 20383
rect 21640 20340 21692 20349
rect 22376 20476 22428 20528
rect 23296 20476 23348 20528
rect 22284 20408 22336 20460
rect 5172 20272 5224 20324
rect 16580 20315 16632 20324
rect 16580 20281 16589 20315
rect 16589 20281 16623 20315
rect 16623 20281 16632 20315
rect 16580 20272 16632 20281
rect 20076 20272 20128 20324
rect 25964 20315 26016 20324
rect 7472 20204 7524 20256
rect 12164 20247 12216 20256
rect 12164 20213 12173 20247
rect 12173 20213 12207 20247
rect 12207 20213 12216 20247
rect 12164 20204 12216 20213
rect 14740 20247 14792 20256
rect 14740 20213 14749 20247
rect 14749 20213 14783 20247
rect 14783 20213 14792 20247
rect 14740 20204 14792 20213
rect 16120 20204 16172 20256
rect 17408 20247 17460 20256
rect 17408 20213 17417 20247
rect 17417 20213 17451 20247
rect 17451 20213 17460 20247
rect 17408 20204 17460 20213
rect 17960 20204 18012 20256
rect 25964 20281 25973 20315
rect 25973 20281 26007 20315
rect 26007 20281 26016 20315
rect 25964 20272 26016 20281
rect 26240 20272 26292 20324
rect 26700 20315 26752 20324
rect 26700 20281 26709 20315
rect 26709 20281 26743 20315
rect 26743 20281 26752 20315
rect 26700 20272 26752 20281
rect 28172 20315 28224 20324
rect 28172 20281 28181 20315
rect 28181 20281 28215 20315
rect 28215 20281 28224 20315
rect 28172 20272 28224 20281
rect 28080 20204 28132 20256
rect 10246 20102 10298 20154
rect 10310 20102 10362 20154
rect 10374 20102 10426 20154
rect 10438 20102 10490 20154
rect 19510 20102 19562 20154
rect 19574 20102 19626 20154
rect 19638 20102 19690 20154
rect 19702 20102 19754 20154
rect 4160 20000 4212 20052
rect 4344 20000 4396 20052
rect 9956 20000 10008 20052
rect 20076 20000 20128 20052
rect 4712 19932 4764 19984
rect 1860 19907 1912 19916
rect 1860 19873 1869 19907
rect 1869 19873 1903 19907
rect 1903 19873 1912 19907
rect 1860 19864 1912 19873
rect 2780 19864 2832 19916
rect 3148 19907 3200 19916
rect 3148 19873 3157 19907
rect 3157 19873 3191 19907
rect 3191 19873 3200 19907
rect 3148 19864 3200 19873
rect 7380 19932 7432 19984
rect 8300 19932 8352 19984
rect 8668 19932 8720 19984
rect 9036 19932 9088 19984
rect 9496 19932 9548 19984
rect 9864 19932 9916 19984
rect 7472 19907 7524 19916
rect 7472 19873 7481 19907
rect 7481 19873 7515 19907
rect 7515 19873 7524 19907
rect 7472 19864 7524 19873
rect 8116 19907 8168 19916
rect 8116 19873 8125 19907
rect 8125 19873 8159 19907
rect 8159 19873 8168 19907
rect 8116 19864 8168 19873
rect 9128 19907 9180 19916
rect 9128 19873 9137 19907
rect 9137 19873 9171 19907
rect 9171 19873 9180 19907
rect 9128 19864 9180 19873
rect 9220 19864 9272 19916
rect 9680 19864 9732 19916
rect 11244 19932 11296 19984
rect 15016 19932 15068 19984
rect 16120 19932 16172 19984
rect 16580 19932 16632 19984
rect 17592 19907 17644 19916
rect 3884 19796 3936 19848
rect 17592 19873 17601 19907
rect 17601 19873 17635 19907
rect 17635 19873 17644 19907
rect 17592 19864 17644 19873
rect 18328 19864 18380 19916
rect 25228 19864 25280 19916
rect 25688 19907 25740 19916
rect 25688 19873 25697 19907
rect 25697 19873 25731 19907
rect 25731 19873 25740 19907
rect 25688 19864 25740 19873
rect 26516 19907 26568 19916
rect 26516 19873 26525 19907
rect 26525 19873 26559 19907
rect 26559 19873 26568 19907
rect 26516 19864 26568 19873
rect 26792 19864 26844 19916
rect 2412 19728 2464 19780
rect 3332 19771 3384 19780
rect 3332 19737 3341 19771
rect 3341 19737 3375 19771
rect 3375 19737 3384 19771
rect 3332 19728 3384 19737
rect 6368 19728 6420 19780
rect 11152 19796 11204 19848
rect 12348 19796 12400 19848
rect 12532 19796 12584 19848
rect 16580 19796 16632 19848
rect 17684 19839 17736 19848
rect 17408 19728 17460 19780
rect 17684 19805 17693 19839
rect 17693 19805 17727 19839
rect 17727 19805 17736 19839
rect 17684 19796 17736 19805
rect 17868 19796 17920 19848
rect 20536 19796 20588 19848
rect 23388 19796 23440 19848
rect 25872 19771 25924 19780
rect 25872 19737 25881 19771
rect 25881 19737 25915 19771
rect 25915 19737 25924 19771
rect 25872 19728 25924 19737
rect 26792 19728 26844 19780
rect 27160 19728 27212 19780
rect 28172 19771 28224 19780
rect 28172 19737 28181 19771
rect 28181 19737 28215 19771
rect 28215 19737 28224 19771
rect 28172 19728 28224 19737
rect 4160 19703 4212 19712
rect 4160 19669 4169 19703
rect 4169 19669 4203 19703
rect 4203 19669 4212 19703
rect 4160 19660 4212 19669
rect 6184 19660 6236 19712
rect 11244 19660 11296 19712
rect 11612 19660 11664 19712
rect 17868 19660 17920 19712
rect 19984 19703 20036 19712
rect 19984 19669 19993 19703
rect 19993 19669 20027 19703
rect 20027 19669 20036 19703
rect 19984 19660 20036 19669
rect 25412 19660 25464 19712
rect 25780 19660 25832 19712
rect 27804 19660 27856 19712
rect 5614 19558 5666 19610
rect 5678 19558 5730 19610
rect 5742 19558 5794 19610
rect 5806 19558 5858 19610
rect 14878 19558 14930 19610
rect 14942 19558 14994 19610
rect 15006 19558 15058 19610
rect 15070 19558 15122 19610
rect 24142 19558 24194 19610
rect 24206 19558 24258 19610
rect 24270 19558 24322 19610
rect 24334 19558 24386 19610
rect 7656 19456 7708 19508
rect 9496 19499 9548 19508
rect 9496 19465 9505 19499
rect 9505 19465 9539 19499
rect 9539 19465 9548 19499
rect 9496 19456 9548 19465
rect 10968 19456 11020 19508
rect 13360 19456 13412 19508
rect 16120 19499 16172 19508
rect 16120 19465 16129 19499
rect 16129 19465 16163 19499
rect 16163 19465 16172 19499
rect 16120 19456 16172 19465
rect 17040 19456 17092 19508
rect 21364 19456 21416 19508
rect 28080 19456 28132 19508
rect 6092 19388 6144 19440
rect 14740 19388 14792 19440
rect 4160 19320 4212 19372
rect 4804 19363 4856 19372
rect 4804 19329 4813 19363
rect 4813 19329 4847 19363
rect 4847 19329 4856 19363
rect 4804 19320 4856 19329
rect 6368 19320 6420 19372
rect 10140 19363 10192 19372
rect 2872 19252 2924 19304
rect 2964 19252 3016 19304
rect 4252 19252 4304 19304
rect 5172 19252 5224 19304
rect 7012 19252 7064 19304
rect 7104 19252 7156 19304
rect 7380 19295 7432 19304
rect 7380 19261 7389 19295
rect 7389 19261 7423 19295
rect 7423 19261 7432 19295
rect 7380 19252 7432 19261
rect 7472 19252 7524 19304
rect 10140 19329 10149 19363
rect 10149 19329 10183 19363
rect 10183 19329 10192 19363
rect 10140 19320 10192 19329
rect 21732 19388 21784 19440
rect 16580 19320 16632 19372
rect 1860 19227 1912 19236
rect 1860 19193 1869 19227
rect 1869 19193 1903 19227
rect 1903 19193 1912 19227
rect 1860 19184 1912 19193
rect 1584 19116 1636 19168
rect 2688 19159 2740 19168
rect 2688 19125 2697 19159
rect 2697 19125 2731 19159
rect 2731 19125 2740 19159
rect 2688 19116 2740 19125
rect 4988 19184 5040 19236
rect 5264 19184 5316 19236
rect 4068 19116 4120 19168
rect 4252 19159 4304 19168
rect 4252 19125 4261 19159
rect 4261 19125 4295 19159
rect 4295 19125 4304 19159
rect 4252 19116 4304 19125
rect 4528 19116 4580 19168
rect 6920 19116 6972 19168
rect 10968 19184 11020 19236
rect 13360 19252 13412 19304
rect 14832 19184 14884 19236
rect 9864 19159 9916 19168
rect 9864 19125 9873 19159
rect 9873 19125 9907 19159
rect 9907 19125 9916 19159
rect 9864 19116 9916 19125
rect 9956 19159 10008 19168
rect 9956 19125 9965 19159
rect 9965 19125 9999 19159
rect 9999 19125 10008 19159
rect 9956 19116 10008 19125
rect 10876 19116 10928 19168
rect 11612 19116 11664 19168
rect 16396 19184 16448 19236
rect 17224 19252 17276 19304
rect 18696 19252 18748 19304
rect 19340 19252 19392 19304
rect 21548 19320 21600 19372
rect 21916 19320 21968 19372
rect 20536 19252 20588 19304
rect 20720 19252 20772 19304
rect 19064 19116 19116 19168
rect 20628 19116 20680 19168
rect 20904 19116 20956 19168
rect 23480 19252 23532 19304
rect 25412 19388 25464 19440
rect 26240 19388 26292 19440
rect 25780 19363 25832 19372
rect 23940 19295 23992 19304
rect 23940 19261 23949 19295
rect 23949 19261 23983 19295
rect 23983 19261 23992 19295
rect 23940 19252 23992 19261
rect 24032 19252 24084 19304
rect 25780 19329 25789 19363
rect 25789 19329 25823 19363
rect 25823 19329 25832 19363
rect 25780 19320 25832 19329
rect 26056 19252 26108 19304
rect 23848 19184 23900 19236
rect 21180 19159 21232 19168
rect 21180 19125 21189 19159
rect 21189 19125 21223 19159
rect 21223 19125 21232 19159
rect 21180 19116 21232 19125
rect 21548 19116 21600 19168
rect 23020 19116 23072 19168
rect 26332 19184 26384 19236
rect 27436 19184 27488 19236
rect 25320 19116 25372 19168
rect 25688 19159 25740 19168
rect 25688 19125 25697 19159
rect 25697 19125 25731 19159
rect 25731 19125 25740 19159
rect 25688 19116 25740 19125
rect 26148 19116 26200 19168
rect 10246 19014 10298 19066
rect 10310 19014 10362 19066
rect 10374 19014 10426 19066
rect 10438 19014 10490 19066
rect 19510 19014 19562 19066
rect 19574 19014 19626 19066
rect 19638 19014 19690 19066
rect 19702 19014 19754 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 2596 18912 2648 18964
rect 2780 18912 2832 18964
rect 1768 18844 1820 18896
rect 2044 18776 2096 18828
rect 2412 18776 2464 18828
rect 4528 18844 4580 18896
rect 5172 18844 5224 18896
rect 5540 18912 5592 18964
rect 6092 18912 6144 18964
rect 6644 18912 6696 18964
rect 3424 18819 3476 18828
rect 3424 18785 3433 18819
rect 3433 18785 3467 18819
rect 3467 18785 3476 18819
rect 3424 18776 3476 18785
rect 1400 18708 1452 18760
rect 5172 18708 5224 18760
rect 9128 18912 9180 18964
rect 9772 18912 9824 18964
rect 9956 18912 10008 18964
rect 10876 18955 10928 18964
rect 10876 18921 10885 18955
rect 10885 18921 10919 18955
rect 10919 18921 10928 18955
rect 10876 18912 10928 18921
rect 12532 18912 12584 18964
rect 13912 18912 13964 18964
rect 14096 18912 14148 18964
rect 14648 18912 14700 18964
rect 14832 18912 14884 18964
rect 8944 18819 8996 18828
rect 8944 18785 8953 18819
rect 8953 18785 8987 18819
rect 8987 18785 8996 18819
rect 8944 18776 8996 18785
rect 11796 18844 11848 18896
rect 12348 18844 12400 18896
rect 14188 18844 14240 18896
rect 9496 18776 9548 18828
rect 12072 18776 12124 18828
rect 12164 18776 12216 18828
rect 13912 18776 13964 18828
rect 15844 18776 15896 18828
rect 17960 18844 18012 18896
rect 18052 18844 18104 18896
rect 19064 18844 19116 18896
rect 17592 18776 17644 18828
rect 19524 18819 19576 18828
rect 9036 18708 9088 18760
rect 9220 18751 9272 18760
rect 9220 18717 9229 18751
rect 9229 18717 9263 18751
rect 9263 18717 9272 18751
rect 9220 18708 9272 18717
rect 9404 18708 9456 18760
rect 11060 18708 11112 18760
rect 11244 18708 11296 18760
rect 11704 18708 11756 18760
rect 12716 18708 12768 18760
rect 14280 18708 14332 18760
rect 11888 18640 11940 18692
rect 12164 18640 12216 18692
rect 13268 18640 13320 18692
rect 14648 18640 14700 18692
rect 15568 18708 15620 18760
rect 17408 18708 17460 18760
rect 17684 18708 17736 18760
rect 15844 18640 15896 18692
rect 19524 18785 19533 18819
rect 19533 18785 19567 18819
rect 19567 18785 19576 18819
rect 19524 18776 19576 18785
rect 19616 18819 19668 18828
rect 19616 18785 19625 18819
rect 19625 18785 19659 18819
rect 19659 18785 19668 18819
rect 19984 18819 20036 18828
rect 19616 18776 19668 18785
rect 19984 18785 19993 18819
rect 19993 18785 20027 18819
rect 20027 18785 20036 18819
rect 19984 18776 20036 18785
rect 18696 18708 18748 18760
rect 20904 18640 20956 18692
rect 6000 18572 6052 18624
rect 6276 18572 6328 18624
rect 8576 18615 8628 18624
rect 8576 18581 8585 18615
rect 8585 18581 8619 18615
rect 8619 18581 8628 18615
rect 8576 18572 8628 18581
rect 11704 18572 11756 18624
rect 15200 18572 15252 18624
rect 16580 18572 16632 18624
rect 19064 18572 19116 18624
rect 21548 18844 21600 18896
rect 22744 18887 22796 18896
rect 21640 18819 21692 18828
rect 21640 18785 21649 18819
rect 21649 18785 21683 18819
rect 21683 18785 21692 18819
rect 21640 18776 21692 18785
rect 22744 18853 22753 18887
rect 22753 18853 22787 18887
rect 22787 18853 22796 18887
rect 22744 18844 22796 18853
rect 23848 18887 23900 18896
rect 23848 18853 23857 18887
rect 23857 18853 23891 18887
rect 23891 18853 23900 18887
rect 23848 18844 23900 18853
rect 23940 18844 23992 18896
rect 25412 18887 25464 18896
rect 25412 18853 25421 18887
rect 25421 18853 25455 18887
rect 25455 18853 25464 18887
rect 25412 18844 25464 18853
rect 25688 18887 25740 18896
rect 23020 18819 23072 18828
rect 21272 18640 21324 18692
rect 21364 18640 21416 18692
rect 21732 18640 21784 18692
rect 23020 18785 23029 18819
rect 23029 18785 23063 18819
rect 23063 18785 23072 18819
rect 23020 18776 23072 18785
rect 23112 18819 23164 18828
rect 23112 18785 23121 18819
rect 23121 18785 23155 18819
rect 23155 18785 23164 18819
rect 23480 18819 23532 18828
rect 23112 18776 23164 18785
rect 23480 18785 23489 18819
rect 23489 18785 23523 18819
rect 23523 18785 23532 18819
rect 23480 18776 23532 18785
rect 24124 18776 24176 18828
rect 25688 18853 25697 18887
rect 25697 18853 25731 18887
rect 25731 18853 25740 18887
rect 25688 18844 25740 18853
rect 22652 18708 22704 18760
rect 24216 18708 24268 18760
rect 25964 18776 26016 18828
rect 26148 18819 26200 18828
rect 26148 18785 26157 18819
rect 26157 18785 26191 18819
rect 26191 18785 26200 18819
rect 26148 18776 26200 18785
rect 26240 18776 26292 18828
rect 25872 18708 25924 18760
rect 24124 18640 24176 18692
rect 28172 18683 28224 18692
rect 28172 18649 28181 18683
rect 28181 18649 28215 18683
rect 28215 18649 28224 18683
rect 28172 18640 28224 18649
rect 22376 18572 22428 18624
rect 25044 18572 25096 18624
rect 25412 18572 25464 18624
rect 26608 18572 26660 18624
rect 5614 18470 5666 18522
rect 5678 18470 5730 18522
rect 5742 18470 5794 18522
rect 5806 18470 5858 18522
rect 14878 18470 14930 18522
rect 14942 18470 14994 18522
rect 15006 18470 15058 18522
rect 15070 18470 15122 18522
rect 24142 18470 24194 18522
rect 24206 18470 24258 18522
rect 24270 18470 24322 18522
rect 24334 18470 24386 18522
rect 2412 18368 2464 18420
rect 5448 18411 5500 18420
rect 5448 18377 5457 18411
rect 5457 18377 5491 18411
rect 5491 18377 5500 18411
rect 5448 18368 5500 18377
rect 2688 18300 2740 18352
rect 11796 18368 11848 18420
rect 11888 18368 11940 18420
rect 15844 18368 15896 18420
rect 17592 18368 17644 18420
rect 18328 18411 18380 18420
rect 18328 18377 18337 18411
rect 18337 18377 18371 18411
rect 18371 18377 18380 18411
rect 18328 18368 18380 18377
rect 9220 18300 9272 18352
rect 2320 18232 2372 18284
rect 2780 18096 2832 18148
rect 1860 18071 1912 18080
rect 1860 18037 1869 18071
rect 1869 18037 1903 18071
rect 1903 18037 1912 18071
rect 1860 18028 1912 18037
rect 2320 18071 2372 18080
rect 2320 18037 2329 18071
rect 2329 18037 2363 18071
rect 2363 18037 2372 18071
rect 3056 18207 3108 18216
rect 3056 18173 3065 18207
rect 3065 18173 3099 18207
rect 3099 18173 3108 18207
rect 4804 18232 4856 18284
rect 5908 18232 5960 18284
rect 11612 18300 11664 18352
rect 3056 18164 3108 18173
rect 4160 18164 4212 18216
rect 5080 18164 5132 18216
rect 13820 18300 13872 18352
rect 13084 18232 13136 18284
rect 13912 18232 13964 18284
rect 17408 18300 17460 18352
rect 19524 18368 19576 18420
rect 20812 18411 20864 18420
rect 15844 18232 15896 18284
rect 19984 18300 20036 18352
rect 20812 18377 20821 18411
rect 20821 18377 20855 18411
rect 20855 18377 20864 18411
rect 20812 18368 20864 18377
rect 21272 18368 21324 18420
rect 21548 18368 21600 18420
rect 23480 18300 23532 18352
rect 24676 18368 24728 18420
rect 25044 18300 25096 18352
rect 19248 18232 19300 18284
rect 8760 18164 8812 18216
rect 9404 18164 9456 18216
rect 10140 18164 10192 18216
rect 11060 18164 11112 18216
rect 11520 18164 11572 18216
rect 11704 18164 11756 18216
rect 14648 18164 14700 18216
rect 16028 18164 16080 18216
rect 16580 18207 16632 18216
rect 16580 18173 16589 18207
rect 16589 18173 16623 18207
rect 16623 18173 16632 18207
rect 16580 18164 16632 18173
rect 6000 18096 6052 18148
rect 16396 18096 16448 18148
rect 16672 18096 16724 18148
rect 17868 18164 17920 18216
rect 21732 18232 21784 18284
rect 22284 18275 22336 18284
rect 22284 18241 22293 18275
rect 22293 18241 22327 18275
rect 22327 18241 22336 18275
rect 22284 18232 22336 18241
rect 23940 18232 23992 18284
rect 25964 18368 26016 18420
rect 26148 18368 26200 18420
rect 27436 18411 27488 18420
rect 27436 18377 27445 18411
rect 27445 18377 27479 18411
rect 27479 18377 27488 18411
rect 27436 18368 27488 18377
rect 28080 18368 28132 18420
rect 20720 18207 20772 18216
rect 20720 18173 20729 18207
rect 20729 18173 20763 18207
rect 20763 18173 20772 18207
rect 20720 18164 20772 18173
rect 20904 18207 20956 18216
rect 20904 18173 20913 18207
rect 20913 18173 20947 18207
rect 20947 18173 20956 18207
rect 20904 18164 20956 18173
rect 21180 18207 21232 18216
rect 21180 18173 21189 18207
rect 21189 18173 21223 18207
rect 21223 18173 21232 18207
rect 21180 18164 21232 18173
rect 22376 18164 22428 18216
rect 28080 18275 28132 18284
rect 28080 18241 28089 18275
rect 28089 18241 28123 18275
rect 28123 18241 28132 18275
rect 28080 18232 28132 18241
rect 25320 18164 25372 18216
rect 27804 18207 27856 18216
rect 27804 18173 27813 18207
rect 27813 18173 27847 18207
rect 27847 18173 27856 18207
rect 27804 18164 27856 18173
rect 4804 18071 4856 18080
rect 2320 18028 2372 18037
rect 4804 18037 4813 18071
rect 4813 18037 4847 18071
rect 4847 18037 4856 18071
rect 4804 18028 4856 18037
rect 8300 18028 8352 18080
rect 12072 18028 12124 18080
rect 15568 18028 15620 18080
rect 15752 18028 15804 18080
rect 21272 18096 21324 18148
rect 17040 18028 17092 18080
rect 23940 18096 23992 18148
rect 27712 18028 27764 18080
rect 10246 17926 10298 17978
rect 10310 17926 10362 17978
rect 10374 17926 10426 17978
rect 10438 17926 10490 17978
rect 19510 17926 19562 17978
rect 19574 17926 19626 17978
rect 19638 17926 19690 17978
rect 19702 17926 19754 17978
rect 2780 17867 2832 17876
rect 2780 17833 2789 17867
rect 2789 17833 2823 17867
rect 2823 17833 2832 17867
rect 2780 17824 2832 17833
rect 4804 17824 4856 17876
rect 8852 17824 8904 17876
rect 8944 17824 8996 17876
rect 9588 17824 9640 17876
rect 10140 17824 10192 17876
rect 10692 17867 10744 17876
rect 10692 17833 10701 17867
rect 10701 17833 10735 17867
rect 10735 17833 10744 17867
rect 10692 17824 10744 17833
rect 14188 17867 14240 17876
rect 1860 17756 1912 17808
rect 4344 17756 4396 17808
rect 5172 17756 5224 17808
rect 6184 17756 6236 17808
rect 8576 17799 8628 17808
rect 8576 17765 8610 17799
rect 8610 17765 8628 17799
rect 8576 17756 8628 17765
rect 8668 17756 8720 17808
rect 14188 17833 14197 17867
rect 14197 17833 14231 17867
rect 14231 17833 14240 17867
rect 14188 17824 14240 17833
rect 15476 17824 15528 17876
rect 16396 17824 16448 17876
rect 18236 17824 18288 17876
rect 21640 17824 21692 17876
rect 26516 17824 26568 17876
rect 3056 17688 3108 17740
rect 4160 17688 4212 17740
rect 3884 17663 3936 17672
rect 3884 17629 3893 17663
rect 3893 17629 3927 17663
rect 3927 17629 3936 17663
rect 3884 17620 3936 17629
rect 2964 17552 3016 17604
rect 7380 17688 7432 17740
rect 7472 17688 7524 17740
rect 12716 17688 12768 17740
rect 14188 17688 14240 17740
rect 14556 17731 14608 17740
rect 14556 17697 14565 17731
rect 14565 17697 14599 17731
rect 14599 17697 14608 17731
rect 14556 17688 14608 17697
rect 17592 17688 17644 17740
rect 17960 17731 18012 17740
rect 17960 17697 17969 17731
rect 17969 17697 18003 17731
rect 18003 17697 18012 17731
rect 17960 17688 18012 17697
rect 23480 17756 23532 17808
rect 25044 17756 25096 17808
rect 23020 17688 23072 17740
rect 26608 17688 26660 17740
rect 26884 17731 26936 17740
rect 5908 17552 5960 17604
rect 7012 17552 7064 17604
rect 6736 17484 6788 17536
rect 7288 17484 7340 17536
rect 11244 17620 11296 17672
rect 12256 17620 12308 17672
rect 14648 17620 14700 17672
rect 17868 17663 17920 17672
rect 17592 17552 17644 17604
rect 17868 17629 17877 17663
rect 17877 17629 17911 17663
rect 17911 17629 17920 17663
rect 17868 17620 17920 17629
rect 25688 17620 25740 17672
rect 26884 17697 26893 17731
rect 26893 17697 26927 17731
rect 26927 17697 26936 17731
rect 26884 17688 26936 17697
rect 28172 17595 28224 17604
rect 28172 17561 28181 17595
rect 28181 17561 28215 17595
rect 28215 17561 28224 17595
rect 28172 17552 28224 17561
rect 8484 17484 8536 17536
rect 11888 17484 11940 17536
rect 5614 17382 5666 17434
rect 5678 17382 5730 17434
rect 5742 17382 5794 17434
rect 5806 17382 5858 17434
rect 14878 17382 14930 17434
rect 14942 17382 14994 17434
rect 15006 17382 15058 17434
rect 15070 17382 15122 17434
rect 24142 17382 24194 17434
rect 24206 17382 24258 17434
rect 24270 17382 24322 17434
rect 24334 17382 24386 17434
rect 3056 17323 3108 17332
rect 3056 17289 3065 17323
rect 3065 17289 3099 17323
rect 3099 17289 3108 17323
rect 3056 17280 3108 17289
rect 5172 17323 5224 17332
rect 5172 17289 5181 17323
rect 5181 17289 5215 17323
rect 5215 17289 5224 17323
rect 5172 17280 5224 17289
rect 9864 17280 9916 17332
rect 20536 17280 20588 17332
rect 20904 17280 20956 17332
rect 26884 17323 26936 17332
rect 26884 17289 26893 17323
rect 26893 17289 26927 17323
rect 26927 17289 26936 17323
rect 26884 17280 26936 17289
rect 4988 17212 5040 17264
rect 1676 17144 1728 17196
rect 14556 17212 14608 17264
rect 20996 17212 21048 17264
rect 21364 17212 21416 17264
rect 21640 17255 21692 17264
rect 21640 17221 21649 17255
rect 21649 17221 21683 17255
rect 21683 17221 21692 17255
rect 21640 17212 21692 17221
rect 6092 17144 6144 17196
rect 6644 17144 6696 17196
rect 7564 17187 7616 17196
rect 7564 17153 7573 17187
rect 7573 17153 7607 17187
rect 7607 17153 7616 17187
rect 7564 17144 7616 17153
rect 19248 17144 19300 17196
rect 20904 17144 20956 17196
rect 21088 17144 21140 17196
rect 28356 17144 28408 17196
rect 1952 17119 2004 17128
rect 1952 17085 1961 17119
rect 1961 17085 1995 17119
rect 1995 17085 2004 17119
rect 1952 17076 2004 17085
rect 2872 17076 2924 17128
rect 3976 17076 4028 17128
rect 4988 17076 5040 17128
rect 7288 17119 7340 17128
rect 7288 17085 7297 17119
rect 7297 17085 7331 17119
rect 7331 17085 7340 17119
rect 7288 17076 7340 17085
rect 9588 17119 9640 17128
rect 9588 17085 9597 17119
rect 9597 17085 9631 17119
rect 9631 17085 9640 17119
rect 9588 17076 9640 17085
rect 2688 17008 2740 17060
rect 6000 17008 6052 17060
rect 9404 17008 9456 17060
rect 11428 17076 11480 17128
rect 11888 17076 11940 17128
rect 15200 17076 15252 17128
rect 20076 17008 20128 17060
rect 26240 17051 26292 17060
rect 26240 17017 26249 17051
rect 26249 17017 26283 17051
rect 26283 17017 26292 17051
rect 26240 17008 26292 17017
rect 26332 17008 26384 17060
rect 5632 16983 5684 16992
rect 5632 16949 5641 16983
rect 5641 16949 5675 16983
rect 5675 16949 5684 16983
rect 6920 16983 6972 16992
rect 5632 16940 5684 16949
rect 6920 16949 6929 16983
rect 6929 16949 6963 16983
rect 6963 16949 6972 16983
rect 6920 16940 6972 16949
rect 8300 16940 8352 16992
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 18328 16983 18380 16992
rect 18328 16949 18337 16983
rect 18337 16949 18371 16983
rect 18371 16949 18380 16983
rect 18328 16940 18380 16949
rect 18420 16940 18472 16992
rect 21180 16940 21232 16992
rect 24400 16940 24452 16992
rect 24768 16940 24820 16992
rect 27436 16983 27488 16992
rect 27436 16949 27445 16983
rect 27445 16949 27479 16983
rect 27479 16949 27488 16983
rect 27436 16940 27488 16949
rect 27804 16983 27856 16992
rect 27804 16949 27813 16983
rect 27813 16949 27847 16983
rect 27847 16949 27856 16983
rect 27804 16940 27856 16949
rect 27896 16983 27948 16992
rect 27896 16949 27905 16983
rect 27905 16949 27939 16983
rect 27939 16949 27948 16983
rect 27896 16940 27948 16949
rect 10246 16838 10298 16890
rect 10310 16838 10362 16890
rect 10374 16838 10426 16890
rect 10438 16838 10490 16890
rect 19510 16838 19562 16890
rect 19574 16838 19626 16890
rect 19638 16838 19690 16890
rect 19702 16838 19754 16890
rect 1768 16779 1820 16788
rect 1768 16745 1777 16779
rect 1777 16745 1811 16779
rect 1811 16745 1820 16779
rect 1768 16736 1820 16745
rect 1952 16643 2004 16652
rect 1952 16609 1961 16643
rect 1961 16609 1995 16643
rect 1995 16609 2004 16643
rect 1952 16600 2004 16609
rect 2688 16668 2740 16720
rect 4620 16736 4672 16788
rect 5632 16736 5684 16788
rect 5908 16736 5960 16788
rect 7472 16736 7524 16788
rect 8300 16779 8352 16788
rect 8300 16745 8309 16779
rect 8309 16745 8343 16779
rect 8343 16745 8352 16779
rect 8300 16736 8352 16745
rect 9496 16736 9548 16788
rect 10048 16736 10100 16788
rect 17132 16736 17184 16788
rect 6920 16668 6972 16720
rect 14464 16668 14516 16720
rect 15936 16668 15988 16720
rect 17960 16668 18012 16720
rect 18328 16668 18380 16720
rect 20812 16668 20864 16720
rect 2780 16600 2832 16652
rect 3240 16643 3292 16652
rect 3240 16609 3249 16643
rect 3249 16609 3283 16643
rect 3283 16609 3292 16643
rect 3240 16600 3292 16609
rect 3332 16600 3384 16652
rect 2596 16464 2648 16516
rect 6828 16600 6880 16652
rect 9404 16600 9456 16652
rect 14280 16600 14332 16652
rect 17592 16643 17644 16652
rect 6736 16532 6788 16584
rect 13084 16532 13136 16584
rect 17592 16609 17601 16643
rect 17601 16609 17635 16643
rect 17635 16609 17644 16643
rect 17592 16600 17644 16609
rect 17868 16600 17920 16652
rect 18420 16600 18472 16652
rect 19984 16600 20036 16652
rect 20996 16643 21048 16652
rect 20996 16609 21005 16643
rect 21005 16609 21039 16643
rect 21039 16609 21048 16643
rect 20996 16600 21048 16609
rect 17224 16396 17276 16448
rect 20168 16532 20220 16584
rect 20904 16575 20956 16584
rect 20904 16541 20913 16575
rect 20913 16541 20947 16575
rect 20947 16541 20956 16575
rect 20904 16532 20956 16541
rect 21180 16668 21232 16720
rect 24676 16668 24728 16720
rect 24768 16668 24820 16720
rect 27712 16668 27764 16720
rect 23572 16600 23624 16652
rect 22652 16532 22704 16584
rect 23112 16532 23164 16584
rect 24032 16600 24084 16652
rect 25228 16600 25280 16652
rect 26884 16643 26936 16652
rect 26884 16609 26893 16643
rect 26893 16609 26927 16643
rect 26927 16609 26936 16643
rect 26884 16600 26936 16609
rect 28172 16643 28224 16652
rect 28172 16609 28181 16643
rect 28181 16609 28215 16643
rect 28215 16609 28224 16643
rect 28172 16600 28224 16609
rect 24216 16575 24268 16584
rect 24216 16541 24225 16575
rect 24225 16541 24259 16575
rect 24259 16541 24268 16575
rect 24216 16532 24268 16541
rect 22284 16464 22336 16516
rect 24400 16464 24452 16516
rect 20076 16396 20128 16448
rect 20720 16439 20772 16448
rect 20720 16405 20729 16439
rect 20729 16405 20763 16439
rect 20763 16405 20772 16439
rect 20720 16396 20772 16405
rect 24860 16396 24912 16448
rect 25688 16396 25740 16448
rect 5614 16294 5666 16346
rect 5678 16294 5730 16346
rect 5742 16294 5794 16346
rect 5806 16294 5858 16346
rect 14878 16294 14930 16346
rect 14942 16294 14994 16346
rect 15006 16294 15058 16346
rect 15070 16294 15122 16346
rect 24142 16294 24194 16346
rect 24206 16294 24258 16346
rect 24270 16294 24322 16346
rect 24334 16294 24386 16346
rect 4988 16235 5040 16244
rect 4988 16201 4997 16235
rect 4997 16201 5031 16235
rect 5031 16201 5040 16235
rect 4988 16192 5040 16201
rect 12164 16192 12216 16244
rect 15568 16192 15620 16244
rect 17592 16192 17644 16244
rect 18420 16192 18472 16244
rect 18972 16192 19024 16244
rect 21640 16235 21692 16244
rect 4252 16124 4304 16176
rect 1860 16031 1912 16040
rect 1860 15997 1869 16031
rect 1869 15997 1903 16031
rect 1903 15997 1912 16031
rect 1860 15988 1912 15997
rect 5908 16124 5960 16176
rect 15108 16124 15160 16176
rect 5172 15988 5224 16040
rect 15200 15988 15252 16040
rect 15844 16056 15896 16108
rect 20168 16124 20220 16176
rect 21640 16201 21649 16235
rect 21649 16201 21683 16235
rect 21683 16201 21692 16235
rect 21640 16192 21692 16201
rect 22284 16192 22336 16244
rect 23572 16235 23624 16244
rect 23572 16201 23581 16235
rect 23581 16201 23615 16235
rect 23615 16201 23624 16235
rect 23572 16192 23624 16201
rect 25228 16235 25280 16244
rect 25228 16201 25237 16235
rect 25237 16201 25271 16235
rect 25271 16201 25280 16235
rect 25228 16192 25280 16201
rect 26792 16192 26844 16244
rect 17224 16056 17276 16108
rect 17132 15988 17184 16040
rect 17960 15988 18012 16040
rect 18328 15988 18380 16040
rect 19984 15988 20036 16040
rect 22560 16056 22612 16108
rect 22652 16031 22704 16040
rect 2964 15920 3016 15972
rect 5080 15920 5132 15972
rect 15936 15963 15988 15972
rect 1952 15895 2004 15904
rect 1952 15861 1961 15895
rect 1961 15861 1995 15895
rect 1995 15861 2004 15895
rect 1952 15852 2004 15861
rect 3700 15852 3752 15904
rect 10876 15895 10928 15904
rect 10876 15861 10885 15895
rect 10885 15861 10919 15895
rect 10919 15861 10928 15895
rect 10876 15852 10928 15861
rect 11428 15852 11480 15904
rect 13084 15852 13136 15904
rect 13268 15895 13320 15904
rect 13268 15861 13277 15895
rect 13277 15861 13311 15895
rect 13311 15861 13320 15895
rect 13268 15852 13320 15861
rect 15568 15852 15620 15904
rect 15936 15929 15945 15963
rect 15945 15929 15979 15963
rect 15979 15929 15988 15963
rect 15936 15920 15988 15929
rect 16120 15920 16172 15972
rect 18972 15920 19024 15972
rect 20720 15920 20772 15972
rect 22652 15997 22661 16031
rect 22661 15997 22695 16031
rect 22695 15997 22704 16031
rect 22652 15988 22704 15997
rect 22928 15988 22980 16040
rect 23112 15988 23164 16040
rect 27988 16124 28040 16176
rect 25780 16099 25832 16108
rect 25780 16065 25789 16099
rect 25789 16065 25823 16099
rect 25823 16065 25832 16099
rect 25780 16056 25832 16065
rect 17224 15852 17276 15904
rect 17500 15852 17552 15904
rect 17960 15852 18012 15904
rect 20260 15852 20312 15904
rect 22284 15895 22336 15904
rect 22284 15861 22293 15895
rect 22293 15861 22327 15895
rect 22327 15861 22336 15895
rect 22284 15852 22336 15861
rect 22744 15920 22796 15972
rect 24952 15988 25004 16040
rect 25688 16031 25740 16040
rect 25688 15997 25697 16031
rect 25697 15997 25731 16031
rect 25731 15997 25740 16031
rect 25688 15988 25740 15997
rect 26240 15988 26292 16040
rect 26516 15988 26568 16040
rect 27252 16031 27304 16040
rect 27252 15997 27261 16031
rect 27261 15997 27295 16031
rect 27295 15997 27304 16031
rect 27252 15988 27304 15997
rect 27528 16031 27580 16040
rect 27528 15997 27537 16031
rect 27537 15997 27571 16031
rect 27571 15997 27580 16031
rect 27528 15988 27580 15997
rect 25504 15920 25556 15972
rect 25872 15920 25924 15972
rect 10246 15750 10298 15802
rect 10310 15750 10362 15802
rect 10374 15750 10426 15802
rect 10438 15750 10490 15802
rect 19510 15750 19562 15802
rect 19574 15750 19626 15802
rect 19638 15750 19690 15802
rect 19702 15750 19754 15802
rect 5080 15648 5132 15700
rect 5448 15648 5500 15700
rect 20168 15648 20220 15700
rect 26424 15691 26476 15700
rect 26424 15657 26433 15691
rect 26433 15657 26467 15691
rect 26467 15657 26476 15691
rect 26424 15648 26476 15657
rect 27528 15648 27580 15700
rect 1860 15623 1912 15632
rect 1860 15589 1869 15623
rect 1869 15589 1903 15623
rect 1903 15589 1912 15623
rect 1860 15580 1912 15589
rect 1584 15512 1636 15564
rect 2596 15580 2648 15632
rect 3884 15580 3936 15632
rect 4436 15580 4488 15632
rect 4620 15580 4672 15632
rect 10692 15580 10744 15632
rect 11060 15623 11112 15632
rect 11060 15589 11069 15623
rect 11069 15589 11103 15623
rect 11103 15589 11112 15623
rect 11060 15580 11112 15589
rect 11980 15580 12032 15632
rect 2964 15555 3016 15564
rect 2964 15521 2973 15555
rect 2973 15521 3007 15555
rect 3007 15521 3016 15555
rect 2964 15512 3016 15521
rect 3976 15555 4028 15564
rect 3976 15521 3985 15555
rect 3985 15521 4019 15555
rect 4019 15521 4028 15555
rect 3976 15512 4028 15521
rect 4252 15512 4304 15564
rect 4436 15444 4488 15496
rect 4620 15444 4672 15496
rect 9496 15512 9548 15564
rect 12164 15512 12216 15564
rect 15568 15580 15620 15632
rect 17960 15580 18012 15632
rect 18972 15623 19024 15632
rect 18972 15589 18981 15623
rect 18981 15589 19015 15623
rect 19015 15589 19024 15623
rect 18972 15580 19024 15589
rect 19064 15580 19116 15632
rect 19340 15623 19392 15632
rect 19340 15589 19371 15623
rect 19371 15589 19392 15623
rect 19340 15580 19392 15589
rect 21640 15580 21692 15632
rect 23112 15580 23164 15632
rect 24768 15580 24820 15632
rect 25228 15580 25280 15632
rect 8300 15487 8352 15496
rect 8300 15453 8309 15487
rect 8309 15453 8343 15487
rect 8343 15453 8352 15487
rect 8300 15444 8352 15453
rect 10968 15487 11020 15496
rect 10968 15453 10977 15487
rect 10977 15453 11011 15487
rect 11011 15453 11020 15487
rect 10968 15444 11020 15453
rect 13820 15512 13872 15564
rect 15476 15512 15528 15564
rect 16304 15512 16356 15564
rect 16672 15512 16724 15564
rect 17132 15512 17184 15564
rect 20076 15512 20128 15564
rect 20260 15512 20312 15564
rect 22744 15512 22796 15564
rect 25596 15580 25648 15632
rect 25688 15580 25740 15632
rect 13912 15487 13964 15496
rect 13912 15453 13921 15487
rect 13921 15453 13955 15487
rect 13955 15453 13964 15487
rect 13912 15444 13964 15453
rect 15200 15444 15252 15496
rect 15936 15444 15988 15496
rect 18696 15444 18748 15496
rect 11428 15376 11480 15428
rect 13084 15376 13136 15428
rect 4160 15308 4212 15360
rect 4344 15351 4396 15360
rect 4344 15317 4353 15351
rect 4353 15317 4387 15351
rect 4387 15317 4396 15351
rect 4344 15308 4396 15317
rect 9680 15351 9732 15360
rect 9680 15317 9689 15351
rect 9689 15317 9723 15351
rect 9723 15317 9732 15351
rect 9680 15308 9732 15317
rect 12348 15308 12400 15360
rect 15200 15308 15252 15360
rect 15568 15376 15620 15428
rect 16120 15376 16172 15428
rect 18328 15376 18380 15428
rect 22284 15444 22336 15496
rect 23848 15444 23900 15496
rect 25504 15444 25556 15496
rect 20536 15376 20588 15428
rect 23480 15376 23532 15428
rect 24492 15376 24544 15428
rect 18972 15308 19024 15360
rect 27528 15308 27580 15360
rect 5614 15206 5666 15258
rect 5678 15206 5730 15258
rect 5742 15206 5794 15258
rect 5806 15206 5858 15258
rect 14878 15206 14930 15258
rect 14942 15206 14994 15258
rect 15006 15206 15058 15258
rect 15070 15206 15122 15258
rect 24142 15206 24194 15258
rect 24206 15206 24258 15258
rect 24270 15206 24322 15258
rect 24334 15206 24386 15258
rect 2780 15104 2832 15156
rect 6828 15104 6880 15156
rect 9496 15147 9548 15156
rect 9496 15113 9505 15147
rect 9505 15113 9539 15147
rect 9539 15113 9548 15147
rect 9496 15104 9548 15113
rect 10692 15147 10744 15156
rect 10692 15113 10701 15147
rect 10701 15113 10735 15147
rect 10735 15113 10744 15147
rect 10692 15104 10744 15113
rect 12164 15104 12216 15156
rect 13820 15104 13872 15156
rect 15844 15104 15896 15156
rect 16120 15104 16172 15156
rect 17684 15147 17736 15156
rect 17684 15113 17693 15147
rect 17693 15113 17727 15147
rect 17727 15113 17736 15147
rect 17684 15104 17736 15113
rect 21916 15147 21968 15156
rect 21916 15113 21925 15147
rect 21925 15113 21959 15147
rect 21959 15113 21968 15147
rect 21916 15104 21968 15113
rect 27804 15104 27856 15156
rect 27896 15104 27948 15156
rect 1400 14968 1452 15020
rect 1768 14900 1820 14952
rect 1584 14875 1636 14884
rect 1584 14841 1593 14875
rect 1593 14841 1627 14875
rect 1627 14841 1636 14875
rect 1584 14832 1636 14841
rect 2504 14900 2556 14952
rect 5080 15036 5132 15088
rect 12532 15036 12584 15088
rect 6644 14968 6696 15020
rect 10048 15011 10100 15020
rect 10048 14977 10057 15011
rect 10057 14977 10091 15011
rect 10091 14977 10100 15011
rect 10048 14968 10100 14977
rect 10876 14968 10928 15020
rect 11244 14968 11296 15020
rect 11704 14968 11756 15020
rect 3700 14900 3752 14952
rect 5080 14900 5132 14952
rect 5264 14900 5316 14952
rect 5448 14943 5500 14952
rect 5448 14909 5457 14943
rect 5457 14909 5491 14943
rect 5491 14909 5500 14943
rect 5448 14900 5500 14909
rect 5908 14943 5960 14952
rect 5908 14909 5917 14943
rect 5917 14909 5951 14943
rect 5951 14909 5960 14943
rect 5908 14900 5960 14909
rect 6276 14900 6328 14952
rect 9680 14900 9732 14952
rect 12348 14943 12400 14952
rect 12348 14909 12357 14943
rect 12357 14909 12391 14943
rect 12391 14909 12400 14943
rect 12348 14900 12400 14909
rect 13360 15036 13412 15088
rect 13544 15036 13596 15088
rect 14648 14968 14700 15020
rect 15200 14968 15252 15020
rect 13820 14943 13872 14952
rect 2872 14832 2924 14884
rect 1768 14764 1820 14816
rect 3516 14764 3568 14816
rect 4068 14764 4120 14816
rect 4436 14764 4488 14816
rect 4804 14764 4856 14816
rect 5172 14807 5224 14816
rect 5172 14773 5181 14807
rect 5181 14773 5215 14807
rect 5215 14773 5224 14807
rect 5172 14764 5224 14773
rect 5816 14832 5868 14884
rect 10600 14832 10652 14884
rect 6460 14807 6512 14816
rect 6460 14773 6469 14807
rect 6469 14773 6503 14807
rect 6503 14773 6512 14807
rect 6460 14764 6512 14773
rect 7380 14807 7432 14816
rect 7380 14773 7389 14807
rect 7389 14773 7423 14807
rect 7423 14773 7432 14807
rect 7380 14764 7432 14773
rect 9128 14764 9180 14816
rect 10140 14764 10192 14816
rect 12256 14764 12308 14816
rect 12808 14832 12860 14884
rect 13084 14832 13136 14884
rect 13820 14909 13829 14943
rect 13829 14909 13863 14943
rect 13863 14909 13872 14943
rect 13820 14900 13872 14909
rect 17500 14968 17552 15020
rect 26056 15011 26108 15020
rect 26056 14977 26065 15011
rect 26065 14977 26099 15011
rect 26099 14977 26108 15011
rect 26056 14968 26108 14977
rect 17592 14900 17644 14952
rect 21548 14900 21600 14952
rect 21732 14900 21784 14952
rect 22652 14900 22704 14952
rect 26424 14900 26476 14952
rect 14280 14832 14332 14884
rect 17132 14875 17184 14884
rect 17132 14841 17141 14875
rect 17141 14841 17175 14875
rect 17175 14841 17184 14875
rect 17132 14832 17184 14841
rect 24860 14832 24912 14884
rect 25872 14832 25924 14884
rect 27436 14900 27488 14952
rect 17592 14764 17644 14816
rect 22468 14764 22520 14816
rect 10246 14662 10298 14714
rect 10310 14662 10362 14714
rect 10374 14662 10426 14714
rect 10438 14662 10490 14714
rect 19510 14662 19562 14714
rect 19574 14662 19626 14714
rect 19638 14662 19690 14714
rect 19702 14662 19754 14714
rect 1768 14603 1820 14612
rect 1768 14569 1777 14603
rect 1777 14569 1811 14603
rect 1811 14569 1820 14603
rect 1768 14560 1820 14569
rect 2504 14560 2556 14612
rect 3884 14560 3936 14612
rect 4436 14560 4488 14612
rect 4804 14560 4856 14612
rect 10140 14603 10192 14612
rect 10140 14569 10149 14603
rect 10149 14569 10183 14603
rect 10183 14569 10192 14603
rect 10140 14560 10192 14569
rect 10968 14603 11020 14612
rect 10968 14569 10977 14603
rect 10977 14569 11011 14603
rect 11011 14569 11020 14603
rect 10968 14560 11020 14569
rect 13820 14560 13872 14612
rect 14188 14560 14240 14612
rect 14648 14560 14700 14612
rect 17592 14560 17644 14612
rect 17868 14603 17920 14612
rect 17868 14569 17877 14603
rect 17877 14569 17911 14603
rect 17911 14569 17920 14603
rect 17868 14560 17920 14569
rect 19064 14560 19116 14612
rect 21088 14603 21140 14612
rect 21088 14569 21097 14603
rect 21097 14569 21131 14603
rect 21131 14569 21140 14603
rect 21088 14560 21140 14569
rect 21916 14560 21968 14612
rect 22652 14603 22704 14612
rect 22652 14569 22661 14603
rect 22661 14569 22695 14603
rect 22695 14569 22704 14603
rect 22652 14560 22704 14569
rect 26056 14560 26108 14612
rect 1952 14467 2004 14476
rect 1952 14433 1961 14467
rect 1961 14433 1995 14467
rect 1995 14433 2004 14467
rect 1952 14424 2004 14433
rect 2780 14424 2832 14476
rect 3792 14492 3844 14544
rect 3700 14467 3752 14476
rect 3700 14433 3709 14467
rect 3709 14433 3743 14467
rect 3743 14433 3752 14467
rect 3700 14424 3752 14433
rect 3976 14424 4028 14476
rect 4436 14424 4488 14476
rect 4804 14288 4856 14340
rect 6460 14424 6512 14476
rect 7104 14424 7156 14476
rect 9680 14492 9732 14544
rect 12440 14535 12492 14544
rect 12440 14501 12449 14535
rect 12449 14501 12483 14535
rect 12483 14501 12492 14535
rect 12440 14492 12492 14501
rect 13084 14492 13136 14544
rect 10968 14424 11020 14476
rect 12348 14424 12400 14476
rect 13360 14467 13412 14476
rect 13360 14433 13369 14467
rect 13369 14433 13403 14467
rect 13403 14433 13412 14467
rect 13360 14424 13412 14433
rect 14188 14424 14240 14476
rect 17500 14467 17552 14476
rect 17500 14433 17509 14467
rect 17509 14433 17543 14467
rect 17543 14433 17552 14467
rect 17500 14424 17552 14433
rect 9680 14356 9732 14408
rect 9956 14356 10008 14408
rect 17868 14356 17920 14408
rect 17684 14288 17736 14340
rect 4988 14220 5040 14272
rect 9128 14220 9180 14272
rect 9864 14220 9916 14272
rect 10600 14220 10652 14272
rect 25688 14492 25740 14544
rect 25964 14535 26016 14544
rect 25964 14501 25973 14535
rect 25973 14501 26007 14535
rect 26007 14501 26016 14535
rect 25964 14492 26016 14501
rect 27988 14535 28040 14544
rect 27988 14501 27997 14535
rect 27997 14501 28031 14535
rect 28031 14501 28040 14535
rect 27988 14492 28040 14501
rect 20720 14424 20772 14476
rect 21180 14467 21232 14476
rect 21180 14433 21189 14467
rect 21189 14433 21223 14467
rect 21223 14433 21232 14467
rect 21180 14424 21232 14433
rect 22652 14424 22704 14476
rect 23020 14424 23072 14476
rect 20904 14356 20956 14408
rect 21916 14356 21968 14408
rect 26424 14399 26476 14408
rect 26424 14365 26433 14399
rect 26433 14365 26467 14399
rect 26467 14365 26476 14399
rect 26424 14356 26476 14365
rect 20812 14331 20864 14340
rect 20812 14297 20821 14331
rect 20821 14297 20855 14331
rect 20855 14297 20864 14331
rect 20812 14288 20864 14297
rect 26700 14288 26752 14340
rect 27252 14288 27304 14340
rect 28172 14331 28224 14340
rect 28172 14297 28181 14331
rect 28181 14297 28215 14331
rect 28215 14297 28224 14331
rect 28172 14288 28224 14297
rect 27988 14220 28040 14272
rect 5614 14118 5666 14170
rect 5678 14118 5730 14170
rect 5742 14118 5794 14170
rect 5806 14118 5858 14170
rect 14878 14118 14930 14170
rect 14942 14118 14994 14170
rect 15006 14118 15058 14170
rect 15070 14118 15122 14170
rect 24142 14118 24194 14170
rect 24206 14118 24258 14170
rect 24270 14118 24322 14170
rect 24334 14118 24386 14170
rect 2320 14059 2372 14068
rect 2320 14025 2329 14059
rect 2329 14025 2363 14059
rect 2363 14025 2372 14059
rect 2320 14016 2372 14025
rect 2872 14059 2924 14068
rect 2872 14025 2881 14059
rect 2881 14025 2915 14059
rect 2915 14025 2924 14059
rect 2872 14016 2924 14025
rect 4712 14059 4764 14068
rect 4712 14025 4721 14059
rect 4721 14025 4755 14059
rect 4755 14025 4764 14059
rect 4712 14016 4764 14025
rect 10968 14059 11020 14068
rect 10968 14025 10977 14059
rect 10977 14025 11011 14059
rect 11011 14025 11020 14059
rect 10968 14016 11020 14025
rect 17132 14059 17184 14068
rect 17132 14025 17141 14059
rect 17141 14025 17175 14059
rect 17175 14025 17184 14059
rect 17132 14016 17184 14025
rect 20996 14016 21048 14068
rect 22652 14016 22704 14068
rect 23296 14016 23348 14068
rect 27436 14016 27488 14068
rect 3332 13948 3384 14000
rect 4620 13991 4672 14000
rect 4620 13957 4629 13991
rect 4629 13957 4663 13991
rect 4663 13957 4672 13991
rect 4620 13948 4672 13957
rect 7196 13948 7248 14000
rect 2596 13880 2648 13932
rect 2504 13812 2556 13864
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 4988 13880 5040 13932
rect 4896 13812 4948 13864
rect 7104 13855 7156 13864
rect 7104 13821 7113 13855
rect 7113 13821 7147 13855
rect 7147 13821 7156 13855
rect 7104 13812 7156 13821
rect 8208 13880 8260 13932
rect 12072 13948 12124 14000
rect 16580 13948 16632 14000
rect 17868 13948 17920 14000
rect 23848 13948 23900 14000
rect 11704 13880 11756 13932
rect 18880 13923 18932 13932
rect 18880 13889 18889 13923
rect 18889 13889 18923 13923
rect 18923 13889 18932 13923
rect 18880 13880 18932 13889
rect 20536 13880 20588 13932
rect 21088 13923 21140 13932
rect 21088 13889 21097 13923
rect 21097 13889 21131 13923
rect 21131 13889 21140 13923
rect 21088 13880 21140 13889
rect 9772 13855 9824 13864
rect 9772 13821 9781 13855
rect 9781 13821 9815 13855
rect 9815 13821 9824 13855
rect 9772 13812 9824 13821
rect 9864 13855 9916 13864
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 11888 13812 11940 13864
rect 14188 13812 14240 13864
rect 17040 13812 17092 13864
rect 17684 13855 17736 13864
rect 17684 13821 17693 13855
rect 17693 13821 17727 13855
rect 17727 13821 17736 13855
rect 17684 13812 17736 13821
rect 19984 13812 20036 13864
rect 20812 13855 20864 13864
rect 20812 13821 20821 13855
rect 20821 13821 20855 13855
rect 20855 13821 20864 13855
rect 20812 13812 20864 13821
rect 20996 13812 21048 13864
rect 21180 13855 21232 13864
rect 21180 13821 21189 13855
rect 21189 13821 21223 13855
rect 21223 13821 21232 13855
rect 21180 13812 21232 13821
rect 1492 13744 1544 13796
rect 4344 13787 4396 13796
rect 4344 13753 4353 13787
rect 4353 13753 4387 13787
rect 4387 13753 4396 13787
rect 4344 13744 4396 13753
rect 9220 13744 9272 13796
rect 9496 13744 9548 13796
rect 15936 13744 15988 13796
rect 21548 13744 21600 13796
rect 22468 13812 22520 13864
rect 24860 13812 24912 13864
rect 25964 13855 26016 13864
rect 25964 13821 25973 13855
rect 25973 13821 26007 13855
rect 26007 13821 26016 13855
rect 25964 13812 26016 13821
rect 26792 13812 26844 13864
rect 25228 13744 25280 13796
rect 27988 13855 28040 13864
rect 27988 13821 27997 13855
rect 27997 13821 28031 13855
rect 28031 13821 28040 13855
rect 27988 13812 28040 13821
rect 28172 13855 28224 13864
rect 28172 13821 28181 13855
rect 28181 13821 28215 13855
rect 28215 13821 28224 13855
rect 28172 13812 28224 13821
rect 27896 13744 27948 13796
rect 3516 13676 3568 13728
rect 12256 13719 12308 13728
rect 12256 13685 12265 13719
rect 12265 13685 12299 13719
rect 12299 13685 12308 13719
rect 12256 13676 12308 13685
rect 18328 13719 18380 13728
rect 18328 13685 18337 13719
rect 18337 13685 18371 13719
rect 18371 13685 18380 13719
rect 18328 13676 18380 13685
rect 18696 13719 18748 13728
rect 18696 13685 18705 13719
rect 18705 13685 18739 13719
rect 18739 13685 18748 13719
rect 18696 13676 18748 13685
rect 20720 13676 20772 13728
rect 10246 13574 10298 13626
rect 10310 13574 10362 13626
rect 10374 13574 10426 13626
rect 10438 13574 10490 13626
rect 19510 13574 19562 13626
rect 19574 13574 19626 13626
rect 19638 13574 19690 13626
rect 19702 13574 19754 13626
rect 2320 13472 2372 13524
rect 3516 13472 3568 13524
rect 3884 13472 3936 13524
rect 4160 13472 4212 13524
rect 9772 13472 9824 13524
rect 10140 13472 10192 13524
rect 12164 13472 12216 13524
rect 12992 13472 13044 13524
rect 13452 13472 13504 13524
rect 14096 13472 14148 13524
rect 17684 13472 17736 13524
rect 18696 13472 18748 13524
rect 19984 13515 20036 13524
rect 19984 13481 19993 13515
rect 19993 13481 20027 13515
rect 20027 13481 20036 13515
rect 19984 13472 20036 13481
rect 20720 13472 20772 13524
rect 21732 13472 21784 13524
rect 1860 13379 1912 13388
rect 1860 13345 1869 13379
rect 1869 13345 1903 13379
rect 1903 13345 1912 13379
rect 1860 13336 1912 13345
rect 2596 13379 2648 13388
rect 2596 13345 2605 13379
rect 2605 13345 2639 13379
rect 2639 13345 2648 13379
rect 2596 13336 2648 13345
rect 3424 13379 3476 13388
rect 3424 13345 3433 13379
rect 3433 13345 3467 13379
rect 3467 13345 3476 13379
rect 3424 13336 3476 13345
rect 3792 13336 3844 13388
rect 7656 13379 7708 13388
rect 7656 13345 7665 13379
rect 7665 13345 7699 13379
rect 7699 13345 7708 13379
rect 7656 13336 7708 13345
rect 7840 13336 7892 13388
rect 8208 13336 8260 13388
rect 9036 13404 9088 13456
rect 11980 13404 12032 13456
rect 12348 13404 12400 13456
rect 9128 13379 9180 13388
rect 9128 13345 9137 13379
rect 9137 13345 9171 13379
rect 9171 13345 9180 13379
rect 9128 13336 9180 13345
rect 10600 13336 10652 13388
rect 11244 13336 11296 13388
rect 13820 13336 13872 13388
rect 17592 13404 17644 13456
rect 18328 13404 18380 13456
rect 19248 13404 19300 13456
rect 25412 13472 25464 13524
rect 25688 13472 25740 13524
rect 16580 13336 16632 13388
rect 17500 13336 17552 13388
rect 20168 13336 20220 13388
rect 21088 13379 21140 13388
rect 5172 13311 5224 13320
rect 5172 13277 5181 13311
rect 5181 13277 5215 13311
rect 5215 13277 5224 13311
rect 5172 13268 5224 13277
rect 6460 13268 6512 13320
rect 6644 13268 6696 13320
rect 7932 13268 7984 13320
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 17684 13311 17736 13320
rect 2320 13200 2372 13252
rect 8208 13243 8260 13252
rect 8208 13209 8217 13243
rect 8217 13209 8251 13243
rect 8251 13209 8260 13243
rect 8208 13200 8260 13209
rect 6000 13132 6052 13184
rect 13912 13132 13964 13184
rect 17684 13277 17693 13311
rect 17693 13277 17727 13311
rect 17727 13277 17736 13311
rect 17684 13268 17736 13277
rect 15200 13200 15252 13252
rect 14740 13132 14792 13184
rect 18328 13132 18380 13184
rect 20444 13132 20496 13184
rect 21088 13345 21097 13379
rect 21097 13345 21131 13379
rect 21131 13345 21140 13379
rect 21088 13336 21140 13345
rect 21548 13336 21600 13388
rect 23848 13379 23900 13388
rect 23848 13345 23857 13379
rect 23857 13345 23891 13379
rect 23891 13345 23900 13379
rect 23848 13336 23900 13345
rect 20812 13200 20864 13252
rect 21180 13268 21232 13320
rect 20996 13132 21048 13184
rect 23572 13268 23624 13320
rect 24032 13336 24084 13388
rect 25044 13336 25096 13388
rect 24860 13268 24912 13320
rect 22928 13200 22980 13252
rect 23112 13200 23164 13252
rect 23940 13243 23992 13252
rect 23940 13209 23949 13243
rect 23949 13209 23983 13243
rect 23983 13209 23992 13243
rect 23940 13200 23992 13209
rect 24860 13132 24912 13184
rect 28172 13243 28224 13252
rect 28172 13209 28181 13243
rect 28181 13209 28215 13243
rect 28215 13209 28224 13243
rect 28172 13200 28224 13209
rect 25872 13132 25924 13184
rect 26148 13132 26200 13184
rect 5614 13030 5666 13082
rect 5678 13030 5730 13082
rect 5742 13030 5794 13082
rect 5806 13030 5858 13082
rect 14878 13030 14930 13082
rect 14942 13030 14994 13082
rect 15006 13030 15058 13082
rect 15070 13030 15122 13082
rect 24142 13030 24194 13082
rect 24206 13030 24258 13082
rect 24270 13030 24322 13082
rect 24334 13030 24386 13082
rect 4160 12928 4212 12980
rect 5172 12928 5224 12980
rect 1584 12792 1636 12844
rect 2780 12724 2832 12776
rect 2964 12724 3016 12776
rect 4160 12724 4212 12776
rect 11612 12928 11664 12980
rect 7012 12860 7064 12912
rect 8208 12835 8260 12844
rect 5908 12767 5960 12776
rect 1860 12699 1912 12708
rect 1860 12665 1869 12699
rect 1869 12665 1903 12699
rect 1903 12665 1912 12699
rect 1860 12656 1912 12665
rect 5908 12733 5917 12767
rect 5917 12733 5951 12767
rect 5951 12733 5960 12767
rect 5908 12724 5960 12733
rect 6000 12767 6052 12776
rect 6000 12733 6009 12767
rect 6009 12733 6043 12767
rect 6043 12733 6052 12767
rect 6184 12767 6236 12776
rect 6000 12724 6052 12733
rect 6184 12733 6193 12767
rect 6193 12733 6227 12767
rect 6227 12733 6236 12767
rect 6184 12724 6236 12733
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 7472 12767 7524 12776
rect 7472 12733 7481 12767
rect 7481 12733 7515 12767
rect 7515 12733 7524 12767
rect 7472 12724 7524 12733
rect 7840 12767 7892 12776
rect 7840 12733 7849 12767
rect 7849 12733 7883 12767
rect 7883 12733 7892 12767
rect 7840 12724 7892 12733
rect 8208 12801 8217 12835
rect 8217 12801 8251 12835
rect 8251 12801 8260 12835
rect 8208 12792 8260 12801
rect 10692 12724 10744 12776
rect 7288 12656 7340 12708
rect 11980 12792 12032 12844
rect 13912 12860 13964 12912
rect 14096 12860 14148 12912
rect 15108 12792 15160 12844
rect 11796 12724 11848 12776
rect 13636 12767 13688 12776
rect 13636 12733 13645 12767
rect 13645 12733 13679 12767
rect 13679 12733 13688 12767
rect 13636 12724 13688 12733
rect 14188 12724 14240 12776
rect 17500 12928 17552 12980
rect 17684 12971 17736 12980
rect 17684 12937 17693 12971
rect 17693 12937 17727 12971
rect 17727 12937 17736 12971
rect 17684 12928 17736 12937
rect 16120 12792 16172 12844
rect 19156 12928 19208 12980
rect 22284 12928 22336 12980
rect 24032 12928 24084 12980
rect 26700 12971 26752 12980
rect 26700 12937 26709 12971
rect 26709 12937 26743 12971
rect 26743 12937 26752 12971
rect 26700 12928 26752 12937
rect 17684 12792 17736 12844
rect 17040 12724 17092 12776
rect 17500 12767 17552 12776
rect 17500 12733 17509 12767
rect 17509 12733 17543 12767
rect 17543 12733 17552 12767
rect 17868 12767 17920 12776
rect 17500 12724 17552 12733
rect 17868 12733 17877 12767
rect 17877 12733 17911 12767
rect 17911 12733 17920 12767
rect 17868 12724 17920 12733
rect 17960 12724 18012 12776
rect 18144 12724 18196 12776
rect 18328 12792 18380 12844
rect 21180 12860 21232 12912
rect 22100 12860 22152 12912
rect 19156 12792 19208 12844
rect 22560 12792 22612 12844
rect 27896 12835 27948 12844
rect 27896 12801 27905 12835
rect 27905 12801 27939 12835
rect 27939 12801 27948 12835
rect 27896 12792 27948 12801
rect 28356 12792 28408 12844
rect 21364 12724 21416 12776
rect 3976 12588 4028 12640
rect 5172 12588 5224 12640
rect 13728 12656 13780 12708
rect 12072 12631 12124 12640
rect 12072 12597 12081 12631
rect 12081 12597 12115 12631
rect 12115 12597 12124 12631
rect 12072 12588 12124 12597
rect 12256 12588 12308 12640
rect 13636 12588 13688 12640
rect 14464 12588 14516 12640
rect 15568 12656 15620 12708
rect 18328 12656 18380 12708
rect 18696 12699 18748 12708
rect 18696 12665 18705 12699
rect 18705 12665 18739 12699
rect 18739 12665 18748 12699
rect 18696 12656 18748 12665
rect 16396 12588 16448 12640
rect 16580 12631 16632 12640
rect 16580 12597 16589 12631
rect 16589 12597 16623 12631
rect 16623 12597 16632 12631
rect 16580 12588 16632 12597
rect 17408 12588 17460 12640
rect 22284 12656 22336 12708
rect 23112 12724 23164 12776
rect 23296 12767 23348 12776
rect 23296 12733 23305 12767
rect 23305 12733 23339 12767
rect 23339 12733 23348 12767
rect 23296 12724 23348 12733
rect 21272 12588 21324 12640
rect 22560 12631 22612 12640
rect 22560 12597 22569 12631
rect 22569 12597 22603 12631
rect 22603 12597 22612 12631
rect 22560 12588 22612 12597
rect 23388 12656 23440 12708
rect 25504 12724 25556 12776
rect 25596 12724 25648 12776
rect 26148 12767 26200 12776
rect 25228 12656 25280 12708
rect 25688 12699 25740 12708
rect 25688 12665 25697 12699
rect 25697 12665 25731 12699
rect 25731 12665 25740 12699
rect 25688 12656 25740 12665
rect 26148 12733 26157 12767
rect 26157 12733 26191 12767
rect 26191 12733 26200 12767
rect 26148 12724 26200 12733
rect 26056 12656 26108 12708
rect 26516 12631 26568 12640
rect 26516 12597 26525 12631
rect 26525 12597 26559 12631
rect 26559 12597 26568 12631
rect 26516 12588 26568 12597
rect 27436 12631 27488 12640
rect 27436 12597 27445 12631
rect 27445 12597 27479 12631
rect 27479 12597 27488 12631
rect 27436 12588 27488 12597
rect 27528 12588 27580 12640
rect 10246 12486 10298 12538
rect 10310 12486 10362 12538
rect 10374 12486 10426 12538
rect 10438 12486 10490 12538
rect 19510 12486 19562 12538
rect 19574 12486 19626 12538
rect 19638 12486 19690 12538
rect 19702 12486 19754 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 2596 12384 2648 12436
rect 3240 12384 3292 12436
rect 4804 12384 4856 12436
rect 5908 12384 5960 12436
rect 8116 12384 8168 12436
rect 2688 12359 2740 12368
rect 2044 12248 2096 12300
rect 2320 12291 2372 12300
rect 2320 12257 2329 12291
rect 2329 12257 2363 12291
rect 2363 12257 2372 12291
rect 2320 12248 2372 12257
rect 2688 12325 2697 12359
rect 2697 12325 2731 12359
rect 2731 12325 2740 12359
rect 2688 12316 2740 12325
rect 4528 12316 4580 12368
rect 9588 12316 9640 12368
rect 1400 12180 1452 12232
rect 3332 12248 3384 12300
rect 3700 12248 3752 12300
rect 6368 12248 6420 12300
rect 7288 12248 7340 12300
rect 8208 12248 8260 12300
rect 9220 12291 9272 12300
rect 9220 12257 9229 12291
rect 9229 12257 9263 12291
rect 9263 12257 9272 12291
rect 9220 12248 9272 12257
rect 9864 12248 9916 12300
rect 11244 12316 11296 12368
rect 11336 12248 11388 12300
rect 2872 12180 2924 12232
rect 7380 12223 7432 12232
rect 3608 12155 3660 12164
rect 3608 12121 3617 12155
rect 3617 12121 3651 12155
rect 3651 12121 3660 12155
rect 3608 12112 3660 12121
rect 7380 12189 7389 12223
rect 7389 12189 7423 12223
rect 7423 12189 7432 12223
rect 7380 12180 7432 12189
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 9404 12180 9456 12232
rect 11612 12180 11664 12232
rect 13452 12384 13504 12436
rect 13820 12427 13872 12436
rect 13820 12393 13829 12427
rect 13829 12393 13863 12427
rect 13863 12393 13872 12427
rect 13820 12384 13872 12393
rect 14280 12384 14332 12436
rect 15752 12384 15804 12436
rect 18328 12384 18380 12436
rect 19248 12384 19300 12436
rect 12440 12180 12492 12232
rect 12808 12291 12860 12300
rect 12808 12257 12817 12291
rect 12817 12257 12851 12291
rect 12851 12257 12860 12291
rect 13636 12316 13688 12368
rect 12808 12248 12860 12257
rect 13084 12248 13136 12300
rect 13820 12248 13872 12300
rect 13912 12248 13964 12300
rect 15292 12316 15344 12368
rect 15844 12316 15896 12368
rect 17224 12316 17276 12368
rect 14464 12291 14516 12300
rect 13636 12180 13688 12232
rect 14464 12257 14473 12291
rect 14473 12257 14507 12291
rect 14507 12257 14516 12291
rect 14464 12248 14516 12257
rect 15384 12291 15436 12300
rect 15384 12257 15393 12291
rect 15393 12257 15427 12291
rect 15427 12257 15436 12291
rect 15384 12248 15436 12257
rect 15660 12248 15712 12300
rect 15292 12223 15344 12232
rect 15292 12189 15301 12223
rect 15301 12189 15335 12223
rect 15335 12189 15344 12223
rect 15292 12180 15344 12189
rect 16212 12180 16264 12232
rect 18604 12316 18656 12368
rect 19340 12316 19392 12368
rect 19984 12384 20036 12436
rect 20260 12359 20312 12368
rect 20260 12325 20269 12359
rect 20269 12325 20303 12359
rect 20303 12325 20312 12359
rect 20260 12316 20312 12325
rect 21088 12384 21140 12436
rect 22560 12384 22612 12436
rect 25412 12427 25464 12436
rect 25412 12393 25421 12427
rect 25421 12393 25455 12427
rect 25455 12393 25464 12427
rect 25412 12384 25464 12393
rect 26148 12384 26200 12436
rect 27528 12384 27580 12436
rect 21364 12316 21416 12368
rect 19248 12248 19300 12300
rect 21916 12248 21968 12300
rect 23388 12316 23440 12368
rect 23940 12248 23992 12300
rect 26700 12248 26752 12300
rect 18604 12180 18656 12232
rect 18972 12180 19024 12232
rect 20812 12180 20864 12232
rect 21180 12223 21232 12232
rect 21180 12189 21189 12223
rect 21189 12189 21223 12223
rect 21223 12189 21232 12223
rect 21180 12180 21232 12189
rect 3792 12044 3844 12096
rect 4988 12044 5040 12096
rect 5908 12044 5960 12096
rect 7288 12044 7340 12096
rect 7472 12044 7524 12096
rect 7748 12044 7800 12096
rect 8116 12044 8168 12096
rect 8208 12044 8260 12096
rect 9128 12044 9180 12096
rect 20536 12112 20588 12164
rect 23388 12180 23440 12232
rect 23848 12180 23900 12232
rect 24768 12180 24820 12232
rect 23296 12112 23348 12164
rect 25044 12112 25096 12164
rect 25228 12112 25280 12164
rect 26240 12180 26292 12232
rect 26424 12223 26476 12232
rect 26424 12189 26433 12223
rect 26433 12189 26467 12223
rect 26467 12189 26476 12223
rect 26424 12180 26476 12189
rect 9956 12044 10008 12096
rect 11244 12044 11296 12096
rect 21364 12044 21416 12096
rect 21456 12044 21508 12096
rect 25964 12044 26016 12096
rect 5614 11942 5666 11994
rect 5678 11942 5730 11994
rect 5742 11942 5794 11994
rect 5806 11942 5858 11994
rect 14878 11942 14930 11994
rect 14942 11942 14994 11994
rect 15006 11942 15058 11994
rect 15070 11942 15122 11994
rect 24142 11942 24194 11994
rect 24206 11942 24258 11994
rect 24270 11942 24322 11994
rect 24334 11942 24386 11994
rect 2872 11840 2924 11892
rect 6368 11883 6420 11892
rect 6368 11849 6377 11883
rect 6377 11849 6411 11883
rect 6411 11849 6420 11883
rect 6368 11840 6420 11849
rect 7656 11840 7708 11892
rect 9128 11840 9180 11892
rect 9588 11883 9640 11892
rect 9588 11849 9597 11883
rect 9597 11849 9631 11883
rect 9631 11849 9640 11883
rect 9588 11840 9640 11849
rect 11796 11840 11848 11892
rect 12072 11840 12124 11892
rect 20536 11883 20588 11892
rect 20536 11849 20545 11883
rect 20545 11849 20579 11883
rect 20579 11849 20588 11883
rect 20536 11840 20588 11849
rect 23388 11840 23440 11892
rect 25044 11840 25096 11892
rect 25228 11840 25280 11892
rect 27896 11840 27948 11892
rect 1492 11636 1544 11688
rect 2412 11679 2464 11688
rect 2412 11645 2421 11679
rect 2421 11645 2455 11679
rect 2455 11645 2464 11679
rect 2412 11636 2464 11645
rect 7472 11772 7524 11824
rect 7932 11772 7984 11824
rect 5080 11704 5132 11756
rect 6276 11704 6328 11756
rect 6460 11704 6512 11756
rect 8208 11704 8260 11756
rect 3976 11568 4028 11620
rect 2320 11500 2372 11552
rect 4528 11543 4580 11552
rect 4528 11509 4537 11543
rect 4537 11509 4571 11543
rect 4571 11509 4580 11543
rect 4528 11500 4580 11509
rect 4988 11568 5040 11620
rect 5172 11568 5224 11620
rect 8116 11636 8168 11688
rect 12624 11772 12676 11824
rect 14096 11772 14148 11824
rect 14740 11815 14792 11824
rect 14740 11781 14749 11815
rect 14749 11781 14783 11815
rect 14783 11781 14792 11815
rect 14740 11772 14792 11781
rect 22744 11772 22796 11824
rect 25596 11815 25648 11824
rect 25596 11781 25605 11815
rect 25605 11781 25639 11815
rect 25639 11781 25648 11815
rect 25596 11772 25648 11781
rect 9680 11704 9732 11756
rect 11244 11747 11296 11756
rect 11244 11713 11253 11747
rect 11253 11713 11287 11747
rect 11287 11713 11296 11747
rect 11244 11704 11296 11713
rect 11796 11704 11848 11756
rect 8484 11636 8536 11688
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 11520 11636 11572 11688
rect 11980 11636 12032 11688
rect 13912 11704 13964 11756
rect 21456 11747 21508 11756
rect 21456 11713 21465 11747
rect 21465 11713 21499 11747
rect 21499 11713 21508 11747
rect 21456 11704 21508 11713
rect 23296 11747 23348 11756
rect 23296 11713 23305 11747
rect 23305 11713 23339 11747
rect 23339 11713 23348 11747
rect 23296 11704 23348 11713
rect 26148 11704 26200 11756
rect 27804 11704 27856 11756
rect 28264 11704 28316 11756
rect 12900 11679 12952 11688
rect 12900 11645 12909 11679
rect 12909 11645 12943 11679
rect 12943 11645 12952 11679
rect 12900 11636 12952 11645
rect 13268 11636 13320 11688
rect 20720 11679 20772 11688
rect 20720 11645 20729 11679
rect 20729 11645 20763 11679
rect 20763 11645 20772 11679
rect 20720 11636 20772 11645
rect 20996 11679 21048 11688
rect 20996 11645 21005 11679
rect 21005 11645 21039 11679
rect 21039 11645 21048 11679
rect 20996 11636 21048 11645
rect 21364 11636 21416 11688
rect 22560 11636 22612 11688
rect 25412 11679 25464 11688
rect 5632 11543 5684 11552
rect 5632 11509 5641 11543
rect 5641 11509 5675 11543
rect 5675 11509 5684 11543
rect 5632 11500 5684 11509
rect 7656 11568 7708 11620
rect 10692 11568 10744 11620
rect 11336 11568 11388 11620
rect 25412 11645 25421 11679
rect 25421 11645 25455 11679
rect 25455 11645 25464 11679
rect 25412 11636 25464 11645
rect 25964 11636 26016 11688
rect 27436 11636 27488 11688
rect 8484 11543 8536 11552
rect 8484 11509 8493 11543
rect 8493 11509 8527 11543
rect 8527 11509 8536 11543
rect 8484 11500 8536 11509
rect 9312 11500 9364 11552
rect 9496 11500 9548 11552
rect 13452 11500 13504 11552
rect 14740 11500 14792 11552
rect 19248 11500 19300 11552
rect 20628 11500 20680 11552
rect 20904 11543 20956 11552
rect 20904 11509 20913 11543
rect 20913 11509 20947 11543
rect 20947 11509 20956 11543
rect 20904 11500 20956 11509
rect 22744 11500 22796 11552
rect 26516 11500 26568 11552
rect 10246 11398 10298 11450
rect 10310 11398 10362 11450
rect 10374 11398 10426 11450
rect 10438 11398 10490 11450
rect 19510 11398 19562 11450
rect 19574 11398 19626 11450
rect 19638 11398 19690 11450
rect 19702 11398 19754 11450
rect 5632 11228 5684 11280
rect 8484 11296 8536 11348
rect 9312 11296 9364 11348
rect 10692 11296 10744 11348
rect 12900 11296 12952 11348
rect 12992 11296 13044 11348
rect 13636 11296 13688 11348
rect 13728 11228 13780 11280
rect 1952 11203 2004 11212
rect 1952 11169 1961 11203
rect 1961 11169 1995 11203
rect 1995 11169 2004 11203
rect 1952 11160 2004 11169
rect 2780 11160 2832 11212
rect 3240 11203 3292 11212
rect 3240 11169 3249 11203
rect 3249 11169 3283 11203
rect 3283 11169 3292 11203
rect 3240 11160 3292 11169
rect 3148 11092 3200 11144
rect 3516 11203 3568 11212
rect 3516 11169 3525 11203
rect 3525 11169 3559 11203
rect 3559 11169 3568 11203
rect 3976 11203 4028 11212
rect 3516 11160 3568 11169
rect 3976 11169 3985 11203
rect 3985 11169 4019 11203
rect 4019 11169 4028 11203
rect 3976 11160 4028 11169
rect 5356 11160 5408 11212
rect 7472 11160 7524 11212
rect 8208 11203 8260 11212
rect 8208 11169 8217 11203
rect 8217 11169 8251 11203
rect 8251 11169 8260 11203
rect 8208 11160 8260 11169
rect 9864 11203 9916 11212
rect 9864 11169 9873 11203
rect 9873 11169 9907 11203
rect 9907 11169 9916 11203
rect 9864 11160 9916 11169
rect 5264 11092 5316 11144
rect 10048 11135 10100 11144
rect 10048 11101 10057 11135
rect 10057 11101 10091 11135
rect 10091 11101 10100 11135
rect 10048 11092 10100 11101
rect 3056 11067 3108 11076
rect 3056 11033 3065 11067
rect 3065 11033 3099 11067
rect 3099 11033 3108 11067
rect 3056 11024 3108 11033
rect 5080 11024 5132 11076
rect 6000 11024 6052 11076
rect 11796 11092 11848 11144
rect 13912 11160 13964 11212
rect 18052 11203 18104 11212
rect 18052 11169 18061 11203
rect 18061 11169 18095 11203
rect 18095 11169 18104 11203
rect 18052 11160 18104 11169
rect 14740 11092 14792 11144
rect 18880 11296 18932 11348
rect 20168 11296 20220 11348
rect 24860 11296 24912 11348
rect 19800 11228 19852 11280
rect 20628 11228 20680 11280
rect 18696 11160 18748 11212
rect 21272 11160 21324 11212
rect 25688 11160 25740 11212
rect 26148 11203 26200 11212
rect 26148 11169 26157 11203
rect 26157 11169 26191 11203
rect 26191 11169 26200 11203
rect 26148 11160 26200 11169
rect 19156 11135 19208 11144
rect 7288 10956 7340 11008
rect 7656 10956 7708 11008
rect 9588 10956 9640 11008
rect 9772 10956 9824 11008
rect 17592 11024 17644 11076
rect 19156 11101 19165 11135
rect 19165 11101 19199 11135
rect 19199 11101 19208 11135
rect 19156 11092 19208 11101
rect 19892 11092 19944 11144
rect 20168 11092 20220 11144
rect 23572 11135 23624 11144
rect 23572 11101 23581 11135
rect 23581 11101 23615 11135
rect 23615 11101 23624 11135
rect 23572 11092 23624 11101
rect 23848 11092 23900 11144
rect 24032 11135 24084 11144
rect 24032 11101 24041 11135
rect 24041 11101 24075 11135
rect 24075 11101 24084 11135
rect 24032 11092 24084 11101
rect 24768 11092 24820 11144
rect 18696 11024 18748 11076
rect 19064 11067 19116 11076
rect 19064 11033 19073 11067
rect 19073 11033 19107 11067
rect 19107 11033 19116 11067
rect 19064 11024 19116 11033
rect 25136 11135 25188 11144
rect 25136 11101 25145 11135
rect 25145 11101 25179 11135
rect 25179 11101 25188 11135
rect 25136 11092 25188 11101
rect 25320 11024 25372 11076
rect 26884 11067 26936 11076
rect 26884 11033 26893 11067
rect 26893 11033 26927 11067
rect 26927 11033 26936 11067
rect 26884 11024 26936 11033
rect 27528 11024 27580 11076
rect 29000 11067 29052 11076
rect 29000 11033 29009 11067
rect 29009 11033 29043 11067
rect 29043 11033 29052 11067
rect 29000 11024 29052 11033
rect 22560 10956 22612 11008
rect 24676 10999 24728 11008
rect 24676 10965 24685 10999
rect 24685 10965 24719 10999
rect 24719 10965 24728 10999
rect 24676 10956 24728 10965
rect 5614 10854 5666 10906
rect 5678 10854 5730 10906
rect 5742 10854 5794 10906
rect 5806 10854 5858 10906
rect 14878 10854 14930 10906
rect 14942 10854 14994 10906
rect 15006 10854 15058 10906
rect 15070 10854 15122 10906
rect 24142 10854 24194 10906
rect 24206 10854 24258 10906
rect 24270 10854 24322 10906
rect 24334 10854 24386 10906
rect 2228 10752 2280 10804
rect 2964 10752 3016 10804
rect 3976 10752 4028 10804
rect 2872 10727 2924 10736
rect 2872 10693 2881 10727
rect 2881 10693 2915 10727
rect 2915 10693 2924 10727
rect 2872 10684 2924 10693
rect 2136 10616 2188 10668
rect 4344 10616 4396 10668
rect 9772 10752 9824 10804
rect 9864 10752 9916 10804
rect 6276 10616 6328 10668
rect 2872 10548 2924 10600
rect 4712 10548 4764 10600
rect 5356 10480 5408 10532
rect 8300 10480 8352 10532
rect 9772 10591 9824 10600
rect 9772 10557 9806 10591
rect 9806 10557 9824 10591
rect 9772 10548 9824 10557
rect 13452 10752 13504 10804
rect 17040 10752 17092 10804
rect 18972 10752 19024 10804
rect 19156 10752 19208 10804
rect 24032 10752 24084 10804
rect 24492 10752 24544 10804
rect 25136 10752 25188 10804
rect 12992 10684 13044 10736
rect 12624 10548 12676 10600
rect 16120 10616 16172 10668
rect 12992 10591 13044 10600
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 12992 10548 13044 10557
rect 13452 10548 13504 10600
rect 15568 10548 15620 10600
rect 17684 10548 17736 10600
rect 22100 10616 22152 10668
rect 23572 10659 23624 10668
rect 23572 10625 23581 10659
rect 23581 10625 23615 10659
rect 23615 10625 23624 10659
rect 23572 10616 23624 10625
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 23940 10616 23992 10625
rect 18420 10548 18472 10600
rect 4804 10455 4856 10464
rect 4804 10421 4813 10455
rect 4813 10421 4847 10455
rect 4847 10421 4856 10455
rect 4804 10412 4856 10421
rect 12072 10480 12124 10532
rect 15200 10480 15252 10532
rect 15936 10480 15988 10532
rect 17132 10523 17184 10532
rect 17132 10489 17141 10523
rect 17141 10489 17175 10523
rect 17175 10489 17184 10523
rect 17132 10480 17184 10489
rect 21180 10480 21232 10532
rect 21548 10480 21600 10532
rect 22284 10548 22336 10600
rect 22928 10548 22980 10600
rect 22652 10480 22704 10532
rect 23940 10480 23992 10532
rect 25872 10684 25924 10736
rect 25320 10616 25372 10668
rect 25504 10616 25556 10668
rect 25964 10616 26016 10668
rect 25412 10548 25464 10600
rect 27988 10480 28040 10532
rect 12532 10455 12584 10464
rect 12532 10421 12541 10455
rect 12541 10421 12575 10455
rect 12575 10421 12584 10455
rect 12532 10412 12584 10421
rect 15568 10412 15620 10464
rect 16212 10455 16264 10464
rect 16212 10421 16221 10455
rect 16221 10421 16255 10455
rect 16255 10421 16264 10455
rect 16212 10412 16264 10421
rect 17684 10412 17736 10464
rect 18236 10455 18288 10464
rect 18236 10421 18245 10455
rect 18245 10421 18279 10455
rect 18279 10421 18288 10455
rect 18236 10412 18288 10421
rect 19800 10412 19852 10464
rect 21916 10412 21968 10464
rect 22560 10455 22612 10464
rect 22560 10421 22569 10455
rect 22569 10421 22603 10455
rect 22603 10421 22612 10455
rect 22560 10412 22612 10421
rect 23848 10455 23900 10464
rect 23848 10421 23857 10455
rect 23857 10421 23891 10455
rect 23891 10421 23900 10455
rect 23848 10412 23900 10421
rect 26240 10455 26292 10464
rect 26240 10421 26249 10455
rect 26249 10421 26283 10455
rect 26283 10421 26292 10455
rect 26240 10412 26292 10421
rect 28264 10412 28316 10464
rect 10246 10310 10298 10362
rect 10310 10310 10362 10362
rect 10374 10310 10426 10362
rect 10438 10310 10490 10362
rect 19510 10310 19562 10362
rect 19574 10310 19626 10362
rect 19638 10310 19690 10362
rect 19702 10310 19754 10362
rect 2688 10208 2740 10260
rect 2780 10208 2832 10260
rect 3700 10208 3752 10260
rect 1584 10115 1636 10124
rect 1584 10081 1593 10115
rect 1593 10081 1627 10115
rect 1627 10081 1636 10115
rect 1584 10072 1636 10081
rect 2136 10140 2188 10192
rect 9220 10251 9272 10260
rect 9220 10217 9229 10251
rect 9229 10217 9263 10251
rect 9263 10217 9272 10251
rect 9220 10208 9272 10217
rect 12072 10208 12124 10260
rect 15200 10208 15252 10260
rect 15568 10208 15620 10260
rect 16028 10208 16080 10260
rect 16580 10208 16632 10260
rect 18052 10208 18104 10260
rect 18144 10208 18196 10260
rect 25872 10208 25924 10260
rect 28080 10251 28132 10260
rect 28080 10217 28089 10251
rect 28089 10217 28123 10251
rect 28123 10217 28132 10251
rect 28080 10208 28132 10217
rect 7104 10183 7156 10192
rect 7104 10149 7113 10183
rect 7113 10149 7147 10183
rect 7147 10149 7156 10183
rect 7104 10140 7156 10149
rect 2228 10115 2280 10124
rect 2228 10081 2237 10115
rect 2237 10081 2271 10115
rect 2271 10081 2280 10115
rect 2228 10072 2280 10081
rect 2964 10115 3016 10124
rect 2964 10081 2973 10115
rect 2973 10081 3007 10115
rect 3007 10081 3016 10115
rect 2964 10072 3016 10081
rect 3240 10072 3292 10124
rect 3516 10072 3568 10124
rect 4804 10072 4856 10124
rect 6184 10072 6236 10124
rect 7288 10072 7340 10124
rect 8208 10140 8260 10192
rect 12532 10140 12584 10192
rect 7840 10072 7892 10124
rect 9036 10115 9088 10124
rect 9036 10081 9045 10115
rect 9045 10081 9079 10115
rect 9079 10081 9088 10115
rect 9036 10072 9088 10081
rect 9312 10072 9364 10124
rect 14096 10072 14148 10124
rect 17040 10072 17092 10124
rect 4252 10004 4304 10056
rect 12164 10004 12216 10056
rect 17868 10004 17920 10056
rect 7472 9936 7524 9988
rect 15108 9936 15160 9988
rect 18420 10140 18472 10192
rect 19156 10140 19208 10192
rect 23388 10140 23440 10192
rect 23940 10140 23992 10192
rect 18880 10115 18932 10124
rect 18880 10081 18889 10115
rect 18889 10081 18923 10115
rect 18923 10081 18932 10115
rect 18880 10072 18932 10081
rect 19248 10072 19300 10124
rect 19800 10072 19852 10124
rect 20720 10115 20772 10124
rect 18604 10004 18656 10056
rect 20720 10081 20729 10115
rect 20729 10081 20763 10115
rect 20763 10081 20772 10115
rect 20720 10072 20772 10081
rect 21088 10115 21140 10124
rect 21088 10081 21097 10115
rect 21097 10081 21131 10115
rect 21131 10081 21140 10115
rect 21088 10072 21140 10081
rect 21180 10072 21232 10124
rect 20812 10047 20864 10056
rect 20812 10013 20821 10047
rect 20821 10013 20855 10047
rect 20855 10013 20864 10047
rect 20812 10004 20864 10013
rect 7656 9868 7708 9920
rect 12624 9868 12676 9920
rect 20444 9868 20496 9920
rect 20812 9868 20864 9920
rect 23572 10072 23624 10124
rect 23848 10072 23900 10124
rect 24676 10140 24728 10192
rect 25504 10072 25556 10124
rect 28356 10072 28408 10124
rect 24768 10047 24820 10056
rect 24768 10013 24777 10047
rect 24777 10013 24811 10047
rect 24811 10013 24820 10047
rect 24768 10004 24820 10013
rect 27896 9868 27948 9920
rect 5614 9766 5666 9818
rect 5678 9766 5730 9818
rect 5742 9766 5794 9818
rect 5806 9766 5858 9818
rect 14878 9766 14930 9818
rect 14942 9766 14994 9818
rect 15006 9766 15058 9818
rect 15070 9766 15122 9818
rect 24142 9766 24194 9818
rect 24206 9766 24258 9818
rect 24270 9766 24322 9818
rect 24334 9766 24386 9818
rect 2872 9707 2924 9716
rect 2872 9673 2881 9707
rect 2881 9673 2915 9707
rect 2915 9673 2924 9707
rect 2872 9664 2924 9673
rect 5356 9664 5408 9716
rect 13452 9664 13504 9716
rect 15568 9664 15620 9716
rect 16212 9664 16264 9716
rect 16580 9664 16632 9716
rect 21916 9707 21968 9716
rect 7472 9596 7524 9648
rect 10600 9596 10652 9648
rect 1400 9528 1452 9580
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 11796 9571 11848 9580
rect 11796 9537 11805 9571
rect 11805 9537 11839 9571
rect 11839 9537 11848 9571
rect 11796 9528 11848 9537
rect 12256 9528 12308 9580
rect 2412 9460 2464 9512
rect 3056 9460 3108 9512
rect 4896 9460 4948 9512
rect 2044 9392 2096 9444
rect 2320 9435 2372 9444
rect 2320 9401 2329 9435
rect 2329 9401 2363 9435
rect 2363 9401 2372 9435
rect 2320 9392 2372 9401
rect 2964 9392 3016 9444
rect 3700 9392 3752 9444
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 3424 9324 3476 9376
rect 4528 9367 4580 9376
rect 4528 9333 4537 9367
rect 4537 9333 4571 9367
rect 4571 9333 4580 9367
rect 4528 9324 4580 9333
rect 4896 9324 4948 9376
rect 6184 9460 6236 9512
rect 6828 9392 6880 9444
rect 7380 9460 7432 9512
rect 10784 9460 10836 9512
rect 11704 9460 11756 9512
rect 14188 9460 14240 9512
rect 11520 9435 11572 9444
rect 6920 9324 6972 9376
rect 7196 9324 7248 9376
rect 11520 9401 11529 9435
rect 11529 9401 11563 9435
rect 11563 9401 11572 9435
rect 11520 9392 11572 9401
rect 12072 9392 12124 9444
rect 14464 9392 14516 9444
rect 14740 9460 14792 9512
rect 16764 9528 16816 9580
rect 21916 9673 21925 9707
rect 21925 9673 21959 9707
rect 21959 9673 21968 9707
rect 21916 9664 21968 9673
rect 23388 9571 23440 9580
rect 17592 9503 17644 9512
rect 17592 9469 17626 9503
rect 17626 9469 17644 9503
rect 16396 9392 16448 9444
rect 17132 9392 17184 9444
rect 17592 9460 17644 9469
rect 19892 9460 19944 9512
rect 23388 9537 23397 9571
rect 23397 9537 23431 9571
rect 23431 9537 23440 9571
rect 23388 9528 23440 9537
rect 23572 9571 23624 9580
rect 23572 9537 23581 9571
rect 23581 9537 23615 9571
rect 23615 9537 23624 9571
rect 23572 9528 23624 9537
rect 25596 9528 25648 9580
rect 26424 9596 26476 9648
rect 26056 9528 26108 9580
rect 21824 9503 21876 9512
rect 21824 9469 21833 9503
rect 21833 9469 21867 9503
rect 21867 9469 21876 9503
rect 21824 9460 21876 9469
rect 22652 9460 22704 9512
rect 26240 9460 26292 9512
rect 26608 9503 26660 9512
rect 26608 9469 26617 9503
rect 26617 9469 26651 9503
rect 26651 9469 26660 9503
rect 26608 9460 26660 9469
rect 27160 9503 27212 9512
rect 27160 9469 27169 9503
rect 27169 9469 27203 9503
rect 27203 9469 27212 9503
rect 27436 9503 27488 9512
rect 27160 9460 27212 9469
rect 27436 9469 27445 9503
rect 27445 9469 27479 9503
rect 27479 9469 27488 9503
rect 27436 9460 27488 9469
rect 19064 9392 19116 9444
rect 20904 9392 20956 9444
rect 11060 9324 11112 9376
rect 11612 9367 11664 9376
rect 11612 9333 11621 9367
rect 11621 9333 11655 9367
rect 11655 9333 11664 9367
rect 11612 9324 11664 9333
rect 11796 9324 11848 9376
rect 14280 9324 14332 9376
rect 15476 9324 15528 9376
rect 15936 9324 15988 9376
rect 18696 9367 18748 9376
rect 18696 9333 18705 9367
rect 18705 9333 18739 9367
rect 18739 9333 18748 9367
rect 18696 9324 18748 9333
rect 19340 9324 19392 9376
rect 21824 9324 21876 9376
rect 10246 9222 10298 9274
rect 10310 9222 10362 9274
rect 10374 9222 10426 9274
rect 10438 9222 10490 9274
rect 19510 9222 19562 9274
rect 19574 9222 19626 9274
rect 19638 9222 19690 9274
rect 19702 9222 19754 9274
rect 3148 9120 3200 9172
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 1860 9095 1912 9104
rect 1860 9061 1869 9095
rect 1869 9061 1903 9095
rect 1903 9061 1912 9095
rect 1860 9052 1912 9061
rect 3056 8984 3108 9036
rect 3424 8984 3476 9036
rect 4436 9120 4488 9172
rect 6828 9163 6880 9172
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 7472 9120 7524 9172
rect 11612 9120 11664 9172
rect 4344 9095 4396 9104
rect 4344 9061 4353 9095
rect 4353 9061 4387 9095
rect 4387 9061 4396 9095
rect 25872 9163 25924 9172
rect 25872 9129 25881 9163
rect 25881 9129 25915 9163
rect 25915 9129 25924 9163
rect 25872 9120 25924 9129
rect 14372 9095 14424 9104
rect 4344 9052 4396 9061
rect 3700 8984 3752 9036
rect 3240 8916 3292 8968
rect 6920 8984 6972 9036
rect 8300 8984 8352 9036
rect 8760 9027 8812 9036
rect 8760 8993 8769 9027
rect 8769 8993 8803 9027
rect 8803 8993 8812 9027
rect 8760 8984 8812 8993
rect 9864 8984 9916 9036
rect 7564 8916 7616 8968
rect 7840 8916 7892 8968
rect 9496 8916 9548 8968
rect 11060 8916 11112 8968
rect 12624 8984 12676 9036
rect 13084 8984 13136 9036
rect 14372 9061 14381 9095
rect 14381 9061 14415 9095
rect 14415 9061 14424 9095
rect 14372 9052 14424 9061
rect 15200 9095 15252 9104
rect 15200 9061 15209 9095
rect 15209 9061 15243 9095
rect 15243 9061 15252 9095
rect 15200 9052 15252 9061
rect 20720 9052 20772 9104
rect 22652 9095 22704 9104
rect 22652 9061 22661 9095
rect 22661 9061 22695 9095
rect 22695 9061 22704 9095
rect 22652 9052 22704 9061
rect 28264 9120 28316 9172
rect 26424 9052 26476 9104
rect 26792 9095 26844 9104
rect 26792 9061 26801 9095
rect 26801 9061 26835 9095
rect 26835 9061 26844 9095
rect 26792 9052 26844 9061
rect 27896 9052 27948 9104
rect 13360 8916 13412 8968
rect 14464 8984 14516 9036
rect 16028 9027 16080 9036
rect 15108 8916 15160 8968
rect 15476 8959 15528 8968
rect 15476 8925 15485 8959
rect 15485 8925 15519 8959
rect 15519 8925 15528 8959
rect 15476 8916 15528 8925
rect 16028 8993 16037 9027
rect 16037 8993 16071 9027
rect 16071 8993 16080 9027
rect 16028 8984 16080 8993
rect 20444 9027 20496 9036
rect 20444 8993 20453 9027
rect 20453 8993 20487 9027
rect 20487 8993 20496 9027
rect 20444 8984 20496 8993
rect 17684 8916 17736 8968
rect 23388 8984 23440 9036
rect 22744 8916 22796 8968
rect 26976 8984 27028 9036
rect 24860 8916 24912 8968
rect 25596 8916 25648 8968
rect 2320 8780 2372 8832
rect 5908 8780 5960 8832
rect 7840 8780 7892 8832
rect 8392 8780 8444 8832
rect 8576 8780 8628 8832
rect 10140 8780 10192 8832
rect 18144 8848 18196 8900
rect 23848 8848 23900 8900
rect 24952 8891 25004 8900
rect 24952 8857 24961 8891
rect 24961 8857 24995 8891
rect 24995 8857 25004 8891
rect 24952 8848 25004 8857
rect 25412 8891 25464 8900
rect 25412 8857 25421 8891
rect 25421 8857 25455 8891
rect 25455 8857 25464 8891
rect 25412 8848 25464 8857
rect 16120 8823 16172 8832
rect 16120 8789 16129 8823
rect 16129 8789 16163 8823
rect 16163 8789 16172 8823
rect 16120 8780 16172 8789
rect 24860 8780 24912 8832
rect 26056 8780 26108 8832
rect 27528 8780 27580 8832
rect 28080 8823 28132 8832
rect 28080 8789 28089 8823
rect 28089 8789 28123 8823
rect 28123 8789 28132 8823
rect 28080 8780 28132 8789
rect 5614 8678 5666 8730
rect 5678 8678 5730 8730
rect 5742 8678 5794 8730
rect 5806 8678 5858 8730
rect 14878 8678 14930 8730
rect 14942 8678 14994 8730
rect 15006 8678 15058 8730
rect 15070 8678 15122 8730
rect 24142 8678 24194 8730
rect 24206 8678 24258 8730
rect 24270 8678 24322 8730
rect 24334 8678 24386 8730
rect 2412 8576 2464 8628
rect 3056 8619 3108 8628
rect 3056 8585 3065 8619
rect 3065 8585 3099 8619
rect 3099 8585 3108 8619
rect 3056 8576 3108 8585
rect 4068 8508 4120 8560
rect 4896 8576 4948 8628
rect 5264 8576 5316 8628
rect 12072 8576 12124 8628
rect 12348 8576 12400 8628
rect 13176 8576 13228 8628
rect 13360 8619 13412 8628
rect 13360 8585 13369 8619
rect 13369 8585 13403 8619
rect 13403 8585 13412 8619
rect 13360 8576 13412 8585
rect 14740 8576 14792 8628
rect 26976 8619 27028 8628
rect 26976 8585 26985 8619
rect 26985 8585 27019 8619
rect 27019 8585 27028 8619
rect 26976 8576 27028 8585
rect 27988 8576 28040 8628
rect 6000 8508 6052 8560
rect 9496 8508 9548 8560
rect 9864 8508 9916 8560
rect 10876 8508 10928 8560
rect 10968 8440 11020 8492
rect 1952 8415 2004 8424
rect 1952 8381 1961 8415
rect 1961 8381 1995 8415
rect 1995 8381 2004 8415
rect 1952 8372 2004 8381
rect 2412 8415 2464 8424
rect 2412 8381 2421 8415
rect 2421 8381 2455 8415
rect 2455 8381 2464 8415
rect 2412 8372 2464 8381
rect 3240 8415 3292 8424
rect 3240 8381 3249 8415
rect 3249 8381 3283 8415
rect 3283 8381 3292 8415
rect 3240 8372 3292 8381
rect 4528 8415 4580 8424
rect 4528 8381 4562 8415
rect 4562 8381 4580 8415
rect 4528 8372 4580 8381
rect 11520 8372 11572 8424
rect 2320 8304 2372 8356
rect 18236 8508 18288 8560
rect 13084 8440 13136 8492
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 21824 8440 21876 8492
rect 12900 8372 12952 8424
rect 14740 8415 14792 8424
rect 14740 8381 14749 8415
rect 14749 8381 14783 8415
rect 14783 8381 14792 8415
rect 14740 8372 14792 8381
rect 16212 8415 16264 8424
rect 16212 8381 16221 8415
rect 16221 8381 16255 8415
rect 16255 8381 16264 8415
rect 16212 8372 16264 8381
rect 16396 8415 16448 8424
rect 16396 8381 16405 8415
rect 16405 8381 16439 8415
rect 16439 8381 16448 8415
rect 16396 8372 16448 8381
rect 24768 8372 24820 8424
rect 26608 8440 26660 8492
rect 27160 8440 27212 8492
rect 27528 8483 27580 8492
rect 27528 8449 27537 8483
rect 27537 8449 27571 8483
rect 27571 8449 27580 8483
rect 27528 8440 27580 8449
rect 28172 8440 28224 8492
rect 25872 8415 25924 8424
rect 25872 8381 25881 8415
rect 25881 8381 25915 8415
rect 25915 8381 25924 8415
rect 25872 8372 25924 8381
rect 26240 8372 26292 8424
rect 27436 8372 27488 8424
rect 28264 8372 28316 8424
rect 12072 8304 12124 8356
rect 12348 8347 12400 8356
rect 12348 8313 12357 8347
rect 12357 8313 12391 8347
rect 12391 8313 12400 8347
rect 12348 8304 12400 8313
rect 15476 8304 15528 8356
rect 6552 8236 6604 8288
rect 9312 8236 9364 8288
rect 9496 8279 9548 8288
rect 9496 8245 9505 8279
rect 9505 8245 9539 8279
rect 9539 8245 9548 8279
rect 9496 8236 9548 8245
rect 9864 8279 9916 8288
rect 9864 8245 9873 8279
rect 9873 8245 9907 8279
rect 9907 8245 9916 8279
rect 9864 8236 9916 8245
rect 9956 8236 10008 8288
rect 13728 8236 13780 8288
rect 19892 8236 19944 8288
rect 20168 8236 20220 8288
rect 25596 8236 25648 8288
rect 26792 8236 26844 8288
rect 10246 8134 10298 8186
rect 10310 8134 10362 8186
rect 10374 8134 10426 8186
rect 10438 8134 10490 8186
rect 19510 8134 19562 8186
rect 19574 8134 19626 8186
rect 19638 8134 19690 8186
rect 19702 8134 19754 8186
rect 2688 8032 2740 8084
rect 2964 8032 3016 8084
rect 4068 8032 4120 8084
rect 8760 8032 8812 8084
rect 9496 8032 9548 8084
rect 12072 8075 12124 8084
rect 12072 8041 12081 8075
rect 12081 8041 12115 8075
rect 12115 8041 12124 8075
rect 12072 8032 12124 8041
rect 12624 8032 12676 8084
rect 13084 8032 13136 8084
rect 14740 8032 14792 8084
rect 16028 8032 16080 8084
rect 16672 8032 16724 8084
rect 16856 8032 16908 8084
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4252 7964 4304 7973
rect 5908 7964 5960 8016
rect 9312 7964 9364 8016
rect 10232 7964 10284 8016
rect 10416 8007 10468 8016
rect 10416 7973 10425 8007
rect 10425 7973 10459 8007
rect 10459 7973 10468 8007
rect 10416 7964 10468 7973
rect 1492 7896 1544 7948
rect 2412 7939 2464 7948
rect 2412 7905 2421 7939
rect 2421 7905 2455 7939
rect 2455 7905 2464 7939
rect 2412 7896 2464 7905
rect 2872 7896 2924 7948
rect 6828 7939 6880 7948
rect 6828 7905 6837 7939
rect 6837 7905 6871 7939
rect 6871 7905 6880 7939
rect 6828 7896 6880 7905
rect 7932 7939 7984 7948
rect 7932 7905 7941 7939
rect 7941 7905 7975 7939
rect 7975 7905 7984 7939
rect 7932 7896 7984 7905
rect 8116 7939 8168 7948
rect 8116 7905 8125 7939
rect 8125 7905 8159 7939
rect 8159 7905 8168 7939
rect 8116 7896 8168 7905
rect 17224 8032 17276 8084
rect 17040 7964 17092 8016
rect 18512 7964 18564 8016
rect 18696 8032 18748 8084
rect 25964 8007 26016 8016
rect 10692 7896 10744 7948
rect 12532 7939 12584 7948
rect 12532 7905 12541 7939
rect 12541 7905 12575 7939
rect 12575 7905 12584 7939
rect 16028 7939 16080 7948
rect 12532 7896 12584 7905
rect 16028 7905 16037 7939
rect 16037 7905 16071 7939
rect 16071 7905 16080 7939
rect 16028 7896 16080 7905
rect 18696 7939 18748 7948
rect 18696 7905 18705 7939
rect 18705 7905 18739 7939
rect 18739 7905 18748 7939
rect 18696 7896 18748 7905
rect 19340 7939 19392 7948
rect 19340 7905 19349 7939
rect 19349 7905 19383 7939
rect 19383 7905 19392 7939
rect 19340 7896 19392 7905
rect 19892 7896 19944 7948
rect 20720 7939 20772 7948
rect 20720 7905 20729 7939
rect 20729 7905 20763 7939
rect 20763 7905 20772 7939
rect 20720 7896 20772 7905
rect 21088 7896 21140 7948
rect 22928 7939 22980 7948
rect 22928 7905 22937 7939
rect 22937 7905 22971 7939
rect 22971 7905 22980 7939
rect 22928 7896 22980 7905
rect 23388 7896 23440 7948
rect 25596 7896 25648 7948
rect 25964 7973 25973 8007
rect 25973 7973 26007 8007
rect 26007 7973 26016 8007
rect 25964 7964 26016 7973
rect 26148 8007 26200 8016
rect 26148 7973 26157 8007
rect 26157 7973 26191 8007
rect 26191 7973 26200 8007
rect 26148 7964 26200 7973
rect 9404 7828 9456 7880
rect 10324 7871 10376 7880
rect 5540 7760 5592 7812
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 13084 7828 13136 7880
rect 14280 7828 14332 7880
rect 16488 7828 16540 7880
rect 17776 7871 17828 7880
rect 17776 7837 17785 7871
rect 17785 7837 17819 7871
rect 17819 7837 17828 7871
rect 17776 7828 17828 7837
rect 18972 7828 19024 7880
rect 23020 7871 23072 7880
rect 6276 7692 6328 7744
rect 7380 7692 7432 7744
rect 8208 7692 8260 7744
rect 9680 7692 9732 7744
rect 15568 7760 15620 7812
rect 17868 7760 17920 7812
rect 20996 7760 21048 7812
rect 23020 7837 23029 7871
rect 23029 7837 23063 7871
rect 23063 7837 23072 7871
rect 23020 7828 23072 7837
rect 23112 7871 23164 7880
rect 23112 7837 23121 7871
rect 23121 7837 23155 7871
rect 23155 7837 23164 7871
rect 23848 7871 23900 7880
rect 23112 7828 23164 7837
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 23848 7828 23900 7837
rect 22468 7760 22520 7812
rect 28356 7828 28408 7880
rect 28172 7803 28224 7812
rect 28172 7769 28181 7803
rect 28181 7769 28215 7803
rect 28215 7769 28224 7803
rect 28172 7760 28224 7769
rect 10784 7692 10836 7744
rect 18696 7692 18748 7744
rect 18880 7692 18932 7744
rect 19340 7692 19392 7744
rect 22560 7735 22612 7744
rect 22560 7701 22569 7735
rect 22569 7701 22603 7735
rect 22603 7701 22612 7735
rect 22560 7692 22612 7701
rect 25964 7692 26016 7744
rect 26792 7735 26844 7744
rect 26792 7701 26801 7735
rect 26801 7701 26835 7735
rect 26835 7701 26844 7735
rect 26792 7692 26844 7701
rect 5614 7590 5666 7642
rect 5678 7590 5730 7642
rect 5742 7590 5794 7642
rect 5806 7590 5858 7642
rect 14878 7590 14930 7642
rect 14942 7590 14994 7642
rect 15006 7590 15058 7642
rect 15070 7590 15122 7642
rect 24142 7590 24194 7642
rect 24206 7590 24258 7642
rect 24270 7590 24322 7642
rect 24334 7590 24386 7642
rect 6828 7488 6880 7540
rect 7932 7488 7984 7540
rect 8392 7488 8444 7540
rect 9864 7488 9916 7540
rect 10416 7531 10468 7540
rect 10416 7497 10425 7531
rect 10425 7497 10459 7531
rect 10459 7497 10468 7531
rect 10416 7488 10468 7497
rect 14004 7488 14056 7540
rect 16212 7488 16264 7540
rect 18512 7531 18564 7540
rect 18512 7497 18521 7531
rect 18521 7497 18555 7531
rect 18555 7497 18564 7531
rect 18512 7488 18564 7497
rect 20812 7488 20864 7540
rect 23388 7488 23440 7540
rect 5356 7420 5408 7472
rect 11612 7420 11664 7472
rect 5816 7352 5868 7404
rect 6000 7352 6052 7404
rect 1860 7284 1912 7336
rect 3056 7327 3108 7336
rect 3056 7293 3065 7327
rect 3065 7293 3099 7327
rect 3099 7293 3108 7327
rect 3056 7284 3108 7293
rect 5264 7284 5316 7336
rect 5908 7284 5960 7336
rect 6644 7284 6696 7336
rect 10784 7352 10836 7404
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 9496 7327 9548 7336
rect 9496 7293 9505 7327
rect 9505 7293 9539 7327
rect 9539 7293 9548 7327
rect 9496 7284 9548 7293
rect 11612 7327 11664 7336
rect 1584 7148 1636 7200
rect 5540 7216 5592 7268
rect 11612 7293 11621 7327
rect 11621 7293 11655 7327
rect 11655 7293 11664 7327
rect 11612 7284 11664 7293
rect 13452 7327 13504 7336
rect 13452 7293 13461 7327
rect 13461 7293 13495 7327
rect 13495 7293 13504 7327
rect 13452 7284 13504 7293
rect 15016 7327 15068 7336
rect 15016 7293 15025 7327
rect 15025 7293 15059 7327
rect 15059 7293 15068 7327
rect 15016 7284 15068 7293
rect 15752 7420 15804 7472
rect 16488 7395 16540 7404
rect 16488 7361 16497 7395
rect 16497 7361 16531 7395
rect 16531 7361 16540 7395
rect 16488 7352 16540 7361
rect 17132 7395 17184 7404
rect 17132 7361 17141 7395
rect 17141 7361 17175 7395
rect 17175 7361 17184 7395
rect 17132 7352 17184 7361
rect 22100 7352 22152 7404
rect 28356 7352 28408 7404
rect 6736 7191 6788 7200
rect 6736 7157 6745 7191
rect 6745 7157 6779 7191
rect 6779 7157 6788 7191
rect 6736 7148 6788 7157
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 7380 7148 7432 7200
rect 9956 7148 10008 7200
rect 11336 7148 11388 7200
rect 14740 7191 14792 7200
rect 14740 7157 14749 7191
rect 14749 7157 14783 7191
rect 14783 7157 14792 7191
rect 14740 7148 14792 7157
rect 14832 7148 14884 7200
rect 15384 7327 15436 7336
rect 15384 7293 15393 7327
rect 15393 7293 15427 7327
rect 15427 7293 15436 7327
rect 20536 7327 20588 7336
rect 15384 7284 15436 7293
rect 20536 7293 20545 7327
rect 20545 7293 20579 7327
rect 20579 7293 20588 7327
rect 20536 7284 20588 7293
rect 20904 7284 20956 7336
rect 22284 7284 22336 7336
rect 24492 7284 24544 7336
rect 25412 7284 25464 7336
rect 15476 7148 15528 7200
rect 17316 7216 17368 7268
rect 19340 7216 19392 7268
rect 23112 7216 23164 7268
rect 25688 7216 25740 7268
rect 20076 7148 20128 7200
rect 22468 7191 22520 7200
rect 22468 7157 22477 7191
rect 22477 7157 22511 7191
rect 22511 7157 22520 7191
rect 22468 7148 22520 7157
rect 23940 7191 23992 7200
rect 23940 7157 23949 7191
rect 23949 7157 23983 7191
rect 23983 7157 23992 7191
rect 23940 7148 23992 7157
rect 26148 7148 26200 7200
rect 27436 7191 27488 7200
rect 27436 7157 27445 7191
rect 27445 7157 27479 7191
rect 27479 7157 27488 7191
rect 27436 7148 27488 7157
rect 27528 7148 27580 7200
rect 28080 7148 28132 7200
rect 10246 7046 10298 7098
rect 10310 7046 10362 7098
rect 10374 7046 10426 7098
rect 10438 7046 10490 7098
rect 19510 7046 19562 7098
rect 19574 7046 19626 7098
rect 19638 7046 19690 7098
rect 19702 7046 19754 7098
rect 2136 6808 2188 6860
rect 2504 6808 2556 6860
rect 4528 6944 4580 6996
rect 8668 6944 8720 6996
rect 9496 6944 9548 6996
rect 10600 6987 10652 6996
rect 10600 6953 10609 6987
rect 10609 6953 10643 6987
rect 10643 6953 10652 6987
rect 10600 6944 10652 6953
rect 11336 6944 11388 6996
rect 15476 6944 15528 6996
rect 15660 6987 15712 6996
rect 15660 6953 15669 6987
rect 15669 6953 15703 6987
rect 15703 6953 15712 6987
rect 15660 6944 15712 6953
rect 17316 6987 17368 6996
rect 17316 6953 17325 6987
rect 17325 6953 17359 6987
rect 17359 6953 17368 6987
rect 17316 6944 17368 6953
rect 5908 6876 5960 6928
rect 8392 6876 8444 6928
rect 10140 6876 10192 6928
rect 3240 6851 3292 6860
rect 3240 6817 3249 6851
rect 3249 6817 3283 6851
rect 3283 6817 3292 6851
rect 3240 6808 3292 6817
rect 3792 6808 3844 6860
rect 3976 6851 4028 6860
rect 3976 6817 3985 6851
rect 3985 6817 4019 6851
rect 4019 6817 4028 6851
rect 3976 6808 4028 6817
rect 4068 6808 4120 6860
rect 6000 6808 6052 6860
rect 6920 6808 6972 6860
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 5540 6740 5592 6792
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 9864 6808 9916 6860
rect 12624 6876 12676 6928
rect 13636 6876 13688 6928
rect 14740 6876 14792 6928
rect 11888 6808 11940 6860
rect 12808 6808 12860 6860
rect 13268 6851 13320 6860
rect 13268 6817 13277 6851
rect 13277 6817 13311 6851
rect 13311 6817 13320 6851
rect 13268 6808 13320 6817
rect 14096 6808 14148 6860
rect 10048 6740 10100 6792
rect 10692 6740 10744 6792
rect 12900 6715 12952 6724
rect 12900 6681 12909 6715
rect 12909 6681 12943 6715
rect 12943 6681 12952 6715
rect 12900 6672 12952 6681
rect 13728 6740 13780 6792
rect 13636 6672 13688 6724
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 3884 6604 3936 6656
rect 5172 6647 5224 6656
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 13452 6604 13504 6656
rect 18512 6944 18564 6996
rect 23112 6987 23164 6996
rect 18420 6876 18472 6928
rect 17960 6851 18012 6860
rect 16580 6740 16632 6792
rect 17960 6817 17969 6851
rect 17969 6817 18003 6851
rect 18003 6817 18012 6851
rect 17960 6808 18012 6817
rect 18052 6672 18104 6724
rect 18788 6808 18840 6860
rect 19064 6851 19116 6860
rect 19064 6817 19073 6851
rect 19073 6817 19107 6851
rect 19107 6817 19116 6851
rect 19340 6876 19392 6928
rect 19800 6919 19852 6928
rect 19800 6885 19809 6919
rect 19809 6885 19843 6919
rect 19843 6885 19852 6919
rect 19800 6876 19852 6885
rect 23112 6953 23121 6987
rect 23121 6953 23155 6987
rect 23155 6953 23164 6987
rect 23112 6944 23164 6953
rect 20076 6876 20128 6928
rect 25688 6987 25740 6996
rect 25688 6953 25697 6987
rect 25697 6953 25731 6987
rect 25731 6953 25740 6987
rect 25688 6944 25740 6953
rect 25964 6944 26016 6996
rect 19064 6808 19116 6817
rect 18604 6740 18656 6792
rect 20536 6808 20588 6860
rect 23020 6851 23072 6860
rect 23020 6817 23029 6851
rect 23029 6817 23063 6851
rect 23063 6817 23072 6851
rect 23020 6808 23072 6817
rect 23940 6808 23992 6860
rect 24860 6876 24912 6928
rect 24584 6851 24636 6860
rect 24584 6817 24593 6851
rect 24593 6817 24627 6851
rect 24627 6817 24636 6851
rect 24584 6808 24636 6817
rect 24676 6808 24728 6860
rect 20996 6740 21048 6792
rect 23572 6740 23624 6792
rect 25872 6740 25924 6792
rect 26148 6783 26200 6792
rect 26148 6749 26157 6783
rect 26157 6749 26191 6783
rect 26191 6749 26200 6783
rect 26148 6740 26200 6749
rect 21088 6672 21140 6724
rect 22928 6672 22980 6724
rect 25044 6672 25096 6724
rect 28172 6715 28224 6724
rect 28172 6681 28181 6715
rect 28181 6681 28215 6715
rect 28215 6681 28224 6715
rect 28172 6672 28224 6681
rect 25136 6647 25188 6656
rect 25136 6613 25145 6647
rect 25145 6613 25179 6647
rect 25179 6613 25188 6647
rect 25136 6604 25188 6613
rect 5614 6502 5666 6554
rect 5678 6502 5730 6554
rect 5742 6502 5794 6554
rect 5806 6502 5858 6554
rect 14878 6502 14930 6554
rect 14942 6502 14994 6554
rect 15006 6502 15058 6554
rect 15070 6502 15122 6554
rect 24142 6502 24194 6554
rect 24206 6502 24258 6554
rect 24270 6502 24322 6554
rect 24334 6502 24386 6554
rect 4160 6400 4212 6452
rect 11244 6443 11296 6452
rect 11244 6409 11253 6443
rect 11253 6409 11287 6443
rect 11287 6409 11296 6443
rect 11244 6400 11296 6409
rect 11336 6443 11388 6452
rect 11336 6409 11345 6443
rect 11345 6409 11379 6443
rect 11379 6409 11388 6443
rect 12164 6443 12216 6452
rect 11336 6400 11388 6409
rect 12164 6409 12173 6443
rect 12173 6409 12207 6443
rect 12207 6409 12216 6443
rect 12164 6400 12216 6409
rect 15384 6400 15436 6452
rect 15752 6400 15804 6452
rect 16212 6400 16264 6452
rect 16488 6400 16540 6452
rect 18604 6400 18656 6452
rect 18788 6443 18840 6452
rect 18788 6409 18797 6443
rect 18797 6409 18831 6443
rect 18831 6409 18840 6443
rect 18788 6400 18840 6409
rect 9864 6332 9916 6384
rect 1400 6264 1452 6316
rect 3424 6264 3476 6316
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 2044 6196 2096 6248
rect 2136 6196 2188 6248
rect 3884 6196 3936 6248
rect 4160 6196 4212 6248
rect 6000 6264 6052 6316
rect 10968 6264 11020 6316
rect 5172 6196 5224 6248
rect 7840 6196 7892 6248
rect 11152 6196 11204 6248
rect 12348 6264 12400 6316
rect 13452 6307 13504 6316
rect 12256 6196 12308 6248
rect 12716 6239 12768 6248
rect 12716 6205 12725 6239
rect 12725 6205 12759 6239
rect 12759 6205 12768 6239
rect 12716 6196 12768 6205
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 14556 6196 14608 6248
rect 15844 6332 15896 6384
rect 17684 6332 17736 6384
rect 15016 6239 15068 6248
rect 15016 6205 15025 6239
rect 15025 6205 15059 6239
rect 15059 6205 15068 6239
rect 15016 6196 15068 6205
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 1768 6060 1820 6112
rect 11060 6171 11112 6180
rect 11060 6137 11069 6171
rect 11069 6137 11103 6171
rect 11103 6137 11112 6171
rect 11060 6128 11112 6137
rect 19800 6264 19852 6316
rect 21088 6400 21140 6452
rect 23940 6400 23992 6452
rect 24584 6400 24636 6452
rect 27528 6400 27580 6452
rect 25504 6332 25556 6384
rect 25964 6332 26016 6384
rect 15936 6239 15988 6248
rect 15936 6205 15945 6239
rect 15945 6205 15979 6239
rect 15979 6205 15988 6239
rect 15936 6196 15988 6205
rect 18696 6239 18748 6248
rect 18696 6205 18705 6239
rect 18705 6205 18739 6239
rect 18739 6205 18748 6239
rect 18696 6196 18748 6205
rect 20076 6196 20128 6248
rect 5448 6060 5500 6112
rect 6736 6060 6788 6112
rect 7196 6060 7248 6112
rect 18328 6128 18380 6180
rect 12992 6060 13044 6112
rect 13452 6060 13504 6112
rect 13820 6103 13872 6112
rect 13820 6069 13829 6103
rect 13829 6069 13863 6103
rect 13863 6069 13872 6103
rect 13820 6060 13872 6069
rect 18052 6060 18104 6112
rect 18420 6060 18472 6112
rect 21364 6103 21416 6112
rect 21364 6069 21373 6103
rect 21373 6069 21407 6103
rect 21407 6069 21416 6103
rect 21364 6060 21416 6069
rect 22560 6196 22612 6248
rect 24676 6264 24728 6316
rect 26240 6264 26292 6316
rect 26516 6264 26568 6316
rect 24768 6196 24820 6248
rect 25136 6196 25188 6248
rect 27436 6196 27488 6248
rect 25872 6128 25924 6180
rect 22744 6060 22796 6112
rect 23020 6060 23072 6112
rect 26148 6060 26200 6112
rect 28172 6103 28224 6112
rect 28172 6069 28181 6103
rect 28181 6069 28215 6103
rect 28215 6069 28224 6103
rect 28172 6060 28224 6069
rect 10246 5958 10298 6010
rect 10310 5958 10362 6010
rect 10374 5958 10426 6010
rect 10438 5958 10490 6010
rect 19510 5958 19562 6010
rect 19574 5958 19626 6010
rect 19638 5958 19690 6010
rect 19702 5958 19754 6010
rect 3700 5856 3752 5908
rect 6368 5856 6420 5908
rect 10968 5899 11020 5908
rect 2228 5831 2280 5840
rect 2228 5797 2237 5831
rect 2237 5797 2271 5831
rect 2271 5797 2280 5831
rect 2228 5788 2280 5797
rect 3792 5788 3844 5840
rect 3608 5720 3660 5772
rect 3332 5695 3384 5704
rect 2504 5627 2556 5636
rect 2504 5593 2513 5627
rect 2513 5593 2547 5627
rect 2547 5593 2556 5627
rect 2504 5584 2556 5593
rect 3332 5661 3341 5695
rect 3341 5661 3375 5695
rect 3375 5661 3384 5695
rect 3332 5652 3384 5661
rect 7196 5788 7248 5840
rect 10968 5865 10977 5899
rect 10977 5865 11011 5899
rect 11011 5865 11020 5899
rect 10968 5856 11020 5865
rect 17960 5856 18012 5908
rect 21364 5856 21416 5908
rect 24492 5856 24544 5908
rect 25320 5899 25372 5908
rect 25320 5865 25329 5899
rect 25329 5865 25363 5899
rect 25363 5865 25372 5899
rect 25320 5856 25372 5865
rect 26056 5899 26108 5908
rect 26056 5865 26065 5899
rect 26065 5865 26099 5899
rect 26099 5865 26108 5899
rect 26056 5856 26108 5865
rect 4252 5763 4304 5772
rect 4252 5729 4261 5763
rect 4261 5729 4295 5763
rect 4295 5729 4304 5763
rect 4252 5720 4304 5729
rect 4344 5720 4396 5772
rect 6552 5720 6604 5772
rect 6828 5763 6880 5772
rect 6828 5729 6837 5763
rect 6837 5729 6871 5763
rect 6871 5729 6880 5763
rect 6828 5720 6880 5729
rect 7656 5720 7708 5772
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 9864 5763 9916 5772
rect 9864 5729 9873 5763
rect 9873 5729 9907 5763
rect 9907 5729 9916 5763
rect 9864 5720 9916 5729
rect 2688 5559 2740 5568
rect 2688 5525 2697 5559
rect 2697 5525 2731 5559
rect 2731 5525 2740 5559
rect 2688 5516 2740 5525
rect 3792 5559 3844 5568
rect 3792 5525 3801 5559
rect 3801 5525 3835 5559
rect 3835 5525 3844 5559
rect 3792 5516 3844 5525
rect 9956 5652 10008 5704
rect 10600 5652 10652 5704
rect 10784 5720 10836 5772
rect 10968 5763 11020 5772
rect 10968 5729 10977 5763
rect 10977 5729 11011 5763
rect 11011 5729 11020 5763
rect 10968 5720 11020 5729
rect 11244 5788 11296 5840
rect 13820 5788 13872 5840
rect 15016 5788 15068 5840
rect 17132 5720 17184 5772
rect 17408 5720 17460 5772
rect 17868 5720 17920 5772
rect 18328 5720 18380 5772
rect 10876 5652 10928 5704
rect 12072 5695 12124 5704
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 13912 5652 13964 5704
rect 18236 5652 18288 5704
rect 18604 5652 18656 5704
rect 24768 5720 24820 5772
rect 28172 5788 28224 5840
rect 25780 5720 25832 5772
rect 25872 5720 25924 5772
rect 26424 5720 26476 5772
rect 26148 5652 26200 5704
rect 6552 5584 6604 5636
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 10692 5516 10744 5568
rect 10784 5559 10836 5568
rect 10784 5525 10793 5559
rect 10793 5525 10827 5559
rect 10827 5525 10836 5559
rect 13636 5584 13688 5636
rect 26700 5584 26752 5636
rect 26884 5627 26936 5636
rect 26884 5593 26893 5627
rect 26893 5593 26927 5627
rect 26927 5593 26936 5627
rect 26884 5584 26936 5593
rect 10784 5516 10836 5525
rect 13268 5516 13320 5568
rect 17960 5516 18012 5568
rect 18696 5516 18748 5568
rect 23940 5516 23992 5568
rect 24492 5559 24544 5568
rect 24492 5525 24501 5559
rect 24501 5525 24535 5559
rect 24535 5525 24544 5559
rect 24492 5516 24544 5525
rect 24584 5516 24636 5568
rect 27436 5516 27488 5568
rect 5614 5414 5666 5466
rect 5678 5414 5730 5466
rect 5742 5414 5794 5466
rect 5806 5414 5858 5466
rect 14878 5414 14930 5466
rect 14942 5414 14994 5466
rect 15006 5414 15058 5466
rect 15070 5414 15122 5466
rect 24142 5414 24194 5466
rect 24206 5414 24258 5466
rect 24270 5414 24322 5466
rect 24334 5414 24386 5466
rect 1768 5355 1820 5364
rect 1768 5321 1777 5355
rect 1777 5321 1811 5355
rect 1811 5321 1820 5355
rect 1768 5312 1820 5321
rect 2688 5355 2740 5364
rect 2688 5321 2697 5355
rect 2697 5321 2731 5355
rect 2731 5321 2740 5355
rect 2688 5312 2740 5321
rect 3332 5312 3384 5364
rect 1584 5244 1636 5296
rect 11060 5312 11112 5364
rect 14740 5312 14792 5364
rect 16580 5312 16632 5364
rect 22836 5312 22888 5364
rect 26516 5312 26568 5364
rect 27344 5312 27396 5364
rect 6000 5244 6052 5296
rect 10784 5244 10836 5296
rect 14188 5244 14240 5296
rect 19892 5244 19944 5296
rect 1952 5151 2004 5160
rect 1952 5117 1961 5151
rect 1961 5117 1995 5151
rect 1995 5117 2004 5151
rect 1952 5108 2004 5117
rect 2780 5108 2832 5160
rect 2964 5151 3016 5160
rect 2964 5117 2973 5151
rect 2973 5117 3007 5151
rect 3007 5117 3016 5151
rect 2964 5108 3016 5117
rect 3240 5108 3292 5160
rect 4988 5108 5040 5160
rect 6920 5176 6972 5228
rect 9680 5176 9732 5228
rect 10692 5219 10744 5228
rect 6368 5151 6420 5160
rect 6368 5117 6377 5151
rect 6377 5117 6411 5151
rect 6411 5117 6420 5151
rect 6368 5108 6420 5117
rect 6460 5108 6512 5160
rect 8208 5151 8260 5160
rect 8208 5117 8217 5151
rect 8217 5117 8251 5151
rect 8251 5117 8260 5151
rect 8208 5108 8260 5117
rect 8392 5151 8444 5160
rect 8392 5117 8401 5151
rect 8401 5117 8435 5151
rect 8435 5117 8444 5151
rect 8392 5108 8444 5117
rect 9864 5108 9916 5160
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 10876 5108 10928 5160
rect 4620 5040 4672 5092
rect 10600 5040 10652 5092
rect 13820 5108 13872 5160
rect 13912 5108 13964 5160
rect 16948 5108 17000 5160
rect 21732 5176 21784 5228
rect 17868 5108 17920 5160
rect 19800 5108 19852 5160
rect 21180 5108 21232 5160
rect 27344 5176 27396 5228
rect 23756 5108 23808 5160
rect 18788 5040 18840 5092
rect 22468 5040 22520 5092
rect 25228 5108 25280 5160
rect 26608 5083 26660 5092
rect 6276 4972 6328 5024
rect 8116 4972 8168 5024
rect 9588 4972 9640 5024
rect 15384 4972 15436 5024
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 18144 4972 18196 5024
rect 19248 4972 19300 5024
rect 19340 4972 19392 5024
rect 20168 4972 20220 5024
rect 23480 5015 23532 5024
rect 23480 4981 23489 5015
rect 23489 4981 23523 5015
rect 23523 4981 23532 5015
rect 23480 4972 23532 4981
rect 25044 4972 25096 5024
rect 26608 5049 26617 5083
rect 26617 5049 26651 5083
rect 26651 5049 26660 5083
rect 26608 5040 26660 5049
rect 27712 5083 27764 5092
rect 27712 5049 27721 5083
rect 27721 5049 27755 5083
rect 27755 5049 27764 5083
rect 27712 5040 27764 5049
rect 27528 4972 27580 5024
rect 10246 4870 10298 4922
rect 10310 4870 10362 4922
rect 10374 4870 10426 4922
rect 10438 4870 10490 4922
rect 19510 4870 19562 4922
rect 19574 4870 19626 4922
rect 19638 4870 19690 4922
rect 19702 4870 19754 4922
rect 3792 4768 3844 4820
rect 5908 4768 5960 4820
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 15200 4811 15252 4820
rect 12440 4768 12492 4777
rect 15200 4777 15209 4811
rect 15209 4777 15243 4811
rect 15243 4777 15252 4811
rect 15200 4768 15252 4777
rect 1400 4632 1452 4684
rect 2780 4632 2832 4684
rect 3240 4675 3292 4684
rect 3240 4641 3249 4675
rect 3249 4641 3283 4675
rect 3283 4641 3292 4675
rect 3240 4632 3292 4641
rect 4436 4632 4488 4684
rect 5908 4632 5960 4684
rect 7288 4632 7340 4684
rect 8116 4675 8168 4684
rect 8116 4641 8125 4675
rect 8125 4641 8159 4675
rect 8159 4641 8168 4675
rect 8116 4632 8168 4641
rect 8760 4675 8812 4684
rect 8760 4641 8769 4675
rect 8769 4641 8803 4675
rect 8803 4641 8812 4675
rect 8760 4632 8812 4641
rect 9036 4675 9088 4684
rect 9036 4641 9045 4675
rect 9045 4641 9079 4675
rect 9079 4641 9088 4675
rect 9036 4632 9088 4641
rect 10692 4700 10744 4752
rect 13820 4743 13872 4752
rect 13820 4709 13829 4743
rect 13829 4709 13863 4743
rect 13863 4709 13872 4743
rect 13820 4700 13872 4709
rect 14188 4700 14240 4752
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 12164 4632 12216 4684
rect 7104 4607 7156 4616
rect 3516 4496 3568 4548
rect 7104 4573 7113 4607
rect 7113 4573 7147 4607
rect 7147 4573 7156 4607
rect 10876 4607 10928 4616
rect 7104 4564 7156 4573
rect 6092 4496 6144 4548
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 14740 4632 14792 4684
rect 16304 4768 16356 4820
rect 16672 4768 16724 4820
rect 17868 4768 17920 4820
rect 16580 4700 16632 4752
rect 17776 4700 17828 4752
rect 16212 4675 16264 4684
rect 16212 4641 16221 4675
rect 16221 4641 16255 4675
rect 16255 4641 16264 4675
rect 16396 4675 16448 4684
rect 16212 4632 16264 4641
rect 16396 4641 16405 4675
rect 16405 4641 16439 4675
rect 16439 4641 16448 4675
rect 16396 4632 16448 4641
rect 18144 4675 18196 4684
rect 18144 4641 18153 4675
rect 18153 4641 18187 4675
rect 18187 4641 18196 4675
rect 18144 4632 18196 4641
rect 9036 4496 9088 4548
rect 13268 4496 13320 4548
rect 15660 4496 15712 4548
rect 16580 4564 16632 4616
rect 18880 4632 18932 4684
rect 20720 4768 20772 4820
rect 23940 4768 23992 4820
rect 19248 4700 19300 4752
rect 20076 4700 20128 4752
rect 18420 4564 18472 4616
rect 19708 4632 19760 4684
rect 22008 4700 22060 4752
rect 22376 4700 22428 4752
rect 23112 4700 23164 4752
rect 23572 4743 23624 4752
rect 23572 4709 23581 4743
rect 23581 4709 23615 4743
rect 23615 4709 23624 4743
rect 23572 4700 23624 4709
rect 23664 4743 23716 4752
rect 23664 4709 23673 4743
rect 23673 4709 23707 4743
rect 23707 4709 23716 4743
rect 23664 4700 23716 4709
rect 24584 4700 24636 4752
rect 25412 4700 25464 4752
rect 21640 4675 21692 4684
rect 19892 4564 19944 4616
rect 20076 4607 20128 4616
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 17684 4496 17736 4548
rect 18880 4496 18932 4548
rect 19984 4496 20036 4548
rect 20996 4564 21048 4616
rect 21640 4641 21649 4675
rect 21649 4641 21683 4675
rect 21683 4641 21692 4675
rect 21640 4632 21692 4641
rect 22744 4632 22796 4684
rect 24492 4675 24544 4684
rect 20628 4496 20680 4548
rect 21548 4564 21600 4616
rect 23388 4564 23440 4616
rect 23940 4564 23992 4616
rect 24492 4641 24501 4675
rect 24501 4641 24535 4675
rect 24535 4641 24544 4675
rect 24492 4632 24544 4641
rect 25320 4632 25372 4684
rect 23020 4496 23072 4548
rect 23848 4496 23900 4548
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 4344 4428 4396 4480
rect 4436 4428 4488 4480
rect 7380 4471 7432 4480
rect 7380 4437 7389 4471
rect 7389 4437 7423 4471
rect 7423 4437 7432 4471
rect 7380 4428 7432 4437
rect 15568 4428 15620 4480
rect 16028 4428 16080 4480
rect 17868 4471 17920 4480
rect 17868 4437 17877 4471
rect 17877 4437 17911 4471
rect 17911 4437 17920 4471
rect 17868 4428 17920 4437
rect 19064 4471 19116 4480
rect 19064 4437 19073 4471
rect 19073 4437 19107 4471
rect 19107 4437 19116 4471
rect 19064 4428 19116 4437
rect 21088 4428 21140 4480
rect 21916 4428 21968 4480
rect 27712 4496 27764 4548
rect 26056 4428 26108 4480
rect 28080 4471 28132 4480
rect 28080 4437 28089 4471
rect 28089 4437 28123 4471
rect 28123 4437 28132 4471
rect 28080 4428 28132 4437
rect 5614 4326 5666 4378
rect 5678 4326 5730 4378
rect 5742 4326 5794 4378
rect 5806 4326 5858 4378
rect 14878 4326 14930 4378
rect 14942 4326 14994 4378
rect 15006 4326 15058 4378
rect 15070 4326 15122 4378
rect 24142 4326 24194 4378
rect 24206 4326 24258 4378
rect 24270 4326 24322 4378
rect 24334 4326 24386 4378
rect 4160 4224 4212 4276
rect 4988 4224 5040 4276
rect 6092 4224 6144 4276
rect 10876 4267 10928 4276
rect 10876 4233 10885 4267
rect 10885 4233 10919 4267
rect 10919 4233 10928 4267
rect 10876 4224 10928 4233
rect 12900 4224 12952 4276
rect 13912 4224 13964 4276
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 4252 4156 4304 4208
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 7564 4088 7616 4140
rect 3056 4020 3108 4072
rect 4160 4020 4212 4072
rect 4344 4020 4396 4072
rect 1676 3952 1728 4004
rect 7472 4020 7524 4072
rect 8392 4088 8444 4140
rect 8484 4088 8536 4140
rect 8760 4088 8812 4140
rect 9864 4088 9916 4140
rect 10968 4156 11020 4208
rect 8208 4063 8260 4072
rect 8208 4029 8217 4063
rect 8217 4029 8251 4063
rect 8251 4029 8260 4063
rect 8208 4020 8260 4029
rect 11612 4088 11664 4140
rect 12164 4088 12216 4140
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 11520 4020 11572 4072
rect 4712 3952 4764 4004
rect 6460 3952 6512 4004
rect 7012 3952 7064 4004
rect 11336 3952 11388 4004
rect 11428 3952 11480 4004
rect 12900 4020 12952 4072
rect 13084 4020 13136 4072
rect 13268 4063 13320 4072
rect 13268 4029 13277 4063
rect 13277 4029 13311 4063
rect 13311 4029 13320 4063
rect 13268 4020 13320 4029
rect 13452 4020 13504 4072
rect 14740 4020 14792 4072
rect 15016 4063 15068 4072
rect 15016 4029 15025 4063
rect 15025 4029 15059 4063
rect 15059 4029 15068 4063
rect 15016 4020 15068 4029
rect 16580 4224 16632 4276
rect 17684 4224 17736 4276
rect 18880 4224 18932 4276
rect 21548 4224 21600 4276
rect 15936 4156 15988 4208
rect 18604 4156 18656 4208
rect 19984 4156 20036 4208
rect 15568 4088 15620 4140
rect 18236 4088 18288 4140
rect 18420 4088 18472 4140
rect 15476 4020 15528 4072
rect 16028 4020 16080 4072
rect 16488 4020 16540 4072
rect 18512 4020 18564 4072
rect 18604 4020 18656 4072
rect 18788 4063 18840 4072
rect 18788 4029 18797 4063
rect 18797 4029 18831 4063
rect 18831 4029 18840 4063
rect 18788 4020 18840 4029
rect 18880 4063 18932 4072
rect 18880 4029 18889 4063
rect 18889 4029 18923 4063
rect 18923 4029 18932 4063
rect 19064 4063 19116 4072
rect 18880 4020 18932 4029
rect 19064 4029 19073 4063
rect 19073 4029 19107 4063
rect 19107 4029 19116 4063
rect 19064 4020 19116 4029
rect 19708 4020 19760 4072
rect 19984 4063 20036 4072
rect 19984 4029 19993 4063
rect 19993 4029 20027 4063
rect 20027 4029 20036 4063
rect 19984 4020 20036 4029
rect 20996 4020 21048 4072
rect 22836 4224 22888 4276
rect 23756 4224 23808 4276
rect 23664 4156 23716 4208
rect 25044 4156 25096 4208
rect 25964 4156 26016 4208
rect 22192 4088 22244 4140
rect 23112 4131 23164 4140
rect 23112 4097 23121 4131
rect 23121 4097 23155 4131
rect 23155 4097 23164 4131
rect 23112 4088 23164 4097
rect 23296 4088 23348 4140
rect 27252 4224 27304 4276
rect 23388 4020 23440 4072
rect 23480 4020 23532 4072
rect 26056 4063 26108 4072
rect 26056 4029 26065 4063
rect 26065 4029 26099 4063
rect 26099 4029 26108 4063
rect 26056 4020 26108 4029
rect 26700 4020 26752 4072
rect 2596 3927 2648 3936
rect 2596 3893 2605 3927
rect 2605 3893 2639 3927
rect 2639 3893 2648 3927
rect 2596 3884 2648 3893
rect 2872 3884 2924 3936
rect 4160 3884 4212 3936
rect 6184 3927 6236 3936
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6184 3884 6236 3893
rect 8668 3884 8720 3936
rect 9588 3927 9640 3936
rect 9588 3893 9597 3927
rect 9597 3893 9631 3927
rect 9631 3893 9640 3927
rect 9588 3884 9640 3893
rect 12256 3884 12308 3936
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 12900 3884 12952 3893
rect 14740 3927 14792 3936
rect 14740 3893 14749 3927
rect 14749 3893 14783 3927
rect 14783 3893 14792 3927
rect 14740 3884 14792 3893
rect 14832 3884 14884 3936
rect 20628 3884 20680 3936
rect 22468 3884 22520 3936
rect 23572 3952 23624 4004
rect 22652 3884 22704 3936
rect 23204 3884 23256 3936
rect 25504 3927 25556 3936
rect 25504 3893 25513 3927
rect 25513 3893 25547 3927
rect 25547 3893 25556 3927
rect 25504 3884 25556 3893
rect 25872 3952 25924 4004
rect 27896 3952 27948 4004
rect 10246 3782 10298 3834
rect 10310 3782 10362 3834
rect 10374 3782 10426 3834
rect 10438 3782 10490 3834
rect 19510 3782 19562 3834
rect 19574 3782 19626 3834
rect 19638 3782 19690 3834
rect 19702 3782 19754 3834
rect 1676 3723 1728 3732
rect 1676 3689 1685 3723
rect 1685 3689 1719 3723
rect 1719 3689 1728 3723
rect 1676 3680 1728 3689
rect 4160 3723 4212 3732
rect 4160 3689 4169 3723
rect 4169 3689 4203 3723
rect 4203 3689 4212 3723
rect 4160 3680 4212 3689
rect 5080 3680 5132 3732
rect 7380 3680 7432 3732
rect 7472 3680 7524 3732
rect 10048 3680 10100 3732
rect 11980 3680 12032 3732
rect 13084 3680 13136 3732
rect 15016 3680 15068 3732
rect 16396 3723 16448 3732
rect 16396 3689 16405 3723
rect 16405 3689 16439 3723
rect 16439 3689 16448 3723
rect 16396 3680 16448 3689
rect 2596 3612 2648 3664
rect 4436 3544 4488 3596
rect 4988 3587 5040 3596
rect 4988 3553 4997 3587
rect 4997 3553 5031 3587
rect 5031 3553 5040 3587
rect 4988 3544 5040 3553
rect 6276 3544 6328 3596
rect 7748 3544 7800 3596
rect 9036 3544 9088 3596
rect 9404 3587 9456 3596
rect 9404 3553 9413 3587
rect 9413 3553 9447 3587
rect 9447 3553 9456 3587
rect 9404 3544 9456 3553
rect 10600 3587 10652 3596
rect 10600 3553 10609 3587
rect 10609 3553 10643 3587
rect 10643 3553 10652 3587
rect 10600 3544 10652 3553
rect 11336 3612 11388 3664
rect 12348 3544 12400 3596
rect 12900 3612 12952 3664
rect 14740 3612 14792 3664
rect 17868 3612 17920 3664
rect 18512 3612 18564 3664
rect 20076 3680 20128 3732
rect 20352 3723 20404 3732
rect 20352 3689 20361 3723
rect 20361 3689 20395 3723
rect 20395 3689 20404 3723
rect 20352 3680 20404 3689
rect 21640 3680 21692 3732
rect 23204 3680 23256 3732
rect 24584 3723 24636 3732
rect 24584 3689 24593 3723
rect 24593 3689 24627 3723
rect 24627 3689 24636 3723
rect 24584 3680 24636 3689
rect 25320 3723 25372 3732
rect 25320 3689 25329 3723
rect 25329 3689 25363 3723
rect 25363 3689 25372 3723
rect 25320 3680 25372 3689
rect 26792 3723 26844 3732
rect 16212 3587 16264 3596
rect 16212 3553 16221 3587
rect 16221 3553 16255 3587
rect 16255 3553 16264 3587
rect 16212 3544 16264 3553
rect 16672 3544 16724 3596
rect 7564 3476 7616 3528
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 5448 3408 5500 3460
rect 11336 3476 11388 3528
rect 11704 3476 11756 3528
rect 11980 3476 12032 3528
rect 12072 3476 12124 3528
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 12440 3476 12492 3485
rect 14096 3476 14148 3528
rect 15660 3476 15712 3528
rect 8668 3408 8720 3460
rect 11428 3408 11480 3460
rect 15844 3408 15896 3460
rect 4896 3340 4948 3392
rect 7104 3340 7156 3392
rect 11152 3340 11204 3392
rect 17224 3340 17276 3392
rect 17868 3476 17920 3528
rect 19984 3544 20036 3596
rect 21916 3612 21968 3664
rect 19248 3476 19300 3528
rect 22560 3587 22612 3596
rect 22560 3553 22569 3587
rect 22569 3553 22603 3587
rect 22603 3553 22612 3587
rect 22560 3544 22612 3553
rect 22468 3476 22520 3528
rect 22928 3544 22980 3596
rect 25412 3544 25464 3596
rect 22836 3476 22888 3528
rect 25136 3476 25188 3528
rect 25780 3587 25832 3596
rect 26792 3689 26801 3723
rect 26801 3689 26835 3723
rect 26835 3689 26844 3723
rect 26792 3680 26844 3689
rect 25780 3553 25794 3587
rect 25794 3553 25828 3587
rect 25828 3553 25832 3587
rect 25780 3544 25832 3553
rect 26148 3476 26200 3528
rect 19248 3340 19300 3392
rect 26424 3408 26476 3460
rect 28172 3451 28224 3460
rect 24492 3340 24544 3392
rect 27896 3340 27948 3392
rect 28172 3417 28181 3451
rect 28181 3417 28215 3451
rect 28215 3417 28224 3451
rect 28172 3408 28224 3417
rect 29276 3340 29328 3392
rect 5614 3238 5666 3290
rect 5678 3238 5730 3290
rect 5742 3238 5794 3290
rect 5806 3238 5858 3290
rect 14878 3238 14930 3290
rect 14942 3238 14994 3290
rect 15006 3238 15058 3290
rect 15070 3238 15122 3290
rect 24142 3238 24194 3290
rect 24206 3238 24258 3290
rect 24270 3238 24322 3290
rect 24334 3238 24386 3290
rect 2872 3179 2924 3188
rect 2872 3145 2881 3179
rect 2881 3145 2915 3179
rect 2915 3145 2924 3179
rect 2872 3136 2924 3145
rect 6644 3068 6696 3120
rect 11612 3136 11664 3188
rect 11796 3136 11848 3188
rect 15568 3136 15620 3188
rect 16304 3136 16356 3188
rect 17040 3179 17092 3188
rect 17040 3145 17049 3179
rect 17049 3145 17083 3179
rect 17083 3145 17092 3179
rect 17040 3136 17092 3145
rect 17224 3136 17276 3188
rect 11152 3068 11204 3120
rect 12624 3068 12676 3120
rect 12900 3068 12952 3120
rect 15752 3068 15804 3120
rect 16212 3068 16264 3120
rect 19156 3068 19208 3120
rect 19892 3068 19944 3120
rect 22376 3111 22428 3120
rect 22376 3077 22385 3111
rect 22385 3077 22419 3111
rect 22419 3077 22428 3111
rect 22376 3068 22428 3077
rect 22928 3111 22980 3120
rect 22928 3077 22937 3111
rect 22937 3077 22971 3111
rect 22971 3077 22980 3111
rect 22928 3068 22980 3077
rect 23020 3068 23072 3120
rect 2964 3000 3016 3052
rect 4896 3000 4948 3052
rect 6920 3000 6972 3052
rect 12164 3043 12216 3052
rect 12164 3009 12173 3043
rect 12173 3009 12207 3043
rect 12207 3009 12216 3043
rect 12164 3000 12216 3009
rect 13360 3000 13412 3052
rect 15200 3000 15252 3052
rect 17684 3043 17736 3052
rect 17684 3009 17693 3043
rect 17693 3009 17727 3043
rect 17727 3009 17736 3043
rect 17684 3000 17736 3009
rect 1676 2975 1728 2984
rect 1676 2941 1685 2975
rect 1685 2941 1719 2975
rect 1719 2941 1728 2975
rect 1676 2932 1728 2941
rect 3148 2932 3200 2984
rect 3516 2932 3568 2984
rect 6184 2932 6236 2984
rect 7104 2932 7156 2984
rect 7564 2932 7616 2984
rect 9588 2932 9640 2984
rect 10048 2932 10100 2984
rect 16212 2932 16264 2984
rect 17316 2932 17368 2984
rect 20168 3000 20220 3052
rect 18420 2932 18472 2984
rect 19340 2932 19392 2984
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 20076 2932 20128 2984
rect 21088 2932 21140 2984
rect 23112 2932 23164 2984
rect 25136 3068 25188 3120
rect 25872 3068 25924 3120
rect 17132 2864 17184 2916
rect 21916 2864 21968 2916
rect 22008 2864 22060 2916
rect 23020 2864 23072 2916
rect 6920 2796 6972 2848
rect 7564 2796 7616 2848
rect 7748 2796 7800 2848
rect 11980 2839 12032 2848
rect 11980 2805 11989 2839
rect 11989 2805 12023 2839
rect 12023 2805 12032 2839
rect 11980 2796 12032 2805
rect 12440 2796 12492 2848
rect 14096 2796 14148 2848
rect 15108 2796 15160 2848
rect 15384 2796 15436 2848
rect 21364 2796 21416 2848
rect 21548 2796 21600 2848
rect 23664 2932 23716 2984
rect 23940 2864 23992 2916
rect 24492 2864 24544 2916
rect 24768 2796 24820 2848
rect 25780 2975 25832 2984
rect 25780 2941 25794 2975
rect 25794 2941 25828 2975
rect 25828 2941 25832 2975
rect 25780 2932 25832 2941
rect 25964 2975 26016 2984
rect 25964 2941 25973 2975
rect 25973 2941 26007 2975
rect 26007 2941 26016 2975
rect 27528 3136 27580 3188
rect 27252 3068 27304 3120
rect 27896 3043 27948 3052
rect 27896 3009 27905 3043
rect 27905 3009 27939 3043
rect 27939 3009 27948 3043
rect 27896 3000 27948 3009
rect 25964 2932 26016 2941
rect 26792 2907 26844 2916
rect 26792 2873 26801 2907
rect 26801 2873 26835 2907
rect 26835 2873 26844 2907
rect 26792 2864 26844 2873
rect 26976 2907 27028 2916
rect 26976 2873 26985 2907
rect 26985 2873 27019 2907
rect 27019 2873 27028 2907
rect 26976 2864 27028 2873
rect 27252 2796 27304 2848
rect 27344 2796 27396 2848
rect 27896 2796 27948 2848
rect 10246 2694 10298 2746
rect 10310 2694 10362 2746
rect 10374 2694 10426 2746
rect 10438 2694 10490 2746
rect 19510 2694 19562 2746
rect 19574 2694 19626 2746
rect 19638 2694 19690 2746
rect 19702 2694 19754 2746
rect 4528 2592 4580 2644
rect 4988 2592 5040 2644
rect 9404 2592 9456 2644
rect 10600 2592 10652 2644
rect 11980 2592 12032 2644
rect 12164 2592 12216 2644
rect 13544 2592 13596 2644
rect 15568 2635 15620 2644
rect 15568 2601 15577 2635
rect 15577 2601 15611 2635
rect 15611 2601 15620 2635
rect 15568 2592 15620 2601
rect 16212 2635 16264 2644
rect 16212 2601 16221 2635
rect 16221 2601 16255 2635
rect 16255 2601 16264 2635
rect 16212 2592 16264 2601
rect 17316 2592 17368 2644
rect 19984 2592 20036 2644
rect 664 2456 716 2508
rect 2596 2499 2648 2508
rect 2596 2465 2605 2499
rect 2605 2465 2639 2499
rect 2639 2465 2648 2499
rect 2596 2456 2648 2465
rect 12716 2524 12768 2576
rect 14280 2524 14332 2576
rect 21364 2592 21416 2644
rect 1952 2388 2004 2440
rect 3332 2388 3384 2440
rect 6092 2456 6144 2508
rect 7472 2456 7524 2508
rect 8576 2499 8628 2508
rect 8576 2465 8585 2499
rect 8585 2465 8619 2499
rect 8619 2465 8628 2499
rect 8576 2456 8628 2465
rect 8760 2456 8812 2508
rect 10140 2456 10192 2508
rect 11152 2499 11204 2508
rect 11152 2465 11161 2499
rect 11161 2465 11195 2499
rect 11195 2465 11204 2499
rect 11152 2456 11204 2465
rect 12256 2499 12308 2508
rect 12256 2465 12265 2499
rect 12265 2465 12299 2499
rect 12299 2465 12308 2499
rect 12256 2456 12308 2465
rect 12532 2456 12584 2508
rect 14648 2456 14700 2508
rect 15752 2499 15804 2508
rect 11888 2388 11940 2440
rect 7932 2320 7984 2372
rect 15752 2465 15761 2499
rect 15761 2465 15795 2499
rect 15795 2465 15804 2499
rect 15752 2456 15804 2465
rect 15660 2388 15712 2440
rect 19340 2499 19392 2508
rect 16948 2388 17000 2440
rect 19340 2465 19349 2499
rect 19349 2465 19383 2499
rect 19383 2465 19392 2499
rect 19340 2456 19392 2465
rect 20444 2499 20496 2508
rect 20444 2465 20453 2499
rect 20453 2465 20487 2499
rect 20487 2465 20496 2499
rect 20444 2456 20496 2465
rect 21640 2567 21692 2576
rect 21640 2533 21649 2567
rect 21649 2533 21683 2567
rect 21683 2533 21692 2567
rect 21640 2524 21692 2533
rect 21364 2388 21416 2440
rect 23020 2499 23072 2508
rect 23020 2465 23029 2499
rect 23029 2465 23063 2499
rect 23063 2465 23072 2499
rect 23020 2456 23072 2465
rect 23388 2456 23440 2508
rect 24492 2499 24544 2508
rect 24492 2465 24501 2499
rect 24501 2465 24535 2499
rect 24535 2465 24544 2499
rect 24492 2456 24544 2465
rect 27160 2499 27212 2508
rect 27160 2465 27169 2499
rect 27169 2465 27203 2499
rect 27203 2465 27212 2499
rect 27160 2456 27212 2465
rect 22468 2388 22520 2440
rect 12992 2295 13044 2304
rect 12992 2261 13001 2295
rect 13001 2261 13035 2295
rect 13035 2261 13044 2295
rect 12992 2252 13044 2261
rect 25228 2388 25280 2440
rect 25044 2320 25096 2372
rect 25872 2363 25924 2372
rect 25872 2329 25881 2363
rect 25881 2329 25915 2363
rect 25915 2329 25924 2363
rect 25872 2320 25924 2329
rect 26056 2320 26108 2372
rect 25412 2252 25464 2304
rect 26148 2252 26200 2304
rect 5614 2150 5666 2202
rect 5678 2150 5730 2202
rect 5742 2150 5794 2202
rect 5806 2150 5858 2202
rect 14878 2150 14930 2202
rect 14942 2150 14994 2202
rect 15006 2150 15058 2202
rect 15070 2150 15122 2202
rect 24142 2150 24194 2202
rect 24206 2150 24258 2202
rect 24270 2150 24322 2202
rect 24334 2150 24386 2202
rect 2596 2048 2648 2100
rect 3516 1980 3568 2032
rect 6828 1980 6880 2032
rect 2780 1912 2832 1964
rect 5908 1912 5960 1964
rect 19340 2048 19392 2100
rect 26516 2048 26568 2100
rect 12992 1980 13044 2032
rect 27160 1980 27212 2032
rect 25596 1912 25648 1964
rect 3424 1844 3476 1896
rect 7656 1844 7708 1896
rect 20444 1232 20496 1284
rect 23756 1232 23808 1284
rect 2964 1028 3016 1080
rect 8576 1028 8628 1080
<< metal2 >>
rect 846 55200 902 56800
rect 2594 55200 2650 56800
rect 2778 55720 2834 55729
rect 2778 55655 2834 55664
rect 860 52426 888 55200
rect 2608 53174 2636 55200
rect 2596 53168 2648 53174
rect 2596 53110 2648 53116
rect 2792 53106 2820 55655
rect 3882 55312 3938 55321
rect 3882 55247 3938 55256
rect 3238 54904 3294 54913
rect 3238 54839 3294 54848
rect 3146 54496 3202 54505
rect 3146 54431 3202 54440
rect 2962 54088 3018 54097
rect 2962 54023 3018 54032
rect 2780 53100 2832 53106
rect 2780 53042 2832 53048
rect 2044 52896 2096 52902
rect 2044 52838 2096 52844
rect 2872 52896 2924 52902
rect 2872 52838 2924 52844
rect 1860 52556 1912 52562
rect 1860 52498 1912 52504
rect 848 52420 900 52426
rect 848 52362 900 52368
rect 1872 51921 1900 52498
rect 1952 52352 2004 52358
rect 1952 52294 2004 52300
rect 1858 51912 1914 51921
rect 1858 51847 1914 51856
rect 1492 51808 1544 51814
rect 1492 51750 1544 51756
rect 1400 51264 1452 51270
rect 1400 51206 1452 51212
rect 1412 50425 1440 51206
rect 1504 50833 1532 51750
rect 1964 51649 1992 52294
rect 1950 51640 2006 51649
rect 1950 51575 2006 51584
rect 1860 51468 1912 51474
rect 1860 51410 1912 51416
rect 1490 50824 1546 50833
rect 1490 50759 1546 50768
rect 1398 50416 1454 50425
rect 1398 50351 1454 50360
rect 1872 50289 1900 51410
rect 1952 50720 2004 50726
rect 1952 50662 2004 50668
rect 1858 50280 1914 50289
rect 1858 50215 1914 50224
rect 1400 50176 1452 50182
rect 1400 50118 1452 50124
rect 1412 49201 1440 50118
rect 1964 50017 1992 50662
rect 1950 50008 2006 50017
rect 1950 49943 2006 49952
rect 1860 49292 1912 49298
rect 1860 49234 1912 49240
rect 1398 49192 1454 49201
rect 1398 49127 1454 49136
rect 1216 48136 1268 48142
rect 1216 48078 1268 48084
rect 1228 46510 1256 48078
rect 1872 47734 1900 49234
rect 1952 49088 2004 49094
rect 1952 49030 2004 49036
rect 1964 47977 1992 49030
rect 1950 47968 2006 47977
rect 1950 47903 2006 47912
rect 1860 47728 1912 47734
rect 1860 47670 1912 47676
rect 1952 47456 2004 47462
rect 1952 47398 2004 47404
rect 1216 46504 1268 46510
rect 1216 46446 1268 46452
rect 1228 42158 1256 46446
rect 1584 46436 1636 46442
rect 1584 46378 1636 46384
rect 1596 45626 1624 46378
rect 1768 46028 1820 46034
rect 1768 45970 1820 45976
rect 1584 45620 1636 45626
rect 1584 45562 1636 45568
rect 1400 43648 1452 43654
rect 1400 43590 1452 43596
rect 1308 43444 1360 43450
rect 1308 43386 1360 43392
rect 1320 42673 1348 43386
rect 1306 42664 1362 42673
rect 1306 42599 1362 42608
rect 1412 42265 1440 43590
rect 1780 43382 1808 45970
rect 1964 45529 1992 47398
rect 1950 45520 2006 45529
rect 1950 45455 2006 45464
rect 1952 44736 2004 44742
rect 1952 44678 2004 44684
rect 1860 44464 1912 44470
rect 1860 44406 1912 44412
rect 1768 43376 1820 43382
rect 1768 43318 1820 43324
rect 1584 42832 1636 42838
rect 1584 42774 1636 42780
rect 1398 42256 1454 42265
rect 1398 42191 1454 42200
rect 1216 42152 1268 42158
rect 1216 42094 1268 42100
rect 1492 42084 1544 42090
rect 1492 42026 1544 42032
rect 1504 41818 1532 42026
rect 1492 41812 1544 41818
rect 1492 41754 1544 41760
rect 1492 41200 1544 41206
rect 1492 41142 1544 41148
rect 1400 39840 1452 39846
rect 1400 39782 1452 39788
rect 1412 38185 1440 39782
rect 1398 38176 1454 38185
rect 1398 38111 1454 38120
rect 1400 37868 1452 37874
rect 1400 37810 1452 37816
rect 1412 36242 1440 37810
rect 1400 36236 1452 36242
rect 1400 36178 1452 36184
rect 1504 35562 1532 41142
rect 1596 38962 1624 42774
rect 1872 39030 1900 44406
rect 1964 43489 1992 44678
rect 1950 43480 2006 43489
rect 1950 43415 2006 43424
rect 1952 42560 2004 42566
rect 1952 42502 2004 42508
rect 1964 41041 1992 42502
rect 1950 41032 2006 41041
rect 1950 40967 2006 40976
rect 1952 40384 2004 40390
rect 1952 40326 2004 40332
rect 1860 39024 1912 39030
rect 1964 39001 1992 40326
rect 2056 39098 2084 52838
rect 2596 52556 2648 52562
rect 2596 52498 2648 52504
rect 2608 52154 2636 52498
rect 2780 52488 2832 52494
rect 2778 52456 2780 52465
rect 2832 52456 2834 52465
rect 2884 52426 2912 52838
rect 2778 52391 2834 52400
rect 2872 52420 2924 52426
rect 2872 52362 2924 52368
rect 2596 52148 2648 52154
rect 2596 52090 2648 52096
rect 2778 52048 2834 52057
rect 2778 51983 2780 51992
rect 2832 51983 2834 51992
rect 2780 51954 2832 51960
rect 2688 51876 2740 51882
rect 2688 51818 2740 51824
rect 2700 50969 2728 51818
rect 2780 51332 2832 51338
rect 2780 51274 2832 51280
rect 2792 51241 2820 51274
rect 2778 51232 2834 51241
rect 2778 51167 2834 51176
rect 2976 50998 3004 54023
rect 2964 50992 3016 50998
rect 2686 50960 2742 50969
rect 2964 50934 3016 50940
rect 2686 50895 2742 50904
rect 2594 50824 2650 50833
rect 2594 50759 2596 50768
rect 2648 50759 2650 50768
rect 2596 50730 2648 50736
rect 3160 50522 3188 54431
rect 3252 51066 3280 54839
rect 3896 54058 3924 55247
rect 4342 55200 4398 56800
rect 6090 55200 6146 56800
rect 7838 55200 7894 56800
rect 9586 55200 9642 56800
rect 11426 55200 11482 56800
rect 13174 55200 13230 56800
rect 14922 55200 14978 56800
rect 16670 55200 16726 56800
rect 18418 55200 18474 56800
rect 20166 55200 20222 56800
rect 22006 55200 22062 56800
rect 23570 55312 23626 55321
rect 23570 55247 23626 55256
rect 3884 54052 3936 54058
rect 3884 53994 3936 54000
rect 4066 53680 4122 53689
rect 4066 53615 4122 53624
rect 3606 53272 3662 53281
rect 3606 53207 3662 53216
rect 3422 52864 3478 52873
rect 3422 52799 3478 52808
rect 3436 51610 3464 52799
rect 3620 52086 3648 53207
rect 4080 53106 4108 53615
rect 4356 53242 4384 55200
rect 5908 54052 5960 54058
rect 5908 53994 5960 54000
rect 5588 53340 5884 53360
rect 5644 53338 5668 53340
rect 5724 53338 5748 53340
rect 5804 53338 5828 53340
rect 5666 53286 5668 53338
rect 5730 53286 5742 53338
rect 5804 53286 5806 53338
rect 5644 53284 5668 53286
rect 5724 53284 5748 53286
rect 5804 53284 5828 53286
rect 5588 53264 5884 53284
rect 4344 53236 4396 53242
rect 4344 53178 4396 53184
rect 4068 53100 4120 53106
rect 4068 53042 4120 53048
rect 5356 53032 5408 53038
rect 5356 52974 5408 52980
rect 5814 53000 5870 53009
rect 3976 52964 4028 52970
rect 3976 52906 4028 52912
rect 3792 52488 3844 52494
rect 3792 52430 3844 52436
rect 3608 52080 3660 52086
rect 3608 52022 3660 52028
rect 3424 51604 3476 51610
rect 3424 51546 3476 51552
rect 3330 51504 3386 51513
rect 3330 51439 3332 51448
rect 3384 51439 3386 51448
rect 3332 51410 3384 51416
rect 3240 51060 3292 51066
rect 3240 51002 3292 51008
rect 3148 50516 3200 50522
rect 3148 50458 3200 50464
rect 2504 50380 2556 50386
rect 2504 50322 2556 50328
rect 2516 49638 2544 50322
rect 2780 50244 2832 50250
rect 2780 50186 2832 50192
rect 2688 49768 2740 49774
rect 2688 49710 2740 49716
rect 2504 49632 2556 49638
rect 2504 49574 2556 49580
rect 2700 49366 2728 49710
rect 2792 49609 2820 50186
rect 2964 49836 3016 49842
rect 2964 49778 3016 49784
rect 2872 49768 2924 49774
rect 2872 49710 2924 49716
rect 2778 49600 2834 49609
rect 2778 49535 2834 49544
rect 2688 49360 2740 49366
rect 2688 49302 2740 49308
rect 2688 49224 2740 49230
rect 2688 49166 2740 49172
rect 2596 48612 2648 48618
rect 2596 48554 2648 48560
rect 2608 47802 2636 48554
rect 2700 48006 2728 49166
rect 2780 49156 2832 49162
rect 2780 49098 2832 49104
rect 2688 48000 2740 48006
rect 2688 47942 2740 47948
rect 2596 47796 2648 47802
rect 2596 47738 2648 47744
rect 2792 47569 2820 49098
rect 2884 48793 2912 49710
rect 2870 48784 2926 48793
rect 2870 48719 2926 48728
rect 2872 48680 2924 48686
rect 2872 48622 2924 48628
rect 2884 48226 2912 48622
rect 2976 48385 3004 49778
rect 3804 49230 3832 52430
rect 3988 51074 4016 52906
rect 4068 52556 4120 52562
rect 4068 52498 4120 52504
rect 5172 52556 5224 52562
rect 5172 52498 5224 52504
rect 4080 51610 4108 52498
rect 5184 52358 5212 52498
rect 5172 52352 5224 52358
rect 5172 52294 5224 52300
rect 5184 51610 5212 52294
rect 4068 51604 4120 51610
rect 4068 51546 4120 51552
rect 5172 51604 5224 51610
rect 5172 51546 5224 51552
rect 5172 51400 5224 51406
rect 5172 51342 5224 51348
rect 3988 51046 4108 51074
rect 3792 49224 3844 49230
rect 3792 49166 3844 49172
rect 3804 48686 3832 49166
rect 3792 48680 3844 48686
rect 3792 48622 3844 48628
rect 2962 48376 3018 48385
rect 2962 48311 3018 48320
rect 2884 48198 3004 48226
rect 2976 48142 3004 48198
rect 2964 48136 3016 48142
rect 2964 48078 3016 48084
rect 2872 48068 2924 48074
rect 2872 48010 2924 48016
rect 2778 47560 2834 47569
rect 2596 47524 2648 47530
rect 2778 47495 2834 47504
rect 2596 47466 2648 47472
rect 2504 47116 2556 47122
rect 2504 47058 2556 47064
rect 2516 45558 2544 47058
rect 2608 46578 2636 47466
rect 2688 47116 2740 47122
rect 2688 47058 2740 47064
rect 2596 46572 2648 46578
rect 2596 46514 2648 46520
rect 2504 45552 2556 45558
rect 2504 45494 2556 45500
rect 2136 45484 2188 45490
rect 2136 45426 2188 45432
rect 2320 45484 2372 45490
rect 2320 45426 2372 45432
rect 2148 45014 2176 45426
rect 2228 45280 2280 45286
rect 2228 45222 2280 45228
rect 2136 45008 2188 45014
rect 2136 44950 2188 44956
rect 2240 44334 2268 45222
rect 2228 44328 2280 44334
rect 2228 44270 2280 44276
rect 2240 41002 2268 44270
rect 2332 41614 2360 45426
rect 2596 44940 2648 44946
rect 2596 44882 2648 44888
rect 2412 44736 2464 44742
rect 2412 44678 2464 44684
rect 2424 44266 2452 44678
rect 2412 44260 2464 44266
rect 2412 44202 2464 44208
rect 2504 43172 2556 43178
rect 2504 43114 2556 43120
rect 2412 42764 2464 42770
rect 2412 42706 2464 42712
rect 2320 41608 2372 41614
rect 2320 41550 2372 41556
rect 2136 40996 2188 41002
rect 2136 40938 2188 40944
rect 2228 40996 2280 41002
rect 2228 40938 2280 40944
rect 2148 40662 2176 40938
rect 2136 40656 2188 40662
rect 2136 40598 2188 40604
rect 2240 40474 2268 40938
rect 2148 40446 2268 40474
rect 2044 39092 2096 39098
rect 2044 39034 2096 39040
rect 1860 38966 1912 38972
rect 1950 38992 2006 39001
rect 1584 38956 1636 38962
rect 1584 38898 1636 38904
rect 1596 38282 1624 38898
rect 1872 38486 1900 38966
rect 1950 38927 2006 38936
rect 2044 38956 2096 38962
rect 2044 38898 2096 38904
rect 1860 38480 1912 38486
rect 1780 38428 1860 38434
rect 1780 38422 1912 38428
rect 1780 38406 1900 38422
rect 1584 38276 1636 38282
rect 1584 38218 1636 38224
rect 1596 37874 1624 38218
rect 1584 37868 1636 37874
rect 1584 37810 1636 37816
rect 1584 37732 1636 37738
rect 1584 37674 1636 37680
rect 1596 36106 1624 37674
rect 1676 37664 1728 37670
rect 1676 37606 1728 37612
rect 1688 36553 1716 37606
rect 1674 36544 1730 36553
rect 1674 36479 1730 36488
rect 1676 36236 1728 36242
rect 1676 36178 1728 36184
rect 1584 36100 1636 36106
rect 1584 36042 1636 36048
rect 1688 35894 1716 36178
rect 1780 36174 1808 38406
rect 1860 36644 1912 36650
rect 1860 36586 1912 36592
rect 1768 36168 1820 36174
rect 1768 36110 1820 36116
rect 1596 35866 1716 35894
rect 1492 35556 1544 35562
rect 1492 35498 1544 35504
rect 1398 33688 1454 33697
rect 1398 33623 1400 33632
rect 1452 33623 1454 33632
rect 1400 33594 1452 33600
rect 1504 32978 1532 35498
rect 1492 32972 1544 32978
rect 1492 32914 1544 32920
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 1412 31482 1440 31826
rect 1400 31476 1452 31482
rect 1400 31418 1452 31424
rect 1400 31136 1452 31142
rect 1400 31078 1452 31084
rect 1412 30433 1440 31078
rect 1398 30424 1454 30433
rect 1398 30359 1454 30368
rect 1400 29572 1452 29578
rect 1400 29514 1452 29520
rect 1412 29170 1440 29514
rect 1400 29164 1452 29170
rect 1400 29106 1452 29112
rect 1596 26234 1624 35866
rect 1768 35760 1820 35766
rect 1768 35702 1820 35708
rect 1676 34944 1728 34950
rect 1674 34912 1676 34921
rect 1728 34912 1730 34921
rect 1674 34847 1730 34856
rect 1780 32978 1808 35702
rect 1872 35562 1900 36586
rect 1952 36576 2004 36582
rect 1952 36518 2004 36524
rect 1860 35556 1912 35562
rect 1860 35498 1912 35504
rect 1964 35329 1992 36518
rect 2056 35630 2084 38898
rect 2044 35624 2096 35630
rect 2044 35566 2096 35572
rect 1950 35320 2006 35329
rect 1950 35255 2006 35264
rect 2044 34536 2096 34542
rect 2042 34504 2044 34513
rect 2096 34504 2098 34513
rect 2042 34439 2098 34448
rect 2042 34096 2098 34105
rect 2042 34031 2044 34040
rect 2096 34031 2098 34040
rect 2044 34002 2096 34008
rect 2148 33130 2176 40446
rect 2228 39500 2280 39506
rect 2228 39442 2280 39448
rect 2240 38321 2268 39442
rect 2226 38312 2282 38321
rect 2226 38247 2282 38256
rect 2228 38208 2280 38214
rect 2228 38150 2280 38156
rect 2240 37806 2268 38150
rect 2228 37800 2280 37806
rect 2228 37742 2280 37748
rect 2228 36168 2280 36174
rect 2228 36110 2280 36116
rect 2240 34950 2268 36110
rect 2228 34944 2280 34950
rect 2228 34886 2280 34892
rect 1964 33102 2176 33130
rect 1768 32972 1820 32978
rect 1768 32914 1820 32920
rect 1676 29504 1728 29510
rect 1676 29446 1728 29452
rect 1688 29102 1716 29446
rect 1676 29096 1728 29102
rect 1676 29038 1728 29044
rect 1780 28506 1808 32914
rect 1860 30796 1912 30802
rect 1860 30738 1912 30744
rect 1872 30326 1900 30738
rect 1964 30734 1992 33102
rect 2044 32972 2096 32978
rect 2044 32914 2096 32920
rect 2056 32026 2084 32914
rect 2240 32366 2268 34886
rect 2228 32360 2280 32366
rect 2228 32302 2280 32308
rect 2136 32292 2188 32298
rect 2136 32234 2188 32240
rect 2044 32020 2096 32026
rect 2044 31962 2096 31968
rect 2148 31210 2176 32234
rect 2136 31204 2188 31210
rect 2136 31146 2188 31152
rect 1952 30728 2004 30734
rect 1952 30670 2004 30676
rect 1952 30592 2004 30598
rect 1952 30534 2004 30540
rect 1860 30320 1912 30326
rect 1860 30262 1912 30268
rect 1860 30116 1912 30122
rect 1860 30058 1912 30064
rect 1872 29209 1900 30058
rect 1964 29617 1992 30534
rect 1950 29608 2006 29617
rect 1950 29543 2006 29552
rect 1858 29200 1914 29209
rect 1858 29135 1914 29144
rect 1858 28792 1914 28801
rect 1858 28727 1914 28736
rect 1872 28694 1900 28727
rect 1860 28688 1912 28694
rect 1860 28630 1912 28636
rect 2148 28626 2176 31146
rect 2332 29646 2360 41550
rect 2424 41274 2452 42706
rect 2516 41750 2544 43114
rect 2608 42906 2636 44882
rect 2700 44470 2728 47058
rect 2780 46980 2832 46986
rect 2780 46922 2832 46928
rect 2792 46016 2820 46922
rect 2884 46345 2912 48010
rect 3056 47456 3108 47462
rect 3056 47398 3108 47404
rect 2964 47184 3016 47190
rect 2964 47126 3016 47132
rect 2870 46336 2926 46345
rect 2870 46271 2926 46280
rect 2792 45988 2912 46016
rect 2780 45892 2832 45898
rect 2780 45834 2832 45840
rect 2688 44464 2740 44470
rect 2688 44406 2740 44412
rect 2792 44305 2820 45834
rect 2884 44713 2912 45988
rect 2976 45121 3004 47126
rect 2962 45112 3018 45121
rect 2962 45047 3018 45056
rect 2870 44704 2926 44713
rect 2870 44639 2926 44648
rect 3068 44538 3096 47398
rect 3792 47252 3844 47258
rect 3792 47194 3844 47200
rect 3804 47161 3832 47194
rect 3790 47152 3846 47161
rect 3332 47116 3384 47122
rect 3790 47087 3846 47096
rect 3332 47058 3384 47064
rect 3344 46646 3372 47058
rect 3424 46912 3476 46918
rect 3424 46854 3476 46860
rect 3516 46912 3568 46918
rect 3516 46854 3568 46860
rect 3332 46640 3384 46646
rect 3332 46582 3384 46588
rect 3148 46368 3200 46374
rect 3148 46310 3200 46316
rect 3160 46034 3188 46310
rect 3148 46028 3200 46034
rect 3148 45970 3200 45976
rect 3332 46028 3384 46034
rect 3332 45970 3384 45976
rect 3148 45824 3200 45830
rect 3148 45766 3200 45772
rect 3056 44532 3108 44538
rect 3056 44474 3108 44480
rect 3056 44328 3108 44334
rect 2778 44296 2834 44305
rect 3056 44270 3108 44276
rect 2778 44231 2834 44240
rect 2688 43852 2740 43858
rect 2688 43794 2740 43800
rect 2596 42900 2648 42906
rect 2596 42842 2648 42848
rect 2596 42764 2648 42770
rect 2596 42706 2648 42712
rect 2608 42362 2636 42706
rect 2596 42356 2648 42362
rect 2596 42298 2648 42304
rect 2700 42090 2728 43794
rect 2780 43716 2832 43722
rect 2780 43658 2832 43664
rect 2792 43081 2820 43658
rect 2964 43104 3016 43110
rect 2778 43072 2834 43081
rect 2964 43046 3016 43052
rect 2778 43007 2834 43016
rect 2780 42628 2832 42634
rect 2780 42570 2832 42576
rect 2688 42084 2740 42090
rect 2688 42026 2740 42032
rect 2792 41857 2820 42570
rect 2872 42288 2924 42294
rect 2872 42230 2924 42236
rect 2778 41848 2834 41857
rect 2884 41818 2912 42230
rect 2778 41783 2834 41792
rect 2872 41812 2924 41818
rect 2872 41754 2924 41760
rect 2504 41744 2556 41750
rect 2504 41686 2556 41692
rect 2976 41449 3004 43046
rect 3068 41682 3096 44270
rect 3056 41676 3108 41682
rect 3056 41618 3108 41624
rect 3160 41614 3188 45766
rect 3344 45626 3372 45970
rect 3436 45937 3464 46854
rect 3528 46753 3556 46854
rect 3514 46744 3570 46753
rect 3514 46679 3570 46688
rect 3976 46504 4028 46510
rect 3976 46446 4028 46452
rect 3516 45960 3568 45966
rect 3422 45928 3478 45937
rect 3516 45902 3568 45908
rect 3608 45960 3660 45966
rect 3608 45902 3660 45908
rect 3422 45863 3478 45872
rect 3332 45620 3384 45626
rect 3332 45562 3384 45568
rect 3528 45558 3556 45902
rect 3516 45552 3568 45558
rect 3516 45494 3568 45500
rect 3240 45416 3292 45422
rect 3240 45358 3292 45364
rect 3252 44878 3280 45358
rect 3620 45354 3648 45902
rect 3608 45348 3660 45354
rect 3608 45290 3660 45296
rect 3332 45280 3384 45286
rect 3332 45222 3384 45228
rect 3240 44872 3292 44878
rect 3240 44814 3292 44820
rect 3344 43178 3372 45222
rect 3620 44878 3648 45290
rect 3988 45286 4016 46446
rect 3976 45280 4028 45286
rect 3976 45222 4028 45228
rect 3516 44872 3568 44878
rect 3516 44814 3568 44820
rect 3608 44872 3660 44878
rect 3608 44814 3660 44820
rect 3424 43988 3476 43994
rect 3424 43930 3476 43936
rect 3436 43897 3464 43930
rect 3422 43888 3478 43897
rect 3422 43823 3478 43832
rect 3332 43172 3384 43178
rect 3332 43114 3384 43120
rect 3528 42514 3556 44814
rect 3608 44736 3660 44742
rect 3608 44678 3660 44684
rect 3620 42702 3648 44678
rect 3976 43784 4028 43790
rect 3976 43726 4028 43732
rect 3608 42696 3660 42702
rect 3608 42638 3660 42644
rect 3884 42560 3936 42566
rect 3528 42486 3648 42514
rect 3884 42502 3936 42508
rect 3148 41608 3200 41614
rect 3148 41550 3200 41556
rect 3516 41540 3568 41546
rect 3516 41482 3568 41488
rect 2962 41440 3018 41449
rect 2962 41375 3018 41384
rect 2412 41268 2464 41274
rect 2412 41210 2464 41216
rect 3056 40996 3108 41002
rect 3056 40938 3108 40944
rect 2504 40928 2556 40934
rect 2504 40870 2556 40876
rect 2516 40730 2544 40870
rect 2504 40724 2556 40730
rect 2504 40666 2556 40672
rect 2688 40588 2740 40594
rect 2688 40530 2740 40536
rect 2412 39908 2464 39914
rect 2412 39850 2464 39856
rect 2596 39908 2648 39914
rect 2596 39850 2648 39856
rect 2424 37466 2452 39850
rect 2504 39500 2556 39506
rect 2504 39442 2556 39448
rect 2516 37670 2544 39442
rect 2608 39030 2636 39850
rect 2700 39438 2728 40530
rect 3068 40186 3096 40938
rect 3148 40928 3200 40934
rect 3148 40870 3200 40876
rect 3160 40633 3188 40870
rect 3146 40624 3202 40633
rect 3146 40559 3202 40568
rect 3332 40520 3384 40526
rect 3332 40462 3384 40468
rect 3056 40180 3108 40186
rect 3056 40122 3108 40128
rect 2780 39908 2832 39914
rect 2780 39850 2832 39856
rect 2688 39432 2740 39438
rect 2792 39409 2820 39850
rect 2688 39374 2740 39380
rect 2778 39400 2834 39409
rect 2778 39335 2834 39344
rect 2872 39364 2924 39370
rect 2872 39306 2924 39312
rect 2688 39092 2740 39098
rect 2688 39034 2740 39040
rect 2596 39024 2648 39030
rect 2596 38966 2648 38972
rect 2596 38412 2648 38418
rect 2596 38354 2648 38360
rect 2608 37806 2636 38354
rect 2596 37800 2648 37806
rect 2596 37742 2648 37748
rect 2504 37664 2556 37670
rect 2504 37606 2556 37612
rect 2412 37460 2464 37466
rect 2412 37402 2464 37408
rect 2412 37324 2464 37330
rect 2412 37266 2464 37272
rect 2596 37324 2648 37330
rect 2596 37266 2648 37272
rect 2424 35834 2452 37266
rect 2608 36854 2636 37266
rect 2596 36848 2648 36854
rect 2596 36790 2648 36796
rect 2700 36786 2728 39034
rect 2884 38593 2912 39306
rect 2964 39296 3016 39302
rect 2964 39238 3016 39244
rect 2870 38584 2926 38593
rect 2870 38519 2926 38528
rect 2780 38208 2832 38214
rect 2780 38150 2832 38156
rect 2792 37777 2820 38150
rect 2872 38004 2924 38010
rect 2872 37946 2924 37952
rect 2778 37768 2834 37777
rect 2778 37703 2834 37712
rect 2884 37670 2912 37946
rect 2872 37664 2924 37670
rect 2872 37606 2924 37612
rect 2872 37392 2924 37398
rect 2976 37369 3004 39238
rect 3240 38888 3292 38894
rect 3240 38830 3292 38836
rect 3056 38820 3108 38826
rect 3056 38762 3108 38768
rect 3068 38486 3096 38762
rect 3056 38480 3108 38486
rect 3056 38422 3108 38428
rect 3252 38010 3280 38830
rect 3240 38004 3292 38010
rect 3240 37946 3292 37952
rect 3148 37800 3200 37806
rect 3148 37742 3200 37748
rect 3056 37732 3108 37738
rect 3056 37674 3108 37680
rect 2872 37334 2924 37340
rect 2962 37360 3018 37369
rect 2780 37188 2832 37194
rect 2780 37130 2832 37136
rect 2792 36961 2820 37130
rect 2778 36952 2834 36961
rect 2778 36887 2834 36896
rect 2688 36780 2740 36786
rect 2688 36722 2740 36728
rect 2596 36644 2648 36650
rect 2596 36586 2648 36592
rect 2780 36644 2832 36650
rect 2780 36586 2832 36592
rect 2412 35828 2464 35834
rect 2412 35770 2464 35776
rect 2412 34944 2464 34950
rect 2412 34886 2464 34892
rect 2424 34746 2452 34886
rect 2412 34740 2464 34746
rect 2412 34682 2464 34688
rect 2608 34678 2636 36586
rect 2792 36145 2820 36586
rect 2778 36136 2834 36145
rect 2778 36071 2834 36080
rect 2884 35737 2912 37334
rect 2962 37295 3018 37304
rect 3068 36242 3096 37674
rect 3160 36242 3188 37742
rect 3056 36236 3108 36242
rect 3056 36178 3108 36184
rect 3148 36236 3200 36242
rect 3148 36178 3200 36184
rect 3160 35766 3188 36178
rect 3344 35766 3372 40462
rect 3424 37664 3476 37670
rect 3424 37606 3476 37612
rect 3148 35760 3200 35766
rect 2870 35728 2926 35737
rect 3148 35702 3200 35708
rect 3332 35760 3384 35766
rect 3332 35702 3384 35708
rect 2870 35663 2926 35672
rect 2872 35488 2924 35494
rect 2872 35430 2924 35436
rect 2596 34672 2648 34678
rect 2596 34614 2648 34620
rect 2780 34536 2832 34542
rect 2780 34478 2832 34484
rect 2596 34468 2648 34474
rect 2596 34410 2648 34416
rect 2412 34060 2464 34066
rect 2412 34002 2464 34008
rect 2424 32502 2452 34002
rect 2504 33448 2556 33454
rect 2504 33390 2556 33396
rect 2412 32496 2464 32502
rect 2412 32438 2464 32444
rect 2516 31890 2544 33390
rect 2608 33046 2636 34410
rect 2688 33448 2740 33454
rect 2688 33390 2740 33396
rect 2596 33040 2648 33046
rect 2596 32982 2648 32988
rect 2700 32842 2728 33390
rect 2688 32836 2740 32842
rect 2688 32778 2740 32784
rect 2700 32450 2728 32778
rect 2792 32473 2820 34478
rect 2608 32422 2728 32450
rect 2778 32464 2834 32473
rect 2608 32366 2636 32422
rect 2778 32399 2834 32408
rect 2596 32360 2648 32366
rect 2596 32302 2648 32308
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2608 31958 2636 32302
rect 2792 32026 2820 32302
rect 2780 32020 2832 32026
rect 2780 31962 2832 31968
rect 2596 31952 2648 31958
rect 2596 31894 2648 31900
rect 2504 31884 2556 31890
rect 2504 31826 2556 31832
rect 2504 31408 2556 31414
rect 2504 31350 2556 31356
rect 2412 30048 2464 30054
rect 2412 29990 2464 29996
rect 2228 29640 2280 29646
rect 2228 29582 2280 29588
rect 2320 29640 2372 29646
rect 2320 29582 2372 29588
rect 2240 28762 2268 29582
rect 2228 28756 2280 28762
rect 2228 28698 2280 28704
rect 2136 28620 2188 28626
rect 2136 28562 2188 28568
rect 1780 28478 1900 28506
rect 1768 28144 1820 28150
rect 1766 28112 1768 28121
rect 1820 28112 1822 28121
rect 1766 28047 1822 28056
rect 1768 27600 1820 27606
rect 1768 27542 1820 27548
rect 1676 27532 1728 27538
rect 1676 27474 1728 27480
rect 1688 27062 1716 27474
rect 1676 27056 1728 27062
rect 1676 26998 1728 27004
rect 1780 26586 1808 27542
rect 1768 26580 1820 26586
rect 1768 26522 1820 26528
rect 1872 26234 1900 28478
rect 2044 28484 2096 28490
rect 2044 28426 2096 28432
rect 1952 28008 2004 28014
rect 1952 27950 2004 27956
rect 1964 27577 1992 27950
rect 2056 27674 2084 28426
rect 2044 27668 2096 27674
rect 2044 27610 2096 27616
rect 1950 27568 2006 27577
rect 1950 27503 2006 27512
rect 2044 27532 2096 27538
rect 2044 27474 2096 27480
rect 1952 26920 2004 26926
rect 1952 26862 2004 26868
rect 1964 26761 1992 26862
rect 1950 26752 2006 26761
rect 1950 26687 2006 26696
rect 1952 26444 2004 26450
rect 1952 26386 2004 26392
rect 1964 26353 1992 26386
rect 1950 26344 2006 26353
rect 1950 26279 2006 26288
rect 1596 26206 1716 26234
rect 1872 26206 1992 26234
rect 1584 25220 1636 25226
rect 1584 25162 1636 25168
rect 1596 24682 1624 25162
rect 1584 24676 1636 24682
rect 1584 24618 1636 24624
rect 1492 24608 1544 24614
rect 1492 24550 1544 24556
rect 1400 23180 1452 23186
rect 1400 23122 1452 23128
rect 1412 22273 1440 23122
rect 1398 22264 1454 22273
rect 1398 22199 1454 22208
rect 1504 22080 1532 24550
rect 1584 23588 1636 23594
rect 1584 23530 1636 23536
rect 1596 22681 1624 23530
rect 1582 22672 1638 22681
rect 1582 22607 1638 22616
rect 1412 22052 1532 22080
rect 1584 22092 1636 22098
rect 1412 21554 1440 22052
rect 1584 22034 1636 22040
rect 1492 21888 1544 21894
rect 1492 21830 1544 21836
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1412 18766 1440 21490
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1412 15026 1440 18702
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 1412 12238 1440 14962
rect 1504 13802 1532 21830
rect 1596 21049 1624 22034
rect 1688 21486 1716 26206
rect 1858 25936 1914 25945
rect 1768 25900 1820 25906
rect 1858 25871 1914 25880
rect 1768 25842 1820 25848
rect 1780 25650 1808 25842
rect 1872 25838 1900 25871
rect 1860 25832 1912 25838
rect 1860 25774 1912 25780
rect 1780 25622 1900 25650
rect 1766 25528 1822 25537
rect 1766 25463 1822 25472
rect 1780 25430 1808 25463
rect 1768 25424 1820 25430
rect 1768 25366 1820 25372
rect 1768 24676 1820 24682
rect 1768 24618 1820 24624
rect 1780 24562 1808 24618
rect 1872 24562 1900 25622
rect 1780 24534 1900 24562
rect 1872 23730 1900 24534
rect 1964 24426 1992 26206
rect 2056 25906 2084 27474
rect 2044 25900 2096 25906
rect 2044 25842 2096 25848
rect 2044 25764 2096 25770
rect 2044 25706 2096 25712
rect 2056 24682 2084 25706
rect 2148 25430 2176 28562
rect 2228 26308 2280 26314
rect 2228 26250 2280 26256
rect 2136 25424 2188 25430
rect 2136 25366 2188 25372
rect 2240 24750 2268 26250
rect 2332 25702 2360 29582
rect 2424 28937 2452 29990
rect 2410 28928 2466 28937
rect 2410 28863 2466 28872
rect 2424 27538 2452 28863
rect 2516 28218 2544 31350
rect 2688 31272 2740 31278
rect 2688 31214 2740 31220
rect 2596 30796 2648 30802
rect 2596 30738 2648 30744
rect 2608 29850 2636 30738
rect 2596 29844 2648 29850
rect 2596 29786 2648 29792
rect 2700 29170 2728 31214
rect 2780 30660 2832 30666
rect 2780 30602 2832 30608
rect 2792 30025 2820 30602
rect 2884 30258 2912 35430
rect 3160 35170 3188 35702
rect 3240 35488 3292 35494
rect 3240 35430 3292 35436
rect 3252 35290 3280 35430
rect 3240 35284 3292 35290
rect 3240 35226 3292 35232
rect 3160 35154 3280 35170
rect 3436 35154 3464 37606
rect 3528 37330 3556 41482
rect 3620 40526 3648 42486
rect 3700 41676 3752 41682
rect 3700 41618 3752 41624
rect 3712 40594 3740 41618
rect 3792 41608 3844 41614
rect 3792 41550 3844 41556
rect 3700 40588 3752 40594
rect 3700 40530 3752 40536
rect 3608 40520 3660 40526
rect 3608 40462 3660 40468
rect 3606 39808 3662 39817
rect 3606 39743 3662 39752
rect 3620 39642 3648 39743
rect 3608 39636 3660 39642
rect 3608 39578 3660 39584
rect 3516 37324 3568 37330
rect 3516 37266 3568 37272
rect 3608 37256 3660 37262
rect 3608 37198 3660 37204
rect 3620 36854 3648 37198
rect 3608 36848 3660 36854
rect 3608 36790 3660 36796
rect 3516 35760 3568 35766
rect 3516 35702 3568 35708
rect 3160 35148 3292 35154
rect 3160 35142 3240 35148
rect 3240 35090 3292 35096
rect 3424 35148 3476 35154
rect 3424 35090 3476 35096
rect 3148 35080 3200 35086
rect 3148 35022 3200 35028
rect 3056 33924 3108 33930
rect 3056 33866 3108 33872
rect 2964 32360 3016 32366
rect 2964 32302 3016 32308
rect 2872 30252 2924 30258
rect 2872 30194 2924 30200
rect 2778 30016 2834 30025
rect 2778 29951 2834 29960
rect 2780 29708 2832 29714
rect 2780 29650 2832 29656
rect 2688 29164 2740 29170
rect 2688 29106 2740 29112
rect 2792 29102 2820 29650
rect 2780 29096 2832 29102
rect 2780 29038 2832 29044
rect 2504 28212 2556 28218
rect 2504 28154 2556 28160
rect 2412 27532 2464 27538
rect 2412 27474 2464 27480
rect 2412 26580 2464 26586
rect 2412 26522 2464 26528
rect 2320 25696 2372 25702
rect 2320 25638 2372 25644
rect 2228 24744 2280 24750
rect 2228 24686 2280 24692
rect 2044 24676 2096 24682
rect 2044 24618 2096 24624
rect 1964 24398 2084 24426
rect 1952 24268 2004 24274
rect 1952 24210 2004 24216
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1768 23248 1820 23254
rect 1768 23190 1820 23196
rect 1676 21480 1728 21486
rect 1676 21422 1728 21428
rect 1780 21418 1808 23190
rect 1872 21978 1900 23666
rect 1964 23497 1992 24210
rect 1950 23488 2006 23497
rect 1950 23423 2006 23432
rect 2056 22778 2084 24398
rect 2136 23588 2188 23594
rect 2136 23530 2188 23536
rect 2044 22772 2096 22778
rect 2044 22714 2096 22720
rect 2044 22500 2096 22506
rect 2044 22442 2096 22448
rect 2056 22234 2084 22442
rect 2044 22228 2096 22234
rect 2044 22170 2096 22176
rect 2148 22166 2176 23530
rect 2136 22160 2188 22166
rect 2136 22102 2188 22108
rect 1872 21950 2084 21978
rect 2056 21418 2084 21950
rect 2148 21418 2176 22102
rect 2332 22098 2360 25638
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2228 22024 2280 22030
rect 2228 21966 2280 21972
rect 1768 21412 1820 21418
rect 1768 21354 1820 21360
rect 2044 21412 2096 21418
rect 2044 21354 2096 21360
rect 2136 21412 2188 21418
rect 2136 21354 2188 21360
rect 1582 21040 1638 21049
rect 1582 20975 1638 20984
rect 1676 21004 1728 21010
rect 1676 20946 1728 20952
rect 1688 20233 1716 20946
rect 1952 20392 2004 20398
rect 1952 20334 2004 20340
rect 1674 20224 1730 20233
rect 1674 20159 1730 20168
rect 1860 19916 1912 19922
rect 1860 19858 1912 19864
rect 1872 19417 1900 19858
rect 1964 19825 1992 20334
rect 1950 19816 2006 19825
rect 1950 19751 2006 19760
rect 1858 19408 1914 19417
rect 1858 19343 1914 19352
rect 1860 19236 1912 19242
rect 1860 19178 1912 19184
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1596 18970 1624 19110
rect 1872 19009 1900 19178
rect 1858 19000 1914 19009
rect 1584 18964 1636 18970
rect 1858 18935 1914 18944
rect 1584 18906 1636 18912
rect 1768 18896 1820 18902
rect 1768 18838 1820 18844
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1596 14890 1624 15506
rect 1584 14884 1636 14890
rect 1584 14826 1636 14832
rect 1492 13796 1544 13802
rect 1492 13738 1544 13744
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1596 12442 1624 12786
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 9586 1440 12174
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1504 10849 1532 11630
rect 1490 10840 1546 10849
rect 1490 10775 1546 10784
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 1596 10033 1624 10066
rect 1582 10024 1638 10033
rect 1582 9959 1638 9968
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 6322 1440 9522
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1504 6769 1532 7890
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1490 6760 1546 6769
rect 1490 6695 1546 6704
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1596 6118 1624 7142
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5302 1624 6054
rect 1584 5296 1636 5302
rect 1584 5238 1636 5244
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 664 2508 716 2514
rect 664 2450 716 2456
rect 676 800 704 2450
rect 662 -800 718 800
rect 1412 241 1440 4626
rect 1688 4146 1716 17138
rect 1780 16794 1808 18838
rect 2056 18834 2084 21354
rect 2136 20800 2188 20806
rect 2136 20742 2188 20748
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 1860 18080 1912 18086
rect 1860 18022 1912 18028
rect 1872 17814 1900 18022
rect 1860 17808 1912 17814
rect 1860 17750 1912 17756
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1964 16969 1992 17070
rect 1950 16960 2006 16969
rect 1950 16895 2006 16904
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1964 16561 1992 16594
rect 1950 16552 2006 16561
rect 1950 16487 2006 16496
rect 1858 16144 1914 16153
rect 1858 16079 1914 16088
rect 1872 16046 1900 16079
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1952 15904 2004 15910
rect 1952 15846 2004 15852
rect 1858 15736 1914 15745
rect 1858 15671 1914 15680
rect 1872 15638 1900 15671
rect 1860 15632 1912 15638
rect 1860 15574 1912 15580
rect 1964 15065 1992 15846
rect 1950 15056 2006 15065
rect 1950 14991 2006 15000
rect 1768 14952 1820 14958
rect 2056 14906 2084 18770
rect 1820 14900 2084 14906
rect 1768 14894 2084 14900
rect 1780 14878 2084 14894
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1780 14618 1808 14758
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 1860 13388 1912 13394
rect 1860 13330 1912 13336
rect 1872 12889 1900 13330
rect 1964 13297 1992 14418
rect 1950 13288 2006 13297
rect 1950 13223 2006 13232
rect 1858 12880 1914 12889
rect 1858 12815 1914 12824
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 1872 12481 1900 12650
rect 1858 12472 1914 12481
rect 1858 12407 1914 12416
rect 2056 12306 2084 14878
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 1964 10441 1992 11154
rect 1950 10432 2006 10441
rect 1950 10367 2006 10376
rect 1858 9616 1914 9625
rect 1858 9551 1914 9560
rect 1872 9110 1900 9551
rect 2056 9450 2084 12242
rect 2148 10674 2176 20742
rect 2240 20330 2268 21966
rect 2228 20324 2280 20330
rect 2228 20266 2280 20272
rect 2240 10810 2268 20266
rect 2332 18290 2360 22034
rect 2424 21894 2452 26522
rect 2516 26450 2544 28154
rect 2688 27464 2740 27470
rect 2688 27406 2740 27412
rect 2504 26444 2556 26450
rect 2504 26386 2556 26392
rect 2516 25362 2544 26386
rect 2504 25356 2556 25362
rect 2504 25298 2556 25304
rect 2596 25356 2648 25362
rect 2596 25298 2648 25304
rect 2504 24744 2556 24750
rect 2504 24686 2556 24692
rect 2516 24614 2544 24686
rect 2504 24608 2556 24614
rect 2504 24550 2556 24556
rect 2504 24336 2556 24342
rect 2504 24278 2556 24284
rect 2516 23866 2544 24278
rect 2504 23860 2556 23866
rect 2504 23802 2556 23808
rect 2608 23746 2636 25298
rect 2700 24750 2728 27406
rect 2778 27160 2834 27169
rect 2778 27095 2834 27104
rect 2792 26926 2820 27095
rect 2780 26920 2832 26926
rect 2780 26862 2832 26868
rect 2976 26586 3004 32302
rect 3068 32065 3096 33866
rect 3160 33658 3188 35022
rect 3148 33652 3200 33658
rect 3148 33594 3200 33600
rect 3436 33454 3464 35090
rect 3148 33448 3200 33454
rect 3148 33390 3200 33396
rect 3424 33448 3476 33454
rect 3424 33390 3476 33396
rect 3054 32056 3110 32065
rect 3160 32026 3188 33390
rect 3436 32910 3464 33390
rect 3424 32904 3476 32910
rect 3424 32846 3476 32852
rect 3054 31991 3110 32000
rect 3148 32020 3200 32026
rect 3148 31962 3200 31968
rect 3056 31884 3108 31890
rect 3056 31826 3108 31832
rect 3068 29578 3096 31826
rect 3240 31136 3292 31142
rect 3240 31078 3292 31084
rect 3332 31136 3384 31142
rect 3332 31078 3384 31084
rect 3252 30841 3280 31078
rect 3238 30832 3294 30841
rect 3238 30767 3294 30776
rect 3240 30728 3292 30734
rect 3344 30682 3372 31078
rect 3528 30802 3556 35702
rect 3608 35624 3660 35630
rect 3608 35566 3660 35572
rect 3620 35290 3648 35566
rect 3608 35284 3660 35290
rect 3608 35226 3660 35232
rect 3608 33312 3660 33318
rect 3606 33280 3608 33289
rect 3660 33280 3662 33289
rect 3606 33215 3662 33224
rect 3608 32020 3660 32026
rect 3608 31962 3660 31968
rect 3516 30796 3568 30802
rect 3516 30738 3568 30744
rect 3292 30676 3372 30682
rect 3240 30670 3372 30676
rect 3252 30654 3372 30670
rect 3056 29572 3108 29578
rect 3056 29514 3108 29520
rect 3148 28416 3200 28422
rect 3148 28358 3200 28364
rect 3160 28082 3188 28358
rect 3148 28076 3200 28082
rect 3148 28018 3200 28024
rect 3054 27976 3110 27985
rect 3252 27946 3280 30654
rect 3332 30048 3384 30054
rect 3332 29990 3384 29996
rect 3344 29782 3372 29990
rect 3332 29776 3384 29782
rect 3332 29718 3384 29724
rect 3054 27911 3110 27920
rect 3240 27940 3292 27946
rect 3068 26926 3096 27911
rect 3240 27882 3292 27888
rect 3148 27872 3200 27878
rect 3148 27814 3200 27820
rect 3160 27674 3188 27814
rect 3148 27668 3200 27674
rect 3148 27610 3200 27616
rect 3056 26920 3108 26926
rect 3056 26862 3108 26868
rect 2964 26580 3016 26586
rect 2964 26522 3016 26528
rect 3056 26444 3108 26450
rect 3056 26386 3108 26392
rect 2688 24744 2740 24750
rect 3068 24721 3096 26386
rect 2688 24686 2740 24692
rect 3054 24712 3110 24721
rect 3054 24647 3110 24656
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2516 23718 2636 23746
rect 2412 21888 2464 21894
rect 2412 21830 2464 21836
rect 2412 19780 2464 19786
rect 2412 19722 2464 19728
rect 2424 18834 2452 19722
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 2332 14074 2360 18022
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2332 13530 2360 14010
rect 2424 13852 2452 18362
rect 2516 15178 2544 23718
rect 2700 23322 2728 24550
rect 3148 24268 3200 24274
rect 3148 24210 3200 24216
rect 2872 24200 2924 24206
rect 2872 24142 2924 24148
rect 2778 23896 2834 23905
rect 2778 23831 2834 23840
rect 2792 23662 2820 23831
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2688 23316 2740 23322
rect 2688 23258 2740 23264
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2792 23089 2820 23122
rect 2778 23080 2834 23089
rect 2778 23015 2834 23024
rect 2884 22982 2912 24142
rect 3160 23322 3188 24210
rect 3148 23316 3200 23322
rect 3148 23258 3200 23264
rect 2872 22976 2924 22982
rect 2872 22918 2924 22924
rect 2596 22772 2648 22778
rect 2596 22714 2648 22720
rect 2608 19258 2636 22714
rect 2884 22574 2912 22918
rect 2872 22568 2924 22574
rect 2872 22510 2924 22516
rect 2780 22432 2832 22438
rect 2780 22374 2832 22380
rect 2792 22234 2820 22374
rect 2780 22228 2832 22234
rect 2780 22170 2832 22176
rect 2792 22098 2820 22170
rect 2780 22092 2832 22098
rect 2780 22034 2832 22040
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 2688 21344 2740 21350
rect 2688 21286 2740 21292
rect 2700 20602 2728 21286
rect 2964 20868 3016 20874
rect 2964 20810 3016 20816
rect 2778 20632 2834 20641
rect 2688 20596 2740 20602
rect 2976 20602 3004 20810
rect 2778 20567 2834 20576
rect 2964 20596 3016 20602
rect 2688 20538 2740 20544
rect 2792 19922 2820 20567
rect 2964 20538 3016 20544
rect 2964 20460 3016 20466
rect 2964 20402 3016 20408
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2976 19310 3004 20402
rect 3160 19922 3188 21383
rect 3252 21010 3280 27882
rect 3528 27402 3556 30738
rect 3516 27396 3568 27402
rect 3516 27338 3568 27344
rect 3424 25288 3476 25294
rect 3424 25230 3476 25236
rect 3330 24304 3386 24313
rect 3330 24239 3386 24248
rect 3344 23662 3372 24239
rect 3332 23656 3384 23662
rect 3332 23598 3384 23604
rect 3332 21412 3384 21418
rect 3332 21354 3384 21360
rect 3240 21004 3292 21010
rect 3240 20946 3292 20952
rect 3148 19916 3200 19922
rect 3148 19858 3200 19864
rect 3344 19786 3372 21354
rect 3332 19780 3384 19786
rect 3332 19722 3384 19728
rect 2872 19304 2924 19310
rect 2608 19230 2820 19258
rect 2872 19246 2924 19252
rect 2964 19304 3016 19310
rect 3016 19252 3096 19258
rect 2964 19246 3096 19252
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2700 18986 2728 19110
rect 2608 18970 2728 18986
rect 2792 18970 2820 19230
rect 2596 18964 2728 18970
rect 2648 18958 2728 18964
rect 2596 18906 2648 18912
rect 2700 18358 2728 18958
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 2688 18352 2740 18358
rect 2688 18294 2740 18300
rect 2884 18193 2912 19246
rect 2976 19230 3096 19246
rect 3068 18222 3096 19230
rect 3436 18952 3464 25230
rect 3528 21010 3556 27338
rect 3516 21004 3568 21010
rect 3516 20946 3568 20952
rect 3436 18924 3556 18952
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3436 18601 3464 18770
rect 3422 18592 3478 18601
rect 3422 18527 3478 18536
rect 3056 18216 3108 18222
rect 2870 18184 2926 18193
rect 2780 18148 2832 18154
rect 3056 18158 3108 18164
rect 2870 18119 2926 18128
rect 2780 18090 2832 18096
rect 2792 17882 2820 18090
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2792 17490 2820 17818
rect 3238 17776 3294 17785
rect 3056 17740 3108 17746
rect 3238 17711 3294 17720
rect 3056 17682 3108 17688
rect 2964 17604 3016 17610
rect 2964 17546 3016 17552
rect 2792 17462 2912 17490
rect 2778 17368 2834 17377
rect 2778 17303 2834 17312
rect 2688 17060 2740 17066
rect 2688 17002 2740 17008
rect 2700 16726 2728 17002
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 2792 16658 2820 17303
rect 2884 17134 2912 17462
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2608 15638 2636 16458
rect 2976 15978 3004 17546
rect 3068 17338 3096 17682
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3252 16658 3280 17711
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2976 15570 3004 15914
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2516 15162 2820 15178
rect 2516 15156 2832 15162
rect 2516 15150 2780 15156
rect 2502 15056 2558 15065
rect 2502 14991 2558 15000
rect 2516 14958 2544 14991
rect 2504 14952 2556 14958
rect 2504 14894 2556 14900
rect 2502 14648 2558 14657
rect 2502 14583 2504 14592
rect 2556 14583 2558 14592
rect 2504 14554 2556 14560
rect 2608 13938 2636 15150
rect 2780 15098 2832 15104
rect 2872 14884 2924 14890
rect 2872 14826 2924 14832
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 14113 2820 14418
rect 2778 14104 2834 14113
rect 2884 14074 2912 14826
rect 2778 14039 2834 14048
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2504 13864 2556 13870
rect 2424 13824 2504 13852
rect 2504 13806 2556 13812
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2332 12306 2360 13194
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2332 11558 2360 12242
rect 2412 11688 2464 11694
rect 2410 11656 2412 11665
rect 2464 11656 2466 11665
rect 2410 11591 2466 11600
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2148 10198 2176 10610
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 2240 10130 2268 10746
rect 2228 10124 2280 10130
rect 2228 10066 2280 10072
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2044 9444 2096 9450
rect 2044 9386 2096 9392
rect 2320 9444 2372 9450
rect 2320 9386 2372 9392
rect 1860 9104 1912 9110
rect 1860 9046 1912 9052
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1964 7585 1992 8366
rect 1950 7576 2006 7585
rect 1950 7511 2006 7520
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1872 6254 1900 7278
rect 2056 6254 2084 9386
rect 2332 8838 2360 9386
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2424 8634 2452 9454
rect 2412 8628 2464 8634
rect 2332 8588 2412 8616
rect 2332 8362 2360 8588
rect 2412 8570 2464 8576
rect 2412 8424 2464 8430
rect 2410 8392 2412 8401
rect 2464 8392 2466 8401
rect 2320 8356 2372 8362
rect 2410 8327 2466 8336
rect 2320 8298 2372 8304
rect 2516 8242 2544 13806
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2608 12442 2636 13330
rect 2976 12782 3004 15506
rect 3344 15337 3372 16594
rect 3330 15328 3386 15337
rect 3330 15263 3386 15272
rect 3528 14822 3556 18924
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3422 14512 3478 14521
rect 3422 14447 3478 14456
rect 3332 14000 3384 14006
rect 3332 13942 3384 13948
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3068 13705 3096 13806
rect 3054 13696 3110 13705
rect 3054 13631 3110 13640
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2240 8214 2544 8242
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2148 6254 2176 6802
rect 2240 6798 2268 8214
rect 2608 8106 2636 12378
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2700 10266 2728 12310
rect 2792 12073 2820 12718
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2778 12064 2834 12073
rect 2778 11999 2834 12008
rect 2884 11898 2912 12174
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2778 11248 2834 11257
rect 3252 11218 3280 12378
rect 3344 12306 3372 13942
rect 3436 13394 3464 14447
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3528 13530 3556 13670
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3620 12170 3648 31962
rect 3712 24614 3740 40530
rect 3804 40390 3832 41550
rect 3792 40384 3844 40390
rect 3792 40326 3844 40332
rect 3790 40216 3846 40225
rect 3790 40151 3846 40160
rect 3804 39438 3832 40151
rect 3896 39506 3924 42502
rect 3988 42158 4016 43726
rect 3976 42152 4028 42158
rect 3976 42094 4028 42100
rect 3988 41138 4016 42094
rect 3976 41132 4028 41138
rect 3976 41074 4028 41080
rect 3884 39500 3936 39506
rect 3884 39442 3936 39448
rect 3976 39500 4028 39506
rect 3976 39442 4028 39448
rect 3792 39432 3844 39438
rect 3792 39374 3844 39380
rect 3896 38894 3924 39442
rect 3988 39098 4016 39442
rect 3976 39092 4028 39098
rect 3976 39034 4028 39040
rect 3884 38888 3936 38894
rect 3884 38830 3936 38836
rect 3884 38752 3936 38758
rect 3884 38694 3936 38700
rect 3896 38350 3924 38694
rect 3884 38344 3936 38350
rect 3884 38286 3936 38292
rect 3976 37188 4028 37194
rect 3976 37130 4028 37136
rect 3884 36032 3936 36038
rect 3884 35974 3936 35980
rect 3896 35698 3924 35974
rect 3884 35692 3936 35698
rect 3884 35634 3936 35640
rect 3988 34610 4016 37130
rect 3976 34604 4028 34610
rect 3976 34546 4028 34552
rect 3884 34196 3936 34202
rect 3884 34138 3936 34144
rect 3896 32842 3924 34138
rect 3884 32836 3936 32842
rect 3884 32778 3936 32784
rect 3792 32768 3844 32774
rect 3792 32710 3844 32716
rect 3804 31958 3832 32710
rect 3792 31952 3844 31958
rect 3792 31894 3844 31900
rect 4080 31754 4108 51046
rect 4712 49292 4764 49298
rect 4712 49234 4764 49240
rect 4160 48816 4212 48822
rect 4160 48758 4212 48764
rect 4172 47530 4200 48758
rect 4436 48612 4488 48618
rect 4436 48554 4488 48560
rect 4252 48544 4304 48550
rect 4252 48486 4304 48492
rect 4264 48278 4292 48486
rect 4252 48272 4304 48278
rect 4252 48214 4304 48220
rect 4160 47524 4212 47530
rect 4160 47466 4212 47472
rect 4448 46510 4476 48554
rect 4620 48544 4672 48550
rect 4620 48486 4672 48492
rect 4632 48346 4660 48486
rect 4724 48346 4752 49234
rect 5184 48890 5212 51342
rect 5264 49088 5316 49094
rect 5264 49030 5316 49036
rect 5172 48884 5224 48890
rect 5172 48826 5224 48832
rect 5172 48748 5224 48754
rect 5172 48690 5224 48696
rect 4620 48340 4672 48346
rect 4620 48282 4672 48288
rect 4712 48340 4764 48346
rect 4712 48282 4764 48288
rect 4632 47598 4660 48282
rect 5184 47666 5212 48690
rect 5276 48686 5304 49030
rect 5264 48680 5316 48686
rect 5264 48622 5316 48628
rect 5276 48346 5304 48622
rect 5264 48340 5316 48346
rect 5264 48282 5316 48288
rect 5172 47660 5224 47666
rect 5172 47602 5224 47608
rect 4620 47592 4672 47598
rect 4620 47534 4672 47540
rect 4896 47524 4948 47530
rect 4896 47466 4948 47472
rect 4620 47456 4672 47462
rect 4620 47398 4672 47404
rect 4436 46504 4488 46510
rect 4436 46446 4488 46452
rect 4344 46368 4396 46374
rect 4344 46310 4396 46316
rect 4252 46096 4304 46102
rect 4252 46038 4304 46044
rect 4160 45892 4212 45898
rect 4160 45834 4212 45840
rect 4172 45082 4200 45834
rect 4160 45076 4212 45082
rect 4160 45018 4212 45024
rect 4160 43240 4212 43246
rect 4160 43182 4212 43188
rect 4172 42702 4200 43182
rect 4160 42696 4212 42702
rect 4160 42638 4212 42644
rect 4264 42566 4292 46038
rect 4356 45082 4384 46310
rect 4344 45076 4396 45082
rect 4344 45018 4396 45024
rect 4344 44396 4396 44402
rect 4344 44338 4396 44344
rect 4252 42560 4304 42566
rect 4252 42502 4304 42508
rect 4356 42226 4384 44338
rect 4448 43450 4476 46446
rect 4632 46170 4660 47398
rect 4908 46510 4936 47466
rect 4896 46504 4948 46510
rect 4896 46446 4948 46452
rect 4988 46368 5040 46374
rect 4988 46310 5040 46316
rect 4620 46164 4672 46170
rect 4620 46106 4672 46112
rect 4804 45960 4856 45966
rect 4804 45902 4856 45908
rect 4528 45824 4580 45830
rect 4528 45766 4580 45772
rect 4540 45082 4568 45766
rect 4620 45552 4672 45558
rect 4620 45494 4672 45500
rect 4528 45076 4580 45082
rect 4528 45018 4580 45024
rect 4632 43450 4660 45494
rect 4816 45490 4844 45902
rect 4804 45484 4856 45490
rect 4804 45426 4856 45432
rect 4712 45280 4764 45286
rect 4712 45222 4764 45228
rect 4436 43444 4488 43450
rect 4436 43386 4488 43392
rect 4620 43444 4672 43450
rect 4620 43386 4672 43392
rect 4632 43330 4660 43386
rect 4540 43302 4660 43330
rect 4436 43172 4488 43178
rect 4436 43114 4488 43120
rect 4448 42702 4476 43114
rect 4436 42696 4488 42702
rect 4436 42638 4488 42644
rect 4344 42220 4396 42226
rect 4344 42162 4396 42168
rect 4252 42152 4304 42158
rect 4448 42106 4476 42638
rect 4540 42158 4568 43302
rect 4620 43240 4672 43246
rect 4620 43182 4672 43188
rect 4304 42100 4476 42106
rect 4252 42094 4476 42100
rect 4528 42152 4580 42158
rect 4528 42094 4580 42100
rect 4264 42078 4476 42094
rect 4264 41818 4292 42078
rect 4252 41812 4304 41818
rect 4252 41754 4304 41760
rect 4632 41614 4660 43182
rect 4620 41608 4672 41614
rect 4620 41550 4672 41556
rect 4252 41472 4304 41478
rect 4252 41414 4304 41420
rect 4264 41070 4292 41414
rect 4252 41064 4304 41070
rect 4252 41006 4304 41012
rect 4344 40928 4396 40934
rect 4344 40870 4396 40876
rect 4252 40452 4304 40458
rect 4252 40394 4304 40400
rect 4160 40384 4212 40390
rect 4160 40326 4212 40332
rect 4172 39574 4200 40326
rect 4160 39568 4212 39574
rect 4160 39510 4212 39516
rect 4172 38486 4200 39510
rect 4160 38480 4212 38486
rect 4160 38422 4212 38428
rect 4160 38208 4212 38214
rect 4160 38150 4212 38156
rect 4172 37874 4200 38150
rect 4264 37890 4292 40394
rect 4356 39982 4384 40870
rect 4632 40458 4660 41550
rect 4620 40452 4672 40458
rect 4620 40394 4672 40400
rect 4344 39976 4396 39982
rect 4344 39918 4396 39924
rect 4356 38758 4384 39918
rect 4528 39908 4580 39914
rect 4528 39850 4580 39856
rect 4540 38894 4568 39850
rect 4528 38888 4580 38894
rect 4528 38830 4580 38836
rect 4344 38752 4396 38758
rect 4344 38694 4396 38700
rect 4540 38486 4568 38830
rect 4528 38480 4580 38486
rect 4528 38422 4580 38428
rect 4620 38412 4672 38418
rect 4620 38354 4672 38360
rect 4528 38208 4580 38214
rect 4528 38150 4580 38156
rect 4160 37868 4212 37874
rect 4264 37862 4384 37890
rect 4160 37810 4212 37816
rect 4172 36718 4200 37810
rect 4252 37800 4304 37806
rect 4252 37742 4304 37748
rect 4160 36712 4212 36718
rect 4160 36654 4212 36660
rect 4264 36378 4292 37742
rect 4252 36372 4304 36378
rect 4252 36314 4304 36320
rect 4356 36258 4384 37862
rect 4540 37330 4568 38150
rect 4528 37324 4580 37330
rect 4528 37266 4580 37272
rect 4436 37188 4488 37194
rect 4436 37130 4488 37136
rect 4264 36230 4384 36258
rect 4448 36242 4476 37130
rect 4632 36718 4660 38354
rect 4724 36768 4752 45222
rect 4816 44810 4844 45426
rect 5000 45422 5028 46310
rect 4988 45416 5040 45422
rect 4988 45358 5040 45364
rect 5080 44940 5132 44946
rect 5080 44882 5132 44888
rect 4804 44804 4856 44810
rect 4804 44746 4856 44752
rect 4988 44532 5040 44538
rect 4988 44474 5040 44480
rect 4804 44192 4856 44198
rect 4804 44134 4856 44140
rect 4816 43926 4844 44134
rect 4804 43920 4856 43926
rect 4804 43862 4856 43868
rect 4896 43240 4948 43246
rect 4896 43182 4948 43188
rect 4908 42838 4936 43182
rect 4896 42832 4948 42838
rect 4896 42774 4948 42780
rect 5000 42770 5028 44474
rect 4988 42764 5040 42770
rect 4988 42706 5040 42712
rect 4896 42628 4948 42634
rect 4896 42570 4948 42576
rect 4908 41546 4936 42570
rect 4988 42016 5040 42022
rect 4988 41958 5040 41964
rect 4896 41540 4948 41546
rect 4896 41482 4948 41488
rect 4908 40662 4936 41482
rect 4896 40656 4948 40662
rect 4896 40598 4948 40604
rect 5000 40594 5028 41958
rect 4988 40588 5040 40594
rect 4988 40530 5040 40536
rect 4896 40520 4948 40526
rect 4896 40462 4948 40468
rect 4804 38752 4856 38758
rect 4804 38694 4856 38700
rect 4816 37330 4844 38694
rect 4908 38457 4936 40462
rect 4988 40452 5040 40458
rect 4988 40394 5040 40400
rect 4894 38448 4950 38457
rect 4894 38383 4950 38392
rect 5000 37890 5028 40394
rect 5092 40066 5120 44882
rect 5184 40202 5212 47602
rect 5368 43840 5396 52974
rect 5814 52935 5816 52944
rect 5868 52935 5870 52944
rect 5816 52906 5868 52912
rect 5588 52252 5884 52272
rect 5644 52250 5668 52252
rect 5724 52250 5748 52252
rect 5804 52250 5828 52252
rect 5666 52198 5668 52250
rect 5730 52198 5742 52250
rect 5804 52198 5806 52250
rect 5644 52196 5668 52198
rect 5724 52196 5748 52198
rect 5804 52196 5828 52198
rect 5588 52176 5884 52196
rect 5920 51610 5948 53994
rect 6104 53242 6132 55200
rect 7852 53242 7880 55200
rect 9600 53242 9628 55200
rect 11440 53242 11468 55200
rect 13188 53242 13216 55200
rect 14936 54074 14964 55200
rect 14936 54046 15148 54074
rect 15120 53802 15148 54046
rect 15120 53774 15240 53802
rect 14852 53340 15148 53360
rect 14908 53338 14932 53340
rect 14988 53338 15012 53340
rect 15068 53338 15092 53340
rect 14930 53286 14932 53338
rect 14994 53286 15006 53338
rect 15068 53286 15070 53338
rect 14908 53284 14932 53286
rect 14988 53284 15012 53286
rect 15068 53284 15092 53286
rect 14852 53264 15148 53284
rect 6092 53236 6144 53242
rect 6092 53178 6144 53184
rect 7840 53236 7892 53242
rect 7840 53178 7892 53184
rect 9588 53236 9640 53242
rect 9588 53178 9640 53184
rect 11428 53236 11480 53242
rect 11428 53178 11480 53184
rect 13176 53236 13228 53242
rect 13176 53178 13228 53184
rect 15212 53174 15240 53774
rect 16684 53174 16712 55200
rect 18432 53242 18460 55200
rect 19156 53712 19208 53718
rect 19156 53654 19208 53660
rect 19168 53242 19196 53654
rect 20180 53242 20208 55200
rect 20258 54496 20314 54505
rect 20258 54431 20314 54440
rect 18420 53236 18472 53242
rect 18420 53178 18472 53184
rect 19156 53236 19208 53242
rect 19156 53178 19208 53184
rect 20168 53236 20220 53242
rect 20168 53178 20220 53184
rect 15200 53168 15252 53174
rect 15200 53110 15252 53116
rect 16672 53168 16724 53174
rect 16672 53110 16724 53116
rect 7012 52964 7064 52970
rect 7012 52906 7064 52912
rect 7840 52964 7892 52970
rect 7840 52906 7892 52912
rect 9956 52964 10008 52970
rect 9956 52906 10008 52912
rect 12072 52964 12124 52970
rect 12072 52906 12124 52912
rect 13268 52964 13320 52970
rect 13268 52906 13320 52912
rect 14372 52964 14424 52970
rect 14372 52906 14424 52912
rect 16488 52964 16540 52970
rect 16488 52906 16540 52912
rect 18512 52964 18564 52970
rect 18512 52906 18564 52912
rect 6552 52352 6604 52358
rect 6552 52294 6604 52300
rect 6000 51944 6052 51950
rect 6000 51886 6052 51892
rect 6368 51944 6420 51950
rect 6368 51886 6420 51892
rect 5908 51604 5960 51610
rect 5908 51546 5960 51552
rect 5908 51264 5960 51270
rect 5908 51206 5960 51212
rect 5588 51164 5884 51184
rect 5644 51162 5668 51164
rect 5724 51162 5748 51164
rect 5804 51162 5828 51164
rect 5666 51110 5668 51162
rect 5730 51110 5742 51162
rect 5804 51110 5806 51162
rect 5644 51108 5668 51110
rect 5724 51108 5748 51110
rect 5804 51108 5828 51110
rect 5588 51088 5884 51108
rect 5920 50998 5948 51206
rect 5908 50992 5960 50998
rect 5908 50934 5960 50940
rect 5816 50856 5868 50862
rect 5868 50816 5948 50844
rect 5816 50798 5868 50804
rect 5540 50788 5592 50794
rect 5540 50730 5592 50736
rect 5552 50386 5580 50730
rect 5540 50380 5592 50386
rect 5540 50322 5592 50328
rect 5588 50076 5884 50096
rect 5644 50074 5668 50076
rect 5724 50074 5748 50076
rect 5804 50074 5828 50076
rect 5666 50022 5668 50074
rect 5730 50022 5742 50074
rect 5804 50022 5806 50074
rect 5644 50020 5668 50022
rect 5724 50020 5748 50022
rect 5804 50020 5828 50022
rect 5588 50000 5884 50020
rect 5920 49434 5948 50816
rect 6012 50794 6040 51886
rect 6380 51474 6408 51886
rect 6564 51610 6592 52294
rect 6552 51604 6604 51610
rect 6552 51546 6604 51552
rect 6368 51468 6420 51474
rect 6368 51410 6420 51416
rect 6000 50788 6052 50794
rect 6000 50730 6052 50736
rect 6380 50386 6408 51410
rect 6828 50856 6880 50862
rect 6828 50798 6880 50804
rect 6460 50788 6512 50794
rect 6460 50730 6512 50736
rect 6092 50380 6144 50386
rect 6092 50322 6144 50328
rect 6368 50380 6420 50386
rect 6368 50322 6420 50328
rect 6000 49768 6052 49774
rect 6000 49710 6052 49716
rect 6012 49434 6040 49710
rect 5908 49428 5960 49434
rect 5908 49370 5960 49376
rect 6000 49428 6052 49434
rect 6000 49370 6052 49376
rect 6104 49230 6132 50322
rect 6184 49292 6236 49298
rect 6184 49234 6236 49240
rect 6092 49224 6144 49230
rect 6092 49166 6144 49172
rect 5588 48988 5884 49008
rect 5644 48986 5668 48988
rect 5724 48986 5748 48988
rect 5804 48986 5828 48988
rect 5666 48934 5668 48986
rect 5730 48934 5742 48986
rect 5804 48934 5806 48986
rect 5644 48932 5668 48934
rect 5724 48932 5748 48934
rect 5804 48932 5828 48934
rect 5588 48912 5884 48932
rect 5448 48884 5500 48890
rect 5448 48826 5500 48832
rect 5460 48754 5488 48826
rect 5448 48748 5500 48754
rect 5448 48690 5500 48696
rect 5460 48142 5488 48690
rect 5448 48136 5500 48142
rect 5448 48078 5500 48084
rect 5460 44402 5488 48078
rect 5908 48068 5960 48074
rect 5908 48010 5960 48016
rect 5588 47900 5884 47920
rect 5644 47898 5668 47900
rect 5724 47898 5748 47900
rect 5804 47898 5828 47900
rect 5666 47846 5668 47898
rect 5730 47846 5742 47898
rect 5804 47846 5806 47898
rect 5644 47844 5668 47846
rect 5724 47844 5748 47846
rect 5804 47844 5828 47846
rect 5588 47824 5884 47844
rect 5920 47784 5948 48010
rect 5828 47756 5948 47784
rect 5828 47598 5856 47756
rect 5816 47592 5868 47598
rect 5816 47534 5868 47540
rect 5724 47524 5776 47530
rect 5724 47466 5776 47472
rect 5736 47122 5764 47466
rect 5724 47116 5776 47122
rect 5724 47058 5776 47064
rect 5828 47036 5856 47534
rect 6196 47410 6224 49234
rect 6276 48816 6328 48822
rect 6276 48758 6328 48764
rect 6288 47530 6316 48758
rect 6472 47598 6500 50730
rect 6644 49224 6696 49230
rect 6644 49166 6696 49172
rect 6552 48612 6604 48618
rect 6552 48554 6604 48560
rect 6460 47592 6512 47598
rect 6460 47534 6512 47540
rect 6276 47524 6328 47530
rect 6276 47466 6328 47472
rect 6196 47382 6316 47410
rect 5908 47048 5960 47054
rect 5828 47008 5908 47036
rect 5908 46990 5960 46996
rect 5588 46812 5884 46832
rect 5644 46810 5668 46812
rect 5724 46810 5748 46812
rect 5804 46810 5828 46812
rect 5666 46758 5668 46810
rect 5730 46758 5742 46810
rect 5804 46758 5806 46810
rect 5644 46756 5668 46758
rect 5724 46756 5748 46758
rect 5804 46756 5828 46758
rect 5588 46736 5884 46756
rect 5920 46510 5948 46990
rect 6288 46510 6316 47382
rect 6564 46714 6592 48554
rect 6656 47598 6684 49166
rect 6840 48600 6868 50798
rect 6920 48612 6972 48618
rect 6840 48572 6920 48600
rect 6920 48554 6972 48560
rect 6736 48544 6788 48550
rect 6736 48486 6788 48492
rect 6748 48074 6776 48486
rect 6736 48068 6788 48074
rect 6736 48010 6788 48016
rect 6644 47592 6696 47598
rect 6644 47534 6696 47540
rect 6828 47592 6880 47598
rect 6828 47534 6880 47540
rect 6552 46708 6604 46714
rect 6552 46650 6604 46656
rect 6656 46594 6684 47534
rect 6840 47054 6868 47534
rect 6828 47048 6880 47054
rect 6828 46990 6880 46996
rect 6564 46566 6684 46594
rect 5908 46504 5960 46510
rect 5908 46446 5960 46452
rect 6276 46504 6328 46510
rect 6276 46446 6328 46452
rect 5588 45724 5884 45744
rect 5644 45722 5668 45724
rect 5724 45722 5748 45724
rect 5804 45722 5828 45724
rect 5666 45670 5668 45722
rect 5730 45670 5742 45722
rect 5804 45670 5806 45722
rect 5644 45668 5668 45670
rect 5724 45668 5748 45670
rect 5804 45668 5828 45670
rect 5588 45648 5884 45668
rect 5920 45540 5948 46446
rect 6288 46374 6316 46446
rect 6276 46368 6328 46374
rect 6276 46310 6328 46316
rect 6092 46164 6144 46170
rect 6092 46106 6144 46112
rect 5828 45512 5948 45540
rect 5724 44940 5776 44946
rect 5724 44882 5776 44888
rect 5736 44724 5764 44882
rect 5828 44826 5856 45512
rect 6000 45280 6052 45286
rect 6000 45222 6052 45228
rect 6012 44946 6040 45222
rect 6000 44940 6052 44946
rect 6000 44882 6052 44888
rect 5828 44798 6040 44826
rect 5736 44696 5948 44724
rect 5588 44636 5884 44656
rect 5644 44634 5668 44636
rect 5724 44634 5748 44636
rect 5804 44634 5828 44636
rect 5666 44582 5668 44634
rect 5730 44582 5742 44634
rect 5804 44582 5806 44634
rect 5644 44580 5668 44582
rect 5724 44580 5748 44582
rect 5804 44580 5828 44582
rect 5588 44560 5884 44580
rect 5448 44396 5500 44402
rect 5448 44338 5500 44344
rect 5276 43812 5396 43840
rect 5276 40526 5304 43812
rect 5460 42634 5488 44338
rect 5920 44266 5948 44696
rect 5908 44260 5960 44266
rect 5908 44202 5960 44208
rect 5920 43994 5948 44202
rect 5908 43988 5960 43994
rect 5908 43930 5960 43936
rect 5588 43548 5884 43568
rect 5644 43546 5668 43548
rect 5724 43546 5748 43548
rect 5804 43546 5828 43548
rect 5666 43494 5668 43546
rect 5730 43494 5742 43546
rect 5804 43494 5806 43546
rect 5644 43492 5668 43494
rect 5724 43492 5748 43494
rect 5804 43492 5828 43494
rect 5588 43472 5884 43492
rect 5448 42628 5500 42634
rect 5448 42570 5500 42576
rect 5588 42460 5884 42480
rect 5644 42458 5668 42460
rect 5724 42458 5748 42460
rect 5804 42458 5828 42460
rect 5666 42406 5668 42458
rect 5730 42406 5742 42458
rect 5804 42406 5806 42458
rect 5644 42404 5668 42406
rect 5724 42404 5748 42406
rect 5804 42404 5828 42406
rect 5588 42384 5884 42404
rect 5356 41812 5408 41818
rect 5356 41754 5408 41760
rect 5368 40594 5396 41754
rect 5908 41472 5960 41478
rect 5908 41414 5960 41420
rect 5588 41372 5884 41392
rect 5644 41370 5668 41372
rect 5724 41370 5748 41372
rect 5804 41370 5828 41372
rect 5666 41318 5668 41370
rect 5730 41318 5742 41370
rect 5804 41318 5806 41370
rect 5644 41316 5668 41318
rect 5724 41316 5748 41318
rect 5804 41316 5828 41318
rect 5588 41296 5884 41316
rect 5538 41168 5594 41177
rect 5538 41103 5594 41112
rect 5552 41070 5580 41103
rect 5540 41064 5592 41070
rect 5540 41006 5592 41012
rect 5356 40588 5408 40594
rect 5356 40530 5408 40536
rect 5264 40520 5316 40526
rect 5264 40462 5316 40468
rect 5184 40174 5304 40202
rect 5092 40038 5212 40066
rect 5080 39976 5132 39982
rect 5080 39918 5132 39924
rect 5092 38486 5120 39918
rect 5080 38480 5132 38486
rect 5080 38422 5132 38428
rect 5000 37862 5120 37890
rect 4804 37324 4856 37330
rect 4804 37266 4856 37272
rect 4896 37256 4948 37262
rect 4896 37198 4948 37204
rect 4724 36740 4844 36768
rect 4620 36712 4672 36718
rect 4620 36654 4672 36660
rect 4436 36236 4488 36242
rect 4160 33856 4212 33862
rect 4160 33798 4212 33804
rect 4172 32881 4200 33798
rect 4264 33046 4292 36230
rect 4436 36178 4488 36184
rect 4344 36168 4396 36174
rect 4344 36110 4396 36116
rect 4356 35494 4384 36110
rect 4344 35488 4396 35494
rect 4344 35430 4396 35436
rect 4252 33040 4304 33046
rect 4252 32982 4304 32988
rect 4252 32904 4304 32910
rect 4158 32872 4214 32881
rect 4252 32846 4304 32852
rect 4158 32807 4214 32816
rect 3988 31726 4108 31754
rect 3790 31240 3846 31249
rect 3790 31175 3846 31184
rect 3804 30938 3832 31175
rect 3792 30932 3844 30938
rect 3792 30874 3844 30880
rect 3884 30592 3936 30598
rect 3884 30534 3936 30540
rect 3790 28384 3846 28393
rect 3790 28319 3846 28328
rect 3804 28082 3832 28319
rect 3792 28076 3844 28082
rect 3792 28018 3844 28024
rect 3896 27962 3924 30534
rect 3988 30054 4016 31726
rect 4066 31648 4122 31657
rect 4066 31583 4122 31592
rect 4080 30734 4108 31583
rect 4264 31482 4292 32846
rect 4356 31754 4384 35430
rect 4448 34474 4476 36178
rect 4528 35148 4580 35154
rect 4528 35090 4580 35096
rect 4540 34649 4568 35090
rect 4526 34640 4582 34649
rect 4526 34575 4582 34584
rect 4528 34536 4580 34542
rect 4528 34478 4580 34484
rect 4436 34468 4488 34474
rect 4436 34410 4488 34416
rect 4436 34060 4488 34066
rect 4540 34048 4568 34478
rect 4488 34020 4568 34048
rect 4436 34002 4488 34008
rect 4436 33040 4488 33046
rect 4436 32982 4488 32988
rect 4448 32434 4476 32982
rect 4436 32428 4488 32434
rect 4436 32370 4488 32376
rect 4356 31726 4476 31754
rect 4252 31476 4304 31482
rect 4252 31418 4304 31424
rect 4160 31272 4212 31278
rect 4160 31214 4212 31220
rect 4068 30728 4120 30734
rect 4068 30670 4120 30676
rect 4068 30116 4120 30122
rect 4068 30058 4120 30064
rect 3976 30048 4028 30054
rect 3976 29990 4028 29996
rect 3976 28960 4028 28966
rect 3974 28928 3976 28937
rect 4028 28928 4030 28937
rect 3974 28863 4030 28872
rect 3804 27934 3924 27962
rect 3700 24608 3752 24614
rect 3700 24550 3752 24556
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 3712 21146 3740 21830
rect 3700 21140 3752 21146
rect 3700 21082 3752 21088
rect 3804 20466 3832 27934
rect 3884 27464 3936 27470
rect 3884 27406 3936 27412
rect 3896 22094 3924 27406
rect 3988 26790 4016 28863
rect 4080 28490 4108 30058
rect 4068 28484 4120 28490
rect 4068 28426 4120 28432
rect 4172 27418 4200 31214
rect 4344 30184 4396 30190
rect 4344 30126 4396 30132
rect 4356 29102 4384 30126
rect 4344 29096 4396 29102
rect 4344 29038 4396 29044
rect 4252 29028 4304 29034
rect 4252 28970 4304 28976
rect 4264 28014 4292 28970
rect 4356 28762 4384 29038
rect 4344 28756 4396 28762
rect 4344 28698 4396 28704
rect 4252 28008 4304 28014
rect 4252 27950 4304 27956
rect 4344 27872 4396 27878
rect 4344 27814 4396 27820
rect 4356 27606 4384 27814
rect 4344 27600 4396 27606
rect 4344 27542 4396 27548
rect 4172 27390 4292 27418
rect 4160 27328 4212 27334
rect 4160 27270 4212 27276
rect 4172 27130 4200 27270
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 3976 26784 4028 26790
rect 3976 26726 4028 26732
rect 4160 26444 4212 26450
rect 4160 26386 4212 26392
rect 4066 25120 4122 25129
rect 4172 25106 4200 26386
rect 4264 25838 4292 27390
rect 4252 25832 4304 25838
rect 4252 25774 4304 25780
rect 4264 25362 4292 25774
rect 4252 25356 4304 25362
rect 4304 25316 4384 25344
rect 4252 25298 4304 25304
rect 4122 25078 4200 25106
rect 4066 25055 4122 25064
rect 4252 24064 4304 24070
rect 4252 24006 4304 24012
rect 4264 23322 4292 24006
rect 4252 23316 4304 23322
rect 4252 23258 4304 23264
rect 4160 23180 4212 23186
rect 4160 23122 4212 23128
rect 4068 22704 4120 22710
rect 4068 22646 4120 22652
rect 4080 22166 4108 22646
rect 4068 22160 4120 22166
rect 4068 22102 4120 22108
rect 3896 22066 4016 22094
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 3792 20460 3844 20466
rect 3792 20402 3844 20408
rect 3896 19854 3924 20878
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3896 17678 3924 19790
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3988 17134 4016 22066
rect 4172 21434 4200 23122
rect 4264 22574 4292 23258
rect 4356 23118 4384 25316
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 4252 22568 4304 22574
rect 4252 22510 4304 22516
rect 4344 22432 4396 22438
rect 4250 22400 4306 22409
rect 4344 22374 4396 22380
rect 4250 22335 4306 22344
rect 4264 21554 4292 22335
rect 4252 21548 4304 21554
rect 4252 21490 4304 21496
rect 4172 21406 4292 21434
rect 4160 21344 4212 21350
rect 4160 21286 4212 21292
rect 4172 20058 4200 21286
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4160 19712 4212 19718
rect 4160 19654 4212 19660
rect 4172 19378 4200 19654
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 4264 19310 4292 21406
rect 4356 20058 4384 22374
rect 4344 20052 4396 20058
rect 4344 19994 4396 20000
rect 4252 19304 4304 19310
rect 4304 19252 4384 19258
rect 4252 19246 4384 19252
rect 4264 19230 4384 19246
rect 4068 19168 4120 19174
rect 4252 19168 4304 19174
rect 4120 19128 4200 19156
rect 4068 19110 4120 19116
rect 4172 18222 4200 19128
rect 4252 19110 4304 19116
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3712 14958 3740 15846
rect 3884 15632 3936 15638
rect 3884 15574 3936 15580
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3712 14482 3740 14894
rect 3896 14618 3924 15574
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3792 14544 3844 14550
rect 3792 14486 3844 14492
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 3804 13394 3832 14486
rect 3896 13530 3924 14554
rect 3988 14482 4016 15506
rect 4172 15450 4200 17682
rect 4264 16182 4292 19110
rect 4356 17814 4384 19230
rect 4344 17808 4396 17814
rect 4344 17750 4396 17756
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 4264 15570 4292 16118
rect 4448 15638 4476 31726
rect 4540 31278 4568 34020
rect 4632 32570 4660 36654
rect 4712 36644 4764 36650
rect 4712 36586 4764 36592
rect 4724 34542 4752 36586
rect 4712 34536 4764 34542
rect 4712 34478 4764 34484
rect 4620 32564 4672 32570
rect 4620 32506 4672 32512
rect 4620 32428 4672 32434
rect 4620 32370 4672 32376
rect 4528 31272 4580 31278
rect 4528 31214 4580 31220
rect 4528 29504 4580 29510
rect 4528 29446 4580 29452
rect 4540 28694 4568 29446
rect 4528 28688 4580 28694
rect 4528 28630 4580 28636
rect 4528 28484 4580 28490
rect 4528 28426 4580 28432
rect 4540 25158 4568 28426
rect 4632 26586 4660 32370
rect 4724 30122 4752 34478
rect 4816 33590 4844 36740
rect 4908 34406 4936 37198
rect 4988 35148 5040 35154
rect 4988 35090 5040 35096
rect 5000 34746 5028 35090
rect 4988 34740 5040 34746
rect 4988 34682 5040 34688
rect 4988 34468 5040 34474
rect 4988 34410 5040 34416
rect 4896 34400 4948 34406
rect 4896 34342 4948 34348
rect 4908 34202 4936 34342
rect 5000 34202 5028 34410
rect 4896 34196 4948 34202
rect 4896 34138 4948 34144
rect 4988 34196 5040 34202
rect 4988 34138 5040 34144
rect 4804 33584 4856 33590
rect 4804 33526 4856 33532
rect 4988 32972 5040 32978
rect 4988 32914 5040 32920
rect 4896 32224 4948 32230
rect 4896 32166 4948 32172
rect 4908 32026 4936 32166
rect 4896 32020 4948 32026
rect 4896 31962 4948 31968
rect 5000 31686 5028 32914
rect 4988 31680 5040 31686
rect 4988 31622 5040 31628
rect 5000 31414 5028 31622
rect 4988 31408 5040 31414
rect 4988 31350 5040 31356
rect 5000 30394 5028 31350
rect 4988 30388 5040 30394
rect 4988 30330 5040 30336
rect 4804 30184 4856 30190
rect 4804 30126 4856 30132
rect 4896 30184 4948 30190
rect 4896 30126 4948 30132
rect 4712 30116 4764 30122
rect 4712 30058 4764 30064
rect 4712 29028 4764 29034
rect 4712 28970 4764 28976
rect 4620 26580 4672 26586
rect 4620 26522 4672 26528
rect 4620 26376 4672 26382
rect 4620 26318 4672 26324
rect 4528 25152 4580 25158
rect 4528 25094 4580 25100
rect 4540 23798 4568 25094
rect 4528 23792 4580 23798
rect 4528 23734 4580 23740
rect 4528 23656 4580 23662
rect 4528 23598 4580 23604
rect 4540 21865 4568 23598
rect 4526 21856 4582 21865
rect 4526 21791 4582 21800
rect 4632 20602 4660 26318
rect 4724 23322 4752 28970
rect 4816 28762 4844 30126
rect 4908 29238 4936 30126
rect 4988 29640 5040 29646
rect 4988 29582 5040 29588
rect 4896 29232 4948 29238
rect 4896 29174 4948 29180
rect 5000 29170 5028 29582
rect 4988 29164 5040 29170
rect 4988 29106 5040 29112
rect 5000 28994 5028 29106
rect 4908 28966 5028 28994
rect 4804 28756 4856 28762
rect 4804 28698 4856 28704
rect 4908 28370 4936 28966
rect 4988 28620 5040 28626
rect 4988 28562 5040 28568
rect 4816 28342 4936 28370
rect 4816 26738 4844 28342
rect 4896 28212 4948 28218
rect 4896 28154 4948 28160
rect 4908 26858 4936 28154
rect 4896 26852 4948 26858
rect 4896 26794 4948 26800
rect 4816 26710 4936 26738
rect 4908 26382 4936 26710
rect 4896 26376 4948 26382
rect 4896 26318 4948 26324
rect 4804 25696 4856 25702
rect 4804 25638 4856 25644
rect 4816 25498 4844 25638
rect 4804 25492 4856 25498
rect 4804 25434 4856 25440
rect 4908 25378 4936 26318
rect 4816 25350 4936 25378
rect 4816 24206 4844 25350
rect 4896 24744 4948 24750
rect 4896 24686 4948 24692
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4908 24138 4936 24686
rect 4896 24132 4948 24138
rect 4896 24074 4948 24080
rect 4896 23792 4948 23798
rect 4896 23734 4948 23740
rect 4804 23520 4856 23526
rect 4804 23462 4856 23468
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 4712 22160 4764 22166
rect 4816 22114 4844 23462
rect 4764 22108 4844 22114
rect 4712 22102 4844 22108
rect 4724 22086 4844 22102
rect 4816 21418 4844 22086
rect 4804 21412 4856 21418
rect 4804 21354 4856 21360
rect 4804 20868 4856 20874
rect 4804 20810 4856 20816
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 4712 19984 4764 19990
rect 4712 19926 4764 19932
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4540 18902 4568 19110
rect 4528 18896 4580 18902
rect 4528 18838 4580 18844
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4632 15638 4660 16730
rect 4436 15632 4488 15638
rect 4436 15574 4488 15580
rect 4620 15632 4672 15638
rect 4620 15574 4672 15580
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4436 15496 4488 15502
rect 4172 15422 4292 15450
rect 4436 15438 4488 15444
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4066 14920 4122 14929
rect 4172 14906 4200 15302
rect 4122 14878 4200 14906
rect 4066 14855 4122 14864
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3608 12164 3660 12170
rect 3608 12106 3660 12112
rect 2778 11183 2780 11192
rect 2832 11183 2834 11192
rect 3240 11212 3292 11218
rect 2780 11154 2832 11160
rect 3240 11154 3292 11160
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2884 10606 2912 10678
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2516 8078 2636 8106
rect 2700 8090 2728 9318
rect 2688 8084 2740 8090
rect 2410 7984 2466 7993
rect 2410 7919 2412 7928
rect 2464 7919 2466 7928
rect 2412 7890 2464 7896
rect 2516 6866 2544 8078
rect 2688 8026 2740 8032
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1780 5370 1808 6054
rect 2240 5846 2268 6734
rect 2228 5840 2280 5846
rect 2228 5782 2280 5788
rect 2516 5642 2544 6802
rect 2504 5636 2556 5642
rect 2504 5578 2556 5584
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2700 5370 2728 5510
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2792 5166 2820 10202
rect 2884 9722 2912 10542
rect 2976 10130 3004 10746
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 3068 9518 3096 11018
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2870 9208 2926 9217
rect 2870 9143 2926 9152
rect 2884 7954 2912 9143
rect 2976 8090 3004 9386
rect 3160 9178 3188 11086
rect 3252 10130 3280 11154
rect 3528 10130 3556 11154
rect 3712 10266 3740 12242
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 3068 8634 3096 8978
rect 3252 8974 3280 10066
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 9178 3464 9318
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3424 9036 3476 9042
rect 3528 9024 3556 10066
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3712 9042 3740 9386
rect 3476 8996 3556 9024
rect 3700 9036 3752 9042
rect 3424 8978 3476 8984
rect 3700 8978 3752 8984
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3238 8800 3294 8809
rect 3238 8735 3294 8744
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 3252 8430 3280 8735
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3068 7177 3096 7278
rect 3054 7168 3110 7177
rect 3054 7103 3110 7112
rect 3804 6866 3832 12038
rect 3988 11626 4016 12582
rect 3976 11620 4028 11626
rect 3976 11562 4028 11568
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3988 10810 4016 11154
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 4080 9058 4108 14758
rect 4264 14362 4292 15422
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4172 14334 4292 14362
rect 4172 13530 4200 14334
rect 4356 13802 4384 15302
rect 4448 14822 4476 15438
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 4448 14482 4476 14554
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4632 14328 4660 15438
rect 4448 14300 4660 14328
rect 4344 13796 4396 13802
rect 4344 13738 4396 13744
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4172 12986 4200 13466
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 3896 9030 4108 9058
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3252 5166 3280 6802
rect 3896 6746 3924 9030
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 4080 8090 4108 8502
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3620 6718 3924 6746
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3344 5370 3372 5646
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 1688 3738 1716 3946
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1964 3505 1992 5102
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2596 3936 2648 3942
rect 2792 3913 2820 4626
rect 2872 3936 2924 3942
rect 2596 3878 2648 3884
rect 2778 3904 2834 3913
rect 2608 3670 2636 3878
rect 2872 3878 2924 3884
rect 2778 3839 2834 3848
rect 2596 3664 2648 3670
rect 2596 3606 2648 3612
rect 1950 3496 2006 3505
rect 1950 3431 2006 3440
rect 2884 3194 2912 3878
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 1674 3088 1730 3097
rect 2976 3058 3004 5102
rect 3252 4842 3280 5102
rect 3160 4814 3280 4842
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3068 4078 3096 4422
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 1674 3023 1730 3032
rect 2964 3052 3016 3058
rect 1688 2990 1716 3023
rect 2964 2994 3016 3000
rect 3160 2990 3188 4814
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 1964 800 1992 2382
rect 2608 2106 2636 2450
rect 2596 2100 2648 2106
rect 2596 2042 2648 2048
rect 2780 1964 2832 1970
rect 2780 1906 2832 1912
rect 2792 1465 2820 1906
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 2964 1080 3016 1086
rect 3252 1057 3280 4626
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 2964 1022 3016 1028
rect 3238 1048 3294 1057
rect 1398 232 1454 241
rect 1398 167 1454 176
rect 1950 -800 2006 800
rect 2976 649 3004 1022
rect 3238 983 3294 992
rect 3344 800 3372 2382
rect 3436 2281 3464 6258
rect 3620 5778 3648 6718
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3698 5944 3754 5953
rect 3698 5879 3700 5888
rect 3752 5879 3754 5888
rect 3700 5850 3752 5856
rect 3804 5846 3832 6598
rect 3896 6254 3924 6598
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3792 5568 3844 5574
rect 3988 5545 4016 6802
rect 4080 6361 4108 6802
rect 4172 6458 4200 12718
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4264 8022 4292 9998
rect 4356 9110 4384 10610
rect 4448 9178 4476 14300
rect 4724 14074 4752 19926
rect 4816 19378 4844 20810
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4816 18290 4844 19314
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4816 17882 4844 18022
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4816 14618 4844 14758
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4528 12368 4580 12374
rect 4528 12310 4580 12316
rect 4540 11558 4568 12310
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4066 6352 4122 6361
rect 4066 6287 4122 6296
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 3792 5510 3844 5516
rect 3974 5536 4030 5545
rect 3804 4826 3832 5510
rect 3974 5471 4030 5480
rect 4066 5128 4122 5137
rect 4172 5114 4200 6190
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4122 5086 4200 5114
rect 4066 5063 4122 5072
rect 3792 4820 3844 4826
rect 4264 4808 4292 5714
rect 3792 4762 3844 4768
rect 3988 4780 4292 4808
rect 3516 4548 3568 4554
rect 3516 4490 3568 4496
rect 3528 2990 3556 4490
rect 3988 4321 4016 4780
rect 4066 4720 4122 4729
rect 4356 4706 4384 5714
rect 4122 4678 4384 4706
rect 4448 4690 4476 9114
rect 4540 8430 4568 9318
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4528 6996 4580 7002
rect 4528 6938 4580 6944
rect 4436 4684 4488 4690
rect 4066 4655 4122 4664
rect 4436 4626 4488 4632
rect 4448 4570 4476 4626
rect 4264 4542 4476 4570
rect 3974 4312 4030 4321
rect 3974 4247 4030 4256
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4172 4078 4200 4218
rect 4264 4214 4292 4542
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4356 4078 4384 4422
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4172 3738 4200 3878
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4448 3602 4476 4422
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3514 2680 3570 2689
rect 4540 2650 4568 6938
rect 4632 5098 4660 13942
rect 4724 10606 4752 14010
rect 4816 12442 4844 14282
rect 4908 13870 4936 23734
rect 5000 21690 5028 28562
rect 5092 27402 5120 37862
rect 5184 36258 5212 40038
rect 5276 39488 5304 40174
rect 5368 39930 5396 40530
rect 5448 40384 5500 40390
rect 5448 40326 5500 40332
rect 5460 40050 5488 40326
rect 5588 40284 5884 40304
rect 5644 40282 5668 40284
rect 5724 40282 5748 40284
rect 5804 40282 5828 40284
rect 5666 40230 5668 40282
rect 5730 40230 5742 40282
rect 5804 40230 5806 40282
rect 5644 40228 5668 40230
rect 5724 40228 5748 40230
rect 5804 40228 5828 40230
rect 5588 40208 5884 40228
rect 5448 40044 5500 40050
rect 5448 39986 5500 39992
rect 5368 39902 5488 39930
rect 5276 39460 5396 39488
rect 5264 39364 5316 39370
rect 5264 39306 5316 39312
rect 5276 38894 5304 39306
rect 5264 38888 5316 38894
rect 5264 38830 5316 38836
rect 5368 38214 5396 39460
rect 5356 38208 5408 38214
rect 5356 38150 5408 38156
rect 5356 37732 5408 37738
rect 5356 37674 5408 37680
rect 5368 37398 5396 37674
rect 5356 37392 5408 37398
rect 5356 37334 5408 37340
rect 5264 37324 5316 37330
rect 5264 37266 5316 37272
rect 5276 36378 5304 37266
rect 5264 36372 5316 36378
rect 5264 36314 5316 36320
rect 5184 36230 5396 36258
rect 5264 34400 5316 34406
rect 5264 34342 5316 34348
rect 5276 34066 5304 34342
rect 5172 34060 5224 34066
rect 5172 34002 5224 34008
rect 5264 34060 5316 34066
rect 5264 34002 5316 34008
rect 5184 33454 5212 34002
rect 5264 33584 5316 33590
rect 5264 33526 5316 33532
rect 5172 33448 5224 33454
rect 5172 33390 5224 33396
rect 5172 33312 5224 33318
rect 5172 33254 5224 33260
rect 5184 28558 5212 33254
rect 5276 32026 5304 33526
rect 5264 32020 5316 32026
rect 5264 31962 5316 31968
rect 5264 30388 5316 30394
rect 5264 30330 5316 30336
rect 5276 28994 5304 30330
rect 5368 29102 5396 36230
rect 5460 33318 5488 39902
rect 5588 39196 5884 39216
rect 5644 39194 5668 39196
rect 5724 39194 5748 39196
rect 5804 39194 5828 39196
rect 5666 39142 5668 39194
rect 5730 39142 5742 39194
rect 5804 39142 5806 39194
rect 5644 39140 5668 39142
rect 5724 39140 5748 39142
rect 5804 39140 5828 39142
rect 5588 39120 5884 39140
rect 5920 38418 5948 41414
rect 5908 38412 5960 38418
rect 5908 38354 5960 38360
rect 5588 38108 5884 38128
rect 5644 38106 5668 38108
rect 5724 38106 5748 38108
rect 5804 38106 5828 38108
rect 5666 38054 5668 38106
rect 5730 38054 5742 38106
rect 5804 38054 5806 38106
rect 5644 38052 5668 38054
rect 5724 38052 5748 38054
rect 5804 38052 5828 38054
rect 5588 38032 5884 38052
rect 5908 37800 5960 37806
rect 5908 37742 5960 37748
rect 5588 37020 5884 37040
rect 5644 37018 5668 37020
rect 5724 37018 5748 37020
rect 5804 37018 5828 37020
rect 5666 36966 5668 37018
rect 5730 36966 5742 37018
rect 5804 36966 5806 37018
rect 5644 36964 5668 36966
rect 5724 36964 5748 36966
rect 5804 36964 5828 36966
rect 5588 36944 5884 36964
rect 5920 36718 5948 37742
rect 5908 36712 5960 36718
rect 5908 36654 5960 36660
rect 5588 35932 5884 35952
rect 5644 35930 5668 35932
rect 5724 35930 5748 35932
rect 5804 35930 5828 35932
rect 5666 35878 5668 35930
rect 5730 35878 5742 35930
rect 5804 35878 5806 35930
rect 5644 35876 5668 35878
rect 5724 35876 5748 35878
rect 5804 35876 5828 35878
rect 5588 35856 5884 35876
rect 5908 34944 5960 34950
rect 5908 34886 5960 34892
rect 5588 34844 5884 34864
rect 5644 34842 5668 34844
rect 5724 34842 5748 34844
rect 5804 34842 5828 34844
rect 5666 34790 5668 34842
rect 5730 34790 5742 34842
rect 5804 34790 5806 34842
rect 5644 34788 5668 34790
rect 5724 34788 5748 34790
rect 5804 34788 5828 34790
rect 5588 34768 5884 34788
rect 5538 34640 5594 34649
rect 5538 34575 5540 34584
rect 5592 34575 5594 34584
rect 5540 34546 5592 34552
rect 5588 33756 5884 33776
rect 5644 33754 5668 33756
rect 5724 33754 5748 33756
rect 5804 33754 5828 33756
rect 5666 33702 5668 33754
rect 5730 33702 5742 33754
rect 5804 33702 5806 33754
rect 5644 33700 5668 33702
rect 5724 33700 5748 33702
rect 5804 33700 5828 33702
rect 5588 33680 5884 33700
rect 5920 33454 5948 34886
rect 5908 33448 5960 33454
rect 5908 33390 5960 33396
rect 5448 33312 5500 33318
rect 5448 33254 5500 33260
rect 5588 32668 5884 32688
rect 5644 32666 5668 32668
rect 5724 32666 5748 32668
rect 5804 32666 5828 32668
rect 5666 32614 5668 32666
rect 5730 32614 5742 32666
rect 5804 32614 5806 32666
rect 5644 32612 5668 32614
rect 5724 32612 5748 32614
rect 5804 32612 5828 32614
rect 5588 32592 5884 32612
rect 5632 32428 5684 32434
rect 5632 32370 5684 32376
rect 5540 32292 5592 32298
rect 5540 32234 5592 32240
rect 5552 32026 5580 32234
rect 5540 32020 5592 32026
rect 5540 31962 5592 31968
rect 5644 31822 5672 32370
rect 5448 31816 5500 31822
rect 5448 31758 5500 31764
rect 5632 31816 5684 31822
rect 5632 31758 5684 31764
rect 5460 29889 5488 31758
rect 5588 31580 5884 31600
rect 5644 31578 5668 31580
rect 5724 31578 5748 31580
rect 5804 31578 5828 31580
rect 5666 31526 5668 31578
rect 5730 31526 5742 31578
rect 5804 31526 5806 31578
rect 5644 31524 5668 31526
rect 5724 31524 5748 31526
rect 5804 31524 5828 31526
rect 5588 31504 5884 31524
rect 5908 31272 5960 31278
rect 5908 31214 5960 31220
rect 5588 30492 5884 30512
rect 5644 30490 5668 30492
rect 5724 30490 5748 30492
rect 5804 30490 5828 30492
rect 5666 30438 5668 30490
rect 5730 30438 5742 30490
rect 5804 30438 5806 30490
rect 5644 30436 5668 30438
rect 5724 30436 5748 30438
rect 5804 30436 5828 30438
rect 5588 30416 5884 30436
rect 5920 30274 5948 31214
rect 5552 30246 5948 30274
rect 5446 29880 5502 29889
rect 5446 29815 5502 29824
rect 5448 29708 5500 29714
rect 5448 29650 5500 29656
rect 5460 29170 5488 29650
rect 5552 29578 5580 30246
rect 5908 30184 5960 30190
rect 6012 30172 6040 44798
rect 6104 36378 6132 46106
rect 6184 45280 6236 45286
rect 6184 45222 6236 45228
rect 6196 43450 6224 45222
rect 6184 43444 6236 43450
rect 6184 43386 6236 43392
rect 6288 43330 6316 46310
rect 6460 45280 6512 45286
rect 6460 45222 6512 45228
rect 6368 44872 6420 44878
rect 6368 44814 6420 44820
rect 6380 44198 6408 44814
rect 6472 44538 6500 45222
rect 6460 44532 6512 44538
rect 6460 44474 6512 44480
rect 6564 44418 6592 46566
rect 6932 45490 6960 48554
rect 6920 45484 6972 45490
rect 6920 45426 6972 45432
rect 6828 44940 6880 44946
rect 6828 44882 6880 44888
rect 6644 44804 6696 44810
rect 6644 44746 6696 44752
rect 6472 44390 6592 44418
rect 6368 44192 6420 44198
rect 6368 44134 6420 44140
rect 6380 43790 6408 44134
rect 6368 43784 6420 43790
rect 6368 43726 6420 43732
rect 6196 43302 6316 43330
rect 6196 43246 6224 43302
rect 6184 43240 6236 43246
rect 6184 43182 6236 43188
rect 6276 43172 6328 43178
rect 6380 43160 6408 43726
rect 6328 43132 6408 43160
rect 6276 43114 6328 43120
rect 6184 41608 6236 41614
rect 6184 41550 6236 41556
rect 6196 40594 6224 41550
rect 6184 40588 6236 40594
rect 6184 40530 6236 40536
rect 6196 39098 6224 40530
rect 6184 39092 6236 39098
rect 6184 39034 6236 39040
rect 6182 38448 6238 38457
rect 6182 38383 6238 38392
rect 6196 38214 6224 38383
rect 6184 38208 6236 38214
rect 6184 38150 6236 38156
rect 6092 36372 6144 36378
rect 6092 36314 6144 36320
rect 6104 32484 6132 36314
rect 6288 32502 6316 43114
rect 6368 39976 6420 39982
rect 6368 39918 6420 39924
rect 6380 39438 6408 39918
rect 6368 39432 6420 39438
rect 6368 39374 6420 39380
rect 6368 36712 6420 36718
rect 6368 36654 6420 36660
rect 6380 36174 6408 36654
rect 6368 36168 6420 36174
rect 6368 36110 6420 36116
rect 6380 34610 6408 36110
rect 6368 34604 6420 34610
rect 6368 34546 6420 34552
rect 6380 33930 6408 34546
rect 6368 33924 6420 33930
rect 6368 33866 6420 33872
rect 6276 32496 6328 32502
rect 6104 32456 6224 32484
rect 6196 32366 6224 32456
rect 6276 32438 6328 32444
rect 6092 32360 6144 32366
rect 6092 32302 6144 32308
rect 6184 32360 6236 32366
rect 6368 32360 6420 32366
rect 6184 32302 6236 32308
rect 6288 32320 6368 32348
rect 6104 30326 6132 32302
rect 6288 32026 6316 32320
rect 6368 32302 6420 32308
rect 6368 32224 6420 32230
rect 6368 32166 6420 32172
rect 6276 32020 6328 32026
rect 6276 31962 6328 31968
rect 6288 31754 6316 31962
rect 6196 31726 6316 31754
rect 6092 30320 6144 30326
rect 6092 30262 6144 30268
rect 5960 30144 6040 30172
rect 6092 30184 6144 30190
rect 5908 30126 5960 30132
rect 6092 30126 6144 30132
rect 5722 29880 5778 29889
rect 6104 29866 6132 30126
rect 6196 30122 6224 31726
rect 6380 31482 6408 32166
rect 6368 31476 6420 31482
rect 6368 31418 6420 31424
rect 6368 31272 6420 31278
rect 6368 31214 6420 31220
rect 6184 30116 6236 30122
rect 6184 30058 6236 30064
rect 5722 29815 5778 29824
rect 6012 29838 6132 29866
rect 5736 29646 5764 29815
rect 5908 29708 5960 29714
rect 5908 29650 5960 29656
rect 5724 29640 5776 29646
rect 5724 29582 5776 29588
rect 5540 29572 5592 29578
rect 5540 29514 5592 29520
rect 5588 29404 5884 29424
rect 5644 29402 5668 29404
rect 5724 29402 5748 29404
rect 5804 29402 5828 29404
rect 5666 29350 5668 29402
rect 5730 29350 5742 29402
rect 5804 29350 5806 29402
rect 5644 29348 5668 29350
rect 5724 29348 5748 29350
rect 5804 29348 5828 29350
rect 5588 29328 5884 29348
rect 5448 29164 5500 29170
rect 5448 29106 5500 29112
rect 5356 29096 5408 29102
rect 5356 29038 5408 29044
rect 5816 29028 5868 29034
rect 5276 28966 5396 28994
rect 5816 28970 5868 28976
rect 5264 28688 5316 28694
rect 5264 28630 5316 28636
rect 5172 28552 5224 28558
rect 5172 28494 5224 28500
rect 5080 27396 5132 27402
rect 5080 27338 5132 27344
rect 5080 26852 5132 26858
rect 5080 26794 5132 26800
rect 5092 24750 5120 26794
rect 5172 26308 5224 26314
rect 5172 26250 5224 26256
rect 5184 25838 5212 26250
rect 5172 25832 5224 25838
rect 5172 25774 5224 25780
rect 5276 25650 5304 28630
rect 5184 25622 5304 25650
rect 5368 25650 5396 28966
rect 5828 28762 5856 28970
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 5448 28552 5500 28558
rect 5448 28494 5500 28500
rect 5460 28218 5488 28494
rect 5588 28316 5884 28336
rect 5644 28314 5668 28316
rect 5724 28314 5748 28316
rect 5804 28314 5828 28316
rect 5666 28262 5668 28314
rect 5730 28262 5742 28314
rect 5804 28262 5806 28314
rect 5644 28260 5668 28262
rect 5724 28260 5748 28262
rect 5804 28260 5828 28262
rect 5588 28240 5884 28260
rect 5448 28212 5500 28218
rect 5448 28154 5500 28160
rect 5920 27334 5948 29650
rect 5908 27328 5960 27334
rect 5908 27270 5960 27276
rect 5588 27228 5884 27248
rect 5644 27226 5668 27228
rect 5724 27226 5748 27228
rect 5804 27226 5828 27228
rect 5666 27174 5668 27226
rect 5730 27174 5742 27226
rect 5804 27174 5806 27226
rect 5644 27172 5668 27174
rect 5724 27172 5748 27174
rect 5804 27172 5828 27174
rect 5588 27152 5884 27172
rect 5908 26580 5960 26586
rect 5908 26522 5960 26528
rect 5588 26140 5884 26160
rect 5644 26138 5668 26140
rect 5724 26138 5748 26140
rect 5804 26138 5828 26140
rect 5666 26086 5668 26138
rect 5730 26086 5742 26138
rect 5804 26086 5806 26138
rect 5644 26084 5668 26086
rect 5724 26084 5748 26086
rect 5804 26084 5828 26086
rect 5588 26064 5884 26084
rect 5368 25622 5488 25650
rect 5080 24744 5132 24750
rect 5080 24686 5132 24692
rect 5092 22234 5120 24686
rect 5080 22228 5132 22234
rect 5080 22170 5132 22176
rect 5184 22098 5212 25622
rect 5460 25498 5488 25622
rect 5356 25492 5408 25498
rect 5356 25434 5408 25440
rect 5448 25492 5500 25498
rect 5448 25434 5500 25440
rect 5264 25152 5316 25158
rect 5264 25094 5316 25100
rect 5276 24818 5304 25094
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 5264 24200 5316 24206
rect 5264 24142 5316 24148
rect 5276 22409 5304 24142
rect 5262 22400 5318 22409
rect 5262 22335 5318 22344
rect 5172 22092 5224 22098
rect 5172 22034 5224 22040
rect 5078 21992 5134 22001
rect 5078 21927 5134 21936
rect 4988 21684 5040 21690
rect 4988 21626 5040 21632
rect 5092 21570 5120 21927
rect 5000 21542 5120 21570
rect 5000 19242 5028 21542
rect 5080 20392 5132 20398
rect 5080 20334 5132 20340
rect 4988 19236 5040 19242
rect 4988 19178 5040 19184
rect 4986 18864 5042 18873
rect 4986 18799 5042 18808
rect 5000 17270 5028 18799
rect 5092 18222 5120 20334
rect 5184 20330 5212 22034
rect 5368 21298 5396 25434
rect 5448 25356 5500 25362
rect 5448 25298 5500 25304
rect 5276 21270 5396 21298
rect 5172 20324 5224 20330
rect 5172 20266 5224 20272
rect 5276 19394 5304 21270
rect 5356 21140 5408 21146
rect 5356 21082 5408 21088
rect 5184 19366 5304 19394
rect 5184 19310 5212 19366
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5184 18902 5212 19246
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5172 18896 5224 18902
rect 5172 18838 5224 18844
rect 5172 18760 5224 18766
rect 5276 18748 5304 19178
rect 5224 18720 5304 18748
rect 5172 18702 5224 18708
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5172 17808 5224 17814
rect 5172 17750 5224 17756
rect 5184 17338 5212 17750
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 4988 17264 5040 17270
rect 4988 17206 5040 17212
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 5000 16250 5028 17070
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5080 15972 5132 15978
rect 5080 15914 5132 15920
rect 5092 15706 5120 15914
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 5092 15094 5120 15642
rect 5080 15088 5132 15094
rect 5184 15065 5212 15982
rect 5080 15030 5132 15036
rect 5170 15056 5226 15065
rect 5170 14991 5226 15000
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 5000 13938 5028 14214
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4816 10130 4844 10406
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4908 9518 4936 13806
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5000 11626 5028 12038
rect 5092 11762 5120 14894
rect 5184 14822 5212 14991
rect 5276 14958 5304 18720
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5184 12986 5212 13262
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 5092 11082 5120 11698
rect 5184 11626 5212 12582
rect 5172 11620 5224 11626
rect 5172 11562 5224 11568
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4908 8634 4936 9318
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5184 7936 5212 11562
rect 5368 11218 5396 21082
rect 5460 18426 5488 25298
rect 5588 25052 5884 25072
rect 5644 25050 5668 25052
rect 5724 25050 5748 25052
rect 5804 25050 5828 25052
rect 5666 24998 5668 25050
rect 5730 24998 5742 25050
rect 5804 24998 5806 25050
rect 5644 24996 5668 24998
rect 5724 24996 5748 24998
rect 5804 24996 5828 24998
rect 5588 24976 5884 24996
rect 5920 24834 5948 26522
rect 5552 24806 5948 24834
rect 5552 24682 5580 24806
rect 5816 24744 5868 24750
rect 5868 24704 5948 24732
rect 5816 24686 5868 24692
rect 5540 24676 5592 24682
rect 5540 24618 5592 24624
rect 5816 24608 5868 24614
rect 5816 24550 5868 24556
rect 5828 24410 5856 24550
rect 5816 24404 5868 24410
rect 5816 24346 5868 24352
rect 5588 23964 5884 23984
rect 5644 23962 5668 23964
rect 5724 23962 5748 23964
rect 5804 23962 5828 23964
rect 5666 23910 5668 23962
rect 5730 23910 5742 23962
rect 5804 23910 5806 23962
rect 5644 23908 5668 23910
rect 5724 23908 5748 23910
rect 5804 23908 5828 23910
rect 5588 23888 5884 23908
rect 5920 23798 5948 24704
rect 6012 24070 6040 29838
rect 6196 29730 6224 30058
rect 6104 29702 6224 29730
rect 6104 28098 6132 29702
rect 6276 29572 6328 29578
rect 6276 29514 6328 29520
rect 6184 28552 6236 28558
rect 6184 28494 6236 28500
rect 6196 28218 6224 28494
rect 6184 28212 6236 28218
rect 6184 28154 6236 28160
rect 6104 28070 6224 28098
rect 6092 26308 6144 26314
rect 6092 26250 6144 26256
rect 6104 24886 6132 26250
rect 6196 25906 6224 28070
rect 6288 27282 6316 29514
rect 6380 28422 6408 31214
rect 6368 28416 6420 28422
rect 6368 28358 6420 28364
rect 6380 27402 6408 28358
rect 6368 27396 6420 27402
rect 6368 27338 6420 27344
rect 6288 27254 6408 27282
rect 6380 27062 6408 27254
rect 6368 27056 6420 27062
rect 6368 26998 6420 27004
rect 6276 26988 6328 26994
rect 6276 26930 6328 26936
rect 6184 25900 6236 25906
rect 6184 25842 6236 25848
rect 6092 24880 6144 24886
rect 6092 24822 6144 24828
rect 6092 24608 6144 24614
rect 6092 24550 6144 24556
rect 6000 24064 6052 24070
rect 6000 24006 6052 24012
rect 6104 23866 6132 24550
rect 6092 23860 6144 23866
rect 6092 23802 6144 23808
rect 5908 23792 5960 23798
rect 5908 23734 5960 23740
rect 6092 23588 6144 23594
rect 6092 23530 6144 23536
rect 6104 23050 6132 23530
rect 6092 23044 6144 23050
rect 6092 22986 6144 22992
rect 5588 22876 5884 22896
rect 5644 22874 5668 22876
rect 5724 22874 5748 22876
rect 5804 22874 5828 22876
rect 5666 22822 5668 22874
rect 5730 22822 5742 22874
rect 5804 22822 5806 22874
rect 5644 22820 5668 22822
rect 5724 22820 5748 22822
rect 5804 22820 5828 22822
rect 5588 22800 5884 22820
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5552 22030 5580 22578
rect 5632 22228 5684 22234
rect 5632 22170 5684 22176
rect 5540 22024 5592 22030
rect 5538 21992 5540 22001
rect 5592 21992 5594 22001
rect 5644 21962 5672 22170
rect 5908 22160 5960 22166
rect 5908 22102 5960 22108
rect 5538 21927 5594 21936
rect 5632 21956 5684 21962
rect 5632 21898 5684 21904
rect 5588 21788 5884 21808
rect 5644 21786 5668 21788
rect 5724 21786 5748 21788
rect 5804 21786 5828 21788
rect 5666 21734 5668 21786
rect 5730 21734 5742 21786
rect 5804 21734 5806 21786
rect 5644 21732 5668 21734
rect 5724 21732 5748 21734
rect 5804 21732 5828 21734
rect 5588 21712 5884 21732
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5828 20788 5856 21490
rect 5920 21078 5948 22102
rect 6000 21956 6052 21962
rect 6000 21898 6052 21904
rect 5908 21072 5960 21078
rect 5908 21014 5960 21020
rect 5828 20760 5948 20788
rect 5588 20700 5884 20720
rect 5644 20698 5668 20700
rect 5724 20698 5748 20700
rect 5804 20698 5828 20700
rect 5666 20646 5668 20698
rect 5730 20646 5742 20698
rect 5804 20646 5806 20698
rect 5644 20644 5668 20646
rect 5724 20644 5748 20646
rect 5804 20644 5828 20646
rect 5588 20624 5884 20644
rect 5588 19612 5884 19632
rect 5644 19610 5668 19612
rect 5724 19610 5748 19612
rect 5804 19610 5828 19612
rect 5666 19558 5668 19610
rect 5730 19558 5742 19610
rect 5804 19558 5806 19610
rect 5644 19556 5668 19558
rect 5724 19556 5748 19558
rect 5804 19556 5828 19558
rect 5588 19536 5884 19556
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5552 18873 5580 18906
rect 5538 18864 5594 18873
rect 5538 18799 5594 18808
rect 5588 18524 5884 18544
rect 5644 18522 5668 18524
rect 5724 18522 5748 18524
rect 5804 18522 5828 18524
rect 5666 18470 5668 18522
rect 5730 18470 5742 18522
rect 5804 18470 5806 18522
rect 5644 18468 5668 18470
rect 5724 18468 5748 18470
rect 5804 18468 5828 18470
rect 5588 18448 5884 18468
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5920 18290 5948 20760
rect 6012 18630 6040 21898
rect 6092 20392 6144 20398
rect 6092 20334 6144 20340
rect 6104 19446 6132 20334
rect 6196 19718 6224 25842
rect 6288 25158 6316 26930
rect 6380 25226 6408 26998
rect 6472 26042 6500 44390
rect 6656 43994 6684 44746
rect 6736 44736 6788 44742
rect 6736 44678 6788 44684
rect 6748 44334 6776 44678
rect 6736 44328 6788 44334
rect 6736 44270 6788 44276
rect 6644 43988 6696 43994
rect 6644 43930 6696 43936
rect 6840 43926 6868 44882
rect 6828 43920 6880 43926
rect 6828 43862 6880 43868
rect 6552 43240 6604 43246
rect 6552 43182 6604 43188
rect 6564 39982 6592 43182
rect 6644 41200 6696 41206
rect 6644 41142 6696 41148
rect 6656 41002 6684 41142
rect 6644 40996 6696 41002
rect 6644 40938 6696 40944
rect 7024 40458 7052 52906
rect 7564 52556 7616 52562
rect 7564 52498 7616 52504
rect 7576 51882 7604 52498
rect 7748 52352 7800 52358
rect 7748 52294 7800 52300
rect 7760 51950 7788 52294
rect 7748 51944 7800 51950
rect 7748 51886 7800 51892
rect 7564 51876 7616 51882
rect 7564 51818 7616 51824
rect 7576 50862 7604 51818
rect 7656 51468 7708 51474
rect 7656 51410 7708 51416
rect 7668 51074 7696 51410
rect 7668 51046 7788 51074
rect 7104 50856 7156 50862
rect 7104 50798 7156 50804
rect 7564 50856 7616 50862
rect 7564 50798 7616 50804
rect 7116 50386 7144 50798
rect 7576 50386 7604 50798
rect 7104 50380 7156 50386
rect 7104 50322 7156 50328
rect 7564 50380 7616 50386
rect 7564 50322 7616 50328
rect 7116 48346 7144 50322
rect 7656 50312 7708 50318
rect 7656 50254 7708 50260
rect 7104 48340 7156 48346
rect 7104 48282 7156 48288
rect 7104 48204 7156 48210
rect 7104 48146 7156 48152
rect 7196 48204 7248 48210
rect 7196 48146 7248 48152
rect 7116 47462 7144 48146
rect 7104 47456 7156 47462
rect 7104 47398 7156 47404
rect 7116 47122 7144 47398
rect 7208 47258 7236 48146
rect 7288 47728 7340 47734
rect 7288 47670 7340 47676
rect 7196 47252 7248 47258
rect 7196 47194 7248 47200
rect 7300 47122 7328 47670
rect 7104 47116 7156 47122
rect 7104 47058 7156 47064
rect 7288 47116 7340 47122
rect 7288 47058 7340 47064
rect 7564 47048 7616 47054
rect 7564 46990 7616 46996
rect 7576 45626 7604 46990
rect 7564 45620 7616 45626
rect 7564 45562 7616 45568
rect 7472 45484 7524 45490
rect 7472 45426 7524 45432
rect 7104 44736 7156 44742
rect 7104 44678 7156 44684
rect 7116 44402 7144 44678
rect 7104 44396 7156 44402
rect 7104 44338 7156 44344
rect 7116 41614 7144 44338
rect 7380 42628 7432 42634
rect 7380 42570 7432 42576
rect 7104 41608 7156 41614
rect 7104 41550 7156 41556
rect 7196 41472 7248 41478
rect 7196 41414 7248 41420
rect 7104 40928 7156 40934
rect 7104 40870 7156 40876
rect 7012 40452 7064 40458
rect 7012 40394 7064 40400
rect 6920 40384 6972 40390
rect 6920 40326 6972 40332
rect 6552 39976 6604 39982
rect 6552 39918 6604 39924
rect 6552 39840 6604 39846
rect 6552 39782 6604 39788
rect 6460 26036 6512 26042
rect 6460 25978 6512 25984
rect 6368 25220 6420 25226
rect 6368 25162 6420 25168
rect 6276 25152 6328 25158
rect 6276 25094 6328 25100
rect 6288 22642 6316 25094
rect 6460 24812 6512 24818
rect 6460 24754 6512 24760
rect 6472 24342 6500 24754
rect 6460 24336 6512 24342
rect 6460 24278 6512 24284
rect 6276 22636 6328 22642
rect 6276 22578 6328 22584
rect 6460 22636 6512 22642
rect 6460 22578 6512 22584
rect 6276 21956 6328 21962
rect 6276 21898 6328 21904
rect 6288 21486 6316 21898
rect 6368 21616 6420 21622
rect 6368 21558 6420 21564
rect 6276 21480 6328 21486
rect 6276 21422 6328 21428
rect 6380 20398 6408 21558
rect 6472 21486 6500 22578
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 6380 19786 6408 20334
rect 6368 19780 6420 19786
rect 6368 19722 6420 19728
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 6092 19440 6144 19446
rect 6092 19382 6144 19388
rect 6104 18970 6132 19382
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 5908 18284 5960 18290
rect 5960 18244 6132 18272
rect 5908 18226 5960 18232
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 5908 17604 5960 17610
rect 5908 17546 5960 17552
rect 5588 17436 5884 17456
rect 5644 17434 5668 17436
rect 5724 17434 5748 17436
rect 5804 17434 5828 17436
rect 5666 17382 5668 17434
rect 5730 17382 5742 17434
rect 5804 17382 5806 17434
rect 5644 17380 5668 17382
rect 5724 17380 5748 17382
rect 5804 17380 5828 17382
rect 5588 17360 5884 17380
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5644 16794 5672 16934
rect 5920 16794 5948 17546
rect 6012 17066 6040 18090
rect 6104 17202 6132 18244
rect 6196 17814 6224 19654
rect 6380 19378 6408 19722
rect 6368 19372 6420 19378
rect 6368 19314 6420 19320
rect 6276 18624 6328 18630
rect 6276 18566 6328 18572
rect 6184 17808 6236 17814
rect 6184 17750 6236 17756
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 6000 17060 6052 17066
rect 6000 17002 6052 17008
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5908 16788 5960 16794
rect 5908 16730 5960 16736
rect 5588 16348 5884 16368
rect 5644 16346 5668 16348
rect 5724 16346 5748 16348
rect 5804 16346 5828 16348
rect 5666 16294 5668 16346
rect 5730 16294 5742 16346
rect 5804 16294 5806 16346
rect 5644 16292 5668 16294
rect 5724 16292 5748 16294
rect 5804 16292 5828 16294
rect 5588 16272 5884 16292
rect 5908 16176 5960 16182
rect 5908 16118 5960 16124
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5460 14958 5488 15642
rect 5588 15260 5884 15280
rect 5644 15258 5668 15260
rect 5724 15258 5748 15260
rect 5804 15258 5828 15260
rect 5666 15206 5668 15258
rect 5730 15206 5742 15258
rect 5804 15206 5806 15258
rect 5644 15204 5668 15206
rect 5724 15204 5748 15206
rect 5804 15204 5828 15206
rect 5588 15184 5884 15204
rect 5920 14958 5948 16118
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5908 14952 5960 14958
rect 5960 14912 6132 14940
rect 5908 14894 5960 14900
rect 5816 14884 5868 14890
rect 5816 14826 5868 14832
rect 5828 14770 5856 14826
rect 5828 14742 5948 14770
rect 5588 14172 5884 14192
rect 5644 14170 5668 14172
rect 5724 14170 5748 14172
rect 5804 14170 5828 14172
rect 5666 14118 5668 14170
rect 5730 14118 5742 14170
rect 5804 14118 5806 14170
rect 5644 14116 5668 14118
rect 5724 14116 5748 14118
rect 5804 14116 5828 14118
rect 5588 14096 5884 14116
rect 5588 13084 5884 13104
rect 5644 13082 5668 13084
rect 5724 13082 5748 13084
rect 5804 13082 5828 13084
rect 5666 13030 5668 13082
rect 5730 13030 5742 13082
rect 5804 13030 5806 13082
rect 5644 13028 5668 13030
rect 5724 13028 5748 13030
rect 5804 13028 5828 13030
rect 5588 13008 5884 13028
rect 5920 12866 5948 14742
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 5828 12838 5948 12866
rect 5828 12186 5856 12838
rect 6012 12782 6040 13126
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 5920 12442 5948 12718
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5828 12158 5948 12186
rect 5920 12102 5948 12158
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5588 11996 5884 12016
rect 5644 11994 5668 11996
rect 5724 11994 5748 11996
rect 5804 11994 5828 11996
rect 5666 11942 5668 11994
rect 5730 11942 5742 11994
rect 5804 11942 5806 11994
rect 5644 11940 5668 11942
rect 5724 11940 5748 11942
rect 5804 11940 5828 11942
rect 5588 11920 5884 11940
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5644 11286 5672 11494
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5276 8634 5304 11086
rect 5368 10538 5396 11154
rect 5588 10908 5884 10928
rect 5644 10906 5668 10908
rect 5724 10906 5748 10908
rect 5804 10906 5828 10908
rect 5666 10854 5668 10906
rect 5730 10854 5742 10906
rect 5804 10854 5806 10906
rect 5644 10852 5668 10854
rect 5724 10852 5748 10854
rect 5804 10852 5828 10854
rect 5588 10832 5884 10852
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5368 9722 5396 10474
rect 5588 9820 5884 9840
rect 5644 9818 5668 9820
rect 5724 9818 5748 9820
rect 5804 9818 5828 9820
rect 5666 9766 5668 9818
rect 5730 9766 5742 9818
rect 5804 9766 5806 9818
rect 5644 9764 5668 9766
rect 5724 9764 5748 9766
rect 5804 9764 5828 9766
rect 5588 9744 5884 9764
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5920 8838 5948 12038
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5588 8732 5884 8752
rect 5644 8730 5668 8732
rect 5724 8730 5748 8732
rect 5804 8730 5828 8732
rect 5666 8678 5668 8730
rect 5730 8678 5742 8730
rect 5804 8678 5806 8730
rect 5644 8676 5668 8678
rect 5724 8676 5748 8678
rect 5804 8676 5828 8678
rect 5588 8656 5884 8676
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5092 7908 5212 7936
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 4620 5092 4672 5098
rect 4620 5034 4672 5040
rect 5000 4282 5028 5102
rect 4988 4276 5040 4282
rect 4908 4236 4988 4264
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 3514 2615 3570 2624
rect 4528 2644 4580 2650
rect 3422 2272 3478 2281
rect 3422 2207 3478 2216
rect 3528 2038 3556 2615
rect 4528 2586 4580 2592
rect 3516 2032 3568 2038
rect 3516 1974 3568 1980
rect 3424 1896 3476 1902
rect 3422 1864 3424 1873
rect 3476 1864 3478 1873
rect 3422 1799 3478 1808
rect 4724 800 4752 3946
rect 4908 3398 4936 4236
rect 4988 4218 5040 4224
rect 5092 3738 5120 7908
rect 5276 7342 5304 8570
rect 6012 8566 6040 11018
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 5368 7818 5580 7834
rect 5368 7812 5592 7818
rect 5368 7806 5540 7812
rect 5368 7478 5396 7806
rect 5540 7754 5592 7760
rect 5588 7644 5884 7664
rect 5644 7642 5668 7644
rect 5724 7642 5748 7644
rect 5804 7642 5828 7644
rect 5666 7590 5668 7642
rect 5730 7590 5742 7642
rect 5804 7590 5806 7642
rect 5644 7588 5668 7590
rect 5724 7588 5748 7590
rect 5804 7588 5828 7590
rect 5588 7568 5884 7588
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5552 6798 5580 7210
rect 5828 6798 5856 7346
rect 5920 7342 5948 7958
rect 6012 7410 6040 8502
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5184 6254 5212 6598
rect 5588 6556 5884 6576
rect 5644 6554 5668 6556
rect 5724 6554 5748 6556
rect 5804 6554 5828 6556
rect 5666 6502 5668 6554
rect 5730 6502 5742 6554
rect 5804 6502 5806 6554
rect 5644 6500 5668 6502
rect 5724 6500 5748 6502
rect 5804 6500 5828 6502
rect 5588 6480 5884 6500
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4908 3058 4936 3334
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 5000 2650 5028 3538
rect 5460 3466 5488 6054
rect 5588 5468 5884 5488
rect 5644 5466 5668 5468
rect 5724 5466 5748 5468
rect 5804 5466 5828 5468
rect 5666 5414 5668 5466
rect 5730 5414 5742 5466
rect 5804 5414 5806 5466
rect 5644 5412 5668 5414
rect 5724 5412 5748 5414
rect 5804 5412 5828 5414
rect 5588 5392 5884 5412
rect 5920 4826 5948 6870
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6012 6322 6040 6802
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6012 5302 6040 6258
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5588 4380 5884 4400
rect 5644 4378 5668 4380
rect 5724 4378 5748 4380
rect 5804 4378 5828 4380
rect 5666 4326 5668 4378
rect 5730 4326 5742 4378
rect 5804 4326 5806 4378
rect 5644 4324 5668 4326
rect 5724 4324 5748 4326
rect 5804 4324 5828 4326
rect 5588 4304 5884 4324
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5588 3292 5884 3312
rect 5644 3290 5668 3292
rect 5724 3290 5748 3292
rect 5804 3290 5828 3292
rect 5666 3238 5668 3290
rect 5730 3238 5742 3290
rect 5804 3238 5806 3290
rect 5644 3236 5668 3238
rect 5724 3236 5748 3238
rect 5804 3236 5828 3238
rect 5588 3216 5884 3236
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5588 2204 5884 2224
rect 5644 2202 5668 2204
rect 5724 2202 5748 2204
rect 5804 2202 5828 2204
rect 5666 2150 5668 2202
rect 5730 2150 5742 2202
rect 5804 2150 5806 2202
rect 5644 2148 5668 2150
rect 5724 2148 5748 2150
rect 5804 2148 5828 2150
rect 5588 2128 5884 2148
rect 5920 1970 5948 4626
rect 6104 4554 6132 14912
rect 6196 12782 6224 17750
rect 6288 14958 6316 18566
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6472 14482 6500 14758
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6196 10130 6224 12718
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6380 11898 6408 12242
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6472 11762 6500 13262
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6288 10674 6316 11698
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6196 9518 6224 10066
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6288 7750 6316 10610
rect 6564 8294 6592 39782
rect 6932 39506 6960 40326
rect 6920 39500 6972 39506
rect 6920 39442 6972 39448
rect 6932 38894 6960 39442
rect 7116 39438 7144 40870
rect 7208 40730 7236 41414
rect 7392 41138 7420 42570
rect 7484 41414 7512 45426
rect 7576 44946 7604 45562
rect 7668 45354 7696 50254
rect 7760 49298 7788 51046
rect 7748 49292 7800 49298
rect 7748 49234 7800 49240
rect 7656 45348 7708 45354
rect 7656 45290 7708 45296
rect 7748 45280 7800 45286
rect 7748 45222 7800 45228
rect 7564 44940 7616 44946
rect 7564 44882 7616 44888
rect 7576 44334 7604 44882
rect 7564 44328 7616 44334
rect 7564 44270 7616 44276
rect 7760 44266 7788 45222
rect 7748 44260 7800 44266
rect 7748 44202 7800 44208
rect 7748 43784 7800 43790
rect 7748 43726 7800 43732
rect 7760 42770 7788 43726
rect 7748 42764 7800 42770
rect 7748 42706 7800 42712
rect 7656 42220 7708 42226
rect 7656 42162 7708 42168
rect 7668 41818 7696 42162
rect 7656 41812 7708 41818
rect 7656 41754 7708 41760
rect 7484 41386 7696 41414
rect 7380 41132 7432 41138
rect 7380 41074 7432 41080
rect 7668 40730 7696 41386
rect 7852 41002 7880 52906
rect 8024 52488 8076 52494
rect 8024 52430 8076 52436
rect 7932 51876 7984 51882
rect 7932 51818 7984 51824
rect 7944 51474 7972 51818
rect 7932 51468 7984 51474
rect 7932 51410 7984 51416
rect 8036 50386 8064 52430
rect 8128 52414 8432 52442
rect 8128 52018 8156 52414
rect 8404 52358 8432 52414
rect 9680 52420 9732 52426
rect 9680 52362 9732 52368
rect 8300 52352 8352 52358
rect 8300 52294 8352 52300
rect 8392 52352 8444 52358
rect 8392 52294 8444 52300
rect 8116 52012 8168 52018
rect 8116 51954 8168 51960
rect 8312 51898 8340 52294
rect 8484 52012 8536 52018
rect 8484 51954 8536 51960
rect 8128 51870 8340 51898
rect 8128 51610 8156 51870
rect 8208 51808 8260 51814
rect 8208 51750 8260 51756
rect 8116 51604 8168 51610
rect 8116 51546 8168 51552
rect 8220 51474 8248 51750
rect 8496 51474 8524 51954
rect 9588 51808 9640 51814
rect 9692 51762 9720 52362
rect 9772 51944 9824 51950
rect 9772 51886 9824 51892
rect 9640 51756 9720 51762
rect 9588 51750 9720 51756
rect 9600 51734 9720 51750
rect 8208 51468 8260 51474
rect 8208 51410 8260 51416
rect 8484 51468 8536 51474
rect 8484 51410 8536 51416
rect 9692 51270 9720 51734
rect 8576 51264 8628 51270
rect 8576 51206 8628 51212
rect 9680 51264 9732 51270
rect 9680 51206 9732 51212
rect 8116 50788 8168 50794
rect 8116 50730 8168 50736
rect 8128 50522 8156 50730
rect 8300 50720 8352 50726
rect 8300 50662 8352 50668
rect 8116 50516 8168 50522
rect 8116 50458 8168 50464
rect 8312 50386 8340 50662
rect 8024 50380 8076 50386
rect 8024 50322 8076 50328
rect 8300 50380 8352 50386
rect 8300 50322 8352 50328
rect 7932 49292 7984 49298
rect 7932 49234 7984 49240
rect 7944 48890 7972 49234
rect 7932 48884 7984 48890
rect 7932 48826 7984 48832
rect 8036 48822 8064 50322
rect 8208 49768 8260 49774
rect 8208 49710 8260 49716
rect 8024 48816 8076 48822
rect 8024 48758 8076 48764
rect 8220 48278 8248 49710
rect 8300 48680 8352 48686
rect 8300 48622 8352 48628
rect 8208 48272 8260 48278
rect 8208 48214 8260 48220
rect 8312 48210 8340 48622
rect 8300 48204 8352 48210
rect 8300 48146 8352 48152
rect 8588 48142 8616 51206
rect 9496 50924 9548 50930
rect 9496 50866 9548 50872
rect 9220 50720 9272 50726
rect 9220 50662 9272 50668
rect 9232 50386 9260 50662
rect 9508 50386 9536 50866
rect 9220 50380 9272 50386
rect 9220 50322 9272 50328
rect 9496 50380 9548 50386
rect 9496 50322 9548 50328
rect 9588 49224 9640 49230
rect 9588 49166 9640 49172
rect 9036 49088 9088 49094
rect 9036 49030 9088 49036
rect 9048 48618 9076 49030
rect 9036 48612 9088 48618
rect 9036 48554 9088 48560
rect 8576 48136 8628 48142
rect 8576 48078 8628 48084
rect 8588 47682 8616 48078
rect 8496 47654 8616 47682
rect 9048 47666 9076 48554
rect 9600 48550 9628 49166
rect 9588 48544 9640 48550
rect 9588 48486 9640 48492
rect 9600 48210 9628 48486
rect 9588 48204 9640 48210
rect 9588 48146 9640 48152
rect 9036 47660 9088 47666
rect 8392 47524 8444 47530
rect 8496 47512 8524 47654
rect 9036 47602 9088 47608
rect 8944 47592 8996 47598
rect 8944 47534 8996 47540
rect 8444 47484 8524 47512
rect 8576 47524 8628 47530
rect 8392 47466 8444 47472
rect 8576 47466 8628 47472
rect 8208 46912 8260 46918
rect 8208 46854 8260 46860
rect 8220 46102 8248 46854
rect 8300 46572 8352 46578
rect 8404 46560 8432 47466
rect 8484 46912 8536 46918
rect 8588 46900 8616 47466
rect 8668 47456 8720 47462
rect 8668 47398 8720 47404
rect 8536 46872 8616 46900
rect 8484 46854 8536 46860
rect 8352 46532 8432 46560
rect 8300 46514 8352 46520
rect 8208 46096 8260 46102
rect 8208 46038 8260 46044
rect 8024 45348 8076 45354
rect 8024 45290 8076 45296
rect 8036 44946 8064 45290
rect 7932 44940 7984 44946
rect 7932 44882 7984 44888
rect 8024 44940 8076 44946
rect 8024 44882 8076 44888
rect 7944 43994 7972 44882
rect 8036 44198 8064 44882
rect 8404 44742 8432 46532
rect 8496 46510 8524 46854
rect 8680 46510 8708 47398
rect 8956 47122 8984 47534
rect 9600 47530 9628 48146
rect 9588 47524 9640 47530
rect 9588 47466 9640 47472
rect 9588 47184 9640 47190
rect 9588 47126 9640 47132
rect 8944 47116 8996 47122
rect 8944 47058 8996 47064
rect 9404 47116 9456 47122
rect 9404 47058 9456 47064
rect 8484 46504 8536 46510
rect 8484 46446 8536 46452
rect 8668 46504 8720 46510
rect 8668 46446 8720 46452
rect 8680 46374 8708 46446
rect 8668 46368 8720 46374
rect 8668 46310 8720 46316
rect 8760 44872 8812 44878
rect 8760 44814 8812 44820
rect 8392 44736 8444 44742
rect 8392 44678 8444 44684
rect 8208 44260 8260 44266
rect 8208 44202 8260 44208
rect 8024 44192 8076 44198
rect 8024 44134 8076 44140
rect 8220 43994 8248 44202
rect 7932 43988 7984 43994
rect 7932 43930 7984 43936
rect 8208 43988 8260 43994
rect 8208 43930 8260 43936
rect 8772 41818 8800 44814
rect 8852 42560 8904 42566
rect 8852 42502 8904 42508
rect 8760 41812 8812 41818
rect 8760 41754 8812 41760
rect 8116 41676 8168 41682
rect 8116 41618 8168 41624
rect 8484 41676 8536 41682
rect 8484 41618 8536 41624
rect 8128 41274 8156 41618
rect 8300 41608 8352 41614
rect 8300 41550 8352 41556
rect 8116 41268 8168 41274
rect 8116 41210 8168 41216
rect 7840 40996 7892 41002
rect 7840 40938 7892 40944
rect 7196 40724 7248 40730
rect 7196 40666 7248 40672
rect 7656 40724 7708 40730
rect 7656 40666 7708 40672
rect 7196 40588 7248 40594
rect 7196 40530 7248 40536
rect 7208 40050 7236 40530
rect 7196 40044 7248 40050
rect 7196 39986 7248 39992
rect 7748 39976 7800 39982
rect 7748 39918 7800 39924
rect 7104 39432 7156 39438
rect 7104 39374 7156 39380
rect 6920 38888 6972 38894
rect 6920 38830 6972 38836
rect 7116 38826 7144 39374
rect 7760 39302 7788 39918
rect 8116 39840 8168 39846
rect 8116 39782 8168 39788
rect 8128 39370 8156 39782
rect 8116 39364 8168 39370
rect 8116 39306 8168 39312
rect 7748 39296 7800 39302
rect 7748 39238 7800 39244
rect 7760 38894 7788 39238
rect 8128 38962 8156 39306
rect 8312 39098 8340 41550
rect 8496 39982 8524 41618
rect 8772 41414 8800 41754
rect 8864 41682 8892 42502
rect 8852 41676 8904 41682
rect 8852 41618 8904 41624
rect 8680 41386 8800 41414
rect 8680 39982 8708 41386
rect 8484 39976 8536 39982
rect 8668 39976 8720 39982
rect 8536 39936 8616 39964
rect 8484 39918 8536 39924
rect 8484 39500 8536 39506
rect 8484 39442 8536 39448
rect 8496 39098 8524 39442
rect 8588 39438 8616 39936
rect 8668 39918 8720 39924
rect 8680 39506 8708 39918
rect 8668 39500 8720 39506
rect 8668 39442 8720 39448
rect 8576 39432 8628 39438
rect 8576 39374 8628 39380
rect 8300 39092 8352 39098
rect 8300 39034 8352 39040
rect 8484 39092 8536 39098
rect 8484 39034 8536 39040
rect 8116 38956 8168 38962
rect 8116 38898 8168 38904
rect 7748 38888 7800 38894
rect 7748 38830 7800 38836
rect 7104 38820 7156 38826
rect 7104 38762 7156 38768
rect 6828 37664 6880 37670
rect 6828 37606 6880 37612
rect 6840 36242 6868 37606
rect 6828 36236 6880 36242
rect 6828 36178 6880 36184
rect 6644 35760 6696 35766
rect 6644 35702 6696 35708
rect 6656 34610 6684 35702
rect 6644 34604 6696 34610
rect 6644 34546 6696 34552
rect 6644 33448 6696 33454
rect 6644 33390 6696 33396
rect 6656 30394 6684 33390
rect 6736 31884 6788 31890
rect 6736 31826 6788 31832
rect 6644 30388 6696 30394
rect 6644 30330 6696 30336
rect 6748 30326 6776 31826
rect 6736 30320 6788 30326
rect 6736 30262 6788 30268
rect 6644 30184 6696 30190
rect 6644 30126 6696 30132
rect 6656 29714 6684 30126
rect 6644 29708 6696 29714
rect 6644 29650 6696 29656
rect 6840 29594 6868 36178
rect 6920 35556 6972 35562
rect 6920 35498 6972 35504
rect 6932 35018 6960 35498
rect 6920 35012 6972 35018
rect 6920 34954 6972 34960
rect 7116 32502 7144 38762
rect 8852 38412 8904 38418
rect 8852 38354 8904 38360
rect 8760 37392 8812 37398
rect 8760 37334 8812 37340
rect 7288 37120 7340 37126
rect 7288 37062 7340 37068
rect 7300 36582 7328 37062
rect 7288 36576 7340 36582
rect 7288 36518 7340 36524
rect 7196 36236 7248 36242
rect 7196 36178 7248 36184
rect 7208 35834 7236 36178
rect 7196 35828 7248 35834
rect 7196 35770 7248 35776
rect 7300 35630 7328 36518
rect 8772 36106 8800 37334
rect 8864 37330 8892 38354
rect 8852 37324 8904 37330
rect 8852 37266 8904 37272
rect 8760 36100 8812 36106
rect 8760 36042 8812 36048
rect 7288 35624 7340 35630
rect 7288 35566 7340 35572
rect 8024 35556 8076 35562
rect 8024 35498 8076 35504
rect 7748 34944 7800 34950
rect 7748 34886 7800 34892
rect 7656 34060 7708 34066
rect 7656 34002 7708 34008
rect 7668 33658 7696 34002
rect 7760 33862 7788 34886
rect 7748 33856 7800 33862
rect 7748 33798 7800 33804
rect 7656 33652 7708 33658
rect 7656 33594 7708 33600
rect 7104 32496 7156 32502
rect 7104 32438 7156 32444
rect 7104 32292 7156 32298
rect 7104 32234 7156 32240
rect 7012 31884 7064 31890
rect 7012 31826 7064 31832
rect 7024 31210 7052 31826
rect 7116 31754 7144 32234
rect 7288 31952 7340 31958
rect 7288 31894 7340 31900
rect 7116 31726 7236 31754
rect 7104 31680 7156 31686
rect 7104 31622 7156 31628
rect 7012 31204 7064 31210
rect 7012 31146 7064 31152
rect 6920 30388 6972 30394
rect 6920 30330 6972 30336
rect 6656 29566 6868 29594
rect 6656 28490 6684 29566
rect 6828 29504 6880 29510
rect 6828 29446 6880 29452
rect 6840 29238 6868 29446
rect 6828 29232 6880 29238
rect 6828 29174 6880 29180
rect 6644 28484 6696 28490
rect 6644 28426 6696 28432
rect 6656 26790 6684 28426
rect 6840 28218 6868 29174
rect 6828 28212 6880 28218
rect 6828 28154 6880 28160
rect 6932 28098 6960 30330
rect 7116 28626 7144 31622
rect 7208 31346 7236 31726
rect 7300 31414 7328 31894
rect 7288 31408 7340 31414
rect 7288 31350 7340 31356
rect 7196 31340 7248 31346
rect 7196 31282 7248 31288
rect 7288 31204 7340 31210
rect 7288 31146 7340 31152
rect 7104 28620 7156 28626
rect 7104 28562 7156 28568
rect 7116 28506 7144 28562
rect 6840 28070 6960 28098
rect 7024 28478 7144 28506
rect 6736 28008 6788 28014
rect 6736 27950 6788 27956
rect 6748 27334 6776 27950
rect 6840 27470 6868 28070
rect 6920 27872 6972 27878
rect 6920 27814 6972 27820
rect 6932 27606 6960 27814
rect 7024 27606 7052 28478
rect 7104 28416 7156 28422
rect 7104 28358 7156 28364
rect 7116 28014 7144 28358
rect 7104 28008 7156 28014
rect 7104 27950 7156 27956
rect 7196 28008 7248 28014
rect 7196 27950 7248 27956
rect 7208 27674 7236 27950
rect 7196 27668 7248 27674
rect 7196 27610 7248 27616
rect 6920 27600 6972 27606
rect 6920 27542 6972 27548
rect 7012 27600 7064 27606
rect 7012 27542 7064 27548
rect 7196 27532 7248 27538
rect 7196 27474 7248 27480
rect 6828 27464 6880 27470
rect 6828 27406 6880 27412
rect 6736 27328 6788 27334
rect 6736 27270 6788 27276
rect 6644 26784 6696 26790
rect 6644 26726 6696 26732
rect 6840 26586 6868 27406
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 7208 26042 7236 27474
rect 7300 27130 7328 31146
rect 7564 30796 7616 30802
rect 7564 30738 7616 30744
rect 7472 30728 7524 30734
rect 7472 30670 7524 30676
rect 7484 28626 7512 30670
rect 7576 29238 7604 30738
rect 7760 29646 7788 33798
rect 7840 32768 7892 32774
rect 7840 32710 7892 32716
rect 7852 31958 7880 32710
rect 7840 31952 7892 31958
rect 7840 31894 7892 31900
rect 7932 31136 7984 31142
rect 7932 31078 7984 31084
rect 7944 30802 7972 31078
rect 7932 30796 7984 30802
rect 7932 30738 7984 30744
rect 7748 29640 7800 29646
rect 7748 29582 7800 29588
rect 7564 29232 7616 29238
rect 7564 29174 7616 29180
rect 7576 28694 7604 29174
rect 7760 29102 7788 29582
rect 7748 29096 7800 29102
rect 7748 29038 7800 29044
rect 7932 29096 7984 29102
rect 7932 29038 7984 29044
rect 7944 28762 7972 29038
rect 7932 28756 7984 28762
rect 7932 28698 7984 28704
rect 7564 28688 7616 28694
rect 7564 28630 7616 28636
rect 7472 28620 7524 28626
rect 7472 28562 7524 28568
rect 7380 28552 7432 28558
rect 7380 28494 7432 28500
rect 7392 28218 7420 28494
rect 7380 28212 7432 28218
rect 7380 28154 7432 28160
rect 7378 28112 7434 28121
rect 7378 28047 7380 28056
rect 7432 28047 7434 28056
rect 7380 28018 7432 28024
rect 7380 27328 7432 27334
rect 7380 27270 7432 27276
rect 7288 27124 7340 27130
rect 7288 27066 7340 27072
rect 7196 26036 7248 26042
rect 7196 25978 7248 25984
rect 7392 25922 7420 27270
rect 7484 26042 7512 28562
rect 7472 26036 7524 26042
rect 7472 25978 7524 25984
rect 7392 25894 7512 25922
rect 6920 25832 6972 25838
rect 6920 25774 6972 25780
rect 7380 25832 7432 25838
rect 7380 25774 7432 25780
rect 6644 25764 6696 25770
rect 6644 25706 6696 25712
rect 6656 24342 6684 25706
rect 6644 24336 6696 24342
rect 6644 24278 6696 24284
rect 6656 23866 6684 24278
rect 6828 24268 6880 24274
rect 6828 24210 6880 24216
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 6736 23792 6788 23798
rect 6736 23734 6788 23740
rect 6748 23186 6776 23734
rect 6840 23322 6868 24210
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6736 23180 6788 23186
rect 6736 23122 6788 23128
rect 6644 23044 6696 23050
rect 6644 22986 6696 22992
rect 6656 22574 6684 22986
rect 6748 22642 6776 23122
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6644 22568 6696 22574
rect 6644 22510 6696 22516
rect 6656 22166 6684 22510
rect 6644 22160 6696 22166
rect 6644 22102 6696 22108
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6656 18970 6684 21490
rect 6840 21010 6868 21626
rect 6932 21146 6960 25774
rect 7392 25430 7420 25774
rect 7380 25424 7432 25430
rect 7380 25366 7432 25372
rect 7392 24410 7420 25366
rect 7484 25242 7512 25894
rect 7576 25770 7604 28630
rect 7944 28218 7972 28698
rect 7932 28212 7984 28218
rect 7932 28154 7984 28160
rect 7656 28008 7708 28014
rect 7656 27950 7708 27956
rect 7668 27674 7696 27950
rect 7748 27872 7800 27878
rect 7748 27814 7800 27820
rect 7656 27668 7708 27674
rect 7656 27610 7708 27616
rect 7564 25764 7616 25770
rect 7564 25706 7616 25712
rect 7576 25362 7604 25706
rect 7564 25356 7616 25362
rect 7564 25298 7616 25304
rect 7484 25214 7604 25242
rect 7380 24404 7432 24410
rect 7380 24346 7432 24352
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 7024 19310 7052 24142
rect 7472 22432 7524 22438
rect 7472 22374 7524 22380
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 7116 21690 7144 22034
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 7104 21004 7156 21010
rect 7104 20946 7156 20952
rect 7288 21004 7340 21010
rect 7288 20946 7340 20952
rect 7116 19310 7144 20946
rect 7300 19394 7328 20946
rect 7484 20398 7512 22374
rect 7472 20392 7524 20398
rect 7392 20340 7472 20346
rect 7392 20334 7524 20340
rect 7392 20318 7512 20334
rect 7392 19990 7420 20318
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7380 19984 7432 19990
rect 7380 19926 7432 19932
rect 7484 19922 7512 20198
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7300 19366 7420 19394
rect 7392 19310 7420 19366
rect 7484 19310 7512 19858
rect 7012 19304 7064 19310
rect 6932 19252 7012 19258
rect 6932 19246 7064 19252
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7472 19304 7524 19310
rect 7472 19246 7524 19252
rect 6932 19230 7052 19246
rect 6932 19174 6960 19230
rect 6920 19168 6972 19174
rect 7116 19156 7144 19246
rect 6920 19110 6972 19116
rect 7024 19128 7144 19156
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 7024 17610 7052 19128
rect 7392 17746 7420 19246
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7472 17740 7524 17746
rect 7472 17682 7524 17688
rect 7012 17604 7064 17610
rect 7012 17546 7064 17552
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6656 15026 6684 17138
rect 6748 16590 6776 17478
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6932 16726 6960 16934
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6840 15162 6868 16594
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6656 13326 6684 14962
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 7024 12918 7052 17546
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7300 17134 7328 17478
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 7484 16794 7512 17682
rect 7576 17202 7604 25214
rect 7668 24682 7696 27610
rect 7760 25838 7788 27814
rect 8036 26568 8064 35498
rect 8116 33312 8168 33318
rect 8116 33254 8168 33260
rect 8128 32570 8156 33254
rect 8668 32972 8720 32978
rect 8668 32914 8720 32920
rect 8484 32836 8536 32842
rect 8484 32778 8536 32784
rect 8116 32564 8168 32570
rect 8116 32506 8168 32512
rect 8128 31958 8156 32506
rect 8300 32360 8352 32366
rect 8300 32302 8352 32308
rect 8116 31952 8168 31958
rect 8116 31894 8168 31900
rect 8312 31890 8340 32302
rect 8300 31884 8352 31890
rect 8300 31826 8352 31832
rect 8300 31680 8352 31686
rect 8300 31622 8352 31628
rect 8312 30802 8340 31622
rect 8300 30796 8352 30802
rect 8300 30738 8352 30744
rect 8392 29504 8444 29510
rect 8392 29446 8444 29452
rect 8404 29102 8432 29446
rect 8496 29152 8524 32778
rect 8680 32026 8708 32914
rect 8760 32904 8812 32910
rect 8760 32846 8812 32852
rect 8772 32230 8800 32846
rect 8760 32224 8812 32230
rect 8760 32166 8812 32172
rect 8668 32020 8720 32026
rect 8668 31962 8720 31968
rect 8760 31884 8812 31890
rect 8760 31826 8812 31832
rect 8576 31748 8628 31754
rect 8576 31690 8628 31696
rect 8588 31482 8616 31690
rect 8576 31476 8628 31482
rect 8576 31418 8628 31424
rect 8668 31476 8720 31482
rect 8668 31418 8720 31424
rect 8680 30870 8708 31418
rect 8668 30864 8720 30870
rect 8668 30806 8720 30812
rect 8496 29124 8616 29152
rect 8392 29096 8444 29102
rect 8444 29056 8524 29084
rect 8392 29038 8444 29044
rect 8300 28620 8352 28626
rect 8300 28562 8352 28568
rect 8208 27872 8260 27878
rect 8208 27814 8260 27820
rect 8220 27538 8248 27814
rect 8312 27674 8340 28562
rect 8300 27668 8352 27674
rect 8300 27610 8352 27616
rect 8496 27606 8524 29056
rect 8588 28558 8616 29124
rect 8576 28552 8628 28558
rect 8576 28494 8628 28500
rect 8484 27600 8536 27606
rect 8484 27542 8536 27548
rect 8208 27532 8260 27538
rect 8208 27474 8260 27480
rect 7944 26540 8064 26568
rect 7748 25832 7800 25838
rect 7748 25774 7800 25780
rect 7760 25344 7788 25774
rect 7840 25356 7892 25362
rect 7760 25316 7840 25344
rect 7840 25298 7892 25304
rect 7656 24676 7708 24682
rect 7656 24618 7708 24624
rect 7944 22094 7972 26540
rect 8024 26444 8076 26450
rect 8024 26386 8076 26392
rect 8036 25498 8064 26386
rect 8116 26376 8168 26382
rect 8116 26318 8168 26324
rect 8128 25498 8156 26318
rect 8300 25832 8352 25838
rect 8300 25774 8352 25780
rect 8024 25492 8076 25498
rect 8024 25434 8076 25440
rect 8116 25492 8168 25498
rect 8116 25434 8168 25440
rect 8312 25294 8340 25774
rect 8300 25288 8352 25294
rect 8300 25230 8352 25236
rect 8116 23180 8168 23186
rect 8116 23122 8168 23128
rect 8128 22234 8156 23122
rect 8116 22228 8168 22234
rect 8116 22170 8168 22176
rect 7944 22066 8064 22094
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7668 19514 7696 20402
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7392 14657 7420 14758
rect 7378 14648 7434 14657
rect 7378 14583 7434 14592
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7116 13870 7144 14418
rect 7196 14000 7248 14006
rect 7196 13942 7248 13948
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 7208 12866 7236 13942
rect 7208 12838 7420 12866
rect 7208 12782 7236 12838
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 7300 12306 7328 12650
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7392 12238 7420 12838
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7484 12238 7512 12718
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7300 11014 7328 12038
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 6828 9444 6880 9450
rect 6828 9386 6880 9392
rect 6840 9178 6868 9386
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6932 9042 6960 9318
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6840 7546 6868 7890
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6380 5166 6408 5850
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6564 5642 6592 5714
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6092 4548 6144 4554
rect 6092 4490 6144 4496
rect 6104 4282 6132 4490
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6196 2990 6224 3878
rect 6288 3602 6316 4966
rect 6472 4010 6500 5102
rect 6656 4146 6684 7278
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6748 6118 6776 7142
rect 6932 6866 6960 8978
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6656 3126 6684 4082
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 5908 1964 5960 1970
rect 5908 1906 5960 1912
rect 6104 800 6132 2450
rect 6840 2038 6868 5714
rect 6932 5234 6960 6802
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6932 3058 6960 5170
rect 7024 4010 7052 5510
rect 7116 4622 7144 10134
rect 7300 10130 7328 10950
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 9178 7236 9318
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7208 6118 7236 7142
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7208 5846 7236 6054
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7300 4690 7328 10066
rect 7392 9518 7420 12174
rect 7484 12102 7512 12174
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7484 11218 7512 11766
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7484 9994 7512 11154
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7484 9178 7512 9590
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7576 8974 7604 17138
rect 7656 13388 7708 13394
rect 7840 13388 7892 13394
rect 7656 13330 7708 13336
rect 7760 13348 7840 13376
rect 7668 11898 7696 13330
rect 7760 12102 7788 13348
rect 7840 13330 7892 13336
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7668 11014 7696 11562
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 10010 7696 10950
rect 7852 10130 7880 12718
rect 7944 11830 7972 13262
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7668 9982 7788 10010
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7668 9586 7696 9862
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7392 7206 7420 7686
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 7392 3738 7420 4422
rect 7576 4146 7604 8910
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7484 3738 7512 4014
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7576 3534 7604 4082
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 6932 2854 6960 2994
rect 7116 2990 7144 3334
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 7576 2854 7604 2926
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 6828 2032 6880 2038
rect 6828 1974 6880 1980
rect 7484 800 7512 2450
rect 7668 1902 7696 5714
rect 7760 3602 7788 9982
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7852 8838 7880 8910
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7852 6254 7880 8774
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7944 7546 7972 7890
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7760 2854 7788 3538
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 8036 2774 8064 22066
rect 8312 19990 8340 25230
rect 8484 23724 8536 23730
rect 8484 23666 8536 23672
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 8404 23322 8432 23462
rect 8392 23316 8444 23322
rect 8392 23258 8444 23264
rect 8496 22778 8524 23666
rect 8588 23594 8616 28494
rect 8772 28098 8800 31826
rect 8956 31754 8984 47058
rect 9416 46714 9444 47058
rect 9600 46714 9628 47126
rect 9404 46708 9456 46714
rect 9404 46650 9456 46656
rect 9588 46708 9640 46714
rect 9588 46650 9640 46656
rect 9692 46186 9720 51206
rect 9784 50522 9812 51886
rect 9864 51468 9916 51474
rect 9864 51410 9916 51416
rect 9772 50516 9824 50522
rect 9772 50458 9824 50464
rect 9876 50386 9904 51410
rect 9864 50380 9916 50386
rect 9864 50322 9916 50328
rect 9864 49292 9916 49298
rect 9864 49234 9916 49240
rect 9876 48210 9904 49234
rect 9864 48204 9916 48210
rect 9864 48146 9916 48152
rect 9876 47598 9904 48146
rect 9864 47592 9916 47598
rect 9784 47540 9864 47546
rect 9784 47534 9916 47540
rect 9784 47518 9904 47534
rect 9784 46986 9812 47518
rect 9864 47456 9916 47462
rect 9864 47398 9916 47404
rect 9876 47190 9904 47398
rect 9864 47184 9916 47190
rect 9864 47126 9916 47132
rect 9772 46980 9824 46986
rect 9772 46922 9824 46928
rect 9692 46158 9904 46186
rect 9312 45416 9364 45422
rect 9312 45358 9364 45364
rect 9324 44742 9352 45358
rect 9496 45280 9548 45286
rect 9496 45222 9548 45228
rect 9508 44946 9536 45222
rect 9496 44940 9548 44946
rect 9496 44882 9548 44888
rect 9680 44940 9732 44946
rect 9680 44882 9732 44888
rect 9312 44736 9364 44742
rect 9312 44678 9364 44684
rect 9220 43784 9272 43790
rect 9220 43726 9272 43732
rect 9036 43648 9088 43654
rect 9232 43636 9260 43726
rect 9088 43608 9260 43636
rect 9036 43590 9088 43596
rect 9232 41177 9260 43608
rect 9324 43110 9352 44678
rect 9692 44470 9720 44882
rect 9772 44736 9824 44742
rect 9772 44678 9824 44684
rect 9680 44464 9732 44470
rect 9680 44406 9732 44412
rect 9784 44402 9812 44678
rect 9772 44396 9824 44402
rect 9772 44338 9824 44344
rect 9404 44328 9456 44334
rect 9404 44270 9456 44276
rect 9312 43104 9364 43110
rect 9312 43046 9364 43052
rect 9324 41682 9352 43046
rect 9416 42702 9444 44270
rect 9772 44192 9824 44198
rect 9772 44134 9824 44140
rect 9784 43926 9812 44134
rect 9772 43920 9824 43926
rect 9772 43862 9824 43868
rect 9496 43240 9548 43246
rect 9496 43182 9548 43188
rect 9508 42770 9536 43182
rect 9496 42764 9548 42770
rect 9496 42706 9548 42712
rect 9404 42696 9456 42702
rect 9404 42638 9456 42644
rect 9416 42158 9444 42638
rect 9404 42152 9456 42158
rect 9404 42094 9456 42100
rect 9312 41676 9364 41682
rect 9312 41618 9364 41624
rect 9508 41478 9536 42706
rect 9680 42220 9732 42226
rect 9680 42162 9732 42168
rect 9692 41818 9720 42162
rect 9772 42016 9824 42022
rect 9772 41958 9824 41964
rect 9680 41812 9732 41818
rect 9680 41754 9732 41760
rect 9588 41676 9640 41682
rect 9588 41618 9640 41624
rect 9496 41472 9548 41478
rect 9496 41414 9548 41420
rect 9218 41168 9274 41177
rect 9218 41103 9220 41112
rect 9272 41103 9274 41112
rect 9220 41074 9272 41080
rect 9232 41043 9260 41074
rect 9496 40384 9548 40390
rect 9496 40326 9548 40332
rect 9220 39500 9272 39506
rect 9220 39442 9272 39448
rect 9232 38350 9260 39442
rect 9312 39364 9364 39370
rect 9312 39306 9364 39312
rect 9036 38344 9088 38350
rect 9036 38286 9088 38292
rect 9220 38344 9272 38350
rect 9220 38286 9272 38292
rect 9048 36854 9076 38286
rect 9232 38185 9260 38286
rect 9218 38176 9274 38185
rect 9218 38111 9274 38120
rect 9036 36848 9088 36854
rect 9036 36790 9088 36796
rect 9128 36236 9180 36242
rect 9128 36178 9180 36184
rect 9140 35562 9168 36178
rect 9128 35556 9180 35562
rect 9128 35498 9180 35504
rect 9128 33516 9180 33522
rect 9128 33458 9180 33464
rect 8680 28070 8800 28098
rect 8864 31726 8984 31754
rect 8680 27538 8708 28070
rect 8760 28008 8812 28014
rect 8760 27950 8812 27956
rect 8668 27532 8720 27538
rect 8668 27474 8720 27480
rect 8576 23588 8628 23594
rect 8576 23530 8628 23536
rect 8484 22772 8536 22778
rect 8484 22714 8536 22720
rect 8680 22642 8708 27474
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8300 19984 8352 19990
rect 8300 19926 8352 19932
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 8128 12442 8156 19858
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8312 16998 8340 18022
rect 8404 17218 8432 22510
rect 8484 22500 8536 22506
rect 8484 22442 8536 22448
rect 8496 22166 8524 22442
rect 8588 22234 8616 22510
rect 8576 22228 8628 22234
rect 8576 22170 8628 22176
rect 8484 22160 8536 22166
rect 8484 22102 8536 22108
rect 8668 22024 8720 22030
rect 8668 21966 8720 21972
rect 8680 21486 8708 21966
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8496 20398 8524 20742
rect 8484 20392 8536 20398
rect 8484 20334 8536 20340
rect 8496 17542 8524 20334
rect 8668 19984 8720 19990
rect 8668 19926 8720 19932
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8588 17814 8616 18566
rect 8680 17814 8708 19926
rect 8772 18222 8800 27950
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8864 17882 8892 31726
rect 8944 30660 8996 30666
rect 8944 30602 8996 30608
rect 8956 25378 8984 30602
rect 9140 29782 9168 33458
rect 9220 31884 9272 31890
rect 9220 31826 9272 31832
rect 9128 29776 9180 29782
rect 9128 29718 9180 29724
rect 9140 29170 9168 29718
rect 9128 29164 9180 29170
rect 9128 29106 9180 29112
rect 9232 27946 9260 31826
rect 9220 27940 9272 27946
rect 9220 27882 9272 27888
rect 9036 26444 9088 26450
rect 9036 26386 9088 26392
rect 9048 25498 9076 26386
rect 9036 25492 9088 25498
rect 9036 25434 9088 25440
rect 8956 25350 9076 25378
rect 8944 23044 8996 23050
rect 8944 22986 8996 22992
rect 8956 20806 8984 22986
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 9048 19990 9076 25350
rect 9220 25356 9272 25362
rect 9220 25298 9272 25304
rect 9232 24818 9260 25298
rect 9220 24812 9272 24818
rect 9220 24754 9272 24760
rect 9128 23588 9180 23594
rect 9128 23530 9180 23536
rect 9140 22094 9168 23530
rect 9220 22976 9272 22982
rect 9220 22918 9272 22924
rect 9232 22506 9260 22918
rect 9220 22500 9272 22506
rect 9220 22442 9272 22448
rect 9140 22066 9260 22094
rect 9036 19984 9088 19990
rect 9036 19926 9088 19932
rect 9232 19922 9260 22066
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 9140 18970 9168 19858
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 9232 18850 9260 19858
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 9140 18822 9260 18850
rect 8956 17882 8984 18770
rect 9036 18760 9088 18766
rect 9036 18702 9088 18708
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8944 17876 8996 17882
rect 8944 17818 8996 17824
rect 8576 17808 8628 17814
rect 8576 17750 8628 17756
rect 8668 17808 8720 17814
rect 8668 17750 8720 17756
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8404 17190 8616 17218
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8312 16794 8340 16934
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8220 13394 8248 13874
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 8220 12850 8248 13194
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 8220 12306 8248 12786
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8128 11694 8156 12038
rect 8220 11762 8248 12038
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8220 11218 8248 11698
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8220 10198 8248 11154
rect 8312 10538 8340 15438
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8496 11694 8524 13262
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8496 11354 8524 11494
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8312 9042 8340 10474
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8588 8922 8616 17190
rect 9048 13462 9076 18702
rect 9140 14906 9168 18822
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9232 18358 9260 18702
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 9140 14878 9260 14906
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9140 14278 9168 14758
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9036 13456 9088 13462
rect 9036 13398 9088 13404
rect 9048 10130 9076 13398
rect 9140 13394 9168 14214
rect 9232 13802 9260 14878
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9140 11898 9168 12038
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9232 10266 9260 12242
rect 9324 11558 9352 39306
rect 9508 38486 9536 40326
rect 9600 40050 9628 41618
rect 9784 41070 9812 41958
rect 9876 41682 9904 46158
rect 9864 41676 9916 41682
rect 9864 41618 9916 41624
rect 9864 41540 9916 41546
rect 9864 41482 9916 41488
rect 9772 41064 9824 41070
rect 9772 41006 9824 41012
rect 9876 40934 9904 41482
rect 9864 40928 9916 40934
rect 9864 40870 9916 40876
rect 9772 40452 9824 40458
rect 9772 40394 9824 40400
rect 9588 40044 9640 40050
rect 9588 39986 9640 39992
rect 9680 39296 9732 39302
rect 9784 39284 9812 40394
rect 9876 40372 9904 40870
rect 9968 40526 9996 52906
rect 11520 52896 11572 52902
rect 11520 52838 11572 52844
rect 10220 52796 10516 52816
rect 10276 52794 10300 52796
rect 10356 52794 10380 52796
rect 10436 52794 10460 52796
rect 10298 52742 10300 52794
rect 10362 52742 10374 52794
rect 10436 52742 10438 52794
rect 10276 52740 10300 52742
rect 10356 52740 10380 52742
rect 10436 52740 10460 52742
rect 10220 52720 10516 52740
rect 10600 52080 10652 52086
rect 10600 52022 10652 52028
rect 10220 51708 10516 51728
rect 10276 51706 10300 51708
rect 10356 51706 10380 51708
rect 10436 51706 10460 51708
rect 10298 51654 10300 51706
rect 10362 51654 10374 51706
rect 10436 51654 10438 51706
rect 10276 51652 10300 51654
rect 10356 51652 10380 51654
rect 10436 51652 10460 51654
rect 10220 51632 10516 51652
rect 10612 51610 10640 52022
rect 11244 51876 11296 51882
rect 11244 51818 11296 51824
rect 10784 51808 10836 51814
rect 10784 51750 10836 51756
rect 10796 51610 10824 51750
rect 10600 51604 10652 51610
rect 10600 51546 10652 51552
rect 10784 51604 10836 51610
rect 10784 51546 10836 51552
rect 10784 51468 10836 51474
rect 10784 51410 10836 51416
rect 10796 51377 10824 51410
rect 10968 51400 11020 51406
rect 10782 51368 10838 51377
rect 10968 51342 11020 51348
rect 10782 51303 10838 51312
rect 10220 50620 10516 50640
rect 10276 50618 10300 50620
rect 10356 50618 10380 50620
rect 10436 50618 10460 50620
rect 10298 50566 10300 50618
rect 10362 50566 10374 50618
rect 10436 50566 10438 50618
rect 10276 50564 10300 50566
rect 10356 50564 10380 50566
rect 10436 50564 10460 50566
rect 10220 50544 10516 50564
rect 10220 49532 10516 49552
rect 10276 49530 10300 49532
rect 10356 49530 10380 49532
rect 10436 49530 10460 49532
rect 10298 49478 10300 49530
rect 10362 49478 10374 49530
rect 10436 49478 10438 49530
rect 10276 49476 10300 49478
rect 10356 49476 10380 49478
rect 10436 49476 10460 49478
rect 10220 49456 10516 49476
rect 10692 49224 10744 49230
rect 10692 49166 10744 49172
rect 10048 49088 10100 49094
rect 10048 49030 10100 49036
rect 10060 48142 10088 49030
rect 10600 48816 10652 48822
rect 10600 48758 10652 48764
rect 10140 48680 10192 48686
rect 10140 48622 10192 48628
rect 10152 48346 10180 48622
rect 10220 48444 10516 48464
rect 10276 48442 10300 48444
rect 10356 48442 10380 48444
rect 10436 48442 10460 48444
rect 10298 48390 10300 48442
rect 10362 48390 10374 48442
rect 10436 48390 10438 48442
rect 10276 48388 10300 48390
rect 10356 48388 10380 48390
rect 10436 48388 10460 48390
rect 10220 48368 10516 48388
rect 10140 48340 10192 48346
rect 10140 48282 10192 48288
rect 10048 48136 10100 48142
rect 10048 48078 10100 48084
rect 10140 47456 10192 47462
rect 10140 47398 10192 47404
rect 10152 47122 10180 47398
rect 10220 47356 10516 47376
rect 10276 47354 10300 47356
rect 10356 47354 10380 47356
rect 10436 47354 10460 47356
rect 10298 47302 10300 47354
rect 10362 47302 10374 47354
rect 10436 47302 10438 47354
rect 10276 47300 10300 47302
rect 10356 47300 10380 47302
rect 10436 47300 10460 47302
rect 10220 47280 10516 47300
rect 10612 47190 10640 48758
rect 10704 48686 10732 49166
rect 10692 48680 10744 48686
rect 10692 48622 10744 48628
rect 10600 47184 10652 47190
rect 10600 47126 10652 47132
rect 10140 47116 10192 47122
rect 10140 47058 10192 47064
rect 10508 47116 10560 47122
rect 10508 47058 10560 47064
rect 10520 46578 10548 47058
rect 10508 46572 10560 46578
rect 10508 46514 10560 46520
rect 10048 46368 10100 46374
rect 10048 46310 10100 46316
rect 10060 46170 10088 46310
rect 10220 46268 10516 46288
rect 10276 46266 10300 46268
rect 10356 46266 10380 46268
rect 10436 46266 10460 46268
rect 10298 46214 10300 46266
rect 10362 46214 10374 46266
rect 10436 46214 10438 46266
rect 10276 46212 10300 46214
rect 10356 46212 10380 46214
rect 10436 46212 10460 46214
rect 10220 46192 10516 46212
rect 10048 46164 10100 46170
rect 10048 46106 10100 46112
rect 10612 46034 10640 47126
rect 10600 46028 10652 46034
rect 10600 45970 10652 45976
rect 10704 45914 10732 48622
rect 10796 46578 10824 51303
rect 10980 50930 11008 51342
rect 11256 51074 11284 51818
rect 11256 51046 11376 51074
rect 11348 50998 11376 51046
rect 11336 50992 11388 50998
rect 11336 50934 11388 50940
rect 10968 50924 11020 50930
rect 10968 50866 11020 50872
rect 11060 50176 11112 50182
rect 11060 50118 11112 50124
rect 11072 49298 11100 50118
rect 11348 49842 11376 50934
rect 11336 49836 11388 49842
rect 11336 49778 11388 49784
rect 11060 49292 11112 49298
rect 11060 49234 11112 49240
rect 10968 49088 11020 49094
rect 10968 49030 11020 49036
rect 10980 48278 11008 49030
rect 11072 48686 11100 49234
rect 11152 48748 11204 48754
rect 11152 48690 11204 48696
rect 11060 48680 11112 48686
rect 11060 48622 11112 48628
rect 11060 48544 11112 48550
rect 11060 48486 11112 48492
rect 11072 48346 11100 48486
rect 11060 48340 11112 48346
rect 11060 48282 11112 48288
rect 10968 48272 11020 48278
rect 10968 48214 11020 48220
rect 11164 48210 11192 48690
rect 11152 48204 11204 48210
rect 11152 48146 11204 48152
rect 10876 48000 10928 48006
rect 10876 47942 10928 47948
rect 10784 46572 10836 46578
rect 10784 46514 10836 46520
rect 10612 45886 10732 45914
rect 10220 45180 10516 45200
rect 10276 45178 10300 45180
rect 10356 45178 10380 45180
rect 10436 45178 10460 45180
rect 10298 45126 10300 45178
rect 10362 45126 10374 45178
rect 10436 45126 10438 45178
rect 10276 45124 10300 45126
rect 10356 45124 10380 45126
rect 10436 45124 10460 45126
rect 10220 45104 10516 45124
rect 10048 44328 10100 44334
rect 10048 44270 10100 44276
rect 10060 43994 10088 44270
rect 10220 44092 10516 44112
rect 10276 44090 10300 44092
rect 10356 44090 10380 44092
rect 10436 44090 10460 44092
rect 10298 44038 10300 44090
rect 10362 44038 10374 44090
rect 10436 44038 10438 44090
rect 10276 44036 10300 44038
rect 10356 44036 10380 44038
rect 10436 44036 10460 44038
rect 10220 44016 10516 44036
rect 10048 43988 10100 43994
rect 10048 43930 10100 43936
rect 9956 40520 10008 40526
rect 9956 40462 10008 40468
rect 9876 40344 9996 40372
rect 9864 40044 9916 40050
rect 9864 39986 9916 39992
rect 9876 39506 9904 39986
rect 9864 39500 9916 39506
rect 9864 39442 9916 39448
rect 9864 39296 9916 39302
rect 9784 39256 9864 39284
rect 9680 39238 9732 39244
rect 9864 39238 9916 39244
rect 9692 38962 9720 39238
rect 9680 38956 9732 38962
rect 9680 38898 9732 38904
rect 9864 38888 9916 38894
rect 9864 38830 9916 38836
rect 9588 38820 9640 38826
rect 9588 38762 9640 38768
rect 9496 38480 9548 38486
rect 9496 38422 9548 38428
rect 9404 38344 9456 38350
rect 9402 38312 9404 38321
rect 9456 38312 9458 38321
rect 9402 38247 9458 38256
rect 9496 36576 9548 36582
rect 9496 36518 9548 36524
rect 9508 36378 9536 36518
rect 9496 36372 9548 36378
rect 9496 36314 9548 36320
rect 9404 35624 9456 35630
rect 9404 35566 9456 35572
rect 9416 34678 9444 35566
rect 9508 35154 9536 36314
rect 9496 35148 9548 35154
rect 9496 35090 9548 35096
rect 9404 34672 9456 34678
rect 9404 34614 9456 34620
rect 9404 34536 9456 34542
rect 9404 34478 9456 34484
rect 9416 32298 9444 34478
rect 9496 33856 9548 33862
rect 9496 33798 9548 33804
rect 9508 33386 9536 33798
rect 9496 33380 9548 33386
rect 9496 33322 9548 33328
rect 9508 32978 9536 33322
rect 9496 32972 9548 32978
rect 9496 32914 9548 32920
rect 9600 32858 9628 38762
rect 9680 38480 9732 38486
rect 9680 38422 9732 38428
rect 9692 36718 9720 38422
rect 9876 38282 9904 38830
rect 9864 38276 9916 38282
rect 9864 38218 9916 38224
rect 9968 37856 9996 40344
rect 9784 37828 9996 37856
rect 9680 36712 9732 36718
rect 9680 36654 9732 36660
rect 9680 36032 9732 36038
rect 9680 35974 9732 35980
rect 9508 32830 9628 32858
rect 9404 32292 9456 32298
rect 9404 32234 9456 32240
rect 9404 29164 9456 29170
rect 9404 29106 9456 29112
rect 9416 25362 9444 29106
rect 9508 28014 9536 32830
rect 9692 32586 9720 35974
rect 9600 32558 9720 32586
rect 9600 32230 9628 32558
rect 9680 32428 9732 32434
rect 9680 32370 9732 32376
rect 9588 32224 9640 32230
rect 9588 32166 9640 32172
rect 9692 31754 9720 32370
rect 9784 31890 9812 37828
rect 9956 37732 10008 37738
rect 9956 37674 10008 37680
rect 9864 37324 9916 37330
rect 9864 37266 9916 37272
rect 9876 36174 9904 37266
rect 9864 36168 9916 36174
rect 9864 36110 9916 36116
rect 9968 36038 9996 37674
rect 9956 36032 10008 36038
rect 9956 35974 10008 35980
rect 9956 35828 10008 35834
rect 9956 35770 10008 35776
rect 9864 35488 9916 35494
rect 9864 35430 9916 35436
rect 9876 35154 9904 35430
rect 9864 35148 9916 35154
rect 9864 35090 9916 35096
rect 9968 35034 9996 35770
rect 9876 35006 9996 35034
rect 9876 32910 9904 35006
rect 9956 33448 10008 33454
rect 9956 33390 10008 33396
rect 9864 32904 9916 32910
rect 9864 32846 9916 32852
rect 9864 32768 9916 32774
rect 9864 32710 9916 32716
rect 9876 32366 9904 32710
rect 9968 32434 9996 33390
rect 9956 32428 10008 32434
rect 9956 32370 10008 32376
rect 9864 32360 9916 32366
rect 9864 32302 9916 32308
rect 9864 32224 9916 32230
rect 9864 32166 9916 32172
rect 9956 32224 10008 32230
rect 9956 32166 10008 32172
rect 9772 31884 9824 31890
rect 9772 31826 9824 31832
rect 9692 31726 9812 31754
rect 9588 30184 9640 30190
rect 9588 30126 9640 30132
rect 9600 29578 9628 30126
rect 9680 30048 9732 30054
rect 9680 29990 9732 29996
rect 9588 29572 9640 29578
rect 9588 29514 9640 29520
rect 9692 28762 9720 29990
rect 9680 28756 9732 28762
rect 9680 28698 9732 28704
rect 9784 28558 9812 31726
rect 9876 29458 9904 32166
rect 9968 30666 9996 32166
rect 10060 31958 10088 43930
rect 10612 43874 10640 45886
rect 10796 45558 10824 46514
rect 10888 45966 10916 47942
rect 11060 47456 11112 47462
rect 11060 47398 11112 47404
rect 10968 47048 11020 47054
rect 10968 46990 11020 46996
rect 10876 45960 10928 45966
rect 10876 45902 10928 45908
rect 10784 45552 10836 45558
rect 10784 45494 10836 45500
rect 10796 44810 10824 45494
rect 10784 44804 10836 44810
rect 10784 44746 10836 44752
rect 10692 44328 10744 44334
rect 10692 44270 10744 44276
rect 10520 43846 10640 43874
rect 10704 43858 10732 44270
rect 10692 43852 10744 43858
rect 10520 43194 10548 43846
rect 10692 43794 10744 43800
rect 10600 43716 10652 43722
rect 10600 43658 10652 43664
rect 10612 43382 10640 43658
rect 10704 43450 10732 43794
rect 10784 43648 10836 43654
rect 10784 43590 10836 43596
rect 10796 43450 10824 43590
rect 10692 43444 10744 43450
rect 10692 43386 10744 43392
rect 10784 43444 10836 43450
rect 10784 43386 10836 43392
rect 10600 43376 10652 43382
rect 10600 43318 10652 43324
rect 10692 43240 10744 43246
rect 10520 43166 10640 43194
rect 10692 43182 10744 43188
rect 10220 43004 10516 43024
rect 10276 43002 10300 43004
rect 10356 43002 10380 43004
rect 10436 43002 10460 43004
rect 10298 42950 10300 43002
rect 10362 42950 10374 43002
rect 10436 42950 10438 43002
rect 10276 42948 10300 42950
rect 10356 42948 10380 42950
rect 10436 42948 10460 42950
rect 10220 42928 10516 42948
rect 10140 42152 10192 42158
rect 10140 42094 10192 42100
rect 10152 41818 10180 42094
rect 10220 41916 10516 41936
rect 10276 41914 10300 41916
rect 10356 41914 10380 41916
rect 10436 41914 10460 41916
rect 10298 41862 10300 41914
rect 10362 41862 10374 41914
rect 10436 41862 10438 41914
rect 10276 41860 10300 41862
rect 10356 41860 10380 41862
rect 10436 41860 10460 41862
rect 10220 41840 10516 41860
rect 10140 41812 10192 41818
rect 10140 41754 10192 41760
rect 10140 41676 10192 41682
rect 10140 41618 10192 41624
rect 10048 31952 10100 31958
rect 10048 31894 10100 31900
rect 10048 30864 10100 30870
rect 10048 30806 10100 30812
rect 9956 30660 10008 30666
rect 9956 30602 10008 30608
rect 9956 29776 10008 29782
rect 9956 29718 10008 29724
rect 9968 29578 9996 29718
rect 9956 29572 10008 29578
rect 9956 29514 10008 29520
rect 9876 29430 9996 29458
rect 9864 28960 9916 28966
rect 9864 28902 9916 28908
rect 9876 28762 9904 28902
rect 9864 28756 9916 28762
rect 9864 28698 9916 28704
rect 9772 28552 9824 28558
rect 9772 28494 9824 28500
rect 9496 28008 9548 28014
rect 9496 27950 9548 27956
rect 9680 27328 9732 27334
rect 9680 27270 9732 27276
rect 9692 26314 9720 27270
rect 9680 26308 9732 26314
rect 9680 26250 9732 26256
rect 9588 26240 9640 26246
rect 9588 26182 9640 26188
rect 9600 25838 9628 26182
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 9588 25832 9640 25838
rect 9588 25774 9640 25780
rect 9404 25356 9456 25362
rect 9404 25298 9456 25304
rect 9416 22030 9444 25298
rect 9508 23050 9536 25774
rect 9588 23180 9640 23186
rect 9588 23122 9640 23128
rect 9496 23044 9548 23050
rect 9496 22986 9548 22992
rect 9600 22778 9628 23122
rect 9588 22772 9640 22778
rect 9588 22714 9640 22720
rect 9692 22250 9720 26250
rect 9784 23050 9812 28494
rect 9864 28484 9916 28490
rect 9864 28426 9916 28432
rect 9876 26586 9904 28426
rect 9968 27334 9996 29430
rect 9956 27328 10008 27334
rect 9956 27270 10008 27276
rect 9956 27056 10008 27062
rect 9956 26998 10008 27004
rect 9864 26580 9916 26586
rect 9864 26522 9916 26528
rect 9968 26466 9996 26998
rect 9876 26438 9996 26466
rect 9772 23044 9824 23050
rect 9772 22986 9824 22992
rect 9600 22222 9720 22250
rect 9772 22228 9824 22234
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 9416 18766 9444 21966
rect 9600 21026 9628 22222
rect 9772 22170 9824 22176
rect 9680 22160 9732 22166
rect 9680 22102 9732 22108
rect 9692 21146 9720 22102
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9600 21010 9720 21026
rect 9600 21004 9732 21010
rect 9600 20998 9680 21004
rect 9680 20946 9732 20952
rect 9496 19984 9548 19990
rect 9496 19926 9548 19932
rect 9508 19514 9536 19926
rect 9692 19922 9720 20946
rect 9784 20806 9812 22170
rect 9876 21622 9904 26438
rect 9954 26344 10010 26353
rect 9954 26279 10010 26288
rect 9968 24818 9996 26279
rect 9956 24812 10008 24818
rect 9956 24754 10008 24760
rect 10060 22094 10088 30806
rect 10152 27656 10180 41618
rect 10220 40828 10516 40848
rect 10276 40826 10300 40828
rect 10356 40826 10380 40828
rect 10436 40826 10460 40828
rect 10298 40774 10300 40826
rect 10362 40774 10374 40826
rect 10436 40774 10438 40826
rect 10276 40772 10300 40774
rect 10356 40772 10380 40774
rect 10436 40772 10460 40774
rect 10220 40752 10516 40772
rect 10220 39740 10516 39760
rect 10276 39738 10300 39740
rect 10356 39738 10380 39740
rect 10436 39738 10460 39740
rect 10298 39686 10300 39738
rect 10362 39686 10374 39738
rect 10436 39686 10438 39738
rect 10276 39684 10300 39686
rect 10356 39684 10380 39686
rect 10436 39684 10460 39686
rect 10220 39664 10516 39684
rect 10232 39568 10284 39574
rect 10230 39536 10232 39545
rect 10284 39536 10286 39545
rect 10230 39471 10286 39480
rect 10324 39500 10376 39506
rect 10324 39442 10376 39448
rect 10508 39500 10560 39506
rect 10508 39442 10560 39448
rect 10232 39432 10284 39438
rect 10232 39374 10284 39380
rect 10244 38894 10272 39374
rect 10232 38888 10284 38894
rect 10336 38865 10364 39442
rect 10520 39409 10548 39442
rect 10506 39400 10562 39409
rect 10506 39335 10562 39344
rect 10506 38992 10562 39001
rect 10506 38927 10562 38936
rect 10232 38830 10284 38836
rect 10322 38856 10378 38865
rect 10520 38826 10548 38927
rect 10322 38791 10378 38800
rect 10508 38820 10560 38826
rect 10508 38762 10560 38768
rect 10220 38652 10516 38672
rect 10276 38650 10300 38652
rect 10356 38650 10380 38652
rect 10436 38650 10460 38652
rect 10298 38598 10300 38650
rect 10362 38598 10374 38650
rect 10436 38598 10438 38650
rect 10276 38596 10300 38598
rect 10356 38596 10380 38598
rect 10436 38596 10460 38598
rect 10220 38576 10516 38596
rect 10230 38448 10286 38457
rect 10230 38383 10286 38392
rect 10508 38412 10560 38418
rect 10244 37738 10272 38383
rect 10508 38354 10560 38360
rect 10520 38321 10548 38354
rect 10506 38312 10562 38321
rect 10506 38247 10562 38256
rect 10232 37732 10284 37738
rect 10232 37674 10284 37680
rect 10220 37564 10516 37584
rect 10276 37562 10300 37564
rect 10356 37562 10380 37564
rect 10436 37562 10460 37564
rect 10298 37510 10300 37562
rect 10362 37510 10374 37562
rect 10436 37510 10438 37562
rect 10276 37508 10300 37510
rect 10356 37508 10380 37510
rect 10436 37508 10460 37510
rect 10220 37488 10516 37508
rect 10220 36476 10516 36496
rect 10276 36474 10300 36476
rect 10356 36474 10380 36476
rect 10436 36474 10460 36476
rect 10298 36422 10300 36474
rect 10362 36422 10374 36474
rect 10436 36422 10438 36474
rect 10276 36420 10300 36422
rect 10356 36420 10380 36422
rect 10436 36420 10460 36422
rect 10220 36400 10516 36420
rect 10416 36236 10468 36242
rect 10416 36178 10468 36184
rect 10428 35834 10456 36178
rect 10508 36032 10560 36038
rect 10508 35974 10560 35980
rect 10416 35828 10468 35834
rect 10416 35770 10468 35776
rect 10520 35698 10548 35974
rect 10508 35692 10560 35698
rect 10508 35634 10560 35640
rect 10220 35388 10516 35408
rect 10276 35386 10300 35388
rect 10356 35386 10380 35388
rect 10436 35386 10460 35388
rect 10298 35334 10300 35386
rect 10362 35334 10374 35386
rect 10436 35334 10438 35386
rect 10276 35332 10300 35334
rect 10356 35332 10380 35334
rect 10436 35332 10460 35334
rect 10220 35312 10516 35332
rect 10324 35216 10376 35222
rect 10324 35158 10376 35164
rect 10336 34513 10364 35158
rect 10508 35148 10560 35154
rect 10508 35090 10560 35096
rect 10416 35080 10468 35086
rect 10414 35048 10416 35057
rect 10468 35048 10470 35057
rect 10414 34983 10470 34992
rect 10416 34944 10468 34950
rect 10416 34886 10468 34892
rect 10428 34610 10456 34886
rect 10520 34678 10548 35090
rect 10508 34672 10560 34678
rect 10508 34614 10560 34620
rect 10416 34604 10468 34610
rect 10416 34546 10468 34552
rect 10322 34504 10378 34513
rect 10322 34439 10378 34448
rect 10220 34300 10516 34320
rect 10276 34298 10300 34300
rect 10356 34298 10380 34300
rect 10436 34298 10460 34300
rect 10298 34246 10300 34298
rect 10362 34246 10374 34298
rect 10436 34246 10438 34298
rect 10276 34244 10300 34246
rect 10356 34244 10380 34246
rect 10436 34244 10460 34246
rect 10220 34224 10516 34244
rect 10220 33212 10516 33232
rect 10276 33210 10300 33212
rect 10356 33210 10380 33212
rect 10436 33210 10460 33212
rect 10298 33158 10300 33210
rect 10362 33158 10374 33210
rect 10436 33158 10438 33210
rect 10276 33156 10300 33158
rect 10356 33156 10380 33158
rect 10436 33156 10460 33158
rect 10220 33136 10516 33156
rect 10220 32124 10516 32144
rect 10276 32122 10300 32124
rect 10356 32122 10380 32124
rect 10436 32122 10460 32124
rect 10298 32070 10300 32122
rect 10362 32070 10374 32122
rect 10436 32070 10438 32122
rect 10276 32068 10300 32070
rect 10356 32068 10380 32070
rect 10436 32068 10460 32070
rect 10220 32048 10516 32068
rect 10324 31952 10376 31958
rect 10324 31894 10376 31900
rect 10336 31686 10364 31894
rect 10324 31680 10376 31686
rect 10324 31622 10376 31628
rect 10220 31036 10516 31056
rect 10276 31034 10300 31036
rect 10356 31034 10380 31036
rect 10436 31034 10460 31036
rect 10298 30982 10300 31034
rect 10362 30982 10374 31034
rect 10436 30982 10438 31034
rect 10276 30980 10300 30982
rect 10356 30980 10380 30982
rect 10436 30980 10460 30982
rect 10220 30960 10516 30980
rect 10220 29948 10516 29968
rect 10276 29946 10300 29948
rect 10356 29946 10380 29948
rect 10436 29946 10460 29948
rect 10298 29894 10300 29946
rect 10362 29894 10374 29946
rect 10436 29894 10438 29946
rect 10276 29892 10300 29894
rect 10356 29892 10380 29894
rect 10436 29892 10460 29894
rect 10220 29872 10516 29892
rect 10230 29608 10286 29617
rect 10230 29543 10286 29552
rect 10244 29034 10272 29543
rect 10508 29232 10560 29238
rect 10508 29174 10560 29180
rect 10520 29073 10548 29174
rect 10506 29064 10562 29073
rect 10232 29028 10284 29034
rect 10506 28999 10562 29008
rect 10232 28970 10284 28976
rect 10220 28860 10516 28880
rect 10276 28858 10300 28860
rect 10356 28858 10380 28860
rect 10436 28858 10460 28860
rect 10298 28806 10300 28858
rect 10362 28806 10374 28858
rect 10436 28806 10438 28858
rect 10276 28804 10300 28806
rect 10356 28804 10380 28806
rect 10436 28804 10460 28806
rect 10220 28784 10516 28804
rect 10220 27772 10516 27792
rect 10276 27770 10300 27772
rect 10356 27770 10380 27772
rect 10436 27770 10460 27772
rect 10298 27718 10300 27770
rect 10362 27718 10374 27770
rect 10436 27718 10438 27770
rect 10276 27716 10300 27718
rect 10356 27716 10380 27718
rect 10436 27716 10460 27718
rect 10220 27696 10516 27716
rect 10152 27628 10548 27656
rect 10520 26908 10548 27628
rect 10612 27062 10640 43166
rect 10704 40390 10732 43182
rect 10784 42764 10836 42770
rect 10784 42706 10836 42712
rect 10692 40384 10744 40390
rect 10692 40326 10744 40332
rect 10796 40066 10824 42706
rect 10980 40730 11008 46990
rect 11072 46510 11100 47398
rect 11152 46980 11204 46986
rect 11152 46922 11204 46928
rect 11060 46504 11112 46510
rect 11060 46446 11112 46452
rect 11164 45490 11192 46922
rect 11152 45484 11204 45490
rect 11152 45426 11204 45432
rect 11164 44470 11192 45426
rect 11152 44464 11204 44470
rect 11072 44424 11152 44452
rect 11072 43110 11100 44424
rect 11152 44406 11204 44412
rect 11152 43172 11204 43178
rect 11152 43114 11204 43120
rect 11060 43104 11112 43110
rect 11060 43046 11112 43052
rect 11164 42838 11192 43114
rect 11152 42832 11204 42838
rect 11152 42774 11204 42780
rect 11244 42832 11296 42838
rect 11244 42774 11296 42780
rect 11060 42560 11112 42566
rect 11060 42502 11112 42508
rect 10968 40724 11020 40730
rect 10968 40666 11020 40672
rect 10704 40038 10824 40066
rect 10704 38978 10732 40038
rect 10784 39976 10836 39982
rect 10836 39936 11008 39964
rect 10784 39918 10836 39924
rect 10876 39500 10928 39506
rect 10876 39442 10928 39448
rect 10704 38950 10824 38978
rect 10690 38856 10746 38865
rect 10690 38791 10746 38800
rect 10704 32314 10732 38791
rect 10796 38593 10824 38950
rect 10888 38865 10916 39442
rect 10874 38856 10930 38865
rect 10874 38791 10930 38800
rect 10782 38584 10838 38593
rect 10782 38519 10838 38528
rect 10888 38418 10916 38791
rect 10980 38570 11008 39936
rect 11072 39846 11100 42502
rect 11060 39840 11112 39846
rect 11060 39782 11112 39788
rect 11256 39506 11284 42774
rect 11060 39500 11112 39506
rect 11060 39442 11112 39448
rect 11244 39500 11296 39506
rect 11244 39442 11296 39448
rect 11072 38654 11100 39442
rect 11242 39264 11298 39273
rect 11242 39199 11298 39208
rect 11256 38962 11284 39199
rect 11244 38956 11296 38962
rect 11244 38898 11296 38904
rect 11256 38808 11284 38898
rect 11348 38876 11376 49778
rect 11428 46368 11480 46374
rect 11428 46310 11480 46316
rect 11440 45490 11468 46310
rect 11428 45484 11480 45490
rect 11428 45426 11480 45432
rect 11428 39500 11480 39506
rect 11428 39442 11480 39448
rect 11440 39030 11468 39442
rect 11428 39024 11480 39030
rect 11532 39012 11560 52838
rect 11612 52420 11664 52426
rect 11612 52362 11664 52368
rect 11624 52018 11652 52362
rect 11612 52012 11664 52018
rect 11612 51954 11664 51960
rect 11888 51468 11940 51474
rect 11888 51410 11940 51416
rect 11796 50720 11848 50726
rect 11796 50662 11848 50668
rect 11808 50522 11836 50662
rect 11796 50516 11848 50522
rect 11796 50458 11848 50464
rect 11900 49774 11928 51410
rect 12084 51074 12112 52906
rect 12716 52488 12768 52494
rect 12544 52448 12716 52476
rect 12164 51944 12216 51950
rect 12164 51886 12216 51892
rect 12176 51406 12204 51886
rect 12544 51610 12572 52448
rect 12716 52430 12768 52436
rect 12992 52488 13044 52494
rect 12992 52430 13044 52436
rect 12714 51640 12770 51649
rect 12532 51604 12584 51610
rect 12714 51575 12770 51584
rect 12532 51546 12584 51552
rect 12348 51536 12400 51542
rect 12348 51478 12400 51484
rect 12164 51400 12216 51406
rect 12164 51342 12216 51348
rect 12360 51241 12388 51478
rect 12728 51338 12756 51575
rect 13004 51406 13032 52430
rect 12808 51400 12860 51406
rect 12808 51342 12860 51348
rect 12992 51400 13044 51406
rect 13176 51400 13228 51406
rect 12992 51342 13044 51348
rect 13174 51368 13176 51377
rect 13228 51368 13230 51377
rect 12716 51332 12768 51338
rect 12716 51274 12768 51280
rect 12440 51264 12492 51270
rect 12346 51232 12402 51241
rect 12440 51206 12492 51212
rect 12346 51167 12402 51176
rect 12084 51046 12204 51074
rect 11980 50312 12032 50318
rect 11980 50254 12032 50260
rect 11992 49978 12020 50254
rect 11980 49972 12032 49978
rect 11980 49914 12032 49920
rect 11888 49768 11940 49774
rect 11888 49710 11940 49716
rect 11900 49298 11928 49710
rect 11888 49292 11940 49298
rect 11888 49234 11940 49240
rect 11796 46436 11848 46442
rect 11796 46378 11848 46384
rect 11612 46368 11664 46374
rect 11612 46310 11664 46316
rect 11704 46368 11756 46374
rect 11704 46310 11756 46316
rect 11624 46170 11652 46310
rect 11612 46164 11664 46170
rect 11612 46106 11664 46112
rect 11716 45898 11744 46310
rect 11808 46170 11836 46378
rect 11796 46164 11848 46170
rect 11796 46106 11848 46112
rect 11704 45892 11756 45898
rect 11704 45834 11756 45840
rect 11716 45268 11744 45834
rect 11796 45280 11848 45286
rect 11716 45240 11796 45268
rect 11796 45222 11848 45228
rect 11612 43104 11664 43110
rect 11612 43046 11664 43052
rect 11624 42634 11652 43046
rect 11612 42628 11664 42634
rect 11612 42570 11664 42576
rect 11704 39636 11756 39642
rect 11704 39578 11756 39584
rect 11612 39024 11664 39030
rect 11532 38984 11612 39012
rect 11428 38966 11480 38972
rect 11612 38966 11664 38972
rect 11520 38888 11572 38894
rect 11348 38848 11468 38876
rect 11256 38780 11376 38808
rect 11242 38720 11298 38729
rect 11242 38655 11298 38664
rect 11072 38626 11192 38654
rect 10980 38542 11100 38570
rect 10784 38412 10836 38418
rect 10784 38354 10836 38360
rect 10876 38412 10928 38418
rect 10876 38354 10928 38360
rect 10796 32434 10824 38354
rect 11072 38298 11100 38542
rect 10888 38270 11100 38298
rect 10888 37398 10916 38270
rect 11164 38162 11192 38626
rect 11072 38134 11192 38162
rect 10968 37732 11020 37738
rect 10968 37674 11020 37680
rect 10876 37392 10928 37398
rect 10876 37334 10928 37340
rect 10980 36854 11008 37674
rect 10968 36848 11020 36854
rect 10968 36790 11020 36796
rect 10876 36576 10928 36582
rect 10876 36518 10928 36524
rect 10888 36242 10916 36518
rect 10876 36236 10928 36242
rect 10928 36196 11008 36224
rect 10876 36178 10928 36184
rect 10876 36100 10928 36106
rect 10876 36042 10928 36048
rect 10888 35154 10916 36042
rect 10980 35222 11008 36196
rect 11072 35834 11100 38134
rect 11152 37800 11204 37806
rect 11152 37742 11204 37748
rect 11164 37194 11192 37742
rect 11152 37188 11204 37194
rect 11152 37130 11204 37136
rect 11152 36236 11204 36242
rect 11152 36178 11204 36184
rect 11060 35828 11112 35834
rect 11060 35770 11112 35776
rect 11164 35290 11192 36178
rect 11152 35284 11204 35290
rect 11152 35226 11204 35232
rect 10968 35216 11020 35222
rect 10968 35158 11020 35164
rect 10876 35148 10928 35154
rect 10876 35090 10928 35096
rect 11060 35148 11112 35154
rect 11060 35090 11112 35096
rect 10968 34468 11020 34474
rect 10968 34410 11020 34416
rect 10876 34400 10928 34406
rect 10876 34342 10928 34348
rect 10888 33454 10916 34342
rect 10980 34066 11008 34410
rect 11072 34202 11100 35090
rect 11152 34672 11204 34678
rect 11152 34614 11204 34620
rect 11060 34196 11112 34202
rect 11060 34138 11112 34144
rect 11164 34066 11192 34614
rect 10968 34060 11020 34066
rect 10968 34002 11020 34008
rect 11152 34060 11204 34066
rect 11152 34002 11204 34008
rect 10876 33448 10928 33454
rect 10876 33390 10928 33396
rect 10784 32428 10836 32434
rect 10836 32388 10916 32416
rect 10784 32370 10836 32376
rect 10704 32286 10824 32314
rect 10692 32224 10744 32230
rect 10692 32166 10744 32172
rect 10704 31346 10732 32166
rect 10692 31340 10744 31346
rect 10692 31282 10744 31288
rect 10692 30660 10744 30666
rect 10692 30602 10744 30608
rect 10704 28937 10732 30602
rect 10796 29696 10824 32286
rect 10888 31414 10916 32388
rect 10876 31408 10928 31414
rect 10876 31350 10928 31356
rect 10888 31142 10916 31350
rect 10876 31136 10928 31142
rect 10876 31078 10928 31084
rect 10796 29668 10916 29696
rect 10784 29096 10836 29102
rect 10784 29038 10836 29044
rect 10690 28928 10746 28937
rect 10690 28863 10746 28872
rect 10704 28694 10732 28863
rect 10692 28688 10744 28694
rect 10692 28630 10744 28636
rect 10796 28490 10824 29038
rect 10784 28484 10836 28490
rect 10784 28426 10836 28432
rect 10888 27606 10916 29668
rect 10876 27600 10928 27606
rect 10876 27542 10928 27548
rect 10600 27056 10652 27062
rect 10600 26998 10652 27004
rect 10784 26920 10836 26926
rect 10520 26880 10732 26908
rect 10220 26684 10516 26704
rect 10276 26682 10300 26684
rect 10356 26682 10380 26684
rect 10436 26682 10460 26684
rect 10298 26630 10300 26682
rect 10362 26630 10374 26682
rect 10436 26630 10438 26682
rect 10276 26628 10300 26630
rect 10356 26628 10380 26630
rect 10436 26628 10460 26630
rect 10220 26608 10516 26628
rect 10598 26616 10654 26625
rect 10598 26551 10654 26560
rect 10140 26444 10192 26450
rect 10140 26386 10192 26392
rect 10152 25430 10180 26386
rect 10416 26376 10468 26382
rect 10416 26318 10468 26324
rect 10428 26217 10456 26318
rect 10414 26208 10470 26217
rect 10414 26143 10470 26152
rect 10220 25596 10516 25616
rect 10276 25594 10300 25596
rect 10356 25594 10380 25596
rect 10436 25594 10460 25596
rect 10298 25542 10300 25594
rect 10362 25542 10374 25594
rect 10436 25542 10438 25594
rect 10276 25540 10300 25542
rect 10356 25540 10380 25542
rect 10436 25540 10460 25542
rect 10220 25520 10516 25540
rect 10612 25480 10640 26551
rect 10520 25452 10640 25480
rect 10140 25424 10192 25430
rect 10140 25366 10192 25372
rect 10520 24750 10548 25452
rect 10600 25356 10652 25362
rect 10600 25298 10652 25304
rect 10612 24954 10640 25298
rect 10600 24948 10652 24954
rect 10600 24890 10652 24896
rect 10508 24744 10560 24750
rect 10508 24686 10560 24692
rect 10220 24508 10516 24528
rect 10276 24506 10300 24508
rect 10356 24506 10380 24508
rect 10436 24506 10460 24508
rect 10298 24454 10300 24506
rect 10362 24454 10374 24506
rect 10436 24454 10438 24506
rect 10276 24452 10300 24454
rect 10356 24452 10380 24454
rect 10436 24452 10460 24454
rect 10220 24432 10516 24452
rect 10220 23420 10516 23440
rect 10276 23418 10300 23420
rect 10356 23418 10380 23420
rect 10436 23418 10460 23420
rect 10298 23366 10300 23418
rect 10362 23366 10374 23418
rect 10436 23366 10438 23418
rect 10276 23364 10300 23366
rect 10356 23364 10380 23366
rect 10436 23364 10460 23366
rect 10220 23344 10516 23364
rect 10600 23180 10652 23186
rect 10600 23122 10652 23128
rect 10140 22976 10192 22982
rect 10140 22918 10192 22924
rect 9968 22066 10088 22094
rect 9864 21616 9916 21622
rect 9864 21558 9916 21564
rect 9968 21026 9996 22066
rect 9876 20998 9996 21026
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9876 20584 9904 20998
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 9784 20556 9904 20584
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9784 18970 9812 20556
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 9876 19990 9904 20402
rect 9968 20058 9996 20878
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 10060 20398 10088 20742
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9864 19984 9916 19990
rect 9864 19926 9916 19932
rect 10152 19378 10180 22918
rect 10612 22642 10640 23122
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 10220 22332 10516 22352
rect 10276 22330 10300 22332
rect 10356 22330 10380 22332
rect 10436 22330 10460 22332
rect 10298 22278 10300 22330
rect 10362 22278 10374 22330
rect 10436 22278 10438 22330
rect 10276 22276 10300 22278
rect 10356 22276 10380 22278
rect 10436 22276 10460 22278
rect 10220 22256 10516 22276
rect 10612 22234 10640 22578
rect 10600 22228 10652 22234
rect 10600 22170 10652 22176
rect 10232 22092 10284 22098
rect 10232 22034 10284 22040
rect 10244 21690 10272 22034
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10600 21616 10652 21622
rect 10600 21558 10652 21564
rect 10220 21244 10516 21264
rect 10276 21242 10300 21244
rect 10356 21242 10380 21244
rect 10436 21242 10460 21244
rect 10298 21190 10300 21242
rect 10362 21190 10374 21242
rect 10436 21190 10438 21242
rect 10276 21188 10300 21190
rect 10356 21188 10380 21190
rect 10436 21188 10460 21190
rect 10220 21168 10516 21188
rect 10220 20156 10516 20176
rect 10276 20154 10300 20156
rect 10356 20154 10380 20156
rect 10436 20154 10460 20156
rect 10298 20102 10300 20154
rect 10362 20102 10374 20154
rect 10436 20102 10438 20154
rect 10276 20100 10300 20102
rect 10356 20100 10380 20102
rect 10436 20100 10460 20102
rect 10220 20080 10516 20100
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9956 19168 10008 19174
rect 9956 19110 10008 19116
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9416 17066 9444 18158
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 9416 16658 9444 17002
rect 9508 16794 9536 18770
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9600 17134 9628 17818
rect 9876 17338 9904 19110
rect 9968 18970 9996 19110
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 10152 18306 10180 19314
rect 10220 19068 10516 19088
rect 10276 19066 10300 19068
rect 10356 19066 10380 19068
rect 10436 19066 10460 19068
rect 10298 19014 10300 19066
rect 10362 19014 10374 19066
rect 10436 19014 10438 19066
rect 10276 19012 10300 19014
rect 10356 19012 10380 19014
rect 10436 19012 10460 19014
rect 10220 18992 10516 19012
rect 9968 18278 10180 18306
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9496 15564 9548 15570
rect 9496 15506 9548 15512
rect 9508 15162 9536 15506
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9692 14958 9720 15302
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9692 14550 9720 14894
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9968 14414 9996 18278
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 10152 17882 10180 18158
rect 10220 17980 10516 18000
rect 10276 17978 10300 17980
rect 10356 17978 10380 17980
rect 10436 17978 10460 17980
rect 10298 17926 10300 17978
rect 10362 17926 10374 17978
rect 10436 17926 10438 17978
rect 10276 17924 10300 17926
rect 10356 17924 10380 17926
rect 10436 17924 10460 17926
rect 10220 17904 10516 17924
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10220 16892 10516 16912
rect 10276 16890 10300 16892
rect 10356 16890 10380 16892
rect 10436 16890 10460 16892
rect 10298 16838 10300 16890
rect 10362 16838 10374 16890
rect 10436 16838 10438 16890
rect 10276 16836 10300 16838
rect 10356 16836 10380 16838
rect 10436 16836 10460 16838
rect 10220 16816 10516 16836
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 10060 15026 10088 16730
rect 10220 15804 10516 15824
rect 10276 15802 10300 15804
rect 10356 15802 10380 15804
rect 10436 15802 10460 15804
rect 10298 15750 10300 15802
rect 10362 15750 10374 15802
rect 10436 15750 10438 15802
rect 10276 15748 10300 15750
rect 10356 15748 10380 15750
rect 10436 15748 10460 15750
rect 10220 15728 10516 15748
rect 10048 15020 10100 15026
rect 10612 15008 10640 21558
rect 10704 17921 10732 26880
rect 10784 26862 10836 26868
rect 10796 26625 10824 26862
rect 10876 26784 10928 26790
rect 10876 26726 10928 26732
rect 10782 26616 10838 26625
rect 10782 26551 10838 26560
rect 10784 26444 10836 26450
rect 10784 26386 10836 26392
rect 10796 25498 10824 26386
rect 10888 25906 10916 26726
rect 10980 26602 11008 34002
rect 11060 33312 11112 33318
rect 11060 33254 11112 33260
rect 11072 30870 11100 33254
rect 11164 32978 11192 34002
rect 11152 32972 11204 32978
rect 11152 32914 11204 32920
rect 11164 31890 11192 32914
rect 11152 31884 11204 31890
rect 11152 31826 11204 31832
rect 11152 31680 11204 31686
rect 11152 31622 11204 31628
rect 11060 30864 11112 30870
rect 11060 30806 11112 30812
rect 11060 29164 11112 29170
rect 11060 29106 11112 29112
rect 11072 28762 11100 29106
rect 11060 28756 11112 28762
rect 11060 28698 11112 28704
rect 11060 28552 11112 28558
rect 11060 28494 11112 28500
rect 11072 28082 11100 28494
rect 11060 28076 11112 28082
rect 11060 28018 11112 28024
rect 11058 27432 11114 27441
rect 11058 27367 11114 27376
rect 11072 27130 11100 27367
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 10980 26574 11100 26602
rect 10968 26512 11020 26518
rect 10968 26454 11020 26460
rect 10980 26042 11008 26454
rect 10968 26036 11020 26042
rect 10968 25978 11020 25984
rect 11072 25922 11100 26574
rect 11164 26489 11192 31622
rect 11150 26480 11206 26489
rect 11150 26415 11206 26424
rect 11152 26376 11204 26382
rect 11152 26318 11204 26324
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10980 25894 11100 25922
rect 10876 25696 10928 25702
rect 10876 25638 10928 25644
rect 10784 25492 10836 25498
rect 10784 25434 10836 25440
rect 10888 25430 10916 25638
rect 10876 25424 10928 25430
rect 10876 25366 10928 25372
rect 10888 24954 10916 25366
rect 10876 24948 10928 24954
rect 10876 24890 10928 24896
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10796 21554 10824 24754
rect 10876 23180 10928 23186
rect 10876 23122 10928 23128
rect 10888 22710 10916 23122
rect 10876 22704 10928 22710
rect 10876 22646 10928 22652
rect 10876 22568 10928 22574
rect 10876 22510 10928 22516
rect 10888 22234 10916 22510
rect 10876 22228 10928 22234
rect 10876 22170 10928 22176
rect 10980 22166 11008 25894
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 11072 24138 11100 25230
rect 11060 24132 11112 24138
rect 11060 24074 11112 24080
rect 11164 22574 11192 26318
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 11072 21894 11100 21966
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11072 21690 11100 21830
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10796 20992 10824 21082
rect 10968 21004 11020 21010
rect 10796 20964 10968 20992
rect 10690 17912 10746 17921
rect 10690 17847 10692 17856
rect 10744 17847 10746 17856
rect 10692 17818 10744 17824
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10704 15162 10732 15574
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10612 14980 10732 15008
rect 10048 14962 10100 14968
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9496 13796 9548 13802
rect 9496 13738 9548 13744
rect 9508 12434 9536 13738
rect 9416 12406 9536 12434
rect 9416 12238 9444 12406
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9324 10130 9352 11290
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8312 8894 8616 8922
rect 8116 7948 8168 7954
rect 8312 7936 8340 8894
rect 8588 8838 8616 8894
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8168 7908 8340 7936
rect 8116 7890 8168 7896
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 5166 8248 7686
rect 8404 7546 8432 8774
rect 8772 8090 8800 8978
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 9324 8022 9352 8230
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 9416 7886 9444 12174
rect 9600 11898 9628 12310
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9692 11762 9720 14350
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 13870 9904 14214
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9784 13530 9812 13806
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9508 10452 9536 11494
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9600 10588 9628 10950
rect 9692 10690 9720 11698
rect 9876 11218 9904 12242
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9968 11694 9996 12038
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9784 10810 9812 10950
rect 9876 10810 9904 11154
rect 10060 11150 10088 14962
rect 10600 14884 10652 14890
rect 10600 14826 10652 14832
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10152 14618 10180 14758
rect 10220 14716 10516 14736
rect 10276 14714 10300 14716
rect 10356 14714 10380 14716
rect 10436 14714 10460 14716
rect 10298 14662 10300 14714
rect 10362 14662 10374 14714
rect 10436 14662 10438 14714
rect 10276 14660 10300 14662
rect 10356 14660 10380 14662
rect 10436 14660 10460 14662
rect 10220 14640 10516 14660
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10152 13530 10180 14554
rect 10612 14278 10640 14826
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10220 13628 10516 13648
rect 10276 13626 10300 13628
rect 10356 13626 10380 13628
rect 10436 13626 10460 13628
rect 10298 13574 10300 13626
rect 10362 13574 10374 13626
rect 10436 13574 10438 13626
rect 10276 13572 10300 13574
rect 10356 13572 10380 13574
rect 10436 13572 10460 13574
rect 10220 13552 10516 13572
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10612 13394 10640 14214
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10220 12540 10516 12560
rect 10276 12538 10300 12540
rect 10356 12538 10380 12540
rect 10436 12538 10460 12540
rect 10298 12486 10300 12538
rect 10362 12486 10374 12538
rect 10436 12486 10438 12538
rect 10276 12484 10300 12486
rect 10356 12484 10380 12486
rect 10436 12484 10460 12486
rect 10220 12464 10516 12484
rect 10220 11452 10516 11472
rect 10276 11450 10300 11452
rect 10356 11450 10380 11452
rect 10436 11450 10460 11452
rect 10298 11398 10300 11450
rect 10362 11398 10374 11450
rect 10436 11398 10438 11450
rect 10276 11396 10300 11398
rect 10356 11396 10380 11398
rect 10436 11396 10460 11398
rect 10220 11376 10516 11396
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9692 10662 9904 10690
rect 9772 10600 9824 10606
rect 9600 10560 9772 10588
rect 9772 10542 9824 10548
rect 9508 10424 9628 10452
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9508 8566 9536 8910
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9508 8090 9536 8230
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8404 6934 8432 7482
rect 9496 7336 9548 7342
rect 8666 7304 8722 7313
rect 9496 7278 9548 7284
rect 8666 7239 8722 7248
rect 8680 7002 8708 7239
rect 9508 7002 9536 7278
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8404 5166 8432 6870
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8128 4690 8156 4966
rect 8116 4684 8168 4690
rect 8116 4626 8168 4632
rect 8220 4078 8248 5102
rect 8404 4146 8432 5102
rect 9600 5030 9628 10424
rect 9876 9042 9904 10662
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9876 8566 9904 8978
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9692 5778 9720 7686
rect 9876 7546 9904 8230
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9968 7206 9996 8230
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9876 6390 9904 6802
rect 10060 6798 10088 11086
rect 10220 10364 10516 10384
rect 10276 10362 10300 10364
rect 10356 10362 10380 10364
rect 10436 10362 10460 10364
rect 10298 10310 10300 10362
rect 10362 10310 10374 10362
rect 10436 10310 10438 10362
rect 10276 10308 10300 10310
rect 10356 10308 10380 10310
rect 10436 10308 10460 10310
rect 10220 10288 10516 10308
rect 10612 9654 10640 13330
rect 10704 12782 10732 14980
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10704 11354 10732 11562
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10796 9518 10824 20964
rect 10968 20946 11020 20952
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 10980 19514 11008 20810
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10876 19168 10928 19174
rect 10980 19145 11008 19178
rect 10876 19110 10928 19116
rect 10966 19136 11022 19145
rect 10888 18970 10916 19110
rect 10966 19071 11022 19080
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 11072 18766 11100 21490
rect 11164 21078 11192 22510
rect 11256 21486 11284 38655
rect 11348 38321 11376 38780
rect 11440 38729 11468 38848
rect 11518 38856 11520 38865
rect 11572 38856 11574 38865
rect 11716 38826 11744 39578
rect 11518 38791 11574 38800
rect 11704 38820 11756 38826
rect 11704 38762 11756 38768
rect 11612 38752 11664 38758
rect 11426 38720 11482 38729
rect 11612 38694 11664 38700
rect 11426 38655 11482 38664
rect 11520 38480 11572 38486
rect 11520 38422 11572 38428
rect 11428 38344 11480 38350
rect 11334 38312 11390 38321
rect 11428 38286 11480 38292
rect 11334 38247 11390 38256
rect 11336 38208 11388 38214
rect 11336 38150 11388 38156
rect 11348 35086 11376 38150
rect 11336 35080 11388 35086
rect 11336 35022 11388 35028
rect 11348 33318 11376 35022
rect 11336 33312 11388 33318
rect 11336 33254 11388 33260
rect 11336 32768 11388 32774
rect 11336 32710 11388 32716
rect 11348 32366 11376 32710
rect 11336 32360 11388 32366
rect 11336 32302 11388 32308
rect 11336 31816 11388 31822
rect 11336 31758 11388 31764
rect 11348 30870 11376 31758
rect 11336 30864 11388 30870
rect 11336 30806 11388 30812
rect 11348 30666 11376 30806
rect 11336 30660 11388 30666
rect 11336 30602 11388 30608
rect 11336 28960 11388 28966
rect 11334 28928 11336 28937
rect 11388 28928 11390 28937
rect 11334 28863 11390 28872
rect 11336 28620 11388 28626
rect 11336 28562 11388 28568
rect 11348 28218 11376 28562
rect 11336 28212 11388 28218
rect 11336 28154 11388 28160
rect 11440 28150 11468 38286
rect 11532 37670 11560 38422
rect 11624 38185 11652 38694
rect 11610 38176 11666 38185
rect 11610 38111 11666 38120
rect 11624 37874 11652 38111
rect 11612 37868 11664 37874
rect 11612 37810 11664 37816
rect 11520 37664 11572 37670
rect 11520 37606 11572 37612
rect 11532 37330 11560 37606
rect 11520 37324 11572 37330
rect 11520 37266 11572 37272
rect 11520 37188 11572 37194
rect 11520 37130 11572 37136
rect 11532 36038 11560 37130
rect 11612 36372 11664 36378
rect 11612 36314 11664 36320
rect 11624 36242 11652 36314
rect 11612 36236 11664 36242
rect 11612 36178 11664 36184
rect 11520 36032 11572 36038
rect 11520 35974 11572 35980
rect 11532 34542 11560 35974
rect 11612 35692 11664 35698
rect 11612 35634 11664 35640
rect 11624 35494 11652 35634
rect 11704 35624 11756 35630
rect 11704 35566 11756 35572
rect 11716 35494 11744 35566
rect 11612 35488 11664 35494
rect 11612 35430 11664 35436
rect 11704 35488 11756 35494
rect 11704 35430 11756 35436
rect 11520 34536 11572 34542
rect 11520 34478 11572 34484
rect 11532 31278 11560 34478
rect 11520 31272 11572 31278
rect 11520 31214 11572 31220
rect 11520 30660 11572 30666
rect 11520 30602 11572 30608
rect 11428 28144 11480 28150
rect 11428 28086 11480 28092
rect 11336 28076 11388 28082
rect 11336 28018 11388 28024
rect 11348 25974 11376 28018
rect 11428 28008 11480 28014
rect 11428 27950 11480 27956
rect 11336 25968 11388 25974
rect 11336 25910 11388 25916
rect 11348 24886 11376 25910
rect 11336 24880 11388 24886
rect 11336 24822 11388 24828
rect 11336 24608 11388 24614
rect 11336 24550 11388 24556
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 11152 21072 11204 21078
rect 11152 21014 11204 21020
rect 11256 20369 11284 21422
rect 11242 20360 11298 20369
rect 11242 20295 11298 20304
rect 11244 19984 11296 19990
rect 11244 19926 11296 19932
rect 11152 19848 11204 19854
rect 11152 19790 11204 19796
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10888 15026 10916 15846
rect 11072 15638 11100 18158
rect 11164 16998 11192 19790
rect 11256 19718 11284 19926
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11256 17678 11284 18702
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10980 14618 11008 15438
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10980 14074 11008 14418
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10220 9276 10516 9296
rect 10276 9274 10300 9276
rect 10356 9274 10380 9276
rect 10436 9274 10460 9276
rect 10298 9222 10300 9274
rect 10362 9222 10374 9274
rect 10436 9222 10438 9274
rect 10276 9220 10300 9222
rect 10356 9220 10380 9222
rect 10436 9220 10460 9222
rect 10220 9200 10516 9220
rect 11072 8974 11100 9318
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 10152 6934 10180 8774
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 10220 8188 10516 8208
rect 10276 8186 10300 8188
rect 10356 8186 10380 8188
rect 10436 8186 10460 8188
rect 10298 8134 10300 8186
rect 10362 8134 10374 8186
rect 10436 8134 10438 8186
rect 10276 8132 10300 8134
rect 10356 8132 10380 8134
rect 10436 8132 10460 8134
rect 10220 8112 10516 8132
rect 10232 8016 10284 8022
rect 10230 7984 10232 7993
rect 10416 8016 10468 8022
rect 10284 7984 10286 7993
rect 10416 7958 10468 7964
rect 10230 7919 10286 7928
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10336 7290 10364 7822
rect 10428 7546 10456 7958
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10704 7313 10732 7890
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10796 7410 10824 7686
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10690 7304 10746 7313
rect 10336 7262 10640 7290
rect 10220 7100 10516 7120
rect 10276 7098 10300 7100
rect 10356 7098 10380 7100
rect 10436 7098 10460 7100
rect 10298 7046 10300 7098
rect 10362 7046 10374 7098
rect 10436 7046 10438 7098
rect 10276 7044 10300 7046
rect 10356 7044 10380 7046
rect 10436 7044 10460 7046
rect 10220 7024 10516 7044
rect 10612 7002 10640 7262
rect 10690 7239 10746 7248
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10140 6928 10192 6934
rect 10140 6870 10192 6876
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9876 5778 9904 6326
rect 10220 6012 10516 6032
rect 10276 6010 10300 6012
rect 10356 6010 10380 6012
rect 10436 6010 10460 6012
rect 10298 5958 10300 6010
rect 10362 5958 10374 6010
rect 10436 5958 10438 6010
rect 10276 5956 10300 5958
rect 10356 5956 10380 5958
rect 10436 5956 10460 5958
rect 10220 5936 10516 5956
rect 9954 5808 10010 5817
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9864 5772 9916 5778
rect 10704 5794 10732 6734
rect 10704 5778 10824 5794
rect 10704 5772 10836 5778
rect 10704 5766 10784 5772
rect 9954 5743 10010 5752
rect 9864 5714 9916 5720
rect 9692 5234 9720 5714
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9876 5166 9904 5714
rect 9968 5710 9996 5743
rect 10784 5714 10836 5720
rect 10888 5710 10916 8502
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10980 7410 11008 8434
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10980 5914 11008 6258
rect 11164 6254 11192 16934
rect 11256 15026 11284 17614
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11256 12374 11284 13330
rect 11348 12434 11376 24550
rect 11440 22234 11468 27950
rect 11532 24614 11560 30602
rect 11624 28014 11652 35430
rect 11704 29232 11756 29238
rect 11704 29174 11756 29180
rect 11716 29102 11744 29174
rect 11704 29096 11756 29102
rect 11704 29038 11756 29044
rect 11612 28008 11664 28014
rect 11612 27950 11664 27956
rect 11612 27872 11664 27878
rect 11612 27814 11664 27820
rect 11624 27130 11652 27814
rect 11704 27532 11756 27538
rect 11704 27474 11756 27480
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 11612 26988 11664 26994
rect 11612 26930 11664 26936
rect 11624 26897 11652 26930
rect 11610 26888 11666 26897
rect 11610 26823 11666 26832
rect 11716 26738 11744 27474
rect 11624 26710 11744 26738
rect 11520 24608 11572 24614
rect 11520 24550 11572 24556
rect 11520 22500 11572 22506
rect 11520 22442 11572 22448
rect 11428 22228 11480 22234
rect 11428 22170 11480 22176
rect 11440 17134 11468 22170
rect 11532 21554 11560 22442
rect 11624 22098 11652 26710
rect 11704 26580 11756 26586
rect 11704 26522 11756 26528
rect 11716 25838 11744 26522
rect 11704 25832 11756 25838
rect 11704 25774 11756 25780
rect 11704 25696 11756 25702
rect 11704 25638 11756 25644
rect 11716 24274 11744 25638
rect 11704 24268 11756 24274
rect 11704 24210 11756 24216
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11716 23730 11744 24006
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11612 22092 11664 22098
rect 11808 22094 11836 45222
rect 11888 40520 11940 40526
rect 11888 40462 11940 40468
rect 11900 34406 11928 40462
rect 11980 39908 12032 39914
rect 11980 39850 12032 39856
rect 11992 39642 12020 39850
rect 12072 39840 12124 39846
rect 12072 39782 12124 39788
rect 11980 39636 12032 39642
rect 11980 39578 12032 39584
rect 12084 39506 12112 39782
rect 12072 39500 12124 39506
rect 12072 39442 12124 39448
rect 12176 39098 12204 51046
rect 12452 50862 12480 51206
rect 12532 50992 12584 50998
rect 12532 50934 12584 50940
rect 12440 50856 12492 50862
rect 12440 50798 12492 50804
rect 12544 50674 12572 50934
rect 12716 50924 12768 50930
rect 12716 50866 12768 50872
rect 12452 50646 12572 50674
rect 12256 49292 12308 49298
rect 12256 49234 12308 49240
rect 12268 48754 12296 49234
rect 12348 49224 12400 49230
rect 12348 49166 12400 49172
rect 12360 48754 12388 49166
rect 12256 48748 12308 48754
rect 12256 48690 12308 48696
rect 12348 48748 12400 48754
rect 12348 48690 12400 48696
rect 12452 47122 12480 50646
rect 12624 50312 12676 50318
rect 12544 50272 12624 50300
rect 12440 47116 12492 47122
rect 12440 47058 12492 47064
rect 12544 47054 12572 50272
rect 12624 50254 12676 50260
rect 12728 49774 12756 50866
rect 12716 49768 12768 49774
rect 12716 49710 12768 49716
rect 12728 49042 12756 49710
rect 12820 49230 12848 51342
rect 13004 50862 13032 51342
rect 13174 51303 13230 51312
rect 12992 50856 13044 50862
rect 12992 50798 13044 50804
rect 13084 50856 13136 50862
rect 13084 50798 13136 50804
rect 12900 49632 12952 49638
rect 12900 49574 12952 49580
rect 12912 49230 12940 49574
rect 12808 49224 12860 49230
rect 12808 49166 12860 49172
rect 12900 49224 12952 49230
rect 12900 49166 12952 49172
rect 12728 49014 12848 49042
rect 12624 47116 12676 47122
rect 12624 47058 12676 47064
rect 12532 47048 12584 47054
rect 12532 46990 12584 46996
rect 12544 46442 12572 46990
rect 12532 46436 12584 46442
rect 12532 46378 12584 46384
rect 12348 45824 12400 45830
rect 12348 45766 12400 45772
rect 12360 45558 12388 45766
rect 12348 45552 12400 45558
rect 12348 45494 12400 45500
rect 12360 44946 12388 45494
rect 12636 45286 12664 47058
rect 12820 47054 12848 49014
rect 12912 48686 12940 49166
rect 12900 48680 12952 48686
rect 12900 48622 12952 48628
rect 12808 47048 12860 47054
rect 12808 46990 12860 46996
rect 12624 45280 12676 45286
rect 12624 45222 12676 45228
rect 12348 44940 12400 44946
rect 12348 44882 12400 44888
rect 12820 44198 12848 46990
rect 12900 44872 12952 44878
rect 12900 44814 12952 44820
rect 12912 44402 12940 44814
rect 12900 44396 12952 44402
rect 12900 44338 12952 44344
rect 12808 44192 12860 44198
rect 12808 44134 12860 44140
rect 12624 43852 12676 43858
rect 12624 43794 12676 43800
rect 12348 43104 12400 43110
rect 12348 43046 12400 43052
rect 12360 42922 12388 43046
rect 12360 42894 12572 42922
rect 12544 42838 12572 42894
rect 12532 42832 12584 42838
rect 12532 42774 12584 42780
rect 12348 42764 12400 42770
rect 12348 42706 12400 42712
rect 12256 42628 12308 42634
rect 12256 42570 12308 42576
rect 12268 42226 12296 42570
rect 12256 42220 12308 42226
rect 12256 42162 12308 42168
rect 12360 42158 12388 42706
rect 12348 42152 12400 42158
rect 12348 42094 12400 42100
rect 12440 42084 12492 42090
rect 12440 42026 12492 42032
rect 12452 40610 12480 42026
rect 12532 41676 12584 41682
rect 12532 41618 12584 41624
rect 12360 40582 12480 40610
rect 12360 40390 12388 40582
rect 12440 40520 12492 40526
rect 12440 40462 12492 40468
rect 12348 40384 12400 40390
rect 12348 40326 12400 40332
rect 12452 39506 12480 40462
rect 12544 39982 12572 41618
rect 12532 39976 12584 39982
rect 12532 39918 12584 39924
rect 12440 39500 12492 39506
rect 12268 39460 12440 39488
rect 12164 39092 12216 39098
rect 12164 39034 12216 39040
rect 11978 38992 12034 39001
rect 11978 38927 12034 38936
rect 11992 38758 12020 38927
rect 12072 38888 12124 38894
rect 12072 38830 12124 38836
rect 11980 38752 12032 38758
rect 11980 38694 12032 38700
rect 11980 38344 12032 38350
rect 11980 38286 12032 38292
rect 11992 37806 12020 38286
rect 12084 38214 12112 38830
rect 12072 38208 12124 38214
rect 12072 38150 12124 38156
rect 11980 37800 12032 37806
rect 11980 37742 12032 37748
rect 12072 37732 12124 37738
rect 12072 37674 12124 37680
rect 11980 37664 12032 37670
rect 11980 37606 12032 37612
rect 11992 36718 12020 37606
rect 12084 37398 12112 37674
rect 12268 37482 12296 39460
rect 12440 39442 12492 39448
rect 12530 39400 12586 39409
rect 12530 39335 12532 39344
rect 12584 39335 12586 39344
rect 12532 39306 12584 39312
rect 12532 38752 12584 38758
rect 12532 38694 12584 38700
rect 12348 37664 12400 37670
rect 12348 37606 12400 37612
rect 12176 37454 12296 37482
rect 12176 37398 12204 37454
rect 12072 37392 12124 37398
rect 12164 37392 12216 37398
rect 12072 37334 12124 37340
rect 12162 37360 12164 37369
rect 12216 37360 12218 37369
rect 12162 37295 12218 37304
rect 12256 37324 12308 37330
rect 12360 37312 12388 37606
rect 12308 37284 12388 37312
rect 12438 37288 12494 37297
rect 12256 37266 12308 37272
rect 12164 37256 12216 37262
rect 12438 37223 12494 37232
rect 12164 37198 12216 37204
rect 12176 36718 12204 37198
rect 12452 36786 12480 37223
rect 12440 36780 12492 36786
rect 12440 36722 12492 36728
rect 11980 36712 12032 36718
rect 11980 36654 12032 36660
rect 12164 36712 12216 36718
rect 12164 36654 12216 36660
rect 11980 36100 12032 36106
rect 11980 36042 12032 36048
rect 11888 34400 11940 34406
rect 11888 34342 11940 34348
rect 11992 32774 12020 36042
rect 12176 36038 12204 36654
rect 12164 36032 12216 36038
rect 12164 35974 12216 35980
rect 12348 35488 12400 35494
rect 12348 35430 12400 35436
rect 12360 35154 12388 35430
rect 12544 35329 12572 38694
rect 12530 35320 12586 35329
rect 12530 35255 12586 35264
rect 12348 35148 12400 35154
rect 12348 35090 12400 35096
rect 12532 35148 12584 35154
rect 12532 35090 12584 35096
rect 12072 35080 12124 35086
rect 12070 35048 12072 35057
rect 12124 35048 12126 35057
rect 12070 34983 12126 34992
rect 12360 34610 12388 35090
rect 12348 34604 12400 34610
rect 12176 34564 12348 34592
rect 12176 32978 12204 34564
rect 12348 34546 12400 34552
rect 12164 32972 12216 32978
rect 12164 32914 12216 32920
rect 12348 32972 12400 32978
rect 12348 32914 12400 32920
rect 12072 32904 12124 32910
rect 12072 32846 12124 32852
rect 11980 32768 12032 32774
rect 11980 32710 12032 32716
rect 11888 32360 11940 32366
rect 11888 32302 11940 32308
rect 11900 31278 11928 32302
rect 11888 31272 11940 31278
rect 11888 31214 11940 31220
rect 11900 30598 11928 31214
rect 11980 31204 12032 31210
rect 11980 31146 12032 31152
rect 11888 30592 11940 30598
rect 11888 30534 11940 30540
rect 11992 30190 12020 31146
rect 11980 30184 12032 30190
rect 11980 30126 12032 30132
rect 11888 29096 11940 29102
rect 11886 29064 11888 29073
rect 11940 29064 11942 29073
rect 11886 28999 11942 29008
rect 11980 28008 12032 28014
rect 11980 27950 12032 27956
rect 11886 27024 11942 27033
rect 11886 26959 11888 26968
rect 11940 26959 11942 26968
rect 11888 26930 11940 26936
rect 11888 26852 11940 26858
rect 11888 26794 11940 26800
rect 11612 22034 11664 22040
rect 11716 22066 11836 22094
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 11532 18222 11560 21014
rect 11624 20602 11652 21830
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 11624 19718 11652 20538
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11612 19168 11664 19174
rect 11612 19110 11664 19116
rect 11624 18358 11652 19110
rect 11716 18766 11744 22066
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11808 20777 11836 21286
rect 11794 20768 11850 20777
rect 11794 20703 11850 20712
rect 11900 20618 11928 26794
rect 11992 25702 12020 27950
rect 11980 25696 12032 25702
rect 11980 25638 12032 25644
rect 11978 24848 12034 24857
rect 12084 24834 12112 32846
rect 12164 32768 12216 32774
rect 12164 32710 12216 32716
rect 12176 31142 12204 32710
rect 12256 31816 12308 31822
rect 12256 31758 12308 31764
rect 12164 31136 12216 31142
rect 12164 31078 12216 31084
rect 12268 30802 12296 31758
rect 12360 30841 12388 32914
rect 12440 32360 12492 32366
rect 12440 32302 12492 32308
rect 12452 32026 12480 32302
rect 12440 32020 12492 32026
rect 12440 31962 12492 31968
rect 12440 31408 12492 31414
rect 12440 31350 12492 31356
rect 12452 31142 12480 31350
rect 12440 31136 12492 31142
rect 12440 31078 12492 31084
rect 12346 30832 12402 30841
rect 12256 30796 12308 30802
rect 12452 30802 12480 31078
rect 12346 30767 12402 30776
rect 12440 30796 12492 30802
rect 12256 30738 12308 30744
rect 12440 30738 12492 30744
rect 12440 30592 12492 30598
rect 12440 30534 12492 30540
rect 12348 30388 12400 30394
rect 12348 30330 12400 30336
rect 12164 29776 12216 29782
rect 12164 29718 12216 29724
rect 12176 27062 12204 29718
rect 12256 29164 12308 29170
rect 12256 29106 12308 29112
rect 12164 27056 12216 27062
rect 12164 26998 12216 27004
rect 12162 26752 12218 26761
rect 12162 26687 12218 26696
rect 12034 24806 12112 24834
rect 11978 24783 12034 24792
rect 11808 20590 11928 20618
rect 11808 18902 11836 20590
rect 11796 18896 11848 18902
rect 11796 18838 11848 18844
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 11888 18692 11940 18698
rect 11888 18634 11940 18640
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11612 18352 11664 18358
rect 11612 18294 11664 18300
rect 11716 18222 11744 18566
rect 11900 18426 11928 18634
rect 11796 18420 11848 18426
rect 11796 18362 11848 18368
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11808 18057 11836 18362
rect 11886 18320 11942 18329
rect 11886 18255 11942 18264
rect 11794 18048 11850 18057
rect 11794 17983 11850 17992
rect 11900 17542 11928 18255
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11992 17218 12020 24783
rect 12072 24268 12124 24274
rect 12072 24210 12124 24216
rect 12084 23730 12112 24210
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 12084 23526 12112 23666
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 12084 21486 12112 22034
rect 12176 21894 12204 26687
rect 12268 26518 12296 29106
rect 12360 28082 12388 30330
rect 12452 30190 12480 30534
rect 12440 30184 12492 30190
rect 12440 30126 12492 30132
rect 12440 29504 12492 29510
rect 12440 29446 12492 29452
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 12360 27470 12388 28018
rect 12348 27464 12400 27470
rect 12348 27406 12400 27412
rect 12360 26586 12388 27406
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 12256 26512 12308 26518
rect 12256 26454 12308 26460
rect 12268 25974 12296 26454
rect 12348 26036 12400 26042
rect 12348 25978 12400 25984
rect 12256 25968 12308 25974
rect 12256 25910 12308 25916
rect 12254 24848 12310 24857
rect 12254 24783 12256 24792
rect 12308 24783 12310 24792
rect 12256 24754 12308 24760
rect 12256 24676 12308 24682
rect 12256 24618 12308 24624
rect 12268 23322 12296 24618
rect 12360 24070 12388 25978
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12256 23316 12308 23322
rect 12256 23258 12308 23264
rect 12268 22098 12296 23258
rect 12256 22092 12308 22098
rect 12256 22034 12308 22040
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12072 21480 12124 21486
rect 12072 21422 12124 21428
rect 12084 21078 12112 21422
rect 12072 21072 12124 21078
rect 12072 21014 12124 21020
rect 12176 21010 12204 21626
rect 12268 21486 12296 22034
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 12268 21146 12296 21422
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 12176 20346 12204 20946
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 12084 20318 12204 20346
rect 12084 19009 12112 20318
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 12070 19000 12126 19009
rect 12070 18935 12126 18944
rect 12176 18834 12204 20198
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12084 18086 12112 18770
rect 12164 18692 12216 18698
rect 12164 18634 12216 18640
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 11532 17190 12020 17218
rect 11428 17128 11480 17134
rect 11428 17070 11480 17076
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11440 15434 11468 15846
rect 11428 15428 11480 15434
rect 11428 15370 11480 15376
rect 11348 12406 11468 12434
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11256 11762 11284 12038
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11348 11626 11376 12242
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 7002 11376 7142
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 11348 6458 11376 6938
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 8772 4146 8800 4626
rect 9048 4554 9076 4626
rect 9036 4548 9088 4554
rect 9036 4490 9088 4496
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8496 3534 8524 4082
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8680 3466 8708 3878
rect 9048 3602 9076 4490
rect 9876 4146 9904 5102
rect 10612 5098 10640 5646
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10704 5234 10732 5510
rect 10796 5302 10824 5510
rect 10784 5296 10836 5302
rect 10784 5238 10836 5244
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10600 5092 10652 5098
rect 10600 5034 10652 5040
rect 10220 4924 10516 4944
rect 10276 4922 10300 4924
rect 10356 4922 10380 4924
rect 10436 4922 10460 4924
rect 10298 4870 10300 4922
rect 10362 4870 10374 4922
rect 10436 4870 10438 4922
rect 10276 4868 10300 4870
rect 10356 4868 10380 4870
rect 10436 4868 10460 4870
rect 10220 4848 10516 4868
rect 10612 4690 10640 5034
rect 10704 4758 10732 5170
rect 10888 5166 10916 5646
rect 10876 5160 10928 5166
rect 10796 5120 10876 5148
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 10796 4078 10824 5120
rect 10876 5102 10928 5108
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10888 4282 10916 4558
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10980 4214 11008 5714
rect 11072 5370 11100 6122
rect 11256 5846 11284 6394
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10968 4208 11020 4214
rect 10968 4150 11020 4156
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 11440 4010 11468 12406
rect 11532 11694 11560 17190
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11716 13938 11744 14962
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11610 13288 11666 13297
rect 11610 13223 11666 13232
rect 11624 12986 11652 13223
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11610 12336 11666 12345
rect 11610 12271 11666 12280
rect 11624 12238 11652 12271
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11716 11778 11744 13874
rect 11900 13870 11928 17070
rect 12176 16250 12204 18634
rect 12268 17678 12296 20742
rect 12360 20398 12388 21830
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12360 19854 12388 20334
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12176 15722 12204 16186
rect 12084 15694 12204 15722
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11808 11898 11836 12718
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11716 11762 11836 11778
rect 11716 11756 11848 11762
rect 11716 11750 11796 11756
rect 11796 11698 11848 11704
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11808 11150 11836 11698
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11808 9586 11836 11086
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11704 9512 11756 9518
rect 11518 9480 11574 9489
rect 11704 9454 11756 9460
rect 11518 9415 11520 9424
rect 11572 9415 11574 9424
rect 11520 9386 11572 9392
rect 11532 8430 11560 9386
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11624 9178 11652 9318
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11610 8936 11666 8945
rect 11610 8871 11666 8880
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11624 7478 11652 8871
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11624 4146 11652 7278
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11336 4004 11388 4010
rect 11336 3946 11388 3952
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 9588 3936 9640 3942
rect 11348 3913 11376 3946
rect 9588 3878 9640 3884
rect 11334 3904 11390 3913
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 7944 2746 8064 2774
rect 7944 2378 7972 2746
rect 9416 2650 9444 3538
rect 9600 2990 9628 3878
rect 10220 3836 10516 3856
rect 11334 3839 11390 3848
rect 10276 3834 10300 3836
rect 10356 3834 10380 3836
rect 10436 3834 10460 3836
rect 10298 3782 10300 3834
rect 10362 3782 10374 3834
rect 10436 3782 10438 3834
rect 10276 3780 10300 3782
rect 10356 3780 10380 3782
rect 10436 3780 10460 3782
rect 10220 3760 10516 3780
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10060 2990 10088 3674
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 10220 2748 10516 2768
rect 10276 2746 10300 2748
rect 10356 2746 10380 2748
rect 10436 2746 10460 2748
rect 10298 2694 10300 2746
rect 10362 2694 10374 2746
rect 10436 2694 10438 2746
rect 10276 2692 10300 2694
rect 10356 2692 10380 2694
rect 10436 2692 10460 2694
rect 10220 2672 10516 2692
rect 10612 2650 10640 3538
rect 11348 3534 11376 3606
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11440 3466 11468 3946
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11164 3126 11192 3334
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 11164 2514 11192 3062
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 11152 2508 11204 2514
rect 11152 2450 11204 2456
rect 7932 2372 7984 2378
rect 7932 2314 7984 2320
rect 7656 1896 7708 1902
rect 7656 1838 7708 1844
rect 8588 1086 8616 2450
rect 8576 1080 8628 1086
rect 8576 1022 8628 1028
rect 8772 800 8800 2450
rect 10152 800 10180 2450
rect 11532 800 11560 4014
rect 11624 3194 11652 4082
rect 11716 3534 11744 9454
rect 11808 9382 11836 9522
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11900 7698 11928 13806
rect 11992 13462 12020 15574
rect 12084 14006 12112 15694
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12176 15162 12204 15506
rect 12360 15366 12388 18838
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12360 14958 12388 15302
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 12268 13818 12296 14758
rect 12360 14482 12388 14894
rect 12452 14550 12480 29446
rect 12544 28082 12572 35090
rect 12532 28076 12584 28082
rect 12532 28018 12584 28024
rect 12532 27872 12584 27878
rect 12532 27814 12584 27820
rect 12544 26994 12572 27814
rect 12532 26988 12584 26994
rect 12532 26930 12584 26936
rect 12532 26852 12584 26858
rect 12532 26794 12584 26800
rect 12544 26625 12572 26794
rect 12530 26616 12586 26625
rect 12530 26551 12586 26560
rect 12532 26444 12584 26450
rect 12532 26386 12584 26392
rect 12544 25922 12572 26386
rect 12636 26042 12664 43794
rect 12900 43376 12952 43382
rect 12900 43318 12952 43324
rect 12808 41064 12860 41070
rect 12808 41006 12860 41012
rect 12716 40996 12768 41002
rect 12716 40938 12768 40944
rect 12728 40594 12756 40938
rect 12716 40588 12768 40594
rect 12716 40530 12768 40536
rect 12716 40452 12768 40458
rect 12716 40394 12768 40400
rect 12728 39642 12756 40394
rect 12820 40390 12848 41006
rect 12808 40384 12860 40390
rect 12808 40326 12860 40332
rect 12716 39636 12768 39642
rect 12716 39578 12768 39584
rect 12728 37505 12756 39578
rect 12808 39500 12860 39506
rect 12808 39442 12860 39448
rect 12714 37496 12770 37505
rect 12714 37431 12770 37440
rect 12716 37324 12768 37330
rect 12716 37266 12768 37272
rect 12728 34678 12756 37266
rect 12820 35834 12848 39442
rect 12808 35828 12860 35834
rect 12808 35770 12860 35776
rect 12808 35148 12860 35154
rect 12808 35090 12860 35096
rect 12820 34950 12848 35090
rect 12808 34944 12860 34950
rect 12808 34886 12860 34892
rect 12716 34672 12768 34678
rect 12716 34614 12768 34620
rect 12820 34542 12848 34886
rect 12808 34536 12860 34542
rect 12808 34478 12860 34484
rect 12808 33992 12860 33998
rect 12808 33934 12860 33940
rect 12820 33522 12848 33934
rect 12808 33516 12860 33522
rect 12808 33458 12860 33464
rect 12808 33380 12860 33386
rect 12808 33322 12860 33328
rect 12820 32978 12848 33322
rect 12808 32972 12860 32978
rect 12808 32914 12860 32920
rect 12716 32836 12768 32842
rect 12716 32778 12768 32784
rect 12728 31686 12756 32778
rect 12820 32434 12848 32914
rect 12808 32428 12860 32434
rect 12808 32370 12860 32376
rect 12808 31748 12860 31754
rect 12808 31690 12860 31696
rect 12716 31680 12768 31686
rect 12716 31622 12768 31628
rect 12728 31278 12756 31622
rect 12716 31272 12768 31278
rect 12820 31249 12848 31690
rect 12716 31214 12768 31220
rect 12806 31240 12862 31249
rect 12806 31175 12862 31184
rect 12716 31136 12768 31142
rect 12716 31078 12768 31084
rect 12728 30734 12756 31078
rect 12716 30728 12768 30734
rect 12716 30670 12768 30676
rect 12728 29714 12756 30670
rect 12808 30184 12860 30190
rect 12808 30126 12860 30132
rect 12716 29708 12768 29714
rect 12716 29650 12768 29656
rect 12820 28694 12848 30126
rect 12808 28688 12860 28694
rect 12808 28630 12860 28636
rect 12808 28416 12860 28422
rect 12808 28358 12860 28364
rect 12820 28218 12848 28358
rect 12808 28212 12860 28218
rect 12808 28154 12860 28160
rect 12714 27704 12770 27713
rect 12714 27639 12770 27648
rect 12728 26790 12756 27639
rect 12808 27532 12860 27538
rect 12808 27474 12860 27480
rect 12820 27033 12848 27474
rect 12806 27024 12862 27033
rect 12806 26959 12862 26968
rect 12808 26920 12860 26926
rect 12808 26862 12860 26868
rect 12716 26784 12768 26790
rect 12716 26726 12768 26732
rect 12716 26580 12768 26586
rect 12716 26522 12768 26528
rect 12728 26042 12756 26522
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12716 26036 12768 26042
rect 12716 25978 12768 25984
rect 12544 25894 12664 25922
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12544 24154 12572 25434
rect 12636 25226 12664 25894
rect 12716 25696 12768 25702
rect 12716 25638 12768 25644
rect 12624 25220 12676 25226
rect 12624 25162 12676 25168
rect 12728 24886 12756 25638
rect 12716 24880 12768 24886
rect 12716 24822 12768 24828
rect 12716 24744 12768 24750
rect 12716 24686 12768 24692
rect 12728 24274 12756 24686
rect 12716 24268 12768 24274
rect 12716 24210 12768 24216
rect 12544 24126 12664 24154
rect 12636 23186 12664 24126
rect 12716 24132 12768 24138
rect 12716 24074 12768 24080
rect 12624 23180 12676 23186
rect 12624 23122 12676 23128
rect 12728 23066 12756 24074
rect 12636 23038 12756 23066
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 12544 22642 12572 22918
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12530 21720 12586 21729
rect 12530 21655 12532 21664
rect 12584 21655 12586 21664
rect 12532 21626 12584 21632
rect 12532 20868 12584 20874
rect 12532 20810 12584 20816
rect 12544 20534 12572 20810
rect 12532 20528 12584 20534
rect 12532 20470 12584 20476
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12544 18970 12572 19790
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12636 17218 12664 23038
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12728 21010 12756 21830
rect 12716 21004 12768 21010
rect 12716 20946 12768 20952
rect 12716 20868 12768 20874
rect 12716 20810 12768 20816
rect 12728 20398 12756 20810
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12728 17746 12756 18702
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12636 17190 12756 17218
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12544 14600 12572 15030
rect 12544 14572 12664 14600
rect 12440 14544 12492 14550
rect 12492 14492 12572 14498
rect 12440 14486 12572 14492
rect 12348 14476 12400 14482
rect 12452 14470 12572 14486
rect 12348 14418 12400 14424
rect 12268 13790 12480 13818
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 11992 12850 12020 13398
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 12084 11898 12112 12582
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11808 7670 11928 7698
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11808 3194 11836 7670
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11900 2446 11928 6802
rect 11992 3738 12020 11630
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 12084 10266 12112 10474
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12084 9674 12112 10202
rect 12176 10062 12204 13466
rect 12268 12646 12296 13670
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12360 10962 12388 13398
rect 12452 12238 12480 13790
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12268 10934 12388 10962
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12084 9646 12204 9674
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 12084 8634 12112 9386
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 12084 8090 12112 8298
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12176 6458 12204 9646
rect 12268 9586 12296 10934
rect 12544 10554 12572 14470
rect 12636 11830 12664 14572
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 12452 10526 12572 10554
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12360 8362 12388 8570
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 12084 3534 12112 5646
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12176 4146 12204 4626
rect 12268 4185 12296 6190
rect 12254 4176 12310 4185
rect 12164 4140 12216 4146
rect 12254 4111 12310 4120
rect 12164 4082 12216 4088
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 11992 3346 12020 3470
rect 11992 3318 12112 3346
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 11992 2650 12020 2790
rect 12084 2774 12112 3318
rect 12176 3058 12204 4082
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 12084 2746 12204 2774
rect 12176 2650 12204 2746
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12268 2514 12296 3878
rect 12360 3602 12388 6258
rect 12452 4826 12480 10526
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12544 10198 12572 10406
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12636 9926 12664 10542
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12636 9042 12664 9862
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12636 8090 12664 8978
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12530 7984 12586 7993
rect 12530 7919 12532 7928
rect 12584 7919 12586 7928
rect 12532 7890 12584 7896
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12452 2854 12480 3470
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12544 2514 12572 7890
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12636 3126 12664 6870
rect 12728 6254 12756 17190
rect 12820 15008 12848 26862
rect 12912 21434 12940 43318
rect 13004 21593 13032 50798
rect 13096 49774 13124 50798
rect 13084 49768 13136 49774
rect 13084 49710 13136 49716
rect 13096 43382 13124 49710
rect 13176 49292 13228 49298
rect 13176 49234 13228 49240
rect 13188 48686 13216 49234
rect 13176 48680 13228 48686
rect 13176 48622 13228 48628
rect 13188 45830 13216 48622
rect 13280 46730 13308 52906
rect 14096 52556 14148 52562
rect 14096 52498 14148 52504
rect 13820 51876 13872 51882
rect 13820 51818 13872 51824
rect 13636 51808 13688 51814
rect 13636 51750 13688 51756
rect 13648 51474 13676 51750
rect 13636 51468 13688 51474
rect 13636 51410 13688 51416
rect 13832 51074 13860 51818
rect 14108 51406 14136 52498
rect 14096 51400 14148 51406
rect 14096 51342 14148 51348
rect 13912 51264 13964 51270
rect 13910 51232 13912 51241
rect 13964 51232 13966 51241
rect 13910 51167 13966 51176
rect 13740 51046 13860 51074
rect 13740 50862 13768 51046
rect 13728 50856 13780 50862
rect 13728 50798 13780 50804
rect 13636 50176 13688 50182
rect 13636 50118 13688 50124
rect 13648 49774 13676 50118
rect 13636 49768 13688 49774
rect 13636 49710 13688 49716
rect 13912 49632 13964 49638
rect 13912 49574 13964 49580
rect 13924 49298 13952 49574
rect 13544 49292 13596 49298
rect 13544 49234 13596 49240
rect 13912 49292 13964 49298
rect 13912 49234 13964 49240
rect 13556 49094 13584 49234
rect 13924 49162 13952 49234
rect 13912 49156 13964 49162
rect 13912 49098 13964 49104
rect 13360 49088 13412 49094
rect 13360 49030 13412 49036
rect 13544 49088 13596 49094
rect 13544 49030 13596 49036
rect 13372 48822 13400 49030
rect 13360 48816 13412 48822
rect 13360 48758 13412 48764
rect 13924 48686 13952 49098
rect 13912 48680 13964 48686
rect 13912 48622 13964 48628
rect 14108 47122 14136 51342
rect 14188 50720 14240 50726
rect 14188 50662 14240 50668
rect 14280 50720 14332 50726
rect 14280 50662 14332 50668
rect 14200 50522 14228 50662
rect 14292 50522 14320 50662
rect 14188 50516 14240 50522
rect 14188 50458 14240 50464
rect 14280 50516 14332 50522
rect 14280 50458 14332 50464
rect 14096 47116 14148 47122
rect 14096 47058 14148 47064
rect 14108 46986 14136 47058
rect 14188 47048 14240 47054
rect 14188 46990 14240 46996
rect 14096 46980 14148 46986
rect 14096 46922 14148 46928
rect 13728 46912 13780 46918
rect 13728 46854 13780 46860
rect 13280 46702 13400 46730
rect 13268 46640 13320 46646
rect 13268 46582 13320 46588
rect 13280 45830 13308 46582
rect 13176 45824 13228 45830
rect 13176 45766 13228 45772
rect 13268 45824 13320 45830
rect 13268 45766 13320 45772
rect 13280 44334 13308 45766
rect 13268 44328 13320 44334
rect 13268 44270 13320 44276
rect 13268 44192 13320 44198
rect 13268 44134 13320 44140
rect 13084 43376 13136 43382
rect 13084 43318 13136 43324
rect 13176 42560 13228 42566
rect 13176 42502 13228 42508
rect 13188 41750 13216 42502
rect 13176 41744 13228 41750
rect 13176 41686 13228 41692
rect 13280 41002 13308 44134
rect 13268 40996 13320 41002
rect 13268 40938 13320 40944
rect 13084 40588 13136 40594
rect 13084 40530 13136 40536
rect 13096 35290 13124 40530
rect 13176 40384 13228 40390
rect 13176 40326 13228 40332
rect 13084 35284 13136 35290
rect 13084 35226 13136 35232
rect 13084 34468 13136 34474
rect 13084 34410 13136 34416
rect 13096 34066 13124 34410
rect 13084 34060 13136 34066
rect 13084 34002 13136 34008
rect 13084 33448 13136 33454
rect 13084 33390 13136 33396
rect 13096 33046 13124 33390
rect 13084 33040 13136 33046
rect 13084 32982 13136 32988
rect 13188 32892 13216 40326
rect 13280 39982 13308 40938
rect 13268 39976 13320 39982
rect 13268 39918 13320 39924
rect 13268 38412 13320 38418
rect 13268 38354 13320 38360
rect 13280 37398 13308 38354
rect 13372 37942 13400 46702
rect 13740 46578 13768 46854
rect 13728 46572 13780 46578
rect 13728 46514 13780 46520
rect 13544 46504 13596 46510
rect 13544 46446 13596 46452
rect 13556 46102 13584 46446
rect 14200 46374 14228 46990
rect 13636 46368 13688 46374
rect 13636 46310 13688 46316
rect 14188 46368 14240 46374
rect 14188 46310 14240 46316
rect 13544 46096 13596 46102
rect 13544 46038 13596 46044
rect 13544 45960 13596 45966
rect 13544 45902 13596 45908
rect 13556 45422 13584 45902
rect 13648 45626 13676 46310
rect 13728 46096 13780 46102
rect 13728 46038 13780 46044
rect 13636 45620 13688 45626
rect 13636 45562 13688 45568
rect 13740 45422 13768 46038
rect 14200 46034 14228 46310
rect 14188 46028 14240 46034
rect 14188 45970 14240 45976
rect 13544 45416 13596 45422
rect 13544 45358 13596 45364
rect 13728 45416 13780 45422
rect 13728 45358 13780 45364
rect 13556 44878 13584 45358
rect 13544 44872 13596 44878
rect 13544 44814 13596 44820
rect 13556 43926 13584 44814
rect 13740 44402 13768 45358
rect 14096 45348 14148 45354
rect 14096 45290 14148 45296
rect 14108 44878 14136 45290
rect 14096 44872 14148 44878
rect 14096 44814 14148 44820
rect 14200 44690 14228 45970
rect 14280 45484 14332 45490
rect 14280 45426 14332 45432
rect 14292 45286 14320 45426
rect 14280 45280 14332 45286
rect 14280 45222 14332 45228
rect 14108 44662 14228 44690
rect 13728 44396 13780 44402
rect 13728 44338 13780 44344
rect 14108 44334 14136 44662
rect 14292 44554 14320 45222
rect 14200 44526 14320 44554
rect 14096 44328 14148 44334
rect 14096 44270 14148 44276
rect 13544 43920 13596 43926
rect 13544 43862 13596 43868
rect 13636 42696 13688 42702
rect 13636 42638 13688 42644
rect 13728 42696 13780 42702
rect 13728 42638 13780 42644
rect 14004 42696 14056 42702
rect 14004 42638 14056 42644
rect 13648 42294 13676 42638
rect 13636 42288 13688 42294
rect 13636 42230 13688 42236
rect 13648 41682 13676 42230
rect 13636 41676 13688 41682
rect 13636 41618 13688 41624
rect 13544 41608 13596 41614
rect 13544 41550 13596 41556
rect 13452 41200 13504 41206
rect 13452 41142 13504 41148
rect 13464 40118 13492 41142
rect 13452 40112 13504 40118
rect 13452 40054 13504 40060
rect 13464 39273 13492 40054
rect 13450 39264 13506 39273
rect 13450 39199 13506 39208
rect 13556 38214 13584 41550
rect 13648 41138 13676 41618
rect 13636 41132 13688 41138
rect 13636 41074 13688 41080
rect 13740 40594 13768 42638
rect 13820 40724 13872 40730
rect 13820 40666 13872 40672
rect 13728 40588 13780 40594
rect 13728 40530 13780 40536
rect 13636 39976 13688 39982
rect 13636 39918 13688 39924
rect 13648 39302 13676 39918
rect 13728 39908 13780 39914
rect 13728 39850 13780 39856
rect 13740 39438 13768 39850
rect 13832 39506 13860 40666
rect 14016 40050 14044 42638
rect 14004 40044 14056 40050
rect 14004 39986 14056 39992
rect 13912 39976 13964 39982
rect 13912 39918 13964 39924
rect 13820 39500 13872 39506
rect 13820 39442 13872 39448
rect 13728 39432 13780 39438
rect 13728 39374 13780 39380
rect 13636 39296 13688 39302
rect 13636 39238 13688 39244
rect 13544 38208 13596 38214
rect 13544 38150 13596 38156
rect 13360 37936 13412 37942
rect 13360 37878 13412 37884
rect 13360 37800 13412 37806
rect 13360 37742 13412 37748
rect 13268 37392 13320 37398
rect 13268 37334 13320 37340
rect 13268 36712 13320 36718
rect 13268 36654 13320 36660
rect 13096 32864 13216 32892
rect 13096 26858 13124 32864
rect 13280 32774 13308 36654
rect 13372 36582 13400 37742
rect 13452 37664 13504 37670
rect 13452 37606 13504 37612
rect 13464 37466 13492 37606
rect 13452 37460 13504 37466
rect 13452 37402 13504 37408
rect 13450 37360 13506 37369
rect 13450 37295 13452 37304
rect 13504 37295 13506 37304
rect 13452 37266 13504 37272
rect 13648 37274 13676 39238
rect 13740 37806 13768 39374
rect 13728 37800 13780 37806
rect 13728 37742 13780 37748
rect 13820 37664 13872 37670
rect 13820 37606 13872 37612
rect 13726 37496 13782 37505
rect 13832 37466 13860 37606
rect 13726 37431 13782 37440
rect 13820 37460 13872 37466
rect 13740 37398 13768 37431
rect 13820 37402 13872 37408
rect 13728 37392 13780 37398
rect 13728 37334 13780 37340
rect 13820 37286 13872 37292
rect 13648 37246 13768 37274
rect 13740 36854 13768 37246
rect 13820 37228 13872 37234
rect 13728 36848 13780 36854
rect 13728 36790 13780 36796
rect 13360 36576 13412 36582
rect 13360 36518 13412 36524
rect 13372 34678 13400 36518
rect 13740 36174 13768 36790
rect 13728 36168 13780 36174
rect 13728 36110 13780 36116
rect 13636 36100 13688 36106
rect 13636 36042 13688 36048
rect 13544 35760 13596 35766
rect 13544 35702 13596 35708
rect 13648 35714 13676 36042
rect 13832 35834 13860 37228
rect 13820 35828 13872 35834
rect 13820 35770 13872 35776
rect 13556 35630 13584 35702
rect 13648 35686 13860 35714
rect 13544 35624 13596 35630
rect 13544 35566 13596 35572
rect 13452 35148 13504 35154
rect 13452 35090 13504 35096
rect 13360 34672 13412 34678
rect 13360 34614 13412 34620
rect 13464 34134 13492 35090
rect 13556 34950 13584 35566
rect 13636 35556 13688 35562
rect 13636 35498 13688 35504
rect 13544 34944 13596 34950
rect 13544 34886 13596 34892
rect 13544 34536 13596 34542
rect 13544 34478 13596 34484
rect 13452 34128 13504 34134
rect 13452 34070 13504 34076
rect 13452 33992 13504 33998
rect 13452 33934 13504 33940
rect 13360 33448 13412 33454
rect 13360 33390 13412 33396
rect 13372 32978 13400 33390
rect 13360 32972 13412 32978
rect 13360 32914 13412 32920
rect 13268 32768 13320 32774
rect 13268 32710 13320 32716
rect 13268 32428 13320 32434
rect 13268 32370 13320 32376
rect 13280 32026 13308 32370
rect 13464 32298 13492 33934
rect 13556 33862 13584 34478
rect 13544 33856 13596 33862
rect 13544 33798 13596 33804
rect 13544 32496 13596 32502
rect 13544 32438 13596 32444
rect 13452 32292 13504 32298
rect 13452 32234 13504 32240
rect 13268 32020 13320 32026
rect 13268 31962 13320 31968
rect 13176 31272 13228 31278
rect 13176 31214 13228 31220
rect 13188 27538 13216 31214
rect 13280 28014 13308 31962
rect 13556 31906 13584 32438
rect 13464 31890 13584 31906
rect 13464 31884 13596 31890
rect 13464 31878 13544 31884
rect 13464 30274 13492 31878
rect 13544 31826 13596 31832
rect 13542 31784 13598 31793
rect 13542 31719 13598 31728
rect 13372 30246 13492 30274
rect 13268 28008 13320 28014
rect 13268 27950 13320 27956
rect 13176 27532 13228 27538
rect 13176 27474 13228 27480
rect 13174 27024 13230 27033
rect 13174 26959 13230 26968
rect 13084 26852 13136 26858
rect 13084 26794 13136 26800
rect 13082 26616 13138 26625
rect 13082 26551 13138 26560
rect 13096 25770 13124 26551
rect 13188 26081 13216 26959
rect 13280 26586 13308 27950
rect 13268 26580 13320 26586
rect 13268 26522 13320 26528
rect 13268 26444 13320 26450
rect 13268 26386 13320 26392
rect 13174 26072 13230 26081
rect 13174 26007 13230 26016
rect 13280 25888 13308 26386
rect 13372 26246 13400 30246
rect 13452 30184 13504 30190
rect 13452 30126 13504 30132
rect 13464 29510 13492 30126
rect 13452 29504 13504 29510
rect 13452 29446 13504 29452
rect 13452 29096 13504 29102
rect 13452 29038 13504 29044
rect 13464 27878 13492 29038
rect 13452 27872 13504 27878
rect 13452 27814 13504 27820
rect 13452 27532 13504 27538
rect 13452 27474 13504 27480
rect 13360 26240 13412 26246
rect 13360 26182 13412 26188
rect 13360 26036 13412 26042
rect 13360 25978 13412 25984
rect 13188 25860 13308 25888
rect 13084 25764 13136 25770
rect 13084 25706 13136 25712
rect 13188 25650 13216 25860
rect 13268 25764 13320 25770
rect 13268 25706 13320 25712
rect 13096 25622 13216 25650
rect 12990 21584 13046 21593
rect 12990 21519 13046 21528
rect 12912 21406 13032 21434
rect 12900 21344 12952 21350
rect 12900 21286 12952 21292
rect 12912 20942 12940 21286
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12912 20398 12940 20742
rect 12900 20392 12952 20398
rect 12900 20334 12952 20340
rect 13004 18986 13032 21406
rect 12912 18958 13032 18986
rect 12912 17660 12940 18958
rect 13096 18290 13124 25622
rect 13280 25362 13308 25706
rect 13268 25356 13320 25362
rect 13268 25298 13320 25304
rect 13176 25220 13228 25226
rect 13176 25162 13228 25168
rect 13188 24274 13216 25162
rect 13280 24410 13308 25298
rect 13372 24886 13400 25978
rect 13360 24880 13412 24886
rect 13360 24822 13412 24828
rect 13268 24404 13320 24410
rect 13268 24346 13320 24352
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 13360 24268 13412 24274
rect 13360 24210 13412 24216
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 12912 17632 13032 17660
rect 12820 14980 12940 15008
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 12820 12306 12848 14826
rect 12912 13410 12940 14980
rect 13004 13530 13032 17632
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 13096 15910 13124 16526
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13084 15428 13136 15434
rect 13084 15370 13136 15376
rect 13096 14890 13124 15370
rect 13084 14884 13136 14890
rect 13084 14826 13136 14832
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12912 13382 13032 13410
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12820 10588 12848 12242
rect 13004 12186 13032 13382
rect 13096 12306 13124 14486
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 13004 12158 13124 12186
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12912 11354 12940 11630
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13004 10742 13032 11290
rect 12992 10736 13044 10742
rect 12992 10678 13044 10684
rect 12992 10600 13044 10606
rect 12820 10560 12992 10588
rect 12992 10542 13044 10548
rect 12806 10432 12862 10441
rect 12806 10367 12862 10376
rect 12820 6866 12848 10367
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12912 6730 12940 8366
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12728 2582 12756 6190
rect 13004 6118 13032 10542
rect 13096 9042 13124 12158
rect 13188 10713 13216 24210
rect 13372 24138 13400 24210
rect 13360 24132 13412 24138
rect 13360 24074 13412 24080
rect 13268 24064 13320 24070
rect 13268 24006 13320 24012
rect 13280 18698 13308 24006
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 13372 21486 13400 23462
rect 13360 21480 13412 21486
rect 13360 21422 13412 21428
rect 13372 20534 13400 21422
rect 13360 20528 13412 20534
rect 13360 20470 13412 20476
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 13372 19514 13400 20334
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 13268 15904 13320 15910
rect 13372 15892 13400 19246
rect 13320 15864 13400 15892
rect 13268 15846 13320 15852
rect 13280 11694 13308 15846
rect 13360 15088 13412 15094
rect 13360 15030 13412 15036
rect 13372 14482 13400 15030
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13266 11520 13322 11529
rect 13266 11455 13322 11464
rect 13174 10704 13230 10713
rect 13174 10639 13230 10648
rect 13280 9602 13308 11455
rect 13188 9574 13308 9602
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13096 8498 13124 8978
rect 13188 8634 13216 9574
rect 13372 9058 13400 14418
rect 13464 13530 13492 27474
rect 13556 27130 13584 31719
rect 13544 27124 13596 27130
rect 13544 27066 13596 27072
rect 13544 26920 13596 26926
rect 13544 26862 13596 26868
rect 13556 26450 13584 26862
rect 13544 26444 13596 26450
rect 13544 26386 13596 26392
rect 13544 26240 13596 26246
rect 13544 26182 13596 26188
rect 13556 24342 13584 26182
rect 13544 24336 13596 24342
rect 13544 24278 13596 24284
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13556 23526 13584 24142
rect 13544 23520 13596 23526
rect 13544 23462 13596 23468
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 13556 21690 13584 21966
rect 13648 21690 13676 35498
rect 13728 35488 13780 35494
rect 13728 35430 13780 35436
rect 13740 34610 13768 35430
rect 13832 35034 13860 35686
rect 13924 35290 13952 39918
rect 14004 39500 14056 39506
rect 14004 39442 14056 39448
rect 14016 37806 14044 39442
rect 14004 37800 14056 37806
rect 14004 37742 14056 37748
rect 14004 37392 14056 37398
rect 14002 37360 14004 37369
rect 14056 37360 14058 37369
rect 14002 37295 14058 37304
rect 14108 36650 14136 44270
rect 14200 42702 14228 44526
rect 14280 42764 14332 42770
rect 14280 42706 14332 42712
rect 14188 42696 14240 42702
rect 14188 42638 14240 42644
rect 14292 42090 14320 42706
rect 14280 42084 14332 42090
rect 14280 42026 14332 42032
rect 14384 41414 14412 52906
rect 16120 52488 16172 52494
rect 16120 52430 16172 52436
rect 14852 52252 15148 52272
rect 14908 52250 14932 52252
rect 14988 52250 15012 52252
rect 15068 52250 15092 52252
rect 14930 52198 14932 52250
rect 14994 52198 15006 52250
rect 15068 52198 15070 52250
rect 14908 52196 14932 52198
rect 14988 52196 15012 52198
rect 15068 52196 15092 52198
rect 14852 52176 15148 52196
rect 16132 52018 16160 52430
rect 14648 52012 14700 52018
rect 14648 51954 14700 51960
rect 15476 52012 15528 52018
rect 15476 51954 15528 51960
rect 16120 52012 16172 52018
rect 16120 51954 16172 51960
rect 14660 51074 14688 51954
rect 14740 51808 14792 51814
rect 14740 51750 14792 51756
rect 15108 51808 15160 51814
rect 15108 51750 15160 51756
rect 14752 51542 14780 51750
rect 15120 51610 15148 51750
rect 15108 51604 15160 51610
rect 15108 51546 15160 51552
rect 14740 51536 14792 51542
rect 14740 51478 14792 51484
rect 14852 51164 15148 51184
rect 14908 51162 14932 51164
rect 14988 51162 15012 51164
rect 15068 51162 15092 51164
rect 14930 51110 14932 51162
rect 14994 51110 15006 51162
rect 15068 51110 15070 51162
rect 14908 51108 14932 51110
rect 14988 51108 15012 51110
rect 15068 51108 15092 51110
rect 14852 51088 15148 51108
rect 14660 51046 14780 51074
rect 14752 49298 14780 51046
rect 15292 50720 15344 50726
rect 15292 50662 15344 50668
rect 14852 50076 15148 50096
rect 14908 50074 14932 50076
rect 14988 50074 15012 50076
rect 15068 50074 15092 50076
rect 14930 50022 14932 50074
rect 14994 50022 15006 50074
rect 15068 50022 15070 50074
rect 14908 50020 14932 50022
rect 14988 50020 15012 50022
rect 15068 50020 15092 50022
rect 14852 50000 15148 50020
rect 15200 49700 15252 49706
rect 15200 49642 15252 49648
rect 14740 49292 14792 49298
rect 14740 49234 14792 49240
rect 14648 49088 14700 49094
rect 14648 49030 14700 49036
rect 14660 48754 14688 49030
rect 14648 48748 14700 48754
rect 14648 48690 14700 48696
rect 14556 48680 14608 48686
rect 14556 48622 14608 48628
rect 14568 44878 14596 48622
rect 14648 47116 14700 47122
rect 14648 47058 14700 47064
rect 14660 46646 14688 47058
rect 14648 46640 14700 46646
rect 14648 46582 14700 46588
rect 14752 46458 14780 49234
rect 14852 48988 15148 49008
rect 14908 48986 14932 48988
rect 14988 48986 15012 48988
rect 15068 48986 15092 48988
rect 14930 48934 14932 48986
rect 14994 48934 15006 48986
rect 15068 48934 15070 48986
rect 14908 48932 14932 48934
rect 14988 48932 15012 48934
rect 15068 48932 15092 48934
rect 14852 48912 15148 48932
rect 15212 48822 15240 49642
rect 15200 48816 15252 48822
rect 15200 48758 15252 48764
rect 15304 48754 15332 50662
rect 15488 49842 15516 51954
rect 16396 51876 16448 51882
rect 16396 51818 16448 51824
rect 15842 51640 15898 51649
rect 15842 51575 15898 51584
rect 15856 51542 15884 51575
rect 15844 51536 15896 51542
rect 15844 51478 15896 51484
rect 16304 51264 16356 51270
rect 16304 51206 16356 51212
rect 16316 50862 16344 51206
rect 16408 50998 16436 51818
rect 16396 50992 16448 50998
rect 16396 50934 16448 50940
rect 16304 50856 16356 50862
rect 16304 50798 16356 50804
rect 16396 50380 16448 50386
rect 16396 50322 16448 50328
rect 16304 50176 16356 50182
rect 16304 50118 16356 50124
rect 15476 49836 15528 49842
rect 15476 49778 15528 49784
rect 15384 49768 15436 49774
rect 15384 49710 15436 49716
rect 15396 48890 15424 49710
rect 15384 48884 15436 48890
rect 15384 48826 15436 48832
rect 15292 48748 15344 48754
rect 15292 48690 15344 48696
rect 14852 47900 15148 47920
rect 14908 47898 14932 47900
rect 14988 47898 15012 47900
rect 15068 47898 15092 47900
rect 14930 47846 14932 47898
rect 14994 47846 15006 47898
rect 15068 47846 15070 47898
rect 14908 47844 14932 47846
rect 14988 47844 15012 47846
rect 15068 47844 15092 47846
rect 14852 47824 15148 47844
rect 15488 47666 15516 49778
rect 16316 49706 16344 50118
rect 16408 49910 16436 50322
rect 16396 49904 16448 49910
rect 16396 49846 16448 49852
rect 16304 49700 16356 49706
rect 16304 49642 16356 49648
rect 16408 49094 16436 49846
rect 16120 49088 16172 49094
rect 16120 49030 16172 49036
rect 16396 49088 16448 49094
rect 16396 49030 16448 49036
rect 16132 48754 16160 49030
rect 16120 48748 16172 48754
rect 16120 48690 16172 48696
rect 15200 47660 15252 47666
rect 15200 47602 15252 47608
rect 15476 47660 15528 47666
rect 15476 47602 15528 47608
rect 14852 46812 15148 46832
rect 14908 46810 14932 46812
rect 14988 46810 15012 46812
rect 15068 46810 15092 46812
rect 14930 46758 14932 46810
rect 14994 46758 15006 46810
rect 15068 46758 15070 46810
rect 14908 46756 14932 46758
rect 14988 46756 15012 46758
rect 15068 46756 15092 46758
rect 14852 46736 15148 46756
rect 14832 46572 14884 46578
rect 14832 46514 14884 46520
rect 14844 46458 14872 46514
rect 14752 46430 14872 46458
rect 14556 44872 14608 44878
rect 14556 44814 14608 44820
rect 14464 44804 14516 44810
rect 14464 44746 14516 44752
rect 14200 41386 14412 41414
rect 14096 36644 14148 36650
rect 14096 36586 14148 36592
rect 14004 36236 14056 36242
rect 14004 36178 14056 36184
rect 14016 35562 14044 36178
rect 14200 35698 14228 41386
rect 14280 40520 14332 40526
rect 14280 40462 14332 40468
rect 14292 39642 14320 40462
rect 14372 39840 14424 39846
rect 14372 39782 14424 39788
rect 14280 39636 14332 39642
rect 14280 39578 14332 39584
rect 14384 38400 14412 39782
rect 14292 38372 14412 38400
rect 14188 35692 14240 35698
rect 14188 35634 14240 35640
rect 14004 35556 14056 35562
rect 14004 35498 14056 35504
rect 13912 35284 13964 35290
rect 13912 35226 13964 35232
rect 14004 35148 14056 35154
rect 14004 35090 14056 35096
rect 13910 35048 13966 35057
rect 13832 35006 13910 35034
rect 13910 34983 13966 34992
rect 13728 34604 13780 34610
rect 13728 34546 13780 34552
rect 13726 34504 13782 34513
rect 13726 34439 13782 34448
rect 13740 32337 13768 34439
rect 13820 34400 13872 34406
rect 13820 34342 13872 34348
rect 13832 32978 13860 34342
rect 13924 33998 13952 34983
rect 14016 34610 14044 35090
rect 14292 35034 14320 38372
rect 14372 38208 14424 38214
rect 14372 38150 14424 38156
rect 14384 37194 14412 38150
rect 14372 37188 14424 37194
rect 14372 37130 14424 37136
rect 14372 36644 14424 36650
rect 14372 36586 14424 36592
rect 14108 35006 14320 35034
rect 14004 34604 14056 34610
rect 14004 34546 14056 34552
rect 14004 34060 14056 34066
rect 14004 34002 14056 34008
rect 13912 33992 13964 33998
rect 13912 33934 13964 33940
rect 13912 33448 13964 33454
rect 13912 33390 13964 33396
rect 13820 32972 13872 32978
rect 13820 32914 13872 32920
rect 13924 32502 13952 33390
rect 14016 33318 14044 34002
rect 14004 33312 14056 33318
rect 14004 33254 14056 33260
rect 14004 33040 14056 33046
rect 14004 32982 14056 32988
rect 13912 32496 13964 32502
rect 13912 32438 13964 32444
rect 13726 32328 13782 32337
rect 13726 32263 13782 32272
rect 13728 31952 13780 31958
rect 13728 31894 13780 31900
rect 13740 30394 13768 31894
rect 13820 31884 13872 31890
rect 13820 31826 13872 31832
rect 13832 31142 13860 31826
rect 13912 31816 13964 31822
rect 13912 31758 13964 31764
rect 13820 31136 13872 31142
rect 13820 31078 13872 31084
rect 13924 30802 13952 31758
rect 13912 30796 13964 30802
rect 13912 30738 13964 30744
rect 13820 30592 13872 30598
rect 13820 30534 13872 30540
rect 13728 30388 13780 30394
rect 13728 30330 13780 30336
rect 13728 30252 13780 30258
rect 13728 30194 13780 30200
rect 13740 28490 13768 30194
rect 13832 30190 13860 30534
rect 13820 30184 13872 30190
rect 13820 30126 13872 30132
rect 13924 30122 13952 30738
rect 13912 30116 13964 30122
rect 13912 30058 13964 30064
rect 13818 29880 13874 29889
rect 13818 29815 13820 29824
rect 13872 29815 13874 29824
rect 13912 29844 13964 29850
rect 13820 29786 13872 29792
rect 13912 29786 13964 29792
rect 13728 28484 13780 28490
rect 13728 28426 13780 28432
rect 13740 27130 13768 28426
rect 13820 27872 13872 27878
rect 13820 27814 13872 27820
rect 13832 27606 13860 27814
rect 13820 27600 13872 27606
rect 13820 27542 13872 27548
rect 13728 27124 13780 27130
rect 13728 27066 13780 27072
rect 13740 26790 13768 27066
rect 13924 27033 13952 29786
rect 13910 27024 13966 27033
rect 13820 26988 13872 26994
rect 13910 26959 13966 26968
rect 13820 26930 13872 26936
rect 13728 26784 13780 26790
rect 13728 26726 13780 26732
rect 13832 26586 13860 26930
rect 14016 26874 14044 32982
rect 14108 28694 14136 35006
rect 14188 34128 14240 34134
rect 14188 34070 14240 34076
rect 14200 33522 14228 34070
rect 14280 34060 14332 34066
rect 14280 34002 14332 34008
rect 14188 33516 14240 33522
rect 14188 33458 14240 33464
rect 14188 32836 14240 32842
rect 14188 32778 14240 32784
rect 14200 31346 14228 32778
rect 14188 31340 14240 31346
rect 14188 31282 14240 31288
rect 14188 31136 14240 31142
rect 14188 31078 14240 31084
rect 14200 29850 14228 31078
rect 14292 30802 14320 34002
rect 14280 30796 14332 30802
rect 14280 30738 14332 30744
rect 14188 29844 14240 29850
rect 14188 29786 14240 29792
rect 14292 29714 14320 30738
rect 14280 29708 14332 29714
rect 14280 29650 14332 29656
rect 14280 28960 14332 28966
rect 14280 28902 14332 28908
rect 14096 28688 14148 28694
rect 14096 28630 14148 28636
rect 14188 28620 14240 28626
rect 14188 28562 14240 28568
rect 14096 28076 14148 28082
rect 14096 28018 14148 28024
rect 13924 26846 14044 26874
rect 13820 26580 13872 26586
rect 13820 26522 13872 26528
rect 13728 26240 13780 26246
rect 13728 26182 13780 26188
rect 13740 25242 13768 26182
rect 13820 25764 13872 25770
rect 13820 25706 13872 25712
rect 13832 25498 13860 25706
rect 13820 25492 13872 25498
rect 13820 25434 13872 25440
rect 13740 25214 13860 25242
rect 13728 25152 13780 25158
rect 13728 25094 13780 25100
rect 13740 24274 13768 25094
rect 13728 24268 13780 24274
rect 13728 24210 13780 24216
rect 13832 22760 13860 25214
rect 13740 22732 13860 22760
rect 13544 21684 13596 21690
rect 13544 21626 13596 21632
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13740 21622 13768 22732
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 13832 21622 13860 22578
rect 13728 21616 13780 21622
rect 13556 21564 13728 21570
rect 13556 21558 13780 21564
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 13556 21542 13768 21558
rect 13556 15094 13584 21542
rect 13726 21448 13782 21457
rect 13726 21383 13728 21392
rect 13780 21383 13782 21392
rect 13728 21354 13780 21360
rect 13728 21004 13780 21010
rect 13648 20964 13728 20992
rect 13544 15088 13596 15094
rect 13544 15030 13596 15036
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13464 12442 13492 13466
rect 13648 12782 13676 20964
rect 13728 20946 13780 20952
rect 13726 20904 13782 20913
rect 13924 20890 13952 26846
rect 14004 26512 14056 26518
rect 14004 26454 14056 26460
rect 13726 20839 13782 20848
rect 13832 20862 13952 20890
rect 13636 12776 13688 12782
rect 13556 12724 13636 12730
rect 13556 12718 13688 12724
rect 13556 12702 13676 12718
rect 13740 12714 13768 20839
rect 13832 20210 13860 20862
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13924 20534 13952 20742
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 13832 20182 13952 20210
rect 13924 18970 13952 20182
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13818 18728 13874 18737
rect 13818 18663 13874 18672
rect 13832 18358 13860 18663
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13924 18290 13952 18770
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13832 15162 13860 15506
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13832 14618 13860 14894
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13728 12708 13780 12714
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13464 11665 13492 12378
rect 13450 11656 13506 11665
rect 13450 11591 13506 11600
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 10810 13492 11494
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13464 9722 13492 10542
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13280 9030 13400 9058
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 13096 7886 13124 8026
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13280 7018 13308 9030
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13372 8634 13400 8910
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13280 6990 13400 7018
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 13280 5574 13308 6802
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 13268 4548 13320 4554
rect 13268 4490 13320 4496
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 12912 4078 12940 4218
rect 13280 4078 13308 4490
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12912 3670 12940 3878
rect 13096 3738 13124 4014
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 12912 800 12940 3062
rect 13372 3058 13400 6990
rect 13464 6662 13492 7278
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13464 6322 13492 6598
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13464 4078 13492 6054
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13556 2650 13584 12702
rect 13728 12650 13780 12656
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13648 12374 13676 12582
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13648 11354 13676 12174
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13740 11286 13768 12650
rect 13832 12442 13860 13330
rect 13924 13190 13952 15438
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13924 12306 13952 12854
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13832 11098 13860 12242
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13924 11218 13952 11698
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13648 11070 13860 11098
rect 13648 6934 13676 11070
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13636 6928 13688 6934
rect 13636 6870 13688 6876
rect 13740 6798 13768 8230
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 13648 5642 13676 6666
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5846 13860 6054
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13636 5636 13688 5642
rect 13636 5578 13688 5584
rect 13832 5166 13860 5782
rect 13924 5710 13952 11154
rect 14016 7546 14044 26454
rect 14108 26246 14136 28018
rect 14096 26240 14148 26246
rect 14096 26182 14148 26188
rect 14094 26072 14150 26081
rect 14094 26007 14150 26016
rect 14108 25265 14136 26007
rect 14200 25498 14228 28562
rect 14292 28558 14320 28902
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 14292 26790 14320 28494
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14278 26616 14334 26625
rect 14278 26551 14334 26560
rect 14292 26246 14320 26551
rect 14280 26240 14332 26246
rect 14280 26182 14332 26188
rect 14188 25492 14240 25498
rect 14188 25434 14240 25440
rect 14094 25256 14150 25265
rect 14094 25191 14150 25200
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14108 24410 14136 25094
rect 14200 24410 14228 25434
rect 14280 25424 14332 25430
rect 14278 25392 14280 25401
rect 14332 25392 14334 25401
rect 14278 25327 14334 25336
rect 14280 25220 14332 25226
rect 14280 25162 14332 25168
rect 14292 24954 14320 25162
rect 14280 24948 14332 24954
rect 14280 24890 14332 24896
rect 14278 24848 14334 24857
rect 14278 24783 14334 24792
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 14108 23322 14136 24346
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 14200 23730 14228 24142
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14108 21350 14136 23258
rect 14200 22098 14228 23666
rect 14292 23662 14320 24783
rect 14280 23656 14332 23662
rect 14280 23598 14332 23604
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 14096 21344 14148 21350
rect 14096 21286 14148 21292
rect 14096 20800 14148 20806
rect 14094 20768 14096 20777
rect 14148 20768 14150 20777
rect 14094 20703 14150 20712
rect 14200 20602 14228 22034
rect 14280 21684 14332 21690
rect 14280 21626 14332 21632
rect 14292 21010 14320 21626
rect 14280 21004 14332 21010
rect 14280 20946 14332 20952
rect 14188 20596 14240 20602
rect 14240 20556 14320 20584
rect 14188 20538 14240 20544
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14108 13530 14136 18906
rect 14188 18896 14240 18902
rect 14188 18838 14240 18844
rect 14200 17882 14228 18838
rect 14292 18766 14320 20556
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 14200 14618 14228 17682
rect 14292 16658 14320 18702
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14200 13870 14228 14418
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14108 12918 14136 13466
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 14200 12782 14228 13806
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14108 10130 14136 11766
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 14108 6866 14136 10066
rect 14200 9518 14228 12718
rect 14292 12442 14320 14826
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13924 5166 13952 5646
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13832 4758 13860 5102
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13924 4282 13952 5102
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 14108 4049 14136 6802
rect 14200 5302 14228 9454
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14292 7886 14320 9318
rect 14384 9110 14412 36586
rect 14476 16726 14504 44746
rect 14568 42090 14596 44814
rect 14752 43926 14780 46430
rect 14852 45724 15148 45744
rect 14908 45722 14932 45724
rect 14988 45722 15012 45724
rect 15068 45722 15092 45724
rect 14930 45670 14932 45722
rect 14994 45670 15006 45722
rect 15068 45670 15070 45722
rect 14908 45668 14932 45670
rect 14988 45668 15012 45670
rect 15068 45668 15092 45670
rect 14852 45648 15148 45668
rect 14852 44636 15148 44656
rect 14908 44634 14932 44636
rect 14988 44634 15012 44636
rect 15068 44634 15092 44636
rect 14930 44582 14932 44634
rect 14994 44582 15006 44634
rect 15068 44582 15070 44634
rect 14908 44580 14932 44582
rect 14988 44580 15012 44582
rect 15068 44580 15092 44582
rect 14852 44560 15148 44580
rect 14740 43920 14792 43926
rect 14740 43862 14792 43868
rect 14648 43852 14700 43858
rect 14648 43794 14700 43800
rect 14556 42084 14608 42090
rect 14556 42026 14608 42032
rect 14660 41478 14688 43794
rect 14852 43548 15148 43568
rect 14908 43546 14932 43548
rect 14988 43546 15012 43548
rect 15068 43546 15092 43548
rect 14930 43494 14932 43546
rect 14994 43494 15006 43546
rect 15068 43494 15070 43546
rect 14908 43492 14932 43494
rect 14988 43492 15012 43494
rect 15068 43492 15092 43494
rect 14852 43472 15148 43492
rect 15108 43240 15160 43246
rect 15212 43228 15240 47602
rect 15752 46912 15804 46918
rect 15752 46854 15804 46860
rect 15764 46442 15792 46854
rect 16132 46458 16160 48690
rect 16212 47524 16264 47530
rect 16212 47466 16264 47472
rect 16224 46646 16252 47466
rect 16212 46640 16264 46646
rect 16212 46582 16264 46588
rect 15752 46436 15804 46442
rect 16132 46430 16252 46458
rect 15752 46378 15804 46384
rect 15764 46034 15792 46378
rect 15752 46028 15804 46034
rect 15752 45970 15804 45976
rect 15752 45824 15804 45830
rect 15752 45766 15804 45772
rect 15764 45422 15792 45766
rect 15752 45416 15804 45422
rect 15752 45358 15804 45364
rect 16028 45416 16080 45422
rect 16028 45358 16080 45364
rect 15568 45280 15620 45286
rect 15568 45222 15620 45228
rect 15660 45280 15712 45286
rect 15660 45222 15712 45228
rect 15580 44946 15608 45222
rect 15568 44940 15620 44946
rect 15568 44882 15620 44888
rect 15476 44396 15528 44402
rect 15476 44338 15528 44344
rect 15160 43200 15240 43228
rect 15108 43182 15160 43188
rect 15212 43110 15240 43200
rect 15292 43172 15344 43178
rect 15292 43114 15344 43120
rect 15200 43104 15252 43110
rect 15200 43046 15252 43052
rect 14852 42460 15148 42480
rect 14908 42458 14932 42460
rect 14988 42458 15012 42460
rect 15068 42458 15092 42460
rect 14930 42406 14932 42458
rect 14994 42406 15006 42458
rect 15068 42406 15070 42458
rect 14908 42404 14932 42406
rect 14988 42404 15012 42406
rect 15068 42404 15092 42406
rect 14852 42384 15148 42404
rect 15304 42294 15332 43114
rect 15384 43104 15436 43110
rect 15384 43046 15436 43052
rect 15292 42288 15344 42294
rect 15292 42230 15344 42236
rect 14648 41472 14700 41478
rect 14648 41414 14700 41420
rect 14852 41372 15148 41392
rect 14908 41370 14932 41372
rect 14988 41370 15012 41372
rect 15068 41370 15092 41372
rect 14930 41318 14932 41370
rect 14994 41318 15006 41370
rect 15068 41318 15070 41370
rect 14908 41316 14932 41318
rect 14988 41316 15012 41318
rect 15068 41316 15092 41318
rect 14852 41296 15148 41316
rect 15200 41132 15252 41138
rect 15200 41074 15252 41080
rect 14648 41064 14700 41070
rect 14648 41006 14700 41012
rect 14556 39500 14608 39506
rect 14556 39442 14608 39448
rect 14568 36378 14596 39442
rect 14660 39438 14688 41006
rect 14740 40588 14792 40594
rect 14740 40530 14792 40536
rect 14752 39574 14780 40530
rect 14852 40284 15148 40304
rect 14908 40282 14932 40284
rect 14988 40282 15012 40284
rect 15068 40282 15092 40284
rect 14930 40230 14932 40282
rect 14994 40230 15006 40282
rect 15068 40230 15070 40282
rect 14908 40228 14932 40230
rect 14988 40228 15012 40230
rect 15068 40228 15092 40230
rect 14852 40208 15148 40228
rect 15108 40112 15160 40118
rect 15108 40054 15160 40060
rect 14832 39840 14884 39846
rect 14832 39782 14884 39788
rect 14740 39568 14792 39574
rect 14740 39510 14792 39516
rect 14648 39432 14700 39438
rect 14648 39374 14700 39380
rect 14648 38888 14700 38894
rect 14648 38830 14700 38836
rect 14556 36372 14608 36378
rect 14556 36314 14608 36320
rect 14556 36168 14608 36174
rect 14556 36110 14608 36116
rect 14568 35630 14596 36110
rect 14556 35624 14608 35630
rect 14556 35566 14608 35572
rect 14556 35488 14608 35494
rect 14556 35430 14608 35436
rect 14568 35290 14596 35430
rect 14556 35284 14608 35290
rect 14556 35226 14608 35232
rect 14568 33522 14596 35226
rect 14556 33516 14608 33522
rect 14556 33458 14608 33464
rect 14556 32972 14608 32978
rect 14556 32914 14608 32920
rect 14568 32026 14596 32914
rect 14556 32020 14608 32026
rect 14556 31962 14608 31968
rect 14556 31680 14608 31686
rect 14556 31622 14608 31628
rect 14568 31414 14596 31622
rect 14556 31408 14608 31414
rect 14556 31350 14608 31356
rect 14556 30184 14608 30190
rect 14556 30126 14608 30132
rect 14568 29714 14596 30126
rect 14556 29708 14608 29714
rect 14556 29650 14608 29656
rect 14568 29102 14596 29650
rect 14556 29096 14608 29102
rect 14556 29038 14608 29044
rect 14660 28150 14688 38830
rect 14752 38758 14780 39510
rect 14844 39506 14872 39782
rect 15120 39506 15148 40054
rect 15212 39846 15240 41074
rect 15396 41070 15424 43046
rect 15384 41064 15436 41070
rect 15384 41006 15436 41012
rect 15384 39976 15436 39982
rect 15384 39918 15436 39924
rect 15200 39840 15252 39846
rect 15200 39782 15252 39788
rect 15292 39840 15344 39846
rect 15292 39782 15344 39788
rect 15304 39506 15332 39782
rect 15396 39642 15424 39918
rect 15488 39914 15516 44338
rect 15580 41414 15608 44882
rect 15672 44810 15700 45222
rect 15660 44804 15712 44810
rect 15660 44746 15712 44752
rect 15580 41386 15792 41414
rect 15476 39908 15528 39914
rect 15476 39850 15528 39856
rect 15384 39636 15436 39642
rect 15384 39578 15436 39584
rect 14832 39500 14884 39506
rect 14832 39442 14884 39448
rect 15108 39500 15160 39506
rect 15292 39500 15344 39506
rect 15160 39460 15240 39488
rect 15108 39442 15160 39448
rect 14852 39196 15148 39216
rect 14908 39194 14932 39196
rect 14988 39194 15012 39196
rect 15068 39194 15092 39196
rect 14930 39142 14932 39194
rect 14994 39142 15006 39194
rect 15068 39142 15070 39194
rect 14908 39140 14932 39142
rect 14988 39140 15012 39142
rect 15068 39140 15092 39142
rect 14852 39120 15148 39140
rect 14740 38752 14792 38758
rect 14740 38694 14792 38700
rect 15212 38214 15240 39460
rect 15292 39442 15344 39448
rect 15384 39500 15436 39506
rect 15488 39488 15516 39850
rect 15436 39460 15516 39488
rect 15384 39442 15436 39448
rect 15476 39364 15528 39370
rect 15476 39306 15528 39312
rect 15488 38865 15516 39306
rect 15660 39296 15712 39302
rect 15660 39238 15712 39244
rect 15672 39098 15700 39238
rect 15660 39092 15712 39098
rect 15660 39034 15712 39040
rect 15474 38856 15530 38865
rect 15474 38791 15530 38800
rect 15292 38412 15344 38418
rect 15292 38354 15344 38360
rect 15200 38208 15252 38214
rect 15200 38150 15252 38156
rect 14852 38108 15148 38128
rect 14908 38106 14932 38108
rect 14988 38106 15012 38108
rect 15068 38106 15092 38108
rect 14930 38054 14932 38106
rect 14994 38054 15006 38106
rect 15068 38054 15070 38106
rect 14908 38052 14932 38054
rect 14988 38052 15012 38054
rect 15068 38052 15092 38054
rect 14852 38032 15148 38052
rect 14740 37800 14792 37806
rect 14740 37742 14792 37748
rect 14752 37330 14780 37742
rect 14832 37732 14884 37738
rect 14832 37674 14884 37680
rect 14844 37398 14872 37674
rect 14832 37392 14884 37398
rect 14832 37334 14884 37340
rect 15304 37330 15332 38354
rect 15384 37800 15436 37806
rect 15384 37742 15436 37748
rect 14740 37324 14792 37330
rect 14740 37266 14792 37272
rect 15292 37324 15344 37330
rect 15292 37266 15344 37272
rect 15200 37188 15252 37194
rect 15200 37130 15252 37136
rect 14740 37120 14792 37126
rect 14740 37062 14792 37068
rect 14752 32978 14780 37062
rect 14852 37020 15148 37040
rect 14908 37018 14932 37020
rect 14988 37018 15012 37020
rect 15068 37018 15092 37020
rect 14930 36966 14932 37018
rect 14994 36966 15006 37018
rect 15068 36966 15070 37018
rect 14908 36964 14932 36966
rect 14988 36964 15012 36966
rect 15068 36964 15092 36966
rect 14852 36944 15148 36964
rect 15212 36802 15240 37130
rect 15120 36774 15240 36802
rect 15120 36174 15148 36774
rect 15200 36644 15252 36650
rect 15200 36586 15252 36592
rect 15108 36168 15160 36174
rect 15108 36110 15160 36116
rect 14852 35932 15148 35952
rect 14908 35930 14932 35932
rect 14988 35930 15012 35932
rect 15068 35930 15092 35932
rect 14930 35878 14932 35930
rect 14994 35878 15006 35930
rect 15068 35878 15070 35930
rect 14908 35876 14932 35878
rect 14988 35876 15012 35878
rect 15068 35876 15092 35878
rect 14852 35856 15148 35876
rect 15212 35630 15240 36586
rect 15200 35624 15252 35630
rect 15200 35566 15252 35572
rect 15304 35154 15332 37266
rect 14832 35148 14884 35154
rect 14832 35090 14884 35096
rect 15292 35148 15344 35154
rect 15292 35090 15344 35096
rect 14844 35057 14872 35090
rect 14830 35048 14886 35057
rect 14830 34983 14886 34992
rect 14852 34844 15148 34864
rect 14908 34842 14932 34844
rect 14988 34842 15012 34844
rect 15068 34842 15092 34844
rect 14930 34790 14932 34842
rect 14994 34790 15006 34842
rect 15068 34790 15070 34842
rect 14908 34788 14932 34790
rect 14988 34788 15012 34790
rect 15068 34788 15092 34790
rect 14852 34768 15148 34788
rect 15200 34604 15252 34610
rect 15200 34546 15252 34552
rect 14852 33756 15148 33776
rect 14908 33754 14932 33756
rect 14988 33754 15012 33756
rect 15068 33754 15092 33756
rect 14930 33702 14932 33754
rect 14994 33702 15006 33754
rect 15068 33702 15070 33754
rect 14908 33700 14932 33702
rect 14988 33700 15012 33702
rect 15068 33700 15092 33702
rect 14852 33680 15148 33700
rect 14832 33516 14884 33522
rect 14832 33458 14884 33464
rect 14740 32972 14792 32978
rect 14740 32914 14792 32920
rect 14844 32858 14872 33458
rect 15016 33448 15068 33454
rect 15016 33390 15068 33396
rect 15028 33046 15056 33390
rect 15016 33040 15068 33046
rect 15016 32982 15068 32988
rect 14752 32830 14872 32858
rect 14648 28144 14700 28150
rect 14648 28086 14700 28092
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14568 26625 14596 27406
rect 14752 26976 14780 32830
rect 14852 32668 15148 32688
rect 14908 32666 14932 32668
rect 14988 32666 15012 32668
rect 15068 32666 15092 32668
rect 14930 32614 14932 32666
rect 14994 32614 15006 32666
rect 15068 32614 15070 32666
rect 14908 32612 14932 32614
rect 14988 32612 15012 32614
rect 15068 32612 15092 32614
rect 14852 32592 15148 32612
rect 15108 32428 15160 32434
rect 15108 32370 15160 32376
rect 14924 32292 14976 32298
rect 14924 32234 14976 32240
rect 14936 31958 14964 32234
rect 14924 31952 14976 31958
rect 14924 31894 14976 31900
rect 15120 31890 15148 32370
rect 15108 31884 15160 31890
rect 15108 31826 15160 31832
rect 14852 31580 15148 31600
rect 14908 31578 14932 31580
rect 14988 31578 15012 31580
rect 15068 31578 15092 31580
rect 14930 31526 14932 31578
rect 14994 31526 15006 31578
rect 15068 31526 15070 31578
rect 14908 31524 14932 31526
rect 14988 31524 15012 31526
rect 15068 31524 15092 31526
rect 14852 31504 15148 31524
rect 15106 31376 15162 31385
rect 15106 31311 15162 31320
rect 15120 30802 15148 31311
rect 15108 30796 15160 30802
rect 15108 30738 15160 30744
rect 14852 30492 15148 30512
rect 14908 30490 14932 30492
rect 14988 30490 15012 30492
rect 15068 30490 15092 30492
rect 14930 30438 14932 30490
rect 14994 30438 15006 30490
rect 15068 30438 15070 30490
rect 14908 30436 14932 30438
rect 14988 30436 15012 30438
rect 15068 30436 15092 30438
rect 14852 30416 15148 30436
rect 15108 30252 15160 30258
rect 15108 30194 15160 30200
rect 15120 29560 15148 30194
rect 15212 29730 15240 34546
rect 15304 33318 15332 35090
rect 15292 33312 15344 33318
rect 15292 33254 15344 33260
rect 15292 32360 15344 32366
rect 15292 32302 15344 32308
rect 15304 31958 15332 32302
rect 15292 31952 15344 31958
rect 15292 31894 15344 31900
rect 15304 29850 15332 31894
rect 15396 29850 15424 37742
rect 15488 37670 15516 38791
rect 15660 37800 15712 37806
rect 15660 37742 15712 37748
rect 15476 37664 15528 37670
rect 15476 37606 15528 37612
rect 15568 37664 15620 37670
rect 15568 37606 15620 37612
rect 15580 37398 15608 37606
rect 15672 37398 15700 37742
rect 15568 37392 15620 37398
rect 15568 37334 15620 37340
rect 15660 37392 15712 37398
rect 15660 37334 15712 37340
rect 15476 36780 15528 36786
rect 15476 36722 15528 36728
rect 15488 36242 15516 36722
rect 15476 36236 15528 36242
rect 15476 36178 15528 36184
rect 15474 36136 15530 36145
rect 15474 36071 15530 36080
rect 15488 33862 15516 36071
rect 15580 36020 15608 37334
rect 15660 37256 15712 37262
rect 15660 37198 15712 37204
rect 15672 36718 15700 37198
rect 15660 36712 15712 36718
rect 15660 36654 15712 36660
rect 15672 36145 15700 36654
rect 15658 36136 15714 36145
rect 15658 36071 15714 36080
rect 15580 35992 15700 36020
rect 15568 35760 15620 35766
rect 15568 35702 15620 35708
rect 15580 35290 15608 35702
rect 15568 35284 15620 35290
rect 15568 35226 15620 35232
rect 15672 34066 15700 35992
rect 15660 34060 15712 34066
rect 15660 34002 15712 34008
rect 15568 33992 15620 33998
rect 15568 33934 15620 33940
rect 15476 33856 15528 33862
rect 15476 33798 15528 33804
rect 15476 31952 15528 31958
rect 15476 31894 15528 31900
rect 15488 31385 15516 31894
rect 15580 31754 15608 33934
rect 15580 31726 15700 31754
rect 15568 31680 15620 31686
rect 15568 31622 15620 31628
rect 15474 31376 15530 31385
rect 15474 31311 15530 31320
rect 15476 31272 15528 31278
rect 15580 31260 15608 31622
rect 15528 31232 15608 31260
rect 15476 31214 15528 31220
rect 15474 30832 15530 30841
rect 15474 30767 15476 30776
rect 15528 30767 15530 30776
rect 15476 30738 15528 30744
rect 15566 29880 15622 29889
rect 15292 29844 15344 29850
rect 15292 29786 15344 29792
rect 15384 29844 15436 29850
rect 15566 29815 15622 29824
rect 15384 29786 15436 29792
rect 15580 29782 15608 29815
rect 15568 29776 15620 29782
rect 15212 29702 15424 29730
rect 15568 29718 15620 29724
rect 15292 29572 15344 29578
rect 15120 29532 15240 29560
rect 14852 29404 15148 29424
rect 14908 29402 14932 29404
rect 14988 29402 15012 29404
rect 15068 29402 15092 29404
rect 14930 29350 14932 29402
rect 14994 29350 15006 29402
rect 15068 29350 15070 29402
rect 14908 29348 14932 29350
rect 14988 29348 15012 29350
rect 15068 29348 15092 29350
rect 14852 29328 15148 29348
rect 15212 29220 15240 29532
rect 15292 29514 15344 29520
rect 15120 29192 15240 29220
rect 15120 28506 15148 29192
rect 15120 28478 15240 28506
rect 14852 28316 15148 28336
rect 14908 28314 14932 28316
rect 14988 28314 15012 28316
rect 15068 28314 15092 28316
rect 14930 28262 14932 28314
rect 14994 28262 15006 28314
rect 15068 28262 15070 28314
rect 14908 28260 14932 28262
rect 14988 28260 15012 28262
rect 15068 28260 15092 28262
rect 14852 28240 15148 28260
rect 14924 28144 14976 28150
rect 15212 28098 15240 28478
rect 14924 28086 14976 28092
rect 14936 27606 14964 28086
rect 15120 28070 15240 28098
rect 14924 27600 14976 27606
rect 14924 27542 14976 27548
rect 15120 27470 15148 28070
rect 15200 28008 15252 28014
rect 15200 27950 15252 27956
rect 15108 27464 15160 27470
rect 15108 27406 15160 27412
rect 14852 27228 15148 27248
rect 14908 27226 14932 27228
rect 14988 27226 15012 27228
rect 15068 27226 15092 27228
rect 14930 27174 14932 27226
rect 14994 27174 15006 27226
rect 15068 27174 15070 27226
rect 14908 27172 14932 27174
rect 14988 27172 15012 27174
rect 15068 27172 15092 27174
rect 14852 27152 15148 27172
rect 14660 26948 14780 26976
rect 14554 26616 14610 26625
rect 14554 26551 14610 26560
rect 14660 26568 14688 26948
rect 14738 26888 14794 26897
rect 14738 26823 14740 26832
rect 14792 26823 14794 26832
rect 14832 26852 14884 26858
rect 14740 26794 14792 26800
rect 14832 26794 14884 26800
rect 14660 26540 14780 26568
rect 14556 26444 14608 26450
rect 14556 26386 14608 26392
rect 14648 26444 14700 26450
rect 14648 26386 14700 26392
rect 14568 25838 14596 26386
rect 14556 25832 14608 25838
rect 14556 25774 14608 25780
rect 14568 23254 14596 25774
rect 14556 23248 14608 23254
rect 14556 23190 14608 23196
rect 14568 20874 14596 23190
rect 14660 22234 14688 26386
rect 14752 23662 14780 26540
rect 14844 26518 14872 26794
rect 14832 26512 14884 26518
rect 14832 26454 14884 26460
rect 14852 26140 15148 26160
rect 14908 26138 14932 26140
rect 14988 26138 15012 26140
rect 15068 26138 15092 26140
rect 14930 26086 14932 26138
rect 14994 26086 15006 26138
rect 15068 26086 15070 26138
rect 14908 26084 14932 26086
rect 14988 26084 15012 26086
rect 15068 26084 15092 26086
rect 14852 26064 15148 26084
rect 14924 25968 14976 25974
rect 14924 25910 14976 25916
rect 14936 25362 14964 25910
rect 14924 25356 14976 25362
rect 14924 25298 14976 25304
rect 15212 25294 15240 27950
rect 15200 25288 15252 25294
rect 15200 25230 15252 25236
rect 15304 25226 15332 29514
rect 15292 25220 15344 25226
rect 15292 25162 15344 25168
rect 15396 25158 15424 29702
rect 15566 29608 15622 29617
rect 15566 29543 15568 29552
rect 15620 29543 15622 29552
rect 15568 29514 15620 29520
rect 15476 29504 15528 29510
rect 15476 29446 15528 29452
rect 15488 29073 15516 29446
rect 15474 29064 15530 29073
rect 15474 28999 15530 29008
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 15488 26586 15516 28494
rect 15568 28008 15620 28014
rect 15568 27950 15620 27956
rect 15476 26580 15528 26586
rect 15476 26522 15528 26528
rect 15476 26444 15528 26450
rect 15476 26386 15528 26392
rect 15488 25906 15516 26386
rect 15476 25900 15528 25906
rect 15476 25842 15528 25848
rect 15580 25498 15608 27950
rect 15568 25492 15620 25498
rect 15568 25434 15620 25440
rect 15476 25288 15528 25294
rect 15476 25230 15528 25236
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 14852 25052 15148 25072
rect 14908 25050 14932 25052
rect 14988 25050 15012 25052
rect 15068 25050 15092 25052
rect 14930 24998 14932 25050
rect 14994 24998 15006 25050
rect 15068 24998 15070 25050
rect 14908 24996 14932 24998
rect 14988 24996 15012 24998
rect 15068 24996 15092 24998
rect 14852 24976 15148 24996
rect 15108 24744 15160 24750
rect 15108 24686 15160 24692
rect 15120 24274 15148 24686
rect 15108 24268 15160 24274
rect 15108 24210 15160 24216
rect 14852 23964 15148 23984
rect 14908 23962 14932 23964
rect 14988 23962 15012 23964
rect 15068 23962 15092 23964
rect 14930 23910 14932 23962
rect 14994 23910 15006 23962
rect 15068 23910 15070 23962
rect 14908 23908 14932 23910
rect 14988 23908 15012 23910
rect 15068 23908 15092 23910
rect 14852 23888 15148 23908
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14752 23186 14780 23598
rect 14740 23180 14792 23186
rect 14740 23122 14792 23128
rect 14852 22876 15148 22896
rect 14908 22874 14932 22876
rect 14988 22874 15012 22876
rect 15068 22874 15092 22876
rect 14930 22822 14932 22874
rect 14994 22822 15006 22874
rect 15068 22822 15070 22874
rect 14908 22820 14932 22822
rect 14988 22820 15012 22822
rect 15068 22820 15092 22822
rect 14852 22800 15148 22820
rect 14740 22500 14792 22506
rect 14740 22442 14792 22448
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 14660 21554 14688 22170
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14752 21078 14780 22442
rect 15212 21894 15240 25094
rect 15488 24834 15516 25230
rect 15568 25220 15620 25226
rect 15568 25162 15620 25168
rect 15304 24806 15516 24834
rect 15304 24206 15332 24806
rect 15384 24744 15436 24750
rect 15384 24686 15436 24692
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 14852 21788 15148 21808
rect 14908 21786 14932 21788
rect 14988 21786 15012 21788
rect 15068 21786 15092 21788
rect 14930 21734 14932 21786
rect 14994 21734 15006 21786
rect 15068 21734 15070 21786
rect 14908 21732 14932 21734
rect 14988 21732 15012 21734
rect 15068 21732 15092 21734
rect 14852 21712 15148 21732
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 15200 21412 15252 21418
rect 15200 21354 15252 21360
rect 14740 21072 14792 21078
rect 14740 21014 14792 21020
rect 14556 20868 14608 20874
rect 14556 20810 14608 20816
rect 14568 18306 14596 20810
rect 14852 20700 15148 20720
rect 14908 20698 14932 20700
rect 14988 20698 15012 20700
rect 15068 20698 15092 20700
rect 14930 20646 14932 20698
rect 14994 20646 15006 20698
rect 15068 20646 15070 20698
rect 14908 20644 14932 20646
rect 14988 20644 15012 20646
rect 15068 20644 15092 20646
rect 14852 20624 15148 20644
rect 15212 20398 15240 21354
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 14752 19446 14780 20198
rect 15028 19990 15056 20334
rect 15016 19984 15068 19990
rect 15016 19926 15068 19932
rect 14852 19612 15148 19632
rect 14908 19610 14932 19612
rect 14988 19610 15012 19612
rect 15068 19610 15092 19612
rect 14930 19558 14932 19610
rect 14994 19558 15006 19610
rect 15068 19558 15070 19610
rect 14908 19556 14932 19558
rect 14988 19556 15012 19558
rect 15068 19556 15092 19558
rect 14852 19536 15148 19556
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 14844 18970 14872 19178
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14832 18964 14884 18970
rect 14832 18906 14884 18912
rect 14660 18698 14688 18906
rect 14648 18692 14700 18698
rect 14648 18634 14700 18640
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 14852 18524 15148 18544
rect 14908 18522 14932 18524
rect 14988 18522 15012 18524
rect 15068 18522 15092 18524
rect 14930 18470 14932 18522
rect 14994 18470 15006 18522
rect 15068 18470 15070 18522
rect 14908 18468 14932 18470
rect 14988 18468 15012 18470
rect 15068 18468 15092 18470
rect 14852 18448 15148 18468
rect 14568 18278 14872 18306
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14568 17270 14596 17682
rect 14660 17678 14688 18158
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 14556 17264 14608 17270
rect 14556 17206 14608 17212
rect 14464 16720 14516 16726
rect 14464 16662 14516 16668
rect 14660 15026 14688 17614
rect 14844 17524 14872 18278
rect 14752 17496 14872 17524
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 14752 14804 14780 17496
rect 14852 17436 15148 17456
rect 14908 17434 14932 17436
rect 14988 17434 15012 17436
rect 15068 17434 15092 17436
rect 14930 17382 14932 17434
rect 14994 17382 15006 17434
rect 15068 17382 15070 17434
rect 14908 17380 14932 17382
rect 14988 17380 15012 17382
rect 15068 17380 15092 17382
rect 14852 17360 15148 17380
rect 15212 17134 15240 18566
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 14852 16348 15148 16368
rect 14908 16346 14932 16348
rect 14988 16346 15012 16348
rect 15068 16346 15092 16348
rect 14930 16294 14932 16346
rect 14994 16294 15006 16346
rect 15068 16294 15070 16346
rect 14908 16292 14932 16294
rect 14988 16292 15012 16294
rect 15068 16292 15092 16294
rect 14852 16272 15148 16292
rect 15108 16176 15160 16182
rect 15108 16118 15160 16124
rect 15120 15892 15148 16118
rect 15212 16046 15240 17070
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15120 15864 15240 15892
rect 15212 15502 15240 15864
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 14852 15260 15148 15280
rect 14908 15258 14932 15260
rect 14988 15258 15012 15260
rect 15068 15258 15092 15260
rect 14930 15206 14932 15258
rect 14994 15206 15006 15258
rect 15068 15206 15070 15258
rect 14908 15204 14932 15206
rect 14988 15204 15012 15206
rect 15068 15204 15092 15206
rect 14852 15184 15148 15204
rect 15212 15026 15240 15302
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 14568 14776 14780 14804
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14476 12306 14504 12582
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14476 9042 14504 9386
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14568 6254 14596 14776
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14188 5296 14240 5302
rect 14188 5238 14240 5244
rect 14200 4758 14228 5238
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14094 4040 14150 4049
rect 14094 3975 14150 3984
rect 14108 3534 14136 3975
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14108 2854 14136 3470
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 14280 2576 14332 2582
rect 14280 2518 14332 2524
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 13004 2038 13032 2246
rect 12992 2032 13044 2038
rect 12992 1974 13044 1980
rect 14292 800 14320 2518
rect 14660 2514 14688 14554
rect 14852 14172 15148 14192
rect 14908 14170 14932 14172
rect 14988 14170 15012 14172
rect 15068 14170 15092 14172
rect 14930 14118 14932 14170
rect 14994 14118 15006 14170
rect 15068 14118 15070 14170
rect 14908 14116 14932 14118
rect 14988 14116 15012 14118
rect 15068 14116 15092 14118
rect 14852 14096 15148 14116
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14752 11830 14780 13126
rect 14852 13084 15148 13104
rect 14908 13082 14932 13084
rect 14988 13082 15012 13084
rect 15068 13082 15092 13084
rect 14930 13030 14932 13082
rect 14994 13030 15006 13082
rect 15068 13030 15070 13082
rect 14908 13028 14932 13030
rect 14988 13028 15012 13030
rect 15068 13028 15092 13030
rect 14852 13008 15148 13028
rect 15108 12844 15160 12850
rect 15212 12832 15240 13194
rect 15160 12804 15240 12832
rect 15108 12786 15160 12792
rect 15304 12594 15332 21626
rect 15120 12566 15332 12594
rect 15120 12434 15148 12566
rect 15396 12434 15424 24686
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15488 23050 15516 24346
rect 15580 23474 15608 25162
rect 15672 24750 15700 31726
rect 15660 24744 15712 24750
rect 15660 24686 15712 24692
rect 15580 23446 15700 23474
rect 15476 23044 15528 23050
rect 15476 22986 15528 22992
rect 15568 23044 15620 23050
rect 15568 22986 15620 22992
rect 15488 22166 15516 22986
rect 15580 22574 15608 22986
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15476 22160 15528 22166
rect 15476 22102 15528 22108
rect 15488 21418 15516 22102
rect 15568 21888 15620 21894
rect 15568 21830 15620 21836
rect 15476 21412 15528 21418
rect 15476 21354 15528 21360
rect 15580 21298 15608 21830
rect 15488 21270 15608 21298
rect 15488 21010 15516 21270
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15568 21004 15620 21010
rect 15568 20946 15620 20952
rect 15488 17882 15516 20946
rect 15580 20874 15608 20946
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15580 18086 15608 18702
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15580 15910 15608 16186
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15580 15638 15608 15846
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15120 12406 15240 12434
rect 14852 11996 15148 12016
rect 14908 11994 14932 11996
rect 14988 11994 15012 11996
rect 15068 11994 15092 11996
rect 14930 11942 14932 11994
rect 14994 11942 15006 11994
rect 15068 11942 15070 11994
rect 14908 11940 14932 11942
rect 14988 11940 15012 11942
rect 15068 11940 15092 11942
rect 14852 11920 15148 11940
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14752 11150 14780 11494
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14852 10908 15148 10928
rect 14908 10906 14932 10908
rect 14988 10906 15012 10908
rect 15068 10906 15092 10908
rect 14930 10854 14932 10906
rect 14994 10854 15006 10906
rect 15068 10854 15070 10906
rect 14908 10852 14932 10854
rect 14988 10852 15012 10854
rect 15068 10852 15092 10854
rect 14852 10832 15148 10852
rect 15212 10656 15240 12406
rect 15304 12406 15424 12434
rect 15304 12374 15332 12406
rect 15292 12368 15344 12374
rect 15292 12310 15344 12316
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15120 10628 15240 10656
rect 15120 9994 15148 10628
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 15212 10266 15240 10474
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15108 9988 15160 9994
rect 15108 9930 15160 9936
rect 14852 9820 15148 9840
rect 14908 9818 14932 9820
rect 14988 9818 15012 9820
rect 15068 9818 15092 9820
rect 14930 9766 14932 9818
rect 14994 9766 15006 9818
rect 15068 9766 15070 9818
rect 14908 9764 14932 9766
rect 14988 9764 15012 9766
rect 15068 9764 15092 9766
rect 14852 9744 15148 9764
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14752 8634 14780 9454
rect 15212 9110 15240 10202
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15108 8968 15160 8974
rect 15106 8936 15108 8945
rect 15160 8936 15162 8945
rect 15304 8922 15332 12174
rect 15106 8871 15162 8880
rect 15212 8894 15332 8922
rect 14852 8732 15148 8752
rect 14908 8730 14932 8732
rect 14988 8730 15012 8732
rect 15068 8730 15092 8732
rect 14930 8678 14932 8730
rect 14994 8678 15006 8730
rect 15068 8678 15070 8730
rect 14908 8676 14932 8678
rect 14988 8676 15012 8678
rect 15068 8676 15092 8678
rect 14852 8656 15148 8676
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14752 8090 14780 8366
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14852 7644 15148 7664
rect 14908 7642 14932 7644
rect 14988 7642 15012 7644
rect 15068 7642 15092 7644
rect 14930 7590 14932 7642
rect 14994 7590 15006 7642
rect 15068 7590 15070 7642
rect 14908 7588 14932 7590
rect 14988 7588 15012 7590
rect 15068 7588 15092 7590
rect 14852 7568 15148 7588
rect 15016 7336 15068 7342
rect 15014 7304 15016 7313
rect 15068 7304 15070 7313
rect 15014 7239 15070 7248
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 14752 6934 14780 7142
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14844 6746 14872 7142
rect 14752 6718 14872 6746
rect 14752 5370 14780 6718
rect 14852 6556 15148 6576
rect 14908 6554 14932 6556
rect 14988 6554 15012 6556
rect 15068 6554 15092 6556
rect 14930 6502 14932 6554
rect 14994 6502 15006 6554
rect 15068 6502 15070 6554
rect 14908 6500 14932 6502
rect 14988 6500 15012 6502
rect 15068 6500 15092 6502
rect 14852 6480 15148 6500
rect 15016 6248 15068 6254
rect 15016 6190 15068 6196
rect 15028 5846 15056 6190
rect 15016 5840 15068 5846
rect 15016 5782 15068 5788
rect 14852 5468 15148 5488
rect 14908 5466 14932 5468
rect 14988 5466 15012 5468
rect 15068 5466 15092 5468
rect 14930 5414 14932 5466
rect 14994 5414 15006 5466
rect 15068 5414 15070 5466
rect 14908 5412 14932 5414
rect 14988 5412 15012 5414
rect 15068 5412 15092 5414
rect 14852 5392 15148 5412
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 15212 4826 15240 8894
rect 15396 7426 15424 12242
rect 15488 9382 15516 15506
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15580 12714 15608 15370
rect 15568 12708 15620 12714
rect 15568 12650 15620 12656
rect 15580 10606 15608 12650
rect 15672 12306 15700 23446
rect 15764 22001 15792 41386
rect 15844 39568 15896 39574
rect 15842 39536 15844 39545
rect 15896 39536 15898 39545
rect 15842 39471 15898 39480
rect 15842 39400 15898 39409
rect 15842 39335 15898 39344
rect 15856 39302 15884 39335
rect 15844 39296 15896 39302
rect 15844 39238 15896 39244
rect 16040 37874 16068 45358
rect 16120 45348 16172 45354
rect 16120 45290 16172 45296
rect 16132 44470 16160 45290
rect 16120 44464 16172 44470
rect 16120 44406 16172 44412
rect 16120 41676 16172 41682
rect 16120 41618 16172 41624
rect 16132 41138 16160 41618
rect 16120 41132 16172 41138
rect 16120 41074 16172 41080
rect 16120 39976 16172 39982
rect 16120 39918 16172 39924
rect 16028 37868 16080 37874
rect 16028 37810 16080 37816
rect 15936 37800 15988 37806
rect 15936 37742 15988 37748
rect 15948 37670 15976 37742
rect 15936 37664 15988 37670
rect 15936 37606 15988 37612
rect 16040 36786 16068 37810
rect 16028 36780 16080 36786
rect 16028 36722 16080 36728
rect 15936 36712 15988 36718
rect 15936 36654 15988 36660
rect 15948 36378 15976 36654
rect 15936 36372 15988 36378
rect 15936 36314 15988 36320
rect 15844 36236 15896 36242
rect 15844 36178 15896 36184
rect 15856 34134 15884 36178
rect 16026 35864 16082 35873
rect 16026 35799 16082 35808
rect 16040 35494 16068 35799
rect 16132 35766 16160 39918
rect 16224 36718 16252 46430
rect 16408 44402 16436 49030
rect 16396 44396 16448 44402
rect 16396 44338 16448 44344
rect 16500 44282 16528 52906
rect 18236 52556 18288 52562
rect 18236 52498 18288 52504
rect 17500 51808 17552 51814
rect 17500 51750 17552 51756
rect 17224 50992 17276 50998
rect 17224 50934 17276 50940
rect 16856 50720 16908 50726
rect 16856 50662 16908 50668
rect 16868 50318 16896 50662
rect 17236 50454 17264 50934
rect 17512 50862 17540 51750
rect 18248 51610 18276 52498
rect 18236 51604 18288 51610
rect 18236 51546 18288 51552
rect 18524 51074 18552 52906
rect 19484 52796 19780 52816
rect 19540 52794 19564 52796
rect 19620 52794 19644 52796
rect 19700 52794 19724 52796
rect 19562 52742 19564 52794
rect 19626 52742 19638 52794
rect 19700 52742 19702 52794
rect 19540 52740 19564 52742
rect 19620 52740 19644 52742
rect 19700 52740 19724 52742
rect 19484 52720 19780 52740
rect 20272 52562 20300 54431
rect 20720 53780 20772 53786
rect 20720 53722 20772 53728
rect 20352 52964 20404 52970
rect 20352 52906 20404 52912
rect 20260 52556 20312 52562
rect 20260 52498 20312 52504
rect 19340 52352 19392 52358
rect 19340 52294 19392 52300
rect 19352 51474 19380 52294
rect 19484 51708 19780 51728
rect 19540 51706 19564 51708
rect 19620 51706 19644 51708
rect 19700 51706 19724 51708
rect 19562 51654 19564 51706
rect 19626 51654 19638 51706
rect 19700 51654 19702 51706
rect 19540 51652 19564 51654
rect 19620 51652 19644 51654
rect 19700 51652 19724 51654
rect 19484 51632 19780 51652
rect 19340 51468 19392 51474
rect 19340 51410 19392 51416
rect 18788 51400 18840 51406
rect 18788 51342 18840 51348
rect 18880 51400 18932 51406
rect 18880 51342 18932 51348
rect 18524 51046 18644 51074
rect 18420 50924 18472 50930
rect 18420 50866 18472 50872
rect 17500 50856 17552 50862
rect 17500 50798 17552 50804
rect 18328 50856 18380 50862
rect 18328 50798 18380 50804
rect 18236 50720 18288 50726
rect 18236 50662 18288 50668
rect 18248 50522 18276 50662
rect 18236 50516 18288 50522
rect 18236 50458 18288 50464
rect 17224 50448 17276 50454
rect 17224 50390 17276 50396
rect 16856 50312 16908 50318
rect 16856 50254 16908 50260
rect 16868 48686 16896 50254
rect 17684 50176 17736 50182
rect 17684 50118 17736 50124
rect 18236 50176 18288 50182
rect 18236 50118 18288 50124
rect 17696 49842 17724 50118
rect 18248 49842 18276 50118
rect 17684 49836 17736 49842
rect 17684 49778 17736 49784
rect 18236 49836 18288 49842
rect 18236 49778 18288 49784
rect 16948 49768 17000 49774
rect 16948 49710 17000 49716
rect 16960 49298 16988 49710
rect 17500 49632 17552 49638
rect 17500 49574 17552 49580
rect 16948 49292 17000 49298
rect 16948 49234 17000 49240
rect 16856 48680 16908 48686
rect 16856 48622 16908 48628
rect 16868 48278 16896 48622
rect 16856 48272 16908 48278
rect 16856 48214 16908 48220
rect 16316 44254 16528 44282
rect 16212 36712 16264 36718
rect 16212 36654 16264 36660
rect 16316 36038 16344 44254
rect 16396 43104 16448 43110
rect 16396 43046 16448 43052
rect 16408 42106 16436 43046
rect 16672 42220 16724 42226
rect 16672 42162 16724 42168
rect 16408 42078 16620 42106
rect 16592 42022 16620 42078
rect 16396 42016 16448 42022
rect 16396 41958 16448 41964
rect 16580 42016 16632 42022
rect 16580 41958 16632 41964
rect 16408 41546 16436 41958
rect 16684 41682 16712 42162
rect 16672 41676 16724 41682
rect 16672 41618 16724 41624
rect 16396 41540 16448 41546
rect 16396 41482 16448 41488
rect 16488 41132 16540 41138
rect 16488 41074 16540 41080
rect 16500 39982 16528 41074
rect 16764 40996 16816 41002
rect 16764 40938 16816 40944
rect 16672 40384 16724 40390
rect 16672 40326 16724 40332
rect 16684 39982 16712 40326
rect 16776 40050 16804 40938
rect 16764 40044 16816 40050
rect 16764 39986 16816 39992
rect 16488 39976 16540 39982
rect 16488 39918 16540 39924
rect 16672 39976 16724 39982
rect 16672 39918 16724 39924
rect 16684 39030 16712 39918
rect 16764 39908 16816 39914
rect 16764 39850 16816 39856
rect 16672 39024 16724 39030
rect 16672 38966 16724 38972
rect 16580 38888 16632 38894
rect 16580 38830 16632 38836
rect 16396 38752 16448 38758
rect 16592 38729 16620 38830
rect 16396 38694 16448 38700
rect 16578 38720 16634 38729
rect 16408 38486 16436 38694
rect 16578 38655 16634 38664
rect 16396 38480 16448 38486
rect 16396 38422 16448 38428
rect 16592 37806 16620 38655
rect 16684 37942 16712 38966
rect 16776 38894 16804 39850
rect 16764 38888 16816 38894
rect 16764 38830 16816 38836
rect 16672 37936 16724 37942
rect 16672 37878 16724 37884
rect 16580 37800 16632 37806
rect 16580 37742 16632 37748
rect 16488 37732 16540 37738
rect 16488 37674 16540 37680
rect 16396 36712 16448 36718
rect 16396 36654 16448 36660
rect 16212 36032 16264 36038
rect 16212 35974 16264 35980
rect 16304 36032 16356 36038
rect 16304 35974 16356 35980
rect 16224 35850 16252 35974
rect 16224 35822 16344 35850
rect 16120 35760 16172 35766
rect 16120 35702 16172 35708
rect 16120 35624 16172 35630
rect 16120 35566 16172 35572
rect 16028 35488 16080 35494
rect 15948 35448 16028 35476
rect 15844 34128 15896 34134
rect 15844 34070 15896 34076
rect 15844 33856 15896 33862
rect 15844 33798 15896 33804
rect 15856 31210 15884 33798
rect 15948 32502 15976 35448
rect 16028 35430 16080 35436
rect 16132 35290 16160 35566
rect 16212 35488 16264 35494
rect 16212 35430 16264 35436
rect 16120 35284 16172 35290
rect 16120 35226 16172 35232
rect 16028 34944 16080 34950
rect 16028 34886 16080 34892
rect 16040 34542 16068 34886
rect 16224 34762 16252 35430
rect 16132 34746 16252 34762
rect 16120 34740 16252 34746
rect 16172 34734 16252 34740
rect 16120 34682 16172 34688
rect 16028 34536 16080 34542
rect 16028 34478 16080 34484
rect 16028 34400 16080 34406
rect 16028 34342 16080 34348
rect 16212 34400 16264 34406
rect 16212 34342 16264 34348
rect 16040 34066 16068 34342
rect 16224 34066 16252 34342
rect 16028 34060 16080 34066
rect 16028 34002 16080 34008
rect 16212 34060 16264 34066
rect 16212 34002 16264 34008
rect 16224 33318 16252 34002
rect 16212 33312 16264 33318
rect 16212 33254 16264 33260
rect 16120 32904 16172 32910
rect 16120 32846 16172 32852
rect 15936 32496 15988 32502
rect 15936 32438 15988 32444
rect 16028 32360 16080 32366
rect 16028 32302 16080 32308
rect 15936 32224 15988 32230
rect 15936 32166 15988 32172
rect 15948 31890 15976 32166
rect 15936 31884 15988 31890
rect 15936 31826 15988 31832
rect 16040 31278 16068 32302
rect 16132 32065 16160 32846
rect 16118 32056 16174 32065
rect 16118 31991 16174 32000
rect 16028 31272 16080 31278
rect 16028 31214 16080 31220
rect 15844 31204 15896 31210
rect 15844 31146 15896 31152
rect 16132 30954 16160 31991
rect 16316 31958 16344 35822
rect 16304 31952 16356 31958
rect 16304 31894 16356 31900
rect 16210 31784 16266 31793
rect 16210 31719 16266 31728
rect 16040 30926 16160 30954
rect 16040 30598 16068 30926
rect 16224 30870 16252 31719
rect 16212 30864 16264 30870
rect 16212 30806 16264 30812
rect 16120 30796 16172 30802
rect 16120 30738 16172 30744
rect 16028 30592 16080 30598
rect 16028 30534 16080 30540
rect 15844 30116 15896 30122
rect 15844 30058 15896 30064
rect 15856 29102 15884 30058
rect 15844 29096 15896 29102
rect 15844 29038 15896 29044
rect 15856 26926 15884 29038
rect 16040 28994 16068 30534
rect 16132 30190 16160 30738
rect 16120 30184 16172 30190
rect 16120 30126 16172 30132
rect 16120 29708 16172 29714
rect 16120 29650 16172 29656
rect 15948 28966 16068 28994
rect 16132 28966 16160 29650
rect 15948 28422 15976 28966
rect 16120 28960 16172 28966
rect 16120 28902 16172 28908
rect 16028 28620 16080 28626
rect 16028 28562 16080 28568
rect 15936 28416 15988 28422
rect 15936 28358 15988 28364
rect 15844 26920 15896 26926
rect 15844 26862 15896 26868
rect 15856 26364 15884 26862
rect 15936 26852 15988 26858
rect 15936 26794 15988 26800
rect 15948 26489 15976 26794
rect 15934 26480 15990 26489
rect 15934 26415 15990 26424
rect 15936 26376 15988 26382
rect 15856 26336 15936 26364
rect 15936 26318 15988 26324
rect 16040 26234 16068 28562
rect 16212 28552 16264 28558
rect 16212 28494 16264 28500
rect 16316 28506 16344 31894
rect 16408 28626 16436 36654
rect 16500 36174 16528 37674
rect 16776 36854 16804 38830
rect 16764 36848 16816 36854
rect 16764 36790 16816 36796
rect 16580 36576 16632 36582
rect 16580 36518 16632 36524
rect 16488 36168 16540 36174
rect 16488 36110 16540 36116
rect 16500 35630 16528 36110
rect 16488 35624 16540 35630
rect 16488 35566 16540 35572
rect 16488 34468 16540 34474
rect 16488 34410 16540 34416
rect 16500 34066 16528 34410
rect 16488 34060 16540 34066
rect 16488 34002 16540 34008
rect 16500 33318 16528 34002
rect 16488 33312 16540 33318
rect 16488 33254 16540 33260
rect 16488 32904 16540 32910
rect 16488 32846 16540 32852
rect 16500 32502 16528 32846
rect 16488 32496 16540 32502
rect 16488 32438 16540 32444
rect 16592 32230 16620 36518
rect 16868 36258 16896 48214
rect 16960 41414 16988 49234
rect 17512 48686 17540 49574
rect 17500 48680 17552 48686
rect 17420 48640 17500 48668
rect 17420 48210 17448 48640
rect 17500 48622 17552 48628
rect 17684 48544 17736 48550
rect 17684 48486 17736 48492
rect 17696 48278 17724 48486
rect 17684 48272 17736 48278
rect 17684 48214 17736 48220
rect 17408 48204 17460 48210
rect 17408 48146 17460 48152
rect 17696 47666 17724 48214
rect 18144 48204 18196 48210
rect 18144 48146 18196 48152
rect 18052 48136 18104 48142
rect 18052 48078 18104 48084
rect 17684 47660 17736 47666
rect 17684 47602 17736 47608
rect 17040 47456 17092 47462
rect 17040 47398 17092 47404
rect 17052 46510 17080 47398
rect 17696 46986 17724 47602
rect 18064 47598 18092 48078
rect 18156 47598 18184 48146
rect 18052 47592 18104 47598
rect 18052 47534 18104 47540
rect 18144 47592 18196 47598
rect 18144 47534 18196 47540
rect 18064 47122 18092 47534
rect 18052 47116 18104 47122
rect 18052 47058 18104 47064
rect 18156 46986 18184 47534
rect 18340 47122 18368 50798
rect 18432 50318 18460 50866
rect 18420 50312 18472 50318
rect 18420 50254 18472 50260
rect 18512 50312 18564 50318
rect 18512 50254 18564 50260
rect 18432 49366 18460 50254
rect 18524 49978 18552 50254
rect 18512 49972 18564 49978
rect 18512 49914 18564 49920
rect 18420 49360 18472 49366
rect 18420 49302 18472 49308
rect 18512 48136 18564 48142
rect 18512 48078 18564 48084
rect 18524 47258 18552 48078
rect 18512 47252 18564 47258
rect 18512 47194 18564 47200
rect 18328 47116 18380 47122
rect 18328 47058 18380 47064
rect 17684 46980 17736 46986
rect 17684 46922 17736 46928
rect 18144 46980 18196 46986
rect 18144 46922 18196 46928
rect 18156 46866 18184 46922
rect 18064 46838 18184 46866
rect 17040 46504 17092 46510
rect 17040 46446 17092 46452
rect 17316 46368 17368 46374
rect 17316 46310 17368 46316
rect 17500 46368 17552 46374
rect 17500 46310 17552 46316
rect 17132 46028 17184 46034
rect 17132 45970 17184 45976
rect 17144 45558 17172 45970
rect 17328 45914 17356 46310
rect 17408 46028 17460 46034
rect 17408 45970 17460 45976
rect 17420 45914 17448 45970
rect 17328 45886 17448 45914
rect 17132 45552 17184 45558
rect 17132 45494 17184 45500
rect 17144 44334 17172 45494
rect 17132 44328 17184 44334
rect 17132 44270 17184 44276
rect 17328 44266 17356 45886
rect 17512 45014 17540 46310
rect 18064 45558 18092 46838
rect 18340 46578 18368 47058
rect 18328 46572 18380 46578
rect 18328 46514 18380 46520
rect 18144 46028 18196 46034
rect 18144 45970 18196 45976
rect 18052 45552 18104 45558
rect 18052 45494 18104 45500
rect 18156 45422 18184 45970
rect 18236 45824 18288 45830
rect 18236 45766 18288 45772
rect 18144 45416 18196 45422
rect 18144 45358 18196 45364
rect 18144 45280 18196 45286
rect 18144 45222 18196 45228
rect 17500 45008 17552 45014
rect 17500 44950 17552 44956
rect 18156 44946 18184 45222
rect 18248 44946 18276 45766
rect 18340 45014 18368 46514
rect 18420 45416 18472 45422
rect 18420 45358 18472 45364
rect 18328 45008 18380 45014
rect 18328 44950 18380 44956
rect 17592 44940 17644 44946
rect 17592 44882 17644 44888
rect 18144 44940 18196 44946
rect 18144 44882 18196 44888
rect 18236 44940 18288 44946
rect 18236 44882 18288 44888
rect 17604 44334 17632 44882
rect 18156 44402 18184 44882
rect 18248 44470 18276 44882
rect 18236 44464 18288 44470
rect 18236 44406 18288 44412
rect 18144 44396 18196 44402
rect 18144 44338 18196 44344
rect 17592 44328 17644 44334
rect 17592 44270 17644 44276
rect 17316 44260 17368 44266
rect 17316 44202 17368 44208
rect 16960 41386 17172 41414
rect 17040 40928 17092 40934
rect 17040 40870 17092 40876
rect 17052 40118 17080 40870
rect 17040 40112 17092 40118
rect 17040 40054 17092 40060
rect 16948 39976 17000 39982
rect 16948 39918 17000 39924
rect 16776 36230 16896 36258
rect 16672 35692 16724 35698
rect 16672 35634 16724 35640
rect 16580 32224 16632 32230
rect 16580 32166 16632 32172
rect 16486 31920 16542 31929
rect 16486 31855 16488 31864
rect 16540 31855 16542 31864
rect 16488 31826 16540 31832
rect 16580 31816 16632 31822
rect 16580 31758 16632 31764
rect 16592 31414 16620 31758
rect 16580 31408 16632 31414
rect 16580 31350 16632 31356
rect 16684 30734 16712 35634
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16580 30592 16632 30598
rect 16580 30534 16632 30540
rect 16592 30326 16620 30534
rect 16580 30320 16632 30326
rect 16580 30262 16632 30268
rect 16672 30116 16724 30122
rect 16672 30058 16724 30064
rect 16396 28620 16448 28626
rect 16396 28562 16448 28568
rect 16224 28370 16252 28494
rect 16316 28478 16528 28506
rect 16224 28342 16344 28370
rect 16212 28076 16264 28082
rect 16212 28018 16264 28024
rect 16120 27328 16172 27334
rect 16120 27270 16172 27276
rect 16132 26926 16160 27270
rect 16120 26920 16172 26926
rect 16120 26862 16172 26868
rect 15948 26206 16068 26234
rect 15844 25356 15896 25362
rect 15844 25298 15896 25304
rect 15856 24682 15884 25298
rect 15844 24676 15896 24682
rect 15844 24618 15896 24624
rect 15856 24410 15884 24618
rect 15844 24404 15896 24410
rect 15844 24346 15896 24352
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 15750 21992 15806 22001
rect 15750 21927 15806 21936
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15764 18272 15792 20402
rect 15856 18834 15884 24142
rect 15948 21690 15976 26206
rect 16132 26042 16160 26862
rect 16120 26036 16172 26042
rect 16120 25978 16172 25984
rect 16224 25974 16252 28018
rect 16212 25968 16264 25974
rect 16212 25910 16264 25916
rect 16120 25764 16172 25770
rect 16120 25706 16172 25712
rect 16028 25356 16080 25362
rect 16028 25298 16080 25304
rect 16040 24954 16068 25298
rect 16028 24948 16080 24954
rect 16028 24890 16080 24896
rect 16132 24818 16160 25706
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 16132 24274 16160 24754
rect 16212 24744 16264 24750
rect 16212 24686 16264 24692
rect 16120 24268 16172 24274
rect 16040 24228 16120 24256
rect 16040 23730 16068 24228
rect 16120 24210 16172 24216
rect 16028 23724 16080 23730
rect 16028 23666 16080 23672
rect 16040 22710 16068 23666
rect 16224 23610 16252 24686
rect 16132 23582 16252 23610
rect 16028 22704 16080 22710
rect 16028 22646 16080 22652
rect 16132 22556 16160 23582
rect 16040 22528 16160 22556
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 15936 21480 15988 21486
rect 15936 21422 15988 21428
rect 15948 21146 15976 21422
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 15934 21040 15990 21049
rect 15934 20975 15990 20984
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15844 18692 15896 18698
rect 15844 18634 15896 18640
rect 15856 18426 15884 18634
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15844 18284 15896 18290
rect 15764 18244 15844 18272
rect 15844 18226 15896 18232
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15764 17921 15792 18022
rect 15750 17912 15806 17921
rect 15750 17847 15806 17856
rect 15856 16114 15884 18226
rect 15948 16726 15976 20975
rect 16040 20534 16068 22528
rect 16316 22522 16344 28342
rect 16396 27600 16448 27606
rect 16396 27542 16448 27548
rect 16408 24206 16436 27542
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 16396 23588 16448 23594
rect 16396 23530 16448 23536
rect 16408 23254 16436 23530
rect 16396 23248 16448 23254
rect 16396 23190 16448 23196
rect 16224 22494 16344 22522
rect 16117 22092 16169 22098
rect 16117 22034 16169 22040
rect 16132 21554 16160 22034
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16120 20868 16172 20874
rect 16120 20810 16172 20816
rect 16028 20528 16080 20534
rect 16028 20470 16080 20476
rect 16028 20392 16080 20398
rect 16132 20369 16160 20810
rect 16028 20334 16080 20340
rect 16118 20360 16174 20369
rect 16040 18222 16068 20334
rect 16118 20295 16174 20304
rect 16132 20262 16160 20295
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16120 19984 16172 19990
rect 16120 19926 16172 19932
rect 16132 19514 16160 19926
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 16028 18216 16080 18222
rect 16080 18176 16160 18204
rect 16028 18158 16080 18164
rect 15936 16720 15988 16726
rect 15988 16680 16068 16708
rect 15936 16662 15988 16668
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15856 15162 15884 16050
rect 15936 15972 15988 15978
rect 15936 15914 15988 15920
rect 15948 15502 15976 15914
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 15948 13802 15976 15438
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15580 10266 15608 10406
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15488 8362 15516 8910
rect 15476 8356 15528 8362
rect 15476 8298 15528 8304
rect 15580 7818 15608 9658
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15304 7398 15424 7426
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14752 4078 14780 4626
rect 14852 4380 15148 4400
rect 14908 4378 14932 4380
rect 14988 4378 15012 4380
rect 15068 4378 15092 4380
rect 14930 4326 14932 4378
rect 14994 4326 15006 4378
rect 15068 4326 15070 4378
rect 14908 4324 14932 4326
rect 14988 4324 15012 4326
rect 15068 4324 15092 4326
rect 14852 4304 15148 4324
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 14740 3936 14792 3942
rect 14832 3936 14884 3942
rect 14740 3878 14792 3884
rect 14830 3904 14832 3913
rect 14884 3904 14886 3913
rect 14752 3670 14780 3878
rect 14830 3839 14886 3848
rect 15028 3738 15056 4014
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 14740 3664 14792 3670
rect 14740 3606 14792 3612
rect 15028 3482 15056 3674
rect 15028 3454 15240 3482
rect 14852 3292 15148 3312
rect 14908 3290 14932 3292
rect 14988 3290 15012 3292
rect 15068 3290 15092 3292
rect 14930 3238 14932 3290
rect 14994 3238 15006 3290
rect 15068 3238 15070 3290
rect 14908 3236 14932 3238
rect 14988 3236 15012 3238
rect 15068 3236 15092 3238
rect 14852 3216 15148 3236
rect 15212 3058 15240 3454
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15108 2848 15160 2854
rect 15304 2836 15332 7398
rect 15384 7336 15436 7342
rect 15672 7313 15700 12242
rect 15764 7478 15792 12378
rect 15844 12368 15896 12374
rect 15844 12310 15896 12316
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15384 7278 15436 7284
rect 15658 7304 15714 7313
rect 15396 6458 15424 7278
rect 15658 7239 15714 7248
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15488 7002 15516 7142
rect 15672 7002 15700 7239
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15764 6458 15792 7414
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15856 6390 15884 12310
rect 15934 10568 15990 10577
rect 15934 10503 15936 10512
rect 15988 10503 15990 10512
rect 15936 10474 15988 10480
rect 16040 10266 16068 16680
rect 16132 15978 16160 18176
rect 16120 15972 16172 15978
rect 16120 15914 16172 15920
rect 16132 15434 16160 15914
rect 16120 15428 16172 15434
rect 16120 15370 16172 15376
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16132 12850 16160 15098
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16132 10674 16160 12786
rect 16224 12238 16252 22494
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16316 21962 16344 22374
rect 16304 21956 16356 21962
rect 16304 21898 16356 21904
rect 16408 21434 16436 23190
rect 16316 21406 16436 21434
rect 16316 15570 16344 21406
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16408 19242 16436 21286
rect 16396 19236 16448 19242
rect 16396 19178 16448 19184
rect 16394 19136 16450 19145
rect 16394 19071 16450 19080
rect 16408 18193 16436 19071
rect 16394 18184 16450 18193
rect 16394 18119 16396 18128
rect 16448 18119 16450 18128
rect 16396 18090 16448 18096
rect 16408 18059 16436 18090
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16408 15450 16436 17818
rect 16316 15422 16436 15450
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16224 9722 16252 10406
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15844 6384 15896 6390
rect 15844 6326 15896 6332
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15396 2854 15424 4966
rect 15660 4548 15712 4554
rect 15660 4490 15712 4496
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15580 4146 15608 4422
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15476 4072 15528 4078
rect 15474 4040 15476 4049
rect 15528 4040 15530 4049
rect 15474 3975 15530 3984
rect 15672 3534 15700 4490
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15856 3466 15884 6326
rect 15948 6254 15976 9318
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 16040 8090 16068 8978
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16132 8498 16160 8774
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 15936 6248 15988 6254
rect 15936 6190 15988 6196
rect 16040 5817 16068 7890
rect 16224 7546 16252 8366
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16026 5808 16082 5817
rect 16026 5743 16082 5752
rect 16224 4690 16252 6394
rect 16316 4826 16344 15422
rect 16396 12640 16448 12646
rect 16394 12608 16396 12617
rect 16448 12608 16450 12617
rect 16394 12543 16450 12552
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16408 8430 16436 9386
rect 16500 9330 16528 28478
rect 16580 25832 16632 25838
rect 16580 25774 16632 25780
rect 16592 24954 16620 25774
rect 16580 24948 16632 24954
rect 16580 24890 16632 24896
rect 16684 24800 16712 30058
rect 16592 24772 16712 24800
rect 16592 24342 16620 24772
rect 16672 24676 16724 24682
rect 16672 24618 16724 24624
rect 16684 24410 16712 24618
rect 16672 24404 16724 24410
rect 16672 24346 16724 24352
rect 16580 24336 16632 24342
rect 16580 24278 16632 24284
rect 16592 23662 16620 24278
rect 16672 24200 16724 24206
rect 16672 24142 16724 24148
rect 16580 23656 16632 23662
rect 16580 23598 16632 23604
rect 16592 23050 16620 23598
rect 16684 23594 16712 24142
rect 16672 23588 16724 23594
rect 16672 23530 16724 23536
rect 16580 23044 16632 23050
rect 16580 22986 16632 22992
rect 16684 22930 16712 23530
rect 16592 22902 16712 22930
rect 16592 21554 16620 22902
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16684 22234 16712 22510
rect 16672 22228 16724 22234
rect 16672 22170 16724 22176
rect 16672 21956 16724 21962
rect 16672 21898 16724 21904
rect 16580 21548 16632 21554
rect 16580 21490 16632 21496
rect 16684 20398 16712 21898
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 16580 20324 16632 20330
rect 16580 20266 16632 20272
rect 16592 19990 16620 20266
rect 16580 19984 16632 19990
rect 16580 19926 16632 19932
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16592 19378 16620 19790
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16592 18222 16620 18566
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16672 18148 16724 18154
rect 16672 18090 16724 18096
rect 16684 18057 16712 18090
rect 16670 18048 16726 18057
rect 16670 17983 16726 17992
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16592 13394 16620 13942
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16592 12345 16620 12582
rect 16578 12336 16634 12345
rect 16578 12271 16634 12280
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16592 9722 16620 10202
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16500 9302 16620 9330
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16500 7410 16528 7822
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16592 7290 16620 9302
rect 16684 8090 16712 15506
rect 16776 9586 16804 36230
rect 16856 36168 16908 36174
rect 16856 36110 16908 36116
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16868 8498 16896 36110
rect 16960 34746 16988 39918
rect 17040 38888 17092 38894
rect 17040 38830 17092 38836
rect 16948 34740 17000 34746
rect 16948 34682 17000 34688
rect 17052 34134 17080 38830
rect 17040 34128 17092 34134
rect 17040 34070 17092 34076
rect 16948 33448 17000 33454
rect 16948 33390 17000 33396
rect 16960 30258 16988 33390
rect 17040 32224 17092 32230
rect 17040 32166 17092 32172
rect 17052 31822 17080 32166
rect 17040 31816 17092 31822
rect 17040 31758 17092 31764
rect 17052 30841 17080 31758
rect 17038 30832 17094 30841
rect 17038 30767 17094 30776
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 17040 30048 17092 30054
rect 17040 29990 17092 29996
rect 16948 29708 17000 29714
rect 16948 29650 17000 29656
rect 16960 23610 16988 29650
rect 17052 29646 17080 29990
rect 17040 29640 17092 29646
rect 17040 29582 17092 29588
rect 17040 26784 17092 26790
rect 17040 26726 17092 26732
rect 17052 26353 17080 26726
rect 17038 26344 17094 26353
rect 17038 26279 17094 26288
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 17052 24818 17080 25230
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 17052 24206 17080 24754
rect 17040 24200 17092 24206
rect 17040 24142 17092 24148
rect 16960 23582 17080 23610
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16500 7262 16620 7290
rect 16500 6458 16528 7262
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16592 5370 16620 6734
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16212 4684 16264 4690
rect 15948 4644 16212 4672
rect 15948 4214 15976 4644
rect 16212 4626 16264 4632
rect 16028 4480 16080 4486
rect 16028 4422 16080 4428
rect 15936 4208 15988 4214
rect 15936 4150 15988 4156
rect 16040 4078 16068 4422
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 15844 3460 15896 3466
rect 15844 3402 15896 3408
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15160 2808 15332 2836
rect 15384 2848 15436 2854
rect 15108 2790 15160 2796
rect 15384 2790 15436 2796
rect 15580 2650 15608 3130
rect 16224 3126 16252 3538
rect 16316 3194 16344 4762
rect 16592 4758 16620 5306
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 16580 4752 16632 4758
rect 16580 4694 16632 4700
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16408 3738 16436 4626
rect 16592 4622 16620 4694
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16592 4282 16620 4558
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16486 4176 16542 4185
rect 16486 4111 16542 4120
rect 16500 4078 16528 4111
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16684 3602 16712 4762
rect 16868 3641 16896 8026
rect 16960 5166 16988 23462
rect 17052 23186 17080 23582
rect 17040 23180 17092 23186
rect 17040 23122 17092 23128
rect 17040 21616 17092 21622
rect 17040 21558 17092 21564
rect 17052 19514 17080 21558
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 17038 18184 17094 18193
rect 17038 18119 17094 18128
rect 17052 18086 17080 18119
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 17144 16946 17172 41386
rect 17224 39432 17276 39438
rect 17224 39374 17276 39380
rect 17236 38894 17264 39374
rect 17224 38888 17276 38894
rect 17224 38830 17276 38836
rect 17236 38350 17264 38830
rect 17224 38344 17276 38350
rect 17224 38286 17276 38292
rect 17236 37262 17264 38286
rect 17224 37256 17276 37262
rect 17224 37198 17276 37204
rect 17224 36780 17276 36786
rect 17224 36722 17276 36728
rect 17236 36242 17264 36722
rect 17224 36236 17276 36242
rect 17224 36178 17276 36184
rect 17236 34950 17264 36178
rect 17328 36174 17356 44202
rect 17604 43858 17632 44270
rect 18432 43926 18460 45358
rect 18420 43920 18472 43926
rect 18420 43862 18472 43868
rect 17592 43852 17644 43858
rect 17592 43794 17644 43800
rect 17500 42084 17552 42090
rect 17500 42026 17552 42032
rect 17512 41818 17540 42026
rect 17500 41812 17552 41818
rect 17500 41754 17552 41760
rect 17408 38820 17460 38826
rect 17408 38762 17460 38768
rect 17420 36174 17448 38762
rect 17500 36848 17552 36854
rect 17500 36790 17552 36796
rect 17316 36168 17368 36174
rect 17316 36110 17368 36116
rect 17408 36168 17460 36174
rect 17408 36110 17460 36116
rect 17512 36106 17540 36790
rect 17500 36100 17552 36106
rect 17500 36042 17552 36048
rect 17406 35728 17462 35737
rect 17512 35698 17540 36042
rect 17406 35663 17462 35672
rect 17500 35692 17552 35698
rect 17420 35154 17448 35663
rect 17500 35634 17552 35640
rect 17512 35222 17540 35634
rect 17500 35216 17552 35222
rect 17500 35158 17552 35164
rect 17408 35148 17460 35154
rect 17408 35090 17460 35096
rect 17224 34944 17276 34950
rect 17224 34886 17276 34892
rect 17224 34604 17276 34610
rect 17224 34546 17276 34552
rect 17236 29714 17264 34546
rect 17316 33992 17368 33998
rect 17316 33934 17368 33940
rect 17224 29708 17276 29714
rect 17224 29650 17276 29656
rect 17224 28076 17276 28082
rect 17224 28018 17276 28024
rect 17236 26994 17264 28018
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 17328 26874 17356 33934
rect 17420 31890 17448 35090
rect 17500 34944 17552 34950
rect 17500 34886 17552 34892
rect 17512 32434 17540 34886
rect 17500 32428 17552 32434
rect 17500 32370 17552 32376
rect 17408 31884 17460 31890
rect 17408 31826 17460 31832
rect 17500 31748 17552 31754
rect 17500 31690 17552 31696
rect 17408 31272 17460 31278
rect 17408 31214 17460 31220
rect 17420 30802 17448 31214
rect 17408 30796 17460 30802
rect 17408 30738 17460 30744
rect 17408 30660 17460 30666
rect 17408 30602 17460 30608
rect 17420 30394 17448 30602
rect 17408 30388 17460 30394
rect 17408 30330 17460 30336
rect 17512 28150 17540 31690
rect 17500 28144 17552 28150
rect 17500 28086 17552 28092
rect 17408 27532 17460 27538
rect 17408 27474 17460 27480
rect 17500 27532 17552 27538
rect 17500 27474 17552 27480
rect 17236 26846 17356 26874
rect 17236 23662 17264 26846
rect 17314 26752 17370 26761
rect 17314 26687 17370 26696
rect 17328 25362 17356 26687
rect 17420 26518 17448 27474
rect 17512 27130 17540 27474
rect 17500 27124 17552 27130
rect 17500 27066 17552 27072
rect 17500 26988 17552 26994
rect 17500 26930 17552 26936
rect 17408 26512 17460 26518
rect 17408 26454 17460 26460
rect 17408 26036 17460 26042
rect 17408 25978 17460 25984
rect 17316 25356 17368 25362
rect 17316 25298 17368 25304
rect 17314 24848 17370 24857
rect 17314 24783 17370 24792
rect 17328 24750 17356 24783
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 17236 23526 17264 23598
rect 17224 23520 17276 23526
rect 17224 23462 17276 23468
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 17236 22234 17264 23258
rect 17420 23186 17448 25978
rect 17512 25974 17540 26930
rect 17500 25968 17552 25974
rect 17500 25910 17552 25916
rect 17512 24886 17540 25910
rect 17500 24880 17552 24886
rect 17500 24822 17552 24828
rect 17316 23180 17368 23186
rect 17316 23122 17368 23128
rect 17408 23180 17460 23186
rect 17408 23122 17460 23128
rect 17328 22642 17356 23122
rect 17316 22636 17368 22642
rect 17316 22578 17368 22584
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17236 18737 17264 19246
rect 17222 18728 17278 18737
rect 17222 18663 17278 18672
rect 17052 16918 17172 16946
rect 17052 13954 17080 16918
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 17144 16046 17172 16730
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17236 16114 17264 16390
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17144 15570 17172 15982
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 17144 14074 17172 14826
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17052 13926 17172 13954
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17052 12782 17080 13806
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 17052 10810 17080 12718
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17052 10130 17080 10746
rect 17144 10538 17172 13926
rect 17236 12374 17264 15846
rect 17224 12368 17276 12374
rect 17224 12310 17276 12316
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 17144 9674 17172 10474
rect 17144 9646 17264 9674
rect 17132 9444 17184 9450
rect 17132 9386 17184 9392
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16854 3632 16910 3641
rect 16672 3596 16724 3602
rect 16854 3567 16910 3576
rect 16672 3538 16724 3544
rect 17052 3194 17080 7958
rect 17144 7410 17172 9386
rect 17236 8090 17264 9646
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17132 7404 17184 7410
rect 17328 7392 17356 22578
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17420 19786 17448 20198
rect 17604 20040 17632 43794
rect 18328 43716 18380 43722
rect 18328 43658 18380 43664
rect 17868 42084 17920 42090
rect 17868 42026 17920 42032
rect 17880 38729 17908 42026
rect 18052 41608 18104 41614
rect 18052 41550 18104 41556
rect 18064 40594 18092 41550
rect 18052 40588 18104 40594
rect 18052 40530 18104 40536
rect 18064 40050 18092 40530
rect 18052 40044 18104 40050
rect 18052 39986 18104 39992
rect 18052 39908 18104 39914
rect 18052 39850 18104 39856
rect 17866 38720 17922 38729
rect 17866 38655 17922 38664
rect 17880 38162 17908 38655
rect 17960 38208 18012 38214
rect 17880 38156 17960 38162
rect 17880 38150 18012 38156
rect 17880 38134 18000 38150
rect 18064 37482 18092 39850
rect 17880 37454 18092 37482
rect 17880 37194 17908 37454
rect 17960 37324 18012 37330
rect 17960 37266 18012 37272
rect 17868 37188 17920 37194
rect 17868 37130 17920 37136
rect 17972 36360 18000 37266
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 18064 36582 18092 37198
rect 18052 36576 18104 36582
rect 18052 36518 18104 36524
rect 17880 36332 18000 36360
rect 17880 36224 17908 36332
rect 18052 36236 18104 36242
rect 17880 36196 18000 36224
rect 17868 36100 17920 36106
rect 17868 36042 17920 36048
rect 17880 35562 17908 36042
rect 17868 35556 17920 35562
rect 17868 35498 17920 35504
rect 17972 35290 18000 36196
rect 18052 36178 18104 36184
rect 17960 35284 18012 35290
rect 17960 35226 18012 35232
rect 18064 34746 18092 36178
rect 18144 36032 18196 36038
rect 18144 35974 18196 35980
rect 18236 36032 18288 36038
rect 18236 35974 18288 35980
rect 18052 34740 18104 34746
rect 18052 34682 18104 34688
rect 18050 34640 18106 34649
rect 18050 34575 18106 34584
rect 17684 34536 17736 34542
rect 17684 34478 17736 34484
rect 17696 34066 17724 34478
rect 17868 34400 17920 34406
rect 17960 34400 18012 34406
rect 17868 34342 17920 34348
rect 17958 34368 17960 34377
rect 18012 34368 18014 34377
rect 17880 34066 17908 34342
rect 17958 34303 18014 34312
rect 18064 34134 18092 34575
rect 18052 34128 18104 34134
rect 18052 34070 18104 34076
rect 17684 34060 17736 34066
rect 17684 34002 17736 34008
rect 17868 34060 17920 34066
rect 17868 34002 17920 34008
rect 17960 33856 18012 33862
rect 17960 33798 18012 33804
rect 17868 32768 17920 32774
rect 17868 32710 17920 32716
rect 17776 32360 17828 32366
rect 17776 32302 17828 32308
rect 17684 32292 17736 32298
rect 17684 32234 17736 32240
rect 17696 27946 17724 32234
rect 17788 31890 17816 32302
rect 17880 32230 17908 32710
rect 17868 32224 17920 32230
rect 17868 32166 17920 32172
rect 17776 31884 17828 31890
rect 17776 31826 17828 31832
rect 17868 31680 17920 31686
rect 17868 31622 17920 31628
rect 17880 30802 17908 31622
rect 17868 30796 17920 30802
rect 17868 30738 17920 30744
rect 17776 30660 17828 30666
rect 17776 30602 17828 30608
rect 17684 27940 17736 27946
rect 17684 27882 17736 27888
rect 17696 26926 17724 27882
rect 17684 26920 17736 26926
rect 17684 26862 17736 26868
rect 17696 22710 17724 26862
rect 17684 22704 17736 22710
rect 17684 22646 17736 22652
rect 17696 21962 17724 22646
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 17512 20012 17632 20040
rect 17408 19780 17460 19786
rect 17408 19722 17460 19728
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17420 18358 17448 18702
rect 17408 18352 17460 18358
rect 17408 18294 17460 18300
rect 17512 15910 17540 20012
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 17604 18834 17632 19858
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17604 18426 17632 18770
rect 17696 18766 17724 19790
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 17604 17746 17632 18362
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17604 16658 17632 17546
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17604 16250 17632 16594
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17500 15904 17552 15910
rect 17500 15846 17552 15852
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17512 14482 17540 14962
rect 17604 14958 17632 16186
rect 17696 15162 17724 18702
rect 17684 15156 17736 15162
rect 17684 15098 17736 15104
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17604 14618 17632 14758
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17512 13394 17540 14418
rect 17604 13462 17632 14554
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17696 13870 17724 14282
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17696 13530 17724 13806
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17512 12986 17540 13330
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17604 12866 17632 13398
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17696 12986 17724 13262
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17512 12838 17632 12866
rect 17696 12850 17724 12922
rect 17684 12844 17736 12850
rect 17512 12782 17540 12838
rect 17684 12786 17736 12792
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17408 12640 17460 12646
rect 17406 12608 17408 12617
rect 17460 12608 17462 12617
rect 17406 12543 17462 12552
rect 17512 12434 17540 12718
rect 17512 12406 17724 12434
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 17604 9518 17632 11018
rect 17696 10606 17724 12406
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17696 8974 17724 10406
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17328 7364 17448 7392
rect 17132 7346 17184 7352
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 17328 7002 17356 7210
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17420 5778 17448 7364
rect 17696 6390 17724 8910
rect 17788 7886 17816 30602
rect 17868 28008 17920 28014
rect 17868 27950 17920 27956
rect 17880 27674 17908 27950
rect 17868 27668 17920 27674
rect 17868 27610 17920 27616
rect 17866 27432 17922 27441
rect 17866 27367 17922 27376
rect 17880 27334 17908 27367
rect 17868 27328 17920 27334
rect 17868 27270 17920 27276
rect 17868 26920 17920 26926
rect 17868 26862 17920 26868
rect 17880 26489 17908 26862
rect 17866 26480 17922 26489
rect 17866 26415 17922 26424
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17880 19854 17908 22034
rect 17972 21078 18000 33798
rect 18052 32292 18104 32298
rect 18052 32234 18104 32240
rect 18064 31754 18092 32234
rect 18156 32026 18184 35974
rect 18248 35766 18276 35974
rect 18236 35760 18288 35766
rect 18236 35702 18288 35708
rect 18236 35556 18288 35562
rect 18236 35498 18288 35504
rect 18248 35154 18276 35498
rect 18236 35148 18288 35154
rect 18236 35090 18288 35096
rect 18236 34604 18288 34610
rect 18236 34546 18288 34552
rect 18144 32020 18196 32026
rect 18144 31962 18196 31968
rect 18064 31726 18184 31754
rect 18050 27432 18106 27441
rect 18050 27367 18106 27376
rect 18064 25702 18092 27367
rect 18052 25696 18104 25702
rect 18052 25638 18104 25644
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 18064 23526 18092 23598
rect 18052 23520 18104 23526
rect 18052 23462 18104 23468
rect 18052 22704 18104 22710
rect 18052 22646 18104 22652
rect 18064 22438 18092 22646
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 18064 22098 18092 22374
rect 18052 22092 18104 22098
rect 18052 22034 18104 22040
rect 17960 21072 18012 21078
rect 17960 21014 18012 21020
rect 18052 21072 18104 21078
rect 18052 21014 18104 21020
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17868 19712 17920 19718
rect 17868 19654 17920 19660
rect 17880 18222 17908 19654
rect 17972 18902 18000 20198
rect 18064 18902 18092 21014
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 18052 18896 18104 18902
rect 18052 18838 18104 18844
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 17972 17746 18000 18838
rect 18050 18728 18106 18737
rect 18050 18663 18106 18672
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17880 16658 17908 17614
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17880 14618 17908 16594
rect 17972 16046 18000 16662
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17972 15638 18000 15846
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17880 14006 17908 14350
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17880 12782 17908 13942
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17880 10062 17908 12718
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 16212 3120 16264 3126
rect 16212 3062 16264 3068
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 15764 2514 15792 3062
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 16224 2650 16252 2926
rect 17144 2922 17172 5714
rect 17788 5114 17816 7822
rect 17880 7818 17908 9998
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17972 7018 18000 12718
rect 18064 12288 18092 18663
rect 18156 12782 18184 31726
rect 18248 24070 18276 34546
rect 18340 31754 18368 43658
rect 18420 43104 18472 43110
rect 18420 43046 18472 43052
rect 18432 42770 18460 43046
rect 18420 42764 18472 42770
rect 18420 42706 18472 42712
rect 18420 42084 18472 42090
rect 18420 42026 18472 42032
rect 18432 39982 18460 42026
rect 18616 41414 18644 51046
rect 18800 49774 18828 51342
rect 18892 50862 18920 51342
rect 19616 51264 19668 51270
rect 19616 51206 19668 51212
rect 19628 50862 19656 51206
rect 18880 50856 18932 50862
rect 18880 50798 18932 50804
rect 19616 50856 19668 50862
rect 19616 50798 19668 50804
rect 19984 50720 20036 50726
rect 19984 50662 20036 50668
rect 20076 50720 20128 50726
rect 20076 50662 20128 50668
rect 19484 50620 19780 50640
rect 19540 50618 19564 50620
rect 19620 50618 19644 50620
rect 19700 50618 19724 50620
rect 19562 50566 19564 50618
rect 19626 50566 19638 50618
rect 19700 50566 19702 50618
rect 19540 50564 19564 50566
rect 19620 50564 19644 50566
rect 19700 50564 19724 50566
rect 19484 50544 19780 50564
rect 19996 50454 20024 50662
rect 19984 50448 20036 50454
rect 19984 50390 20036 50396
rect 19248 50380 19300 50386
rect 19248 50322 19300 50328
rect 18788 49768 18840 49774
rect 18788 49710 18840 49716
rect 18880 48204 18932 48210
rect 18880 48146 18932 48152
rect 18788 48000 18840 48006
rect 18788 47942 18840 47948
rect 18800 47530 18828 47942
rect 18788 47524 18840 47530
rect 18788 47466 18840 47472
rect 18788 44804 18840 44810
rect 18788 44746 18840 44752
rect 18696 44464 18748 44470
rect 18696 44406 18748 44412
rect 18708 43246 18736 44406
rect 18800 43858 18828 44746
rect 18788 43852 18840 43858
rect 18788 43794 18840 43800
rect 18892 43790 18920 48146
rect 19260 48006 19288 50322
rect 20088 49978 20116 50662
rect 20260 50312 20312 50318
rect 20260 50254 20312 50260
rect 20168 50176 20220 50182
rect 20168 50118 20220 50124
rect 20076 49972 20128 49978
rect 20076 49914 20128 49920
rect 19340 49768 19392 49774
rect 19340 49710 19392 49716
rect 19352 49366 19380 49710
rect 19484 49532 19780 49552
rect 19540 49530 19564 49532
rect 19620 49530 19644 49532
rect 19700 49530 19724 49532
rect 19562 49478 19564 49530
rect 19626 49478 19638 49530
rect 19700 49478 19702 49530
rect 19540 49476 19564 49478
rect 19620 49476 19644 49478
rect 19700 49476 19724 49478
rect 19484 49456 19780 49476
rect 19340 49360 19392 49366
rect 19340 49302 19392 49308
rect 19484 48444 19780 48464
rect 19540 48442 19564 48444
rect 19620 48442 19644 48444
rect 19700 48442 19724 48444
rect 19562 48390 19564 48442
rect 19626 48390 19638 48442
rect 19700 48390 19702 48442
rect 19540 48388 19564 48390
rect 19620 48388 19644 48390
rect 19700 48388 19724 48390
rect 19484 48368 19780 48388
rect 19984 48136 20036 48142
rect 19984 48078 20036 48084
rect 19064 48000 19116 48006
rect 19064 47942 19116 47948
rect 19248 48000 19300 48006
rect 19248 47942 19300 47948
rect 19076 45014 19104 47942
rect 19064 45008 19116 45014
rect 19064 44950 19116 44956
rect 18972 44940 19024 44946
rect 18972 44882 19024 44888
rect 18984 44198 19012 44882
rect 19156 44736 19208 44742
rect 19156 44678 19208 44684
rect 18972 44192 19024 44198
rect 18972 44134 19024 44140
rect 19168 43858 19196 44678
rect 19064 43852 19116 43858
rect 19064 43794 19116 43800
rect 19156 43852 19208 43858
rect 19156 43794 19208 43800
rect 18880 43784 18932 43790
rect 18880 43726 18932 43732
rect 18696 43240 18748 43246
rect 18696 43182 18748 43188
rect 18788 43240 18840 43246
rect 18788 43182 18840 43188
rect 18800 42226 18828 43182
rect 18892 43110 18920 43726
rect 18972 43172 19024 43178
rect 18972 43114 19024 43120
rect 18880 43104 18932 43110
rect 18880 43046 18932 43052
rect 18984 42838 19012 43114
rect 18972 42832 19024 42838
rect 18972 42774 19024 42780
rect 18788 42220 18840 42226
rect 18788 42162 18840 42168
rect 18524 41386 18644 41414
rect 18420 39976 18472 39982
rect 18420 39918 18472 39924
rect 18420 39840 18472 39846
rect 18420 39782 18472 39788
rect 18432 38350 18460 39782
rect 18420 38344 18472 38350
rect 18420 38286 18472 38292
rect 18432 33862 18460 38286
rect 18524 36310 18552 41386
rect 18604 39908 18656 39914
rect 18604 39850 18656 39856
rect 18616 39506 18644 39850
rect 18604 39500 18656 39506
rect 18604 39442 18656 39448
rect 18800 38282 18828 42162
rect 18880 41472 18932 41478
rect 18880 41414 18932 41420
rect 18892 40594 18920 41414
rect 18880 40588 18932 40594
rect 18880 40530 18932 40536
rect 18972 40588 19024 40594
rect 18972 40530 19024 40536
rect 18984 39030 19012 40530
rect 18972 39024 19024 39030
rect 18972 38966 19024 38972
rect 18788 38276 18840 38282
rect 18788 38218 18840 38224
rect 18604 37868 18656 37874
rect 18604 37810 18656 37816
rect 18616 36582 18644 37810
rect 18984 36786 19012 38966
rect 18972 36780 19024 36786
rect 18972 36722 19024 36728
rect 18604 36576 18656 36582
rect 18604 36518 18656 36524
rect 18696 36576 18748 36582
rect 18696 36518 18748 36524
rect 18512 36304 18564 36310
rect 18512 36246 18564 36252
rect 18616 36242 18644 36518
rect 18604 36236 18656 36242
rect 18604 36178 18656 36184
rect 18512 35624 18564 35630
rect 18512 35566 18564 35572
rect 18524 35290 18552 35566
rect 18512 35284 18564 35290
rect 18512 35226 18564 35232
rect 18420 33856 18472 33862
rect 18420 33798 18472 33804
rect 18420 33380 18472 33386
rect 18420 33322 18472 33328
rect 18432 33046 18460 33322
rect 18420 33040 18472 33046
rect 18420 32982 18472 32988
rect 18524 32978 18552 35226
rect 18708 35154 18736 36518
rect 18880 36304 18932 36310
rect 18880 36246 18932 36252
rect 18788 35760 18840 35766
rect 18786 35728 18788 35737
rect 18840 35728 18842 35737
rect 18786 35663 18842 35672
rect 18892 35578 18920 36246
rect 18972 36236 19024 36242
rect 18972 36178 19024 36184
rect 18984 36038 19012 36178
rect 18972 36032 19024 36038
rect 18972 35974 19024 35980
rect 18800 35550 18920 35578
rect 18604 35148 18656 35154
rect 18604 35090 18656 35096
rect 18696 35148 18748 35154
rect 18696 35090 18748 35096
rect 18616 34746 18644 35090
rect 18604 34740 18656 34746
rect 18604 34682 18656 34688
rect 18800 34354 18828 35550
rect 18616 34326 18828 34354
rect 18512 32972 18564 32978
rect 18512 32914 18564 32920
rect 18616 32570 18644 34326
rect 18696 34128 18748 34134
rect 18696 34070 18748 34076
rect 18708 33130 18736 34070
rect 18788 34060 18840 34066
rect 18788 34002 18840 34008
rect 18800 33318 18828 34002
rect 18788 33312 18840 33318
rect 18788 33254 18840 33260
rect 18708 33102 18920 33130
rect 18696 33040 18748 33046
rect 18696 32982 18748 32988
rect 18708 32774 18736 32982
rect 18696 32768 18748 32774
rect 18696 32710 18748 32716
rect 18604 32564 18656 32570
rect 18604 32506 18656 32512
rect 18788 32564 18840 32570
rect 18788 32506 18840 32512
rect 18512 32428 18564 32434
rect 18512 32370 18564 32376
rect 18524 32026 18552 32370
rect 18800 32366 18828 32506
rect 18788 32360 18840 32366
rect 18708 32320 18788 32348
rect 18512 32020 18564 32026
rect 18512 31962 18564 31968
rect 18524 31890 18552 31962
rect 18512 31884 18564 31890
rect 18512 31826 18564 31832
rect 18340 31726 18460 31754
rect 18328 31272 18380 31278
rect 18328 31214 18380 31220
rect 18340 27577 18368 31214
rect 18326 27568 18382 27577
rect 18326 27503 18382 27512
rect 18326 27432 18382 27441
rect 18326 27367 18382 27376
rect 18340 26450 18368 27367
rect 18328 26444 18380 26450
rect 18328 26386 18380 26392
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 18236 24064 18288 24070
rect 18236 24006 18288 24012
rect 18248 22094 18276 24006
rect 18340 23866 18368 24142
rect 18328 23860 18380 23866
rect 18328 23802 18380 23808
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 18340 23254 18368 23598
rect 18328 23248 18380 23254
rect 18328 23190 18380 23196
rect 18248 22066 18368 22094
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 18248 21146 18276 21286
rect 18236 21140 18288 21146
rect 18236 21082 18288 21088
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18248 17882 18276 20946
rect 18340 20097 18368 22066
rect 18326 20088 18382 20097
rect 18326 20023 18382 20032
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18340 18426 18368 19858
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 18432 17218 18460 31726
rect 18524 31346 18552 31826
rect 18604 31816 18656 31822
rect 18708 31804 18736 32320
rect 18788 32302 18840 32308
rect 18786 32056 18842 32065
rect 18786 31991 18842 32000
rect 18800 31958 18828 31991
rect 18788 31952 18840 31958
rect 18788 31894 18840 31900
rect 18656 31776 18736 31804
rect 18604 31758 18656 31764
rect 18604 31680 18656 31686
rect 18604 31622 18656 31628
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18512 31136 18564 31142
rect 18512 31078 18564 31084
rect 18524 30870 18552 31078
rect 18512 30864 18564 30870
rect 18512 30806 18564 30812
rect 18512 27872 18564 27878
rect 18512 27814 18564 27820
rect 18524 27713 18552 27814
rect 18510 27704 18566 27713
rect 18510 27639 18566 27648
rect 18616 27554 18644 31622
rect 18708 30598 18736 31776
rect 18892 31754 18920 33102
rect 18972 32768 19024 32774
rect 18972 32710 19024 32716
rect 18984 32434 19012 32710
rect 18972 32428 19024 32434
rect 18972 32370 19024 32376
rect 18972 31816 19024 31822
rect 18972 31758 19024 31764
rect 18800 31726 18920 31754
rect 18696 30592 18748 30598
rect 18696 30534 18748 30540
rect 18800 30190 18828 31726
rect 18880 31680 18932 31686
rect 18880 31622 18932 31628
rect 18892 31249 18920 31622
rect 18984 31278 19012 31758
rect 18972 31272 19024 31278
rect 18878 31240 18934 31249
rect 18972 31214 19024 31220
rect 18878 31175 18934 31184
rect 18972 31136 19024 31142
rect 18972 31078 19024 31084
rect 18788 30184 18840 30190
rect 18788 30126 18840 30132
rect 18800 27614 18828 30126
rect 18984 30122 19012 31078
rect 18972 30116 19024 30122
rect 18972 30058 19024 30064
rect 18972 28620 19024 28626
rect 18972 28562 19024 28568
rect 18880 27872 18932 27878
rect 18880 27814 18932 27820
rect 18248 17190 18460 17218
rect 18524 27526 18644 27554
rect 18708 27586 18828 27614
rect 18892 27606 18920 27814
rect 18880 27600 18932 27606
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 18064 12260 18184 12288
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 18064 10266 18092 11154
rect 18156 10441 18184 12260
rect 18248 10554 18276 17190
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18340 16726 18368 16934
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18432 16658 18460 16934
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 18340 15434 18368 15982
rect 18328 15428 18380 15434
rect 18328 15370 18380 15376
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 18340 13462 18368 13670
rect 18328 13456 18380 13462
rect 18328 13398 18380 13404
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18340 12850 18368 13126
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18328 12708 18380 12714
rect 18328 12650 18380 12656
rect 18340 12442 18368 12650
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18432 10713 18460 16186
rect 18418 10704 18474 10713
rect 18418 10639 18474 10648
rect 18420 10600 18472 10606
rect 18248 10526 18368 10554
rect 18420 10542 18472 10548
rect 18236 10464 18288 10470
rect 18142 10432 18198 10441
rect 18236 10406 18288 10412
rect 18142 10367 18198 10376
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 18156 8906 18184 10202
rect 18144 8900 18196 8906
rect 18144 8842 18196 8848
rect 18248 8566 18276 10406
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 17972 6990 18184 7018
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17972 5914 18000 6802
rect 18052 6724 18104 6730
rect 18052 6666 18104 6672
rect 18064 6118 18092 6666
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17880 5166 17908 5714
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17696 5086 17816 5114
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17696 4554 17724 5086
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17788 4758 17816 4966
rect 17880 4826 17908 5102
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17684 4548 17736 4554
rect 17684 4490 17736 4496
rect 17696 4282 17724 4490
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17236 3194 17264 3334
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17696 3058 17724 4218
rect 17880 3670 17908 4422
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17868 3528 17920 3534
rect 17972 3516 18000 5510
rect 18156 5030 18184 6990
rect 18340 6186 18368 10526
rect 18432 10198 18460 10542
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 18418 10024 18474 10033
rect 18418 9959 18474 9968
rect 18432 6934 18460 9959
rect 18524 8022 18552 27526
rect 18604 27464 18656 27470
rect 18604 27406 18656 27412
rect 18616 26450 18644 27406
rect 18604 26444 18656 26450
rect 18604 26386 18656 26392
rect 18616 25838 18644 26386
rect 18604 25832 18656 25838
rect 18604 25774 18656 25780
rect 18708 22094 18736 27586
rect 18880 27542 18932 27548
rect 18788 27532 18840 27538
rect 18788 27474 18840 27480
rect 18800 27441 18828 27474
rect 18786 27432 18842 27441
rect 18786 27367 18842 27376
rect 18892 26926 18920 27542
rect 18984 27062 19012 28562
rect 18972 27056 19024 27062
rect 18972 26998 19024 27004
rect 18788 26920 18840 26926
rect 18788 26862 18840 26868
rect 18880 26920 18932 26926
rect 18880 26862 18932 26868
rect 18800 26586 18828 26862
rect 18984 26772 19012 26998
rect 18892 26744 19012 26772
rect 18788 26580 18840 26586
rect 18788 26522 18840 26528
rect 18788 26376 18840 26382
rect 18788 26318 18840 26324
rect 18800 25906 18828 26318
rect 18788 25900 18840 25906
rect 18788 25842 18840 25848
rect 18616 22066 18736 22094
rect 18616 12617 18644 22066
rect 18800 21078 18828 25842
rect 18788 21072 18840 21078
rect 18788 21014 18840 21020
rect 18788 20936 18840 20942
rect 18788 20878 18840 20884
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 18708 18766 18736 19246
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18708 15502 18736 18702
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18708 13530 18736 13670
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18800 13410 18828 20878
rect 18892 13938 18920 26744
rect 18972 25900 19024 25906
rect 18972 25842 19024 25848
rect 18984 25498 19012 25842
rect 18972 25492 19024 25498
rect 18972 25434 19024 25440
rect 19076 25378 19104 43794
rect 19156 35624 19208 35630
rect 19156 35566 19208 35572
rect 19168 34649 19196 35566
rect 19154 34640 19210 34649
rect 19154 34575 19210 34584
rect 19156 34536 19208 34542
rect 19156 34478 19208 34484
rect 19168 34066 19196 34478
rect 19156 34060 19208 34066
rect 19156 34002 19208 34008
rect 19156 32836 19208 32842
rect 19156 32778 19208 32784
rect 19168 32502 19196 32778
rect 19156 32496 19208 32502
rect 19156 32438 19208 32444
rect 19156 32292 19208 32298
rect 19156 32234 19208 32240
rect 19168 31890 19196 32234
rect 19156 31884 19208 31890
rect 19156 31826 19208 31832
rect 19260 31754 19288 47942
rect 19996 47734 20024 48078
rect 20180 47734 20208 50118
rect 20272 49298 20300 50254
rect 20260 49292 20312 49298
rect 20260 49234 20312 49240
rect 20272 48346 20300 49234
rect 20260 48340 20312 48346
rect 20260 48282 20312 48288
rect 20272 48006 20300 48282
rect 20260 48000 20312 48006
rect 20260 47942 20312 47948
rect 19984 47728 20036 47734
rect 19984 47670 20036 47676
rect 20168 47728 20220 47734
rect 20168 47670 20220 47676
rect 19800 47660 19852 47666
rect 19800 47602 19852 47608
rect 19484 47356 19780 47376
rect 19540 47354 19564 47356
rect 19620 47354 19644 47356
rect 19700 47354 19724 47356
rect 19562 47302 19564 47354
rect 19626 47302 19638 47354
rect 19700 47302 19702 47354
rect 19540 47300 19564 47302
rect 19620 47300 19644 47302
rect 19700 47300 19724 47302
rect 19484 47280 19780 47300
rect 19812 47258 19840 47602
rect 20076 47592 20128 47598
rect 20076 47534 20128 47540
rect 19800 47252 19852 47258
rect 19800 47194 19852 47200
rect 20088 47138 20116 47534
rect 20180 47258 20208 47670
rect 20168 47252 20220 47258
rect 20168 47194 20220 47200
rect 19904 47122 20116 47138
rect 19892 47116 20128 47122
rect 19944 47110 20076 47116
rect 19892 47058 19944 47064
rect 19892 46504 19944 46510
rect 19892 46446 19944 46452
rect 19484 46268 19780 46288
rect 19540 46266 19564 46268
rect 19620 46266 19644 46268
rect 19700 46266 19724 46268
rect 19562 46214 19564 46266
rect 19626 46214 19638 46266
rect 19700 46214 19702 46266
rect 19540 46212 19564 46214
rect 19620 46212 19644 46214
rect 19700 46212 19724 46214
rect 19484 46192 19780 46212
rect 19904 46034 19932 46446
rect 19996 46102 20024 47110
rect 20076 47058 20128 47064
rect 20180 46510 20208 47194
rect 20260 47116 20312 47122
rect 20260 47058 20312 47064
rect 20272 46918 20300 47058
rect 20260 46912 20312 46918
rect 20260 46854 20312 46860
rect 20168 46504 20220 46510
rect 20168 46446 20220 46452
rect 19984 46096 20036 46102
rect 19984 46038 20036 46044
rect 19892 46028 19944 46034
rect 19892 45970 19944 45976
rect 19484 45180 19780 45200
rect 19540 45178 19564 45180
rect 19620 45178 19644 45180
rect 19700 45178 19724 45180
rect 19562 45126 19564 45178
rect 19626 45126 19638 45178
rect 19700 45126 19702 45178
rect 19540 45124 19564 45126
rect 19620 45124 19644 45126
rect 19700 45124 19724 45126
rect 19484 45104 19780 45124
rect 19800 44328 19852 44334
rect 19800 44270 19852 44276
rect 19340 44260 19392 44266
rect 19340 44202 19392 44208
rect 19352 43790 19380 44202
rect 19812 44198 19840 44270
rect 19800 44192 19852 44198
rect 19800 44134 19852 44140
rect 19484 44092 19780 44112
rect 19540 44090 19564 44092
rect 19620 44090 19644 44092
rect 19700 44090 19724 44092
rect 19562 44038 19564 44090
rect 19626 44038 19638 44090
rect 19700 44038 19702 44090
rect 19540 44036 19564 44038
rect 19620 44036 19644 44038
rect 19700 44036 19724 44038
rect 19484 44016 19780 44036
rect 19340 43784 19392 43790
rect 19340 43726 19392 43732
rect 19484 43004 19780 43024
rect 19540 43002 19564 43004
rect 19620 43002 19644 43004
rect 19700 43002 19724 43004
rect 19562 42950 19564 43002
rect 19626 42950 19638 43002
rect 19700 42950 19702 43002
rect 19540 42948 19564 42950
rect 19620 42948 19644 42950
rect 19700 42948 19724 42950
rect 19484 42928 19780 42948
rect 19812 42888 19840 44134
rect 19720 42860 19840 42888
rect 19720 42294 19748 42860
rect 19800 42560 19852 42566
rect 19800 42502 19852 42508
rect 19340 42288 19392 42294
rect 19340 42230 19392 42236
rect 19708 42288 19760 42294
rect 19708 42230 19760 42236
rect 19352 41818 19380 42230
rect 19484 41916 19780 41936
rect 19540 41914 19564 41916
rect 19620 41914 19644 41916
rect 19700 41914 19724 41916
rect 19562 41862 19564 41914
rect 19626 41862 19638 41914
rect 19700 41862 19702 41914
rect 19540 41860 19564 41862
rect 19620 41860 19644 41862
rect 19700 41860 19724 41862
rect 19484 41840 19780 41860
rect 19812 41818 19840 42502
rect 19340 41812 19392 41818
rect 19340 41754 19392 41760
rect 19800 41812 19852 41818
rect 19800 41754 19852 41760
rect 19340 41608 19392 41614
rect 19340 41550 19392 41556
rect 19352 40644 19380 41550
rect 19904 41414 19932 45970
rect 20076 45008 20128 45014
rect 20076 44950 20128 44956
rect 20088 44470 20116 44950
rect 20076 44464 20128 44470
rect 20076 44406 20128 44412
rect 20088 43246 20116 44406
rect 20260 43648 20312 43654
rect 20260 43590 20312 43596
rect 20272 43246 20300 43590
rect 20076 43240 20128 43246
rect 20076 43182 20128 43188
rect 20260 43240 20312 43246
rect 20260 43182 20312 43188
rect 19812 41386 19932 41414
rect 19484 40828 19780 40848
rect 19540 40826 19564 40828
rect 19620 40826 19644 40828
rect 19700 40826 19724 40828
rect 19562 40774 19564 40826
rect 19626 40774 19638 40826
rect 19700 40774 19702 40826
rect 19540 40772 19564 40774
rect 19620 40772 19644 40774
rect 19700 40772 19724 40774
rect 19484 40752 19780 40772
rect 19432 40656 19484 40662
rect 19352 40616 19432 40644
rect 19432 40598 19484 40604
rect 19444 39828 19472 40598
rect 19524 40520 19576 40526
rect 19524 40462 19576 40468
rect 19536 39914 19564 40462
rect 19524 39908 19576 39914
rect 19524 39850 19576 39856
rect 19352 39800 19472 39828
rect 19352 37126 19380 39800
rect 19484 39740 19780 39760
rect 19540 39738 19564 39740
rect 19620 39738 19644 39740
rect 19700 39738 19724 39740
rect 19562 39686 19564 39738
rect 19626 39686 19638 39738
rect 19700 39686 19702 39738
rect 19540 39684 19564 39686
rect 19620 39684 19644 39686
rect 19700 39684 19724 39686
rect 19484 39664 19780 39684
rect 19484 38652 19780 38672
rect 19540 38650 19564 38652
rect 19620 38650 19644 38652
rect 19700 38650 19724 38652
rect 19562 38598 19564 38650
rect 19626 38598 19638 38650
rect 19700 38598 19702 38650
rect 19540 38596 19564 38598
rect 19620 38596 19644 38598
rect 19700 38596 19724 38598
rect 19484 38576 19780 38596
rect 19484 37564 19780 37584
rect 19540 37562 19564 37564
rect 19620 37562 19644 37564
rect 19700 37562 19724 37564
rect 19562 37510 19564 37562
rect 19626 37510 19638 37562
rect 19700 37510 19702 37562
rect 19540 37508 19564 37510
rect 19620 37508 19644 37510
rect 19700 37508 19724 37510
rect 19484 37488 19780 37508
rect 19340 37120 19392 37126
rect 19340 37062 19392 37068
rect 19352 36258 19380 37062
rect 19484 36476 19780 36496
rect 19540 36474 19564 36476
rect 19620 36474 19644 36476
rect 19700 36474 19724 36476
rect 19562 36422 19564 36474
rect 19626 36422 19638 36474
rect 19700 36422 19702 36474
rect 19540 36420 19564 36422
rect 19620 36420 19644 36422
rect 19700 36420 19724 36422
rect 19484 36400 19780 36420
rect 19352 36230 19472 36258
rect 19444 35766 19472 36230
rect 19432 35760 19484 35766
rect 19432 35702 19484 35708
rect 19484 35388 19780 35408
rect 19540 35386 19564 35388
rect 19620 35386 19644 35388
rect 19700 35386 19724 35388
rect 19562 35334 19564 35386
rect 19626 35334 19638 35386
rect 19700 35334 19702 35386
rect 19540 35332 19564 35334
rect 19620 35332 19644 35334
rect 19700 35332 19724 35334
rect 19484 35312 19780 35332
rect 19708 35148 19760 35154
rect 19708 35090 19760 35096
rect 19616 34944 19668 34950
rect 19616 34886 19668 34892
rect 19628 34678 19656 34886
rect 19720 34746 19748 35090
rect 19708 34740 19760 34746
rect 19708 34682 19760 34688
rect 19616 34672 19668 34678
rect 19616 34614 19668 34620
rect 19484 34300 19780 34320
rect 19540 34298 19564 34300
rect 19620 34298 19644 34300
rect 19700 34298 19724 34300
rect 19562 34246 19564 34298
rect 19626 34246 19638 34298
rect 19700 34246 19702 34298
rect 19540 34244 19564 34246
rect 19620 34244 19644 34246
rect 19700 34244 19724 34246
rect 19484 34224 19780 34244
rect 19484 33212 19780 33232
rect 19540 33210 19564 33212
rect 19620 33210 19644 33212
rect 19700 33210 19724 33212
rect 19562 33158 19564 33210
rect 19626 33158 19638 33210
rect 19700 33158 19702 33210
rect 19540 33156 19564 33158
rect 19620 33156 19644 33158
rect 19700 33156 19724 33158
rect 19484 33136 19780 33156
rect 19484 32124 19780 32144
rect 19540 32122 19564 32124
rect 19620 32122 19644 32124
rect 19700 32122 19724 32124
rect 19562 32070 19564 32122
rect 19626 32070 19638 32122
rect 19700 32070 19702 32122
rect 19540 32068 19564 32070
rect 19620 32068 19644 32070
rect 19700 32068 19724 32070
rect 19484 32048 19780 32068
rect 18984 25350 19104 25378
rect 19168 31726 19288 31754
rect 18984 16250 19012 25350
rect 19064 25220 19116 25226
rect 19064 25162 19116 25168
rect 19076 24274 19104 25162
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 19076 22710 19104 24210
rect 19064 22704 19116 22710
rect 19064 22646 19116 22652
rect 19064 22092 19116 22098
rect 19064 22034 19116 22040
rect 19076 21690 19104 22034
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 19076 21078 19104 21286
rect 19064 21072 19116 21078
rect 19064 21014 19116 21020
rect 19076 20398 19104 21014
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 19076 18902 19104 19110
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 19076 18630 19104 18838
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 18972 15972 19024 15978
rect 18972 15914 19024 15920
rect 18984 15638 19012 15914
rect 18972 15632 19024 15638
rect 18970 15600 18972 15609
rect 19064 15632 19116 15638
rect 19024 15600 19026 15609
rect 19064 15574 19116 15580
rect 18970 15535 19026 15544
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18708 13382 18828 13410
rect 18708 12714 18736 13382
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18602 12608 18658 12617
rect 18602 12543 18658 12552
rect 18604 12368 18656 12374
rect 18602 12336 18604 12345
rect 18656 12336 18658 12345
rect 18602 12271 18658 12280
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18616 10062 18644 12174
rect 18708 11218 18736 12650
rect 18786 12608 18842 12617
rect 18786 12543 18842 12552
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18512 8016 18564 8022
rect 18512 7958 18564 7964
rect 18524 7546 18552 7958
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18524 7002 18552 7482
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18420 6928 18472 6934
rect 18420 6870 18472 6876
rect 18616 6798 18644 9998
rect 18708 9382 18736 11018
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18708 7954 18736 8026
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18708 7750 18736 7890
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18800 7018 18828 12543
rect 18892 11354 18920 13874
rect 18984 12238 19012 15302
rect 19076 14618 19104 15574
rect 19064 14612 19116 14618
rect 19064 14554 19116 14560
rect 19168 14464 19196 31726
rect 19484 31036 19780 31056
rect 19540 31034 19564 31036
rect 19620 31034 19644 31036
rect 19700 31034 19724 31036
rect 19562 30982 19564 31034
rect 19626 30982 19638 31034
rect 19700 30982 19702 31034
rect 19540 30980 19564 30982
rect 19620 30980 19644 30982
rect 19700 30980 19724 30982
rect 19484 30960 19780 30980
rect 19432 30796 19484 30802
rect 19432 30738 19484 30744
rect 19708 30796 19760 30802
rect 19708 30738 19760 30744
rect 19444 30598 19472 30738
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19720 30326 19748 30738
rect 19708 30320 19760 30326
rect 19708 30262 19760 30268
rect 19484 29948 19780 29968
rect 19540 29946 19564 29948
rect 19620 29946 19644 29948
rect 19700 29946 19724 29948
rect 19562 29894 19564 29946
rect 19626 29894 19638 29946
rect 19700 29894 19702 29946
rect 19540 29892 19564 29894
rect 19620 29892 19644 29894
rect 19700 29892 19724 29894
rect 19484 29872 19780 29892
rect 19484 28860 19780 28880
rect 19540 28858 19564 28860
rect 19620 28858 19644 28860
rect 19700 28858 19724 28860
rect 19562 28806 19564 28858
rect 19626 28806 19638 28858
rect 19700 28806 19702 28858
rect 19540 28804 19564 28806
rect 19620 28804 19644 28806
rect 19700 28804 19724 28806
rect 19484 28784 19780 28804
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 19248 28484 19300 28490
rect 19248 28426 19300 28432
rect 19260 27538 19288 28426
rect 19248 27532 19300 27538
rect 19248 27474 19300 27480
rect 19260 25294 19288 27474
rect 19352 27418 19380 28494
rect 19484 27772 19780 27792
rect 19540 27770 19564 27772
rect 19620 27770 19644 27772
rect 19700 27770 19724 27772
rect 19562 27718 19564 27770
rect 19626 27718 19638 27770
rect 19700 27718 19702 27770
rect 19540 27716 19564 27718
rect 19620 27716 19644 27718
rect 19700 27716 19724 27718
rect 19484 27696 19780 27716
rect 19352 27390 19472 27418
rect 19444 26840 19472 27390
rect 19524 27328 19576 27334
rect 19524 27270 19576 27276
rect 19536 26926 19564 27270
rect 19524 26920 19576 26926
rect 19524 26862 19576 26868
rect 19352 26812 19472 26840
rect 19352 25974 19380 26812
rect 19484 26684 19780 26704
rect 19540 26682 19564 26684
rect 19620 26682 19644 26684
rect 19700 26682 19724 26684
rect 19562 26630 19564 26682
rect 19626 26630 19638 26682
rect 19700 26630 19702 26682
rect 19540 26628 19564 26630
rect 19620 26628 19644 26630
rect 19700 26628 19724 26630
rect 19484 26608 19780 26628
rect 19340 25968 19392 25974
rect 19340 25910 19392 25916
rect 19352 25838 19380 25910
rect 19340 25832 19392 25838
rect 19340 25774 19392 25780
rect 19352 25294 19380 25774
rect 19484 25596 19780 25616
rect 19540 25594 19564 25596
rect 19620 25594 19644 25596
rect 19700 25594 19724 25596
rect 19562 25542 19564 25594
rect 19626 25542 19638 25594
rect 19700 25542 19702 25594
rect 19540 25540 19564 25542
rect 19620 25540 19644 25542
rect 19700 25540 19724 25542
rect 19484 25520 19780 25540
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 19260 21554 19288 25230
rect 19484 24508 19780 24528
rect 19540 24506 19564 24508
rect 19620 24506 19644 24508
rect 19700 24506 19724 24508
rect 19562 24454 19564 24506
rect 19626 24454 19638 24506
rect 19700 24454 19702 24506
rect 19540 24452 19564 24454
rect 19620 24452 19644 24454
rect 19700 24452 19724 24454
rect 19484 24432 19780 24452
rect 19484 23420 19780 23440
rect 19540 23418 19564 23420
rect 19620 23418 19644 23420
rect 19700 23418 19724 23420
rect 19562 23366 19564 23418
rect 19626 23366 19638 23418
rect 19700 23366 19702 23418
rect 19540 23364 19564 23366
rect 19620 23364 19644 23366
rect 19700 23364 19724 23366
rect 19484 23344 19780 23364
rect 19484 22332 19780 22352
rect 19540 22330 19564 22332
rect 19620 22330 19644 22332
rect 19700 22330 19724 22332
rect 19562 22278 19564 22330
rect 19626 22278 19638 22330
rect 19700 22278 19702 22330
rect 19540 22276 19564 22278
rect 19620 22276 19644 22278
rect 19700 22276 19724 22278
rect 19484 22256 19780 22276
rect 19812 21690 19840 41386
rect 20088 40594 20116 43182
rect 20364 41414 20392 52906
rect 20732 52358 20760 53722
rect 20904 53644 20956 53650
rect 20904 53586 20956 53592
rect 20916 52562 20944 53586
rect 21180 53440 21232 53446
rect 21180 53382 21232 53388
rect 21192 53242 21220 53382
rect 21180 53236 21232 53242
rect 21180 53178 21232 53184
rect 22020 53174 22048 55200
rect 23204 53576 23256 53582
rect 23204 53518 23256 53524
rect 22836 53508 22888 53514
rect 22836 53450 22888 53456
rect 22008 53168 22060 53174
rect 22008 53110 22060 53116
rect 21640 52964 21692 52970
rect 21640 52906 21692 52912
rect 22100 52964 22152 52970
rect 22100 52906 22152 52912
rect 20904 52556 20956 52562
rect 20904 52498 20956 52504
rect 21364 52556 21416 52562
rect 21364 52498 21416 52504
rect 20720 52352 20772 52358
rect 20720 52294 20772 52300
rect 20444 51876 20496 51882
rect 20444 51818 20496 51824
rect 20456 51610 20484 51818
rect 21376 51814 21404 52498
rect 21456 52488 21508 52494
rect 21456 52430 21508 52436
rect 20812 51808 20864 51814
rect 20812 51750 20864 51756
rect 21364 51808 21416 51814
rect 21364 51750 21416 51756
rect 20824 51610 20852 51750
rect 20444 51604 20496 51610
rect 20444 51546 20496 51552
rect 20812 51604 20864 51610
rect 20812 51546 20864 51552
rect 20904 51400 20956 51406
rect 20904 51342 20956 51348
rect 21364 51400 21416 51406
rect 21364 51342 21416 51348
rect 20916 49842 20944 51342
rect 21272 50720 21324 50726
rect 21272 50662 21324 50668
rect 21284 50522 21312 50662
rect 21272 50516 21324 50522
rect 21272 50458 21324 50464
rect 21180 50312 21232 50318
rect 21180 50254 21232 50260
rect 20996 50176 21048 50182
rect 20996 50118 21048 50124
rect 20904 49836 20956 49842
rect 20904 49778 20956 49784
rect 20444 49360 20496 49366
rect 20444 49302 20496 49308
rect 20456 48210 20484 49302
rect 20444 48204 20496 48210
rect 20444 48146 20496 48152
rect 20628 48204 20680 48210
rect 20628 48146 20680 48152
rect 20444 48000 20496 48006
rect 20444 47942 20496 47948
rect 20456 47122 20484 47942
rect 20444 47116 20496 47122
rect 20444 47058 20496 47064
rect 20640 46918 20668 48146
rect 20916 47598 20944 49778
rect 21008 49774 21036 50118
rect 21192 49978 21220 50254
rect 21180 49972 21232 49978
rect 21180 49914 21232 49920
rect 20996 49768 21048 49774
rect 20996 49710 21048 49716
rect 21376 49314 21404 51342
rect 21468 50862 21496 52430
rect 21456 50856 21508 50862
rect 21456 50798 21508 50804
rect 21376 49286 21588 49314
rect 21364 49224 21416 49230
rect 21364 49166 21416 49172
rect 21180 48748 21232 48754
rect 21180 48690 21232 48696
rect 21088 48204 21140 48210
rect 21088 48146 21140 48152
rect 20904 47592 20956 47598
rect 20904 47534 20956 47540
rect 20996 47592 21048 47598
rect 20996 47534 21048 47540
rect 21008 47122 21036 47534
rect 21100 47122 21128 48146
rect 21192 48142 21220 48690
rect 21376 48686 21404 49166
rect 21364 48680 21416 48686
rect 21364 48622 21416 48628
rect 21376 48210 21404 48622
rect 21364 48204 21416 48210
rect 21364 48146 21416 48152
rect 21180 48136 21232 48142
rect 21180 48078 21232 48084
rect 20996 47116 21048 47122
rect 20996 47058 21048 47064
rect 21088 47116 21140 47122
rect 21088 47058 21140 47064
rect 20904 47048 20956 47054
rect 20904 46990 20956 46996
rect 20628 46912 20680 46918
rect 20628 46854 20680 46860
rect 20272 41386 20392 41414
rect 20076 40588 20128 40594
rect 20076 40530 20128 40536
rect 20168 39908 20220 39914
rect 20168 39850 20220 39856
rect 20076 39296 20128 39302
rect 20076 39238 20128 39244
rect 20088 38554 20116 39238
rect 20180 38758 20208 39850
rect 20168 38752 20220 38758
rect 20168 38694 20220 38700
rect 20076 38548 20128 38554
rect 20076 38490 20128 38496
rect 20076 37936 20128 37942
rect 20076 37878 20128 37884
rect 20088 37806 20116 37878
rect 20180 37806 20208 38694
rect 20076 37800 20128 37806
rect 20076 37742 20128 37748
rect 20168 37800 20220 37806
rect 20168 37742 20220 37748
rect 20088 36038 20116 37742
rect 19892 36032 19944 36038
rect 19892 35974 19944 35980
rect 20076 36032 20128 36038
rect 20076 35974 20128 35980
rect 19904 35290 19932 35974
rect 20076 35556 20128 35562
rect 20076 35498 20128 35504
rect 19892 35284 19944 35290
rect 19892 35226 19944 35232
rect 20088 35154 20116 35498
rect 20076 35148 20128 35154
rect 20076 35090 20128 35096
rect 19984 35012 20036 35018
rect 19984 34954 20036 34960
rect 19996 34626 20024 34954
rect 19904 34610 20024 34626
rect 19892 34604 20024 34610
rect 19944 34598 20024 34604
rect 19892 34546 19944 34552
rect 19984 33040 20036 33046
rect 19984 32982 20036 32988
rect 19892 32972 19944 32978
rect 19892 32914 19944 32920
rect 19800 21684 19852 21690
rect 19800 21626 19852 21632
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 19260 18290 19288 21490
rect 19352 19310 19380 21490
rect 19484 21244 19780 21264
rect 19540 21242 19564 21244
rect 19620 21242 19644 21244
rect 19700 21242 19724 21244
rect 19562 21190 19564 21242
rect 19626 21190 19638 21242
rect 19700 21190 19702 21242
rect 19540 21188 19564 21190
rect 19620 21188 19644 21190
rect 19700 21188 19724 21190
rect 19484 21168 19780 21188
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 19484 20156 19780 20176
rect 19540 20154 19564 20156
rect 19620 20154 19644 20156
rect 19700 20154 19724 20156
rect 19562 20102 19564 20154
rect 19626 20102 19638 20154
rect 19700 20102 19702 20154
rect 19540 20100 19564 20102
rect 19620 20100 19644 20102
rect 19700 20100 19724 20102
rect 19484 20080 19780 20100
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19484 19068 19780 19088
rect 19540 19066 19564 19068
rect 19620 19066 19644 19068
rect 19700 19066 19724 19068
rect 19562 19014 19564 19066
rect 19626 19014 19638 19066
rect 19700 19014 19702 19066
rect 19540 19012 19564 19014
rect 19620 19012 19644 19014
rect 19700 19012 19724 19014
rect 19484 18992 19780 19012
rect 19524 18828 19576 18834
rect 19524 18770 19576 18776
rect 19616 18828 19668 18834
rect 19812 18816 19840 21082
rect 19668 18788 19840 18816
rect 19616 18770 19668 18776
rect 19536 18426 19564 18770
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19628 18306 19656 18770
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19352 18278 19656 18306
rect 19260 17202 19288 18226
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 19352 15638 19380 18278
rect 19484 17980 19780 18000
rect 19540 17978 19564 17980
rect 19620 17978 19644 17980
rect 19700 17978 19724 17980
rect 19562 17926 19564 17978
rect 19626 17926 19638 17978
rect 19700 17926 19702 17978
rect 19540 17924 19564 17926
rect 19620 17924 19644 17926
rect 19700 17924 19724 17926
rect 19484 17904 19780 17924
rect 19484 16892 19780 16912
rect 19540 16890 19564 16892
rect 19620 16890 19644 16892
rect 19700 16890 19724 16892
rect 19562 16838 19564 16890
rect 19626 16838 19638 16890
rect 19700 16838 19702 16890
rect 19540 16836 19564 16838
rect 19620 16836 19644 16838
rect 19700 16836 19724 16838
rect 19484 16816 19780 16836
rect 19484 15804 19780 15824
rect 19540 15802 19564 15804
rect 19620 15802 19644 15804
rect 19700 15802 19724 15804
rect 19562 15750 19564 15802
rect 19626 15750 19638 15802
rect 19700 15750 19702 15802
rect 19540 15748 19564 15750
rect 19620 15748 19644 15750
rect 19700 15748 19724 15750
rect 19484 15728 19780 15748
rect 19340 15632 19392 15638
rect 19340 15574 19392 15580
rect 19076 14436 19196 14464
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 19076 11234 19104 14436
rect 19248 13456 19300 13462
rect 19248 13398 19300 13404
rect 19154 13288 19210 13297
rect 19154 13223 19210 13232
rect 19168 12986 19196 13223
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 18984 11206 19104 11234
rect 18984 10810 19012 11206
rect 19168 11150 19196 12786
rect 19260 12442 19288 13398
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19352 12374 19380 15574
rect 19484 14716 19780 14736
rect 19540 14714 19564 14716
rect 19620 14714 19644 14716
rect 19700 14714 19724 14716
rect 19562 14662 19564 14714
rect 19626 14662 19638 14714
rect 19700 14662 19702 14714
rect 19540 14660 19564 14662
rect 19620 14660 19644 14662
rect 19700 14660 19724 14662
rect 19484 14640 19780 14660
rect 19484 13628 19780 13648
rect 19540 13626 19564 13628
rect 19620 13626 19644 13628
rect 19700 13626 19724 13628
rect 19562 13574 19564 13626
rect 19626 13574 19638 13626
rect 19700 13574 19702 13626
rect 19540 13572 19564 13574
rect 19620 13572 19644 13574
rect 19700 13572 19724 13574
rect 19484 13552 19780 13572
rect 19484 12540 19780 12560
rect 19540 12538 19564 12540
rect 19620 12538 19644 12540
rect 19700 12538 19724 12540
rect 19562 12486 19564 12538
rect 19626 12486 19638 12538
rect 19700 12486 19702 12538
rect 19540 12484 19564 12486
rect 19620 12484 19644 12486
rect 19700 12484 19724 12486
rect 19484 12464 19780 12484
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19260 11558 19288 12242
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 18972 10804 19024 10810
rect 18972 10746 19024 10752
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18892 9489 18920 10066
rect 18878 9480 18934 9489
rect 19076 9450 19104 11018
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19168 10198 19196 10746
rect 19156 10192 19208 10198
rect 19156 10134 19208 10140
rect 19248 10124 19300 10130
rect 19352 10112 19380 12310
rect 19904 11642 19932 32914
rect 19996 28082 20024 32982
rect 20272 32910 20300 41386
rect 20536 40928 20588 40934
rect 20536 40870 20588 40876
rect 20548 40662 20576 40870
rect 20536 40656 20588 40662
rect 20536 40598 20588 40604
rect 20352 38344 20404 38350
rect 20352 38286 20404 38292
rect 20364 37942 20392 38286
rect 20444 38208 20496 38214
rect 20444 38150 20496 38156
rect 20352 37936 20404 37942
rect 20352 37878 20404 37884
rect 20352 37664 20404 37670
rect 20352 37606 20404 37612
rect 20364 37398 20392 37606
rect 20456 37398 20484 38150
rect 20352 37392 20404 37398
rect 20352 37334 20404 37340
rect 20444 37392 20496 37398
rect 20444 37334 20496 37340
rect 20352 37256 20404 37262
rect 20352 37198 20404 37204
rect 20364 34746 20392 37198
rect 20536 36576 20588 36582
rect 20536 36518 20588 36524
rect 20548 35698 20576 36518
rect 20536 35692 20588 35698
rect 20536 35634 20588 35640
rect 20444 35148 20496 35154
rect 20444 35090 20496 35096
rect 20352 34740 20404 34746
rect 20352 34682 20404 34688
rect 20364 34406 20392 34682
rect 20352 34400 20404 34406
rect 20352 34342 20404 34348
rect 20260 32904 20312 32910
rect 20260 32846 20312 32852
rect 20364 32434 20392 34342
rect 20456 34134 20484 35090
rect 20444 34128 20496 34134
rect 20444 34070 20496 34076
rect 20444 33380 20496 33386
rect 20444 33322 20496 33328
rect 20352 32428 20404 32434
rect 20352 32370 20404 32376
rect 20456 32366 20484 33322
rect 20536 32904 20588 32910
rect 20536 32846 20588 32852
rect 20548 32570 20576 32846
rect 20536 32564 20588 32570
rect 20536 32506 20588 32512
rect 20548 32434 20576 32506
rect 20536 32428 20588 32434
rect 20536 32370 20588 32376
rect 20444 32360 20496 32366
rect 20444 32302 20496 32308
rect 20536 32292 20588 32298
rect 20536 32234 20588 32240
rect 20444 31884 20496 31890
rect 20444 31826 20496 31832
rect 20260 31272 20312 31278
rect 20260 31214 20312 31220
rect 20272 30870 20300 31214
rect 20260 30864 20312 30870
rect 20260 30806 20312 30812
rect 20456 30802 20484 31826
rect 20548 31278 20576 32234
rect 20536 31272 20588 31278
rect 20536 31214 20588 31220
rect 20444 30796 20496 30802
rect 20444 30738 20496 30744
rect 20076 30728 20128 30734
rect 20076 30670 20128 30676
rect 20088 29850 20116 30670
rect 20456 30258 20484 30738
rect 20548 30598 20576 31214
rect 20536 30592 20588 30598
rect 20536 30534 20588 30540
rect 20444 30252 20496 30258
rect 20444 30194 20496 30200
rect 20350 30152 20406 30161
rect 20350 30087 20352 30096
rect 20404 30087 20406 30096
rect 20352 30058 20404 30064
rect 20076 29844 20128 29850
rect 20076 29786 20128 29792
rect 20088 28121 20116 29786
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 20168 28960 20220 28966
rect 20168 28902 20220 28908
rect 20180 28218 20208 28902
rect 20260 28620 20312 28626
rect 20260 28562 20312 28568
rect 20168 28212 20220 28218
rect 20168 28154 20220 28160
rect 20074 28112 20130 28121
rect 19984 28076 20036 28082
rect 20074 28047 20130 28056
rect 19984 28018 20036 28024
rect 19996 24818 20024 28018
rect 20076 28008 20128 28014
rect 20076 27950 20128 27956
rect 20088 27674 20116 27950
rect 20180 27946 20208 28154
rect 20168 27940 20220 27946
rect 20168 27882 20220 27888
rect 20166 27840 20222 27849
rect 20166 27775 20222 27784
rect 20076 27668 20128 27674
rect 20076 27610 20128 27616
rect 20180 27554 20208 27775
rect 20272 27674 20300 28562
rect 20456 27962 20484 29446
rect 20364 27946 20484 27962
rect 20548 27946 20576 30534
rect 20364 27940 20496 27946
rect 20364 27934 20444 27940
rect 20260 27668 20312 27674
rect 20260 27610 20312 27616
rect 20364 27554 20392 27934
rect 20444 27882 20496 27888
rect 20536 27940 20588 27946
rect 20536 27882 20588 27888
rect 20548 27826 20576 27882
rect 20088 27526 20208 27554
rect 20272 27526 20392 27554
rect 20456 27798 20576 27826
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19996 24342 20024 24754
rect 19984 24336 20036 24342
rect 19984 24278 20036 24284
rect 19996 23526 20024 24278
rect 20088 23594 20116 27526
rect 20168 26784 20220 26790
rect 20168 26726 20220 26732
rect 20180 26042 20208 26726
rect 20272 26586 20300 27526
rect 20352 27464 20404 27470
rect 20352 27406 20404 27412
rect 20260 26580 20312 26586
rect 20260 26522 20312 26528
rect 20168 26036 20220 26042
rect 20168 25978 20220 25984
rect 20180 24682 20208 25978
rect 20168 24676 20220 24682
rect 20168 24618 20220 24624
rect 20076 23588 20128 23594
rect 20076 23530 20128 23536
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19996 22094 20024 23462
rect 19996 22066 20116 22094
rect 20088 21622 20116 22066
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 20076 21616 20128 21622
rect 20076 21558 20128 21564
rect 20076 21412 20128 21418
rect 20076 21354 20128 21360
rect 20088 20330 20116 21354
rect 20076 20324 20128 20330
rect 20076 20266 20128 20272
rect 20088 20058 20116 20266
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19996 18834 20024 19654
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19996 18358 20024 18770
rect 19984 18352 20036 18358
rect 19984 18294 20036 18300
rect 20076 17060 20128 17066
rect 20076 17002 20128 17008
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19996 16046 20024 16594
rect 20088 16454 20116 17002
rect 20180 16590 20208 21626
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20272 20806 20300 21286
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19996 15450 20024 15982
rect 20088 15570 20116 16390
rect 20168 16176 20220 16182
rect 20168 16118 20220 16124
rect 20180 15706 20208 16118
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 20272 15570 20300 15846
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 19996 15422 20208 15450
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 19996 13530 20024 13806
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19996 12442 20024 13466
rect 20180 13394 20208 15422
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19904 11614 20024 11642
rect 19484 11452 19780 11472
rect 19540 11450 19564 11452
rect 19620 11450 19644 11452
rect 19700 11450 19724 11452
rect 19562 11398 19564 11450
rect 19626 11398 19638 11450
rect 19700 11398 19702 11450
rect 19540 11396 19564 11398
rect 19620 11396 19644 11398
rect 19700 11396 19724 11398
rect 19484 11376 19780 11396
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 19812 10470 19840 11222
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19800 10464 19852 10470
rect 19800 10406 19852 10412
rect 19484 10364 19780 10384
rect 19540 10362 19564 10364
rect 19620 10362 19644 10364
rect 19700 10362 19724 10364
rect 19562 10310 19564 10362
rect 19626 10310 19638 10362
rect 19700 10310 19702 10362
rect 19540 10308 19564 10310
rect 19620 10308 19644 10310
rect 19700 10308 19724 10310
rect 19484 10288 19780 10308
rect 19812 10130 19840 10406
rect 19300 10084 19380 10112
rect 19800 10124 19852 10130
rect 19248 10066 19300 10072
rect 19800 10066 19852 10072
rect 19260 10010 19288 10066
rect 19168 9982 19288 10010
rect 18878 9415 18934 9424
rect 19064 9444 19116 9450
rect 18892 7750 18920 9415
rect 19064 9386 19116 9392
rect 18970 8936 19026 8945
rect 18970 8871 19026 8880
rect 18984 7886 19012 8871
rect 19168 8294 19196 9982
rect 19246 9888 19302 9897
rect 19246 9823 19302 9832
rect 19076 8266 19196 8294
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18800 6990 18920 7018
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18800 6458 18828 6802
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 18328 6180 18380 6186
rect 18328 6122 18380 6128
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18156 4690 18184 4966
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 18248 4146 18276 5646
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 17920 3488 18000 3516
rect 17868 3470 17920 3476
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 17328 2650 17356 2926
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 14852 2204 15148 2224
rect 14908 2202 14932 2204
rect 14988 2202 15012 2204
rect 15068 2202 15092 2204
rect 14930 2150 14932 2202
rect 14994 2150 15006 2202
rect 15068 2150 15070 2202
rect 14908 2148 14932 2150
rect 14988 2148 15012 2150
rect 15068 2148 15092 2150
rect 14852 2128 15148 2148
rect 15672 800 15700 2382
rect 16960 800 16988 2382
rect 18340 800 18368 5714
rect 18432 4622 18460 6054
rect 18616 5710 18644 6394
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 18708 5574 18736 6190
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18788 5092 18840 5098
rect 18788 5034 18840 5040
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18604 4208 18656 4214
rect 18604 4150 18656 4156
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 18432 2990 18460 4082
rect 18616 4078 18644 4150
rect 18800 4078 18828 5034
rect 18892 4690 18920 6990
rect 19076 6866 19104 8266
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 19260 5114 19288 9823
rect 19904 9518 19932 11086
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19352 7954 19380 9318
rect 19484 9276 19780 9296
rect 19540 9274 19564 9276
rect 19620 9274 19644 9276
rect 19700 9274 19724 9276
rect 19562 9222 19564 9274
rect 19626 9222 19638 9274
rect 19700 9222 19702 9274
rect 19540 9220 19564 9222
rect 19620 9220 19644 9222
rect 19700 9220 19724 9222
rect 19484 9200 19780 9220
rect 19904 8294 19932 9454
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 19484 8188 19780 8208
rect 19540 8186 19564 8188
rect 19620 8186 19644 8188
rect 19700 8186 19724 8188
rect 19562 8134 19564 8186
rect 19626 8134 19638 8186
rect 19700 8134 19702 8186
rect 19540 8132 19564 8134
rect 19620 8132 19644 8134
rect 19700 8132 19724 8134
rect 19484 8112 19780 8132
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19352 7274 19380 7686
rect 19340 7268 19392 7274
rect 19340 7210 19392 7216
rect 19352 6934 19380 7210
rect 19484 7100 19780 7120
rect 19540 7098 19564 7100
rect 19620 7098 19644 7100
rect 19700 7098 19724 7100
rect 19562 7046 19564 7098
rect 19626 7046 19638 7098
rect 19700 7046 19702 7098
rect 19540 7044 19564 7046
rect 19620 7044 19644 7046
rect 19700 7044 19724 7046
rect 19484 7024 19780 7044
rect 19340 6928 19392 6934
rect 19340 6870 19392 6876
rect 19800 6928 19852 6934
rect 19800 6870 19852 6876
rect 19812 6322 19840 6870
rect 19800 6316 19852 6322
rect 19800 6258 19852 6264
rect 19484 6012 19780 6032
rect 19540 6010 19564 6012
rect 19620 6010 19644 6012
rect 19700 6010 19724 6012
rect 19562 5958 19564 6010
rect 19626 5958 19638 6010
rect 19700 5958 19702 6010
rect 19540 5956 19564 5958
rect 19620 5956 19644 5958
rect 19700 5956 19724 5958
rect 19484 5936 19780 5956
rect 19904 5302 19932 7890
rect 19892 5296 19944 5302
rect 19892 5238 19944 5244
rect 19168 5086 19288 5114
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18880 4548 18932 4554
rect 18880 4490 18932 4496
rect 18892 4282 18920 4490
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 18880 4276 18932 4282
rect 18880 4218 18932 4224
rect 18892 4078 18920 4218
rect 19076 4078 19104 4422
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 18524 3670 18552 4014
rect 18512 3664 18564 3670
rect 18512 3606 18564 3612
rect 19168 3126 19196 5086
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19260 4758 19288 4966
rect 19248 4752 19300 4758
rect 19248 4694 19300 4700
rect 19260 3534 19288 4694
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19260 3398 19288 3470
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19156 3120 19208 3126
rect 19156 3062 19208 3068
rect 19352 2990 19380 4966
rect 19484 4924 19780 4944
rect 19540 4922 19564 4924
rect 19620 4922 19644 4924
rect 19700 4922 19724 4924
rect 19562 4870 19564 4922
rect 19626 4870 19638 4922
rect 19700 4870 19702 4922
rect 19540 4868 19564 4870
rect 19620 4868 19644 4870
rect 19700 4868 19724 4870
rect 19484 4848 19780 4868
rect 19708 4684 19760 4690
rect 19708 4626 19760 4632
rect 19720 4078 19748 4626
rect 19708 4072 19760 4078
rect 19708 4014 19760 4020
rect 19484 3836 19780 3856
rect 19540 3834 19564 3836
rect 19620 3834 19644 3836
rect 19700 3834 19724 3836
rect 19562 3782 19564 3834
rect 19626 3782 19638 3834
rect 19700 3782 19702 3834
rect 19540 3780 19564 3782
rect 19620 3780 19644 3782
rect 19700 3780 19724 3782
rect 19484 3760 19780 3780
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19484 2748 19780 2768
rect 19540 2746 19564 2748
rect 19620 2746 19644 2748
rect 19700 2746 19724 2748
rect 19562 2694 19564 2746
rect 19626 2694 19638 2746
rect 19700 2694 19702 2746
rect 19540 2692 19564 2694
rect 19620 2692 19644 2694
rect 19700 2692 19724 2694
rect 19484 2672 19780 2692
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 19352 2106 19380 2450
rect 19340 2100 19392 2106
rect 19340 2042 19392 2048
rect 19812 1442 19840 5102
rect 19892 4616 19944 4622
rect 19892 4558 19944 4564
rect 19904 3126 19932 4558
rect 19996 4554 20024 11614
rect 20180 11354 20208 13330
rect 20260 12368 20312 12374
rect 20258 12336 20260 12345
rect 20312 12336 20314 12345
rect 20258 12271 20314 12280
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20180 11150 20208 11290
rect 20168 11144 20220 11150
rect 20168 11086 20220 11092
rect 20168 8288 20220 8294
rect 20168 8230 20220 8236
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 20088 6934 20116 7142
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 20076 6248 20128 6254
rect 20180 6236 20208 8230
rect 20128 6208 20208 6236
rect 20076 6190 20128 6196
rect 20088 4758 20116 6190
rect 20168 5024 20220 5030
rect 20168 4966 20220 4972
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 19996 4214 20024 4490
rect 19984 4208 20036 4214
rect 19984 4150 20036 4156
rect 19984 4072 20036 4078
rect 19984 4014 20036 4020
rect 19996 3602 20024 4014
rect 20088 3738 20116 4558
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 19984 3596 20036 3602
rect 20036 3556 20116 3584
rect 19984 3538 20036 3544
rect 19892 3120 19944 3126
rect 19892 3062 19944 3068
rect 20088 2990 20116 3556
rect 20180 3058 20208 4966
rect 20364 3738 20392 27406
rect 20456 27010 20484 27798
rect 20536 27328 20588 27334
rect 20536 27270 20588 27276
rect 20548 27130 20576 27270
rect 20536 27124 20588 27130
rect 20536 27066 20588 27072
rect 20456 26982 20576 27010
rect 20444 24744 20496 24750
rect 20444 24686 20496 24692
rect 20456 24342 20484 24686
rect 20548 24682 20576 26982
rect 20536 24676 20588 24682
rect 20536 24618 20588 24624
rect 20444 24336 20496 24342
rect 20444 24278 20496 24284
rect 20444 22568 20496 22574
rect 20444 22510 20496 22516
rect 20456 20602 20484 22510
rect 20548 21418 20576 24618
rect 20536 21412 20588 21418
rect 20536 21354 20588 21360
rect 20548 21146 20576 21354
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20640 19938 20668 46854
rect 20916 46510 20944 46990
rect 21008 46646 21036 47058
rect 21192 47054 21220 48078
rect 21364 48068 21416 48074
rect 21364 48010 21416 48016
rect 21272 48000 21324 48006
rect 21272 47942 21324 47948
rect 21284 47666 21312 47942
rect 21272 47660 21324 47666
rect 21272 47602 21324 47608
rect 21272 47456 21324 47462
rect 21272 47398 21324 47404
rect 21284 47122 21312 47398
rect 21272 47116 21324 47122
rect 21272 47058 21324 47064
rect 21180 47048 21232 47054
rect 21180 46990 21232 46996
rect 21376 46986 21404 48010
rect 21364 46980 21416 46986
rect 21364 46922 21416 46928
rect 20996 46640 21048 46646
rect 20996 46582 21048 46588
rect 20904 46504 20956 46510
rect 20904 46446 20956 46452
rect 21456 45620 21508 45626
rect 21456 45562 21508 45568
rect 21180 45416 21232 45422
rect 21180 45358 21232 45364
rect 21192 44470 21220 45358
rect 21468 45354 21496 45562
rect 21456 45348 21508 45354
rect 21456 45290 21508 45296
rect 21560 45286 21588 49286
rect 21652 46186 21680 52906
rect 22008 52896 22060 52902
rect 22008 52838 22060 52844
rect 21824 51944 21876 51950
rect 21824 51886 21876 51892
rect 21836 51338 21864 51886
rect 21824 51332 21876 51338
rect 21824 51274 21876 51280
rect 21824 50720 21876 50726
rect 21824 50662 21876 50668
rect 21836 49978 21864 50662
rect 21916 50448 21968 50454
rect 21916 50390 21968 50396
rect 21928 49978 21956 50390
rect 21824 49972 21876 49978
rect 21824 49914 21876 49920
rect 21916 49972 21968 49978
rect 21916 49914 21968 49920
rect 21732 47456 21784 47462
rect 21732 47398 21784 47404
rect 21744 47190 21772 47398
rect 21732 47184 21784 47190
rect 21732 47126 21784 47132
rect 21652 46158 21772 46186
rect 21548 45280 21600 45286
rect 21548 45222 21600 45228
rect 21180 44464 21232 44470
rect 21180 44406 21232 44412
rect 20720 44328 20772 44334
rect 20720 44270 20772 44276
rect 21272 44328 21324 44334
rect 21272 44270 21324 44276
rect 20732 39642 20760 44270
rect 21284 44198 21312 44270
rect 21560 44198 21588 45222
rect 21640 44736 21692 44742
rect 21640 44678 21692 44684
rect 21272 44192 21324 44198
rect 21272 44134 21324 44140
rect 21548 44192 21600 44198
rect 21548 44134 21600 44140
rect 21364 43920 21416 43926
rect 21364 43862 21416 43868
rect 21456 43920 21508 43926
rect 21456 43862 21508 43868
rect 20996 43784 21048 43790
rect 20996 43726 21048 43732
rect 21008 41138 21036 43726
rect 21376 43450 21404 43862
rect 21364 43444 21416 43450
rect 21364 43386 21416 43392
rect 21468 43110 21496 43862
rect 21560 43790 21588 44134
rect 21548 43784 21600 43790
rect 21548 43726 21600 43732
rect 21456 43104 21508 43110
rect 21456 43046 21508 43052
rect 21456 41676 21508 41682
rect 21456 41618 21508 41624
rect 21088 41472 21140 41478
rect 21088 41414 21140 41420
rect 20996 41132 21048 41138
rect 20996 41074 21048 41080
rect 21100 39982 21128 41414
rect 21468 40934 21496 41618
rect 21456 40928 21508 40934
rect 21456 40870 21508 40876
rect 21468 40730 21496 40870
rect 21456 40724 21508 40730
rect 21456 40666 21508 40672
rect 21088 39976 21140 39982
rect 21088 39918 21140 39924
rect 20720 39636 20772 39642
rect 20720 39578 20772 39584
rect 20732 36718 20760 39578
rect 20904 38412 20956 38418
rect 21272 38412 21324 38418
rect 20956 38372 21036 38400
rect 20904 38354 20956 38360
rect 20812 37868 20864 37874
rect 20812 37810 20864 37816
rect 20720 36712 20772 36718
rect 20720 36654 20772 36660
rect 20824 35630 20852 37810
rect 20904 37392 20956 37398
rect 20904 37334 20956 37340
rect 20916 37126 20944 37334
rect 21008 37126 21036 38372
rect 21272 38354 21324 38360
rect 21088 38208 21140 38214
rect 21088 38150 21140 38156
rect 21100 37806 21128 38150
rect 21088 37800 21140 37806
rect 21088 37742 21140 37748
rect 21284 37398 21312 38354
rect 21364 38276 21416 38282
rect 21364 38218 21416 38224
rect 21376 37398 21404 38218
rect 21272 37392 21324 37398
rect 21272 37334 21324 37340
rect 21364 37392 21416 37398
rect 21364 37334 21416 37340
rect 21088 37324 21140 37330
rect 21088 37266 21140 37272
rect 20904 37120 20956 37126
rect 20904 37062 20956 37068
rect 20996 37120 21048 37126
rect 20996 37062 21048 37068
rect 20812 35624 20864 35630
rect 20812 35566 20864 35572
rect 20720 35556 20772 35562
rect 20720 35498 20772 35504
rect 20732 35222 20760 35498
rect 20720 35216 20772 35222
rect 21008 35170 21036 37062
rect 20720 35158 20772 35164
rect 20916 35142 21036 35170
rect 20720 33516 20772 33522
rect 20720 33458 20772 33464
rect 20732 32774 20760 33458
rect 20812 32904 20864 32910
rect 20812 32846 20864 32852
rect 20720 32768 20772 32774
rect 20720 32710 20772 32716
rect 20732 32366 20760 32710
rect 20824 32570 20852 32846
rect 20812 32564 20864 32570
rect 20812 32506 20864 32512
rect 20720 32360 20772 32366
rect 20720 32302 20772 32308
rect 20916 32212 20944 35142
rect 20996 35080 21048 35086
rect 20994 35048 20996 35057
rect 21048 35048 21050 35057
rect 20994 34983 21050 34992
rect 21100 34066 21128 37266
rect 21284 36718 21312 37334
rect 21272 36712 21324 36718
rect 21272 36654 21324 36660
rect 21180 36032 21232 36038
rect 21180 35974 21232 35980
rect 21192 35154 21220 35974
rect 21180 35148 21232 35154
rect 21180 35090 21232 35096
rect 21548 35148 21600 35154
rect 21548 35090 21600 35096
rect 20996 34060 21048 34066
rect 20996 34002 21048 34008
rect 21088 34060 21140 34066
rect 21088 34002 21140 34008
rect 20732 32184 20944 32212
rect 20732 26874 20760 32184
rect 21008 30802 21036 34002
rect 21192 33454 21220 35090
rect 21560 34134 21588 35090
rect 21548 34128 21600 34134
rect 21548 34070 21600 34076
rect 21180 33448 21232 33454
rect 21180 33390 21232 33396
rect 21548 33448 21600 33454
rect 21548 33390 21600 33396
rect 21088 32836 21140 32842
rect 21088 32778 21140 32784
rect 21100 32366 21128 32778
rect 21088 32360 21140 32366
rect 21088 32302 21140 32308
rect 21100 32026 21128 32302
rect 21088 32020 21140 32026
rect 21088 31962 21140 31968
rect 21180 32020 21232 32026
rect 21180 31962 21232 31968
rect 21192 31890 21220 31962
rect 21180 31884 21232 31890
rect 21180 31826 21232 31832
rect 21364 31884 21416 31890
rect 21560 31872 21588 33390
rect 21364 31826 21416 31832
rect 21468 31844 21588 31872
rect 21088 31816 21140 31822
rect 21086 31784 21088 31793
rect 21140 31784 21142 31793
rect 21086 31719 21142 31728
rect 21272 31680 21324 31686
rect 21272 31622 21324 31628
rect 20996 30796 21048 30802
rect 20996 30738 21048 30744
rect 21180 30796 21232 30802
rect 21180 30738 21232 30744
rect 20812 30660 20864 30666
rect 20812 30602 20864 30608
rect 20904 30660 20956 30666
rect 20904 30602 20956 30608
rect 20824 30326 20852 30602
rect 20812 30320 20864 30326
rect 20812 30262 20864 30268
rect 20812 30184 20864 30190
rect 20916 30172 20944 30602
rect 20996 30592 21048 30598
rect 20996 30534 21048 30540
rect 21008 30190 21036 30534
rect 20864 30144 20944 30172
rect 20996 30184 21048 30190
rect 20812 30126 20864 30132
rect 20996 30126 21048 30132
rect 20824 29850 20852 30126
rect 20812 29844 20864 29850
rect 20812 29786 20864 29792
rect 21088 27872 21140 27878
rect 21088 27814 21140 27820
rect 21192 27826 21220 30738
rect 21284 30598 21312 31622
rect 21376 31142 21404 31826
rect 21364 31136 21416 31142
rect 21364 31078 21416 31084
rect 21376 30870 21404 31078
rect 21364 30864 21416 30870
rect 21364 30806 21416 30812
rect 21272 30592 21324 30598
rect 21272 30534 21324 30540
rect 21468 30054 21496 31844
rect 21652 31754 21680 44678
rect 21744 32570 21772 46158
rect 21824 44328 21876 44334
rect 21824 44270 21876 44276
rect 21836 43790 21864 44270
rect 21824 43784 21876 43790
rect 21824 43726 21876 43732
rect 21824 43104 21876 43110
rect 21824 43046 21876 43052
rect 21836 42838 21864 43046
rect 21824 42832 21876 42838
rect 21824 42774 21876 42780
rect 21916 36576 21968 36582
rect 21916 36518 21968 36524
rect 21732 32564 21784 32570
rect 21732 32506 21784 32512
rect 21928 31754 21956 36518
rect 22020 33862 22048 52838
rect 22008 33856 22060 33862
rect 22008 33798 22060 33804
rect 22008 33312 22060 33318
rect 22008 33254 22060 33260
rect 22020 32434 22048 33254
rect 22112 32978 22140 52906
rect 22652 52896 22704 52902
rect 22652 52838 22704 52844
rect 22664 52698 22692 52838
rect 22652 52692 22704 52698
rect 22652 52634 22704 52640
rect 22848 52562 22876 53450
rect 23216 53242 23244 53518
rect 23204 53236 23256 53242
rect 23204 53178 23256 53184
rect 23296 53032 23348 53038
rect 23296 52974 23348 52980
rect 23308 52698 23336 52974
rect 23296 52692 23348 52698
rect 23296 52634 23348 52640
rect 22836 52556 22888 52562
rect 22836 52498 22888 52504
rect 22928 52080 22980 52086
rect 22928 52022 22980 52028
rect 22560 51876 22612 51882
rect 22560 51818 22612 51824
rect 22572 51610 22600 51818
rect 22940 51610 22968 52022
rect 23388 51808 23440 51814
rect 23388 51750 23440 51756
rect 22560 51604 22612 51610
rect 22560 51546 22612 51552
rect 22928 51604 22980 51610
rect 22928 51546 22980 51552
rect 23112 51604 23164 51610
rect 23112 51546 23164 51552
rect 22376 51468 22428 51474
rect 22376 51410 22428 51416
rect 22388 51270 22416 51410
rect 23020 51400 23072 51406
rect 22466 51368 22522 51377
rect 23020 51342 23072 51348
rect 22466 51303 22522 51312
rect 22376 51264 22428 51270
rect 22376 51206 22428 51212
rect 22480 50998 22508 51303
rect 23032 51074 23060 51342
rect 22664 51046 23060 51074
rect 23124 51066 23152 51546
rect 23112 51060 23164 51066
rect 22468 50992 22520 50998
rect 22468 50934 22520 50940
rect 22192 50856 22244 50862
rect 22192 50798 22244 50804
rect 22204 50522 22232 50798
rect 22284 50788 22336 50794
rect 22284 50730 22336 50736
rect 22192 50516 22244 50522
rect 22192 50458 22244 50464
rect 22204 48618 22232 50458
rect 22296 50250 22324 50730
rect 22560 50380 22612 50386
rect 22560 50322 22612 50328
rect 22284 50244 22336 50250
rect 22284 50186 22336 50192
rect 22572 49230 22600 50322
rect 22664 49994 22692 51046
rect 23112 51002 23164 51008
rect 23204 51060 23256 51066
rect 23204 51002 23256 51008
rect 23216 50810 23244 51002
rect 23400 50862 23428 51750
rect 23584 50998 23612 55247
rect 23754 55200 23810 56800
rect 25226 55720 25282 55729
rect 25226 55655 25282 55664
rect 23768 53242 23796 55200
rect 25134 54904 25190 54913
rect 25134 54839 25190 54848
rect 25042 54088 25098 54097
rect 25042 54023 25098 54032
rect 25056 53922 25084 54023
rect 24032 53916 24084 53922
rect 24032 53858 24084 53864
rect 25044 53916 25096 53922
rect 25044 53858 25096 53864
rect 23756 53236 23808 53242
rect 23756 53178 23808 53184
rect 24044 53106 24072 53858
rect 24860 53508 24912 53514
rect 24860 53450 24912 53456
rect 24116 53340 24412 53360
rect 24172 53338 24196 53340
rect 24252 53338 24276 53340
rect 24332 53338 24356 53340
rect 24194 53286 24196 53338
rect 24258 53286 24270 53338
rect 24332 53286 24334 53338
rect 24172 53284 24196 53286
rect 24252 53284 24276 53286
rect 24332 53284 24356 53286
rect 24116 53264 24412 53284
rect 24872 53281 24900 53450
rect 24858 53272 24914 53281
rect 24858 53207 24914 53216
rect 24032 53100 24084 53106
rect 24032 53042 24084 53048
rect 24860 53100 24912 53106
rect 24860 53042 24912 53048
rect 24584 53032 24636 53038
rect 24872 52986 24900 53042
rect 24584 52974 24636 52980
rect 23756 52964 23808 52970
rect 23756 52906 23808 52912
rect 23572 50992 23624 50998
rect 23572 50934 23624 50940
rect 23480 50924 23532 50930
rect 23480 50866 23532 50872
rect 22940 50782 23244 50810
rect 23388 50856 23440 50862
rect 23388 50798 23440 50804
rect 22940 50726 22968 50782
rect 22928 50720 22980 50726
rect 22928 50662 22980 50668
rect 23112 50720 23164 50726
rect 23492 50708 23520 50866
rect 23112 50662 23164 50668
rect 23216 50680 23520 50708
rect 22756 50238 22968 50266
rect 22756 50182 22784 50238
rect 22744 50176 22796 50182
rect 22744 50118 22796 50124
rect 22664 49966 22876 49994
rect 22652 49768 22704 49774
rect 22652 49710 22704 49716
rect 22664 49314 22692 49710
rect 22848 49706 22876 49966
rect 22940 49774 22968 50238
rect 23020 50176 23072 50182
rect 23020 50118 23072 50124
rect 23032 49842 23060 50118
rect 23020 49836 23072 49842
rect 23020 49778 23072 49784
rect 22928 49768 22980 49774
rect 22928 49710 22980 49716
rect 22836 49700 22888 49706
rect 22836 49642 22888 49648
rect 22744 49632 22796 49638
rect 22744 49574 22796 49580
rect 22756 49434 22784 49574
rect 22744 49428 22796 49434
rect 22744 49370 22796 49376
rect 22664 49286 22784 49314
rect 22560 49224 22612 49230
rect 22560 49166 22612 49172
rect 22756 48618 22784 49286
rect 22848 48686 22876 49642
rect 23124 49434 23152 50662
rect 23216 50522 23244 50680
rect 23204 50516 23256 50522
rect 23204 50458 23256 50464
rect 23572 50380 23624 50386
rect 23572 50322 23624 50328
rect 23112 49428 23164 49434
rect 23112 49370 23164 49376
rect 22928 49224 22980 49230
rect 22928 49166 22980 49172
rect 22836 48680 22888 48686
rect 22836 48622 22888 48628
rect 22192 48612 22244 48618
rect 22192 48554 22244 48560
rect 22744 48612 22796 48618
rect 22744 48554 22796 48560
rect 22204 45898 22232 48554
rect 22560 47116 22612 47122
rect 22560 47058 22612 47064
rect 22192 45892 22244 45898
rect 22192 45834 22244 45840
rect 22204 44810 22232 45834
rect 22572 45558 22600 47058
rect 22560 45552 22612 45558
rect 22560 45494 22612 45500
rect 22572 45422 22600 45494
rect 22560 45416 22612 45422
rect 22560 45358 22612 45364
rect 22756 44946 22784 48554
rect 22848 48142 22876 48622
rect 22836 48136 22888 48142
rect 22836 48078 22888 48084
rect 22560 44940 22612 44946
rect 22560 44882 22612 44888
rect 22744 44940 22796 44946
rect 22744 44882 22796 44888
rect 22192 44804 22244 44810
rect 22192 44746 22244 44752
rect 22204 43738 22232 44746
rect 22204 43710 22508 43738
rect 22296 43314 22324 43710
rect 22376 43648 22428 43654
rect 22376 43590 22428 43596
rect 22284 43308 22336 43314
rect 22284 43250 22336 43256
rect 22284 43104 22336 43110
rect 22284 43046 22336 43052
rect 22296 42770 22324 43046
rect 22284 42764 22336 42770
rect 22284 42706 22336 42712
rect 22192 42696 22244 42702
rect 22192 42638 22244 42644
rect 22204 42362 22232 42638
rect 22192 42356 22244 42362
rect 22192 42298 22244 42304
rect 22388 42226 22416 43590
rect 22376 42220 22428 42226
rect 22376 42162 22428 42168
rect 22192 42152 22244 42158
rect 22192 42094 22244 42100
rect 22204 41070 22232 42094
rect 22192 41064 22244 41070
rect 22192 41006 22244 41012
rect 22192 40928 22244 40934
rect 22192 40870 22244 40876
rect 22204 40050 22232 40870
rect 22480 40118 22508 43710
rect 22468 40112 22520 40118
rect 22468 40054 22520 40060
rect 22192 40044 22244 40050
rect 22192 39986 22244 39992
rect 22284 39092 22336 39098
rect 22336 39052 22508 39080
rect 22284 39034 22336 39040
rect 22480 38962 22508 39052
rect 22468 38956 22520 38962
rect 22468 38898 22520 38904
rect 22192 38344 22244 38350
rect 22192 38286 22244 38292
rect 22204 38010 22232 38286
rect 22192 38004 22244 38010
rect 22192 37946 22244 37952
rect 22572 36564 22600 44882
rect 22756 42158 22784 44882
rect 22744 42152 22796 42158
rect 22744 42094 22796 42100
rect 22652 39840 22704 39846
rect 22652 39782 22704 39788
rect 22664 39642 22692 39782
rect 22652 39636 22704 39642
rect 22652 39578 22704 39584
rect 22652 38888 22704 38894
rect 22652 38830 22704 38836
rect 22664 38282 22692 38830
rect 22744 38752 22796 38758
rect 22744 38694 22796 38700
rect 22652 38276 22704 38282
rect 22652 38218 22704 38224
rect 22296 36536 22600 36564
rect 22192 34468 22244 34474
rect 22192 34410 22244 34416
rect 22100 32972 22152 32978
rect 22100 32914 22152 32920
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 22100 32360 22152 32366
rect 21560 31726 21680 31754
rect 21836 31726 21956 31754
rect 22020 32308 22100 32314
rect 22020 32302 22152 32308
rect 22020 32286 22140 32302
rect 21456 30048 21508 30054
rect 21456 29990 21508 29996
rect 21272 28756 21324 28762
rect 21272 28698 21324 28704
rect 21284 27946 21312 28698
rect 21364 28416 21416 28422
rect 21364 28358 21416 28364
rect 21376 28014 21404 28358
rect 21364 28008 21416 28014
rect 21364 27950 21416 27956
rect 21272 27940 21324 27946
rect 21272 27882 21324 27888
rect 21100 27538 21128 27814
rect 21192 27798 21404 27826
rect 21088 27532 21140 27538
rect 21088 27474 21140 27480
rect 20732 26846 21128 26874
rect 20904 25152 20956 25158
rect 20904 25094 20956 25100
rect 20916 24750 20944 25094
rect 20904 24744 20956 24750
rect 20904 24686 20956 24692
rect 20720 24608 20772 24614
rect 20720 24550 20772 24556
rect 20732 23798 20760 24550
rect 20720 23792 20772 23798
rect 20720 23734 20772 23740
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20732 22098 20760 22374
rect 20720 22092 20772 22098
rect 20720 22034 20772 22040
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20732 21146 20760 22034
rect 20720 21140 20772 21146
rect 20720 21082 20772 21088
rect 20824 21026 20852 22034
rect 21008 22030 21036 23598
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20916 21418 20944 21830
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 20904 21412 20956 21418
rect 20904 21354 20956 21360
rect 21008 21078 21036 21422
rect 20996 21072 21048 21078
rect 20824 21010 20944 21026
rect 20996 21014 21048 21020
rect 20824 21004 20956 21010
rect 20824 20998 20904 21004
rect 20904 20946 20956 20952
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20456 19910 20668 19938
rect 20456 13190 20484 19910
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20548 19310 20576 19790
rect 20536 19304 20588 19310
rect 20720 19304 20772 19310
rect 20536 19246 20588 19252
rect 20626 19272 20682 19281
rect 20720 19246 20772 19252
rect 20626 19207 20682 19216
rect 20640 19174 20668 19207
rect 20628 19168 20680 19174
rect 20628 19110 20680 19116
rect 20732 18222 20760 19246
rect 20824 18426 20852 20878
rect 20916 19174 20944 20946
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20916 18698 20944 19110
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20902 18592 20958 18601
rect 20902 18527 20958 18536
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20536 17332 20588 17338
rect 20536 17274 20588 17280
rect 20548 15434 20576 17274
rect 20824 16726 20852 18362
rect 20916 18222 20944 18527
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 20916 17338 20944 18158
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 21008 17270 21036 20334
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 21100 17202 21128 26846
rect 21272 25764 21324 25770
rect 21272 25706 21324 25712
rect 21180 24268 21232 24274
rect 21180 24210 21232 24216
rect 21192 23662 21220 24210
rect 21284 23866 21312 25706
rect 21376 24206 21404 27798
rect 21454 27568 21510 27577
rect 21454 27503 21510 27512
rect 21468 27402 21496 27503
rect 21456 27396 21508 27402
rect 21456 27338 21508 27344
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 21364 24200 21416 24206
rect 21364 24142 21416 24148
rect 21272 23860 21324 23866
rect 21272 23802 21324 23808
rect 21272 23724 21324 23730
rect 21272 23666 21324 23672
rect 21180 23656 21232 23662
rect 21180 23598 21232 23604
rect 21192 21146 21220 23598
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21192 18222 21220 19110
rect 21284 18698 21312 23666
rect 21468 22506 21496 24550
rect 21364 22500 21416 22506
rect 21364 22442 21416 22448
rect 21456 22500 21508 22506
rect 21456 22442 21508 22448
rect 21376 20466 21404 22442
rect 21560 22094 21588 31726
rect 21640 31680 21692 31686
rect 21640 31622 21692 31628
rect 21732 31680 21784 31686
rect 21732 31622 21784 31628
rect 21652 31346 21680 31622
rect 21744 31414 21772 31622
rect 21732 31408 21784 31414
rect 21732 31350 21784 31356
rect 21640 31340 21692 31346
rect 21640 31282 21692 31288
rect 21732 30184 21784 30190
rect 21730 30152 21732 30161
rect 21784 30152 21786 30161
rect 21730 30087 21786 30096
rect 21640 27872 21692 27878
rect 21640 27814 21692 27820
rect 21732 27872 21784 27878
rect 21732 27814 21784 27820
rect 21652 24274 21680 27814
rect 21744 27674 21772 27814
rect 21732 27668 21784 27674
rect 21732 27610 21784 27616
rect 21836 25430 21864 31726
rect 21916 31204 21968 31210
rect 21916 31146 21968 31152
rect 21928 30734 21956 31146
rect 21916 30728 21968 30734
rect 21916 30670 21968 30676
rect 21916 26784 21968 26790
rect 21916 26726 21968 26732
rect 21824 25424 21876 25430
rect 21824 25366 21876 25372
rect 21836 24818 21864 25366
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21928 24750 21956 26726
rect 21916 24744 21968 24750
rect 21916 24686 21968 24692
rect 21732 24676 21784 24682
rect 21732 24618 21784 24624
rect 21640 24268 21692 24274
rect 21640 24210 21692 24216
rect 21652 22574 21680 24210
rect 21744 23730 21772 24618
rect 21928 24206 21956 24686
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21916 24200 21968 24206
rect 21916 24142 21968 24148
rect 21732 23724 21784 23730
rect 21732 23666 21784 23672
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21732 22432 21784 22438
rect 21732 22374 21784 22380
rect 21744 22166 21772 22374
rect 21732 22160 21784 22166
rect 21732 22102 21784 22108
rect 21468 22066 21588 22094
rect 21640 22092 21692 22098
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21376 19514 21404 20402
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21376 18698 21404 19450
rect 21272 18692 21324 18698
rect 21272 18634 21324 18640
rect 21364 18692 21416 18698
rect 21364 18634 21416 18640
rect 21284 18426 21312 18634
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21180 18216 21232 18222
rect 21180 18158 21232 18164
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20916 16590 20944 17138
rect 21192 17082 21220 18158
rect 21272 18148 21324 18154
rect 21272 18090 21324 18096
rect 21100 17054 21220 17082
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20732 15978 20760 16390
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20548 13938 20576 15370
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20732 13734 20760 14418
rect 20916 14414 20944 16526
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 20824 13870 20852 14282
rect 21008 14074 21036 16594
rect 21100 14618 21128 17054
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21192 16726 21220 16934
rect 21180 16720 21232 16726
rect 21180 16662 21232 16668
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 21100 13938 21128 14554
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20732 13530 20760 13670
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20444 13184 20496 13190
rect 20444 13126 20496 13132
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20548 11898 20576 12106
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20732 11694 20760 13466
rect 20824 13258 20852 13806
rect 20812 13252 20864 13258
rect 20812 13194 20864 13200
rect 20824 12434 20852 13194
rect 21008 13190 21036 13806
rect 21100 13394 21128 13874
rect 21192 13870 21220 14418
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 20824 12406 20944 12434
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20640 11286 20668 11494
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20732 10130 20760 11630
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20456 9042 20484 9862
rect 20732 9110 20760 10066
rect 20824 10062 20852 12174
rect 20916 11558 20944 12406
rect 21008 11694 21036 13126
rect 21100 12442 21128 13330
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21192 12918 21220 13262
rect 21180 12912 21232 12918
rect 21180 12854 21232 12860
rect 21284 12730 21312 18090
rect 21364 17264 21416 17270
rect 21364 17206 21416 17212
rect 21376 12782 21404 17206
rect 21192 12702 21312 12730
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 21192 12238 21220 12702
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21284 12356 21312 12582
rect 21468 12434 21496 22066
rect 21640 22034 21692 22040
rect 21652 20482 21680 22034
rect 21744 21690 21772 22102
rect 21732 21684 21784 21690
rect 21732 21626 21784 21632
rect 21744 21078 21772 21626
rect 21732 21072 21784 21078
rect 21732 21014 21784 21020
rect 21560 20454 21680 20482
rect 21560 19378 21588 20454
rect 21640 20392 21692 20398
rect 21744 20380 21772 21014
rect 21692 20352 21772 20380
rect 21640 20334 21692 20340
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21548 19372 21600 19378
rect 21548 19314 21600 19320
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 21560 18902 21588 19110
rect 21548 18896 21600 18902
rect 21744 18873 21772 19382
rect 21548 18838 21600 18844
rect 21730 18864 21786 18873
rect 21640 18828 21692 18834
rect 21730 18799 21786 18808
rect 21640 18770 21692 18776
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21560 14958 21588 18362
rect 21652 17882 21680 18770
rect 21732 18692 21784 18698
rect 21732 18634 21784 18640
rect 21744 18290 21772 18634
rect 21732 18284 21784 18290
rect 21732 18226 21784 18232
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 21640 17264 21692 17270
rect 21640 17206 21692 17212
rect 21652 16250 21680 17206
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 21652 15638 21680 16186
rect 21640 15632 21692 15638
rect 21640 15574 21692 15580
rect 21548 14952 21600 14958
rect 21548 14894 21600 14900
rect 21732 14952 21784 14958
rect 21732 14894 21784 14900
rect 21548 13796 21600 13802
rect 21548 13738 21600 13744
rect 21560 13394 21588 13738
rect 21744 13530 21772 14894
rect 21732 13524 21784 13530
rect 21732 13466 21784 13472
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21468 12406 21588 12434
rect 21364 12368 21416 12374
rect 21284 12328 21364 12356
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20812 9920 20864 9926
rect 20916 9908 20944 11494
rect 20864 9880 20944 9908
rect 20812 9862 20864 9868
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20536 7336 20588 7342
rect 20536 7278 20588 7284
rect 20548 6866 20576 7278
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 20732 4826 20760 7890
rect 20824 7546 20852 9862
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20916 7342 20944 9386
rect 21008 7818 21036 11630
rect 21284 11218 21312 12328
rect 21364 12310 21416 12316
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21376 11694 21404 12038
rect 21468 11762 21496 12038
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21560 10538 21588 12406
rect 21180 10532 21232 10538
rect 21180 10474 21232 10480
rect 21548 10532 21600 10538
rect 21548 10474 21600 10480
rect 21192 10130 21220 10474
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 21180 10124 21232 10130
rect 21180 10066 21232 10072
rect 21100 7954 21128 10066
rect 21836 9602 21864 24142
rect 21916 22024 21968 22030
rect 21916 21966 21968 21972
rect 21928 19378 21956 21966
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 21928 15162 21956 19314
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 21928 14618 21956 15098
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 21916 14408 21968 14414
rect 21916 14350 21968 14356
rect 21928 12306 21956 14350
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 21928 9722 21956 10406
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 21836 9574 21956 9602
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 21836 9382 21864 9454
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21836 8498 21864 9318
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21088 7948 21140 7954
rect 21088 7890 21140 7896
rect 20996 7812 21048 7818
rect 20996 7754 21048 7760
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 21008 6798 21036 7754
rect 20996 6792 21048 6798
rect 20996 6734 21048 6740
rect 21088 6724 21140 6730
rect 21088 6666 21140 6672
rect 21100 6458 21128 6666
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21376 5914 21404 6054
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21732 5228 21784 5234
rect 21732 5170 21784 5176
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 20628 4548 20680 4554
rect 20628 4490 20680 4496
rect 20640 3942 20668 4490
rect 21008 4078 21036 4558
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 20996 4072 21048 4078
rect 20996 4014 21048 4020
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 19996 2650 20024 2926
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 20364 2553 20392 3674
rect 21100 2990 21128 4422
rect 21088 2984 21140 2990
rect 21088 2926 21140 2932
rect 21192 2774 21220 5102
rect 21640 4684 21692 4690
rect 21640 4626 21692 4632
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 21560 4282 21588 4558
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21560 2854 21588 4218
rect 21652 3738 21680 4626
rect 21640 3732 21692 3738
rect 21640 3674 21692 3680
rect 21364 2848 21416 2854
rect 21100 2746 21220 2774
rect 21362 2816 21364 2825
rect 21548 2848 21600 2854
rect 21416 2816 21418 2825
rect 21548 2790 21600 2796
rect 21744 2774 21772 5170
rect 21928 4486 21956 9574
rect 22020 4758 22048 32286
rect 22204 31890 22232 34410
rect 22192 31884 22244 31890
rect 22192 31826 22244 31832
rect 22100 31680 22152 31686
rect 22100 31622 22152 31628
rect 22112 30394 22140 31622
rect 22100 30388 22152 30394
rect 22100 30330 22152 30336
rect 22296 26314 22324 36536
rect 22664 36038 22692 38218
rect 22756 37874 22784 38694
rect 22744 37868 22796 37874
rect 22744 37810 22796 37816
rect 22744 37324 22796 37330
rect 22744 37266 22796 37272
rect 22756 36378 22784 37266
rect 22744 36372 22796 36378
rect 22744 36314 22796 36320
rect 22652 36032 22704 36038
rect 22652 35974 22704 35980
rect 22744 36032 22796 36038
rect 22744 35974 22796 35980
rect 22664 35766 22692 35974
rect 22652 35760 22704 35766
rect 22652 35702 22704 35708
rect 22468 35148 22520 35154
rect 22468 35090 22520 35096
rect 22376 35012 22428 35018
rect 22376 34954 22428 34960
rect 22388 32910 22416 34954
rect 22480 34542 22508 35090
rect 22756 34746 22784 35974
rect 22744 34740 22796 34746
rect 22744 34682 22796 34688
rect 22468 34536 22520 34542
rect 22468 34478 22520 34484
rect 22480 34406 22508 34478
rect 22468 34400 22520 34406
rect 22468 34342 22520 34348
rect 22480 33998 22508 34342
rect 22468 33992 22520 33998
rect 22468 33934 22520 33940
rect 22848 32994 22876 48078
rect 22940 46560 22968 49166
rect 23204 49088 23256 49094
rect 23204 49030 23256 49036
rect 23216 48686 23244 49030
rect 23204 48680 23256 48686
rect 23204 48622 23256 48628
rect 23216 48210 23244 48622
rect 23204 48204 23256 48210
rect 23204 48146 23256 48152
rect 23388 46912 23440 46918
rect 23388 46854 23440 46860
rect 23204 46640 23256 46646
rect 23204 46582 23256 46588
rect 23020 46572 23072 46578
rect 22940 46532 23020 46560
rect 23020 46514 23072 46520
rect 23032 45354 23060 46514
rect 23216 46458 23244 46582
rect 23216 46430 23336 46458
rect 23112 46368 23164 46374
rect 23112 46310 23164 46316
rect 23204 46368 23256 46374
rect 23204 46310 23256 46316
rect 23020 45348 23072 45354
rect 23020 45290 23072 45296
rect 23032 44962 23060 45290
rect 23124 45082 23152 46310
rect 23216 46170 23244 46310
rect 23204 46164 23256 46170
rect 23204 46106 23256 46112
rect 23112 45076 23164 45082
rect 23112 45018 23164 45024
rect 23032 44934 23244 44962
rect 23308 44946 23336 46430
rect 23400 46170 23428 46854
rect 23388 46164 23440 46170
rect 23388 46106 23440 46112
rect 23480 45960 23532 45966
rect 23480 45902 23532 45908
rect 23388 45280 23440 45286
rect 23388 45222 23440 45228
rect 23020 43444 23072 43450
rect 23020 43386 23072 43392
rect 23032 43246 23060 43386
rect 23020 43240 23072 43246
rect 23020 43182 23072 43188
rect 23216 42702 23244 44934
rect 23296 44940 23348 44946
rect 23296 44882 23348 44888
rect 23400 44878 23428 45222
rect 23388 44872 23440 44878
rect 23388 44814 23440 44820
rect 23492 44470 23520 45902
rect 23480 44464 23532 44470
rect 23480 44406 23532 44412
rect 23388 43852 23440 43858
rect 23388 43794 23440 43800
rect 23400 42838 23428 43794
rect 23492 43790 23520 44406
rect 23584 44402 23612 50322
rect 23664 47252 23716 47258
rect 23664 47194 23716 47200
rect 23572 44396 23624 44402
rect 23572 44338 23624 44344
rect 23572 44260 23624 44266
rect 23572 44202 23624 44208
rect 23480 43784 23532 43790
rect 23480 43726 23532 43732
rect 23584 43330 23612 44202
rect 23492 43302 23612 43330
rect 23388 42832 23440 42838
rect 23388 42774 23440 42780
rect 23204 42696 23256 42702
rect 23204 42638 23256 42644
rect 23020 42220 23072 42226
rect 23020 42162 23072 42168
rect 23032 41070 23060 42162
rect 23020 41064 23072 41070
rect 23020 41006 23072 41012
rect 23032 38026 23060 41006
rect 23216 39982 23244 42638
rect 23296 42560 23348 42566
rect 23296 42502 23348 42508
rect 23308 42158 23336 42502
rect 23296 42152 23348 42158
rect 23296 42094 23348 42100
rect 23308 41138 23336 42094
rect 23296 41132 23348 41138
rect 23296 41074 23348 41080
rect 23204 39976 23256 39982
rect 23204 39918 23256 39924
rect 23492 38654 23520 43302
rect 23676 41682 23704 47194
rect 23664 41676 23716 41682
rect 23664 41618 23716 41624
rect 23676 41414 23704 41618
rect 23584 41386 23704 41414
rect 23584 39846 23612 41386
rect 23664 41132 23716 41138
rect 23664 41074 23716 41080
rect 23676 41002 23704 41074
rect 23664 40996 23716 41002
rect 23664 40938 23716 40944
rect 23676 40594 23704 40938
rect 23664 40588 23716 40594
rect 23664 40530 23716 40536
rect 23676 39982 23704 40530
rect 23664 39976 23716 39982
rect 23664 39918 23716 39924
rect 23572 39840 23624 39846
rect 23572 39782 23624 39788
rect 23676 39658 23704 39918
rect 23308 38626 23520 38654
rect 23584 39630 23704 39658
rect 23112 38208 23164 38214
rect 23112 38150 23164 38156
rect 23204 38208 23256 38214
rect 23204 38150 23256 38156
rect 22480 32966 22876 32994
rect 22940 37998 23060 38026
rect 22376 32904 22428 32910
rect 22376 32846 22428 32852
rect 22388 32570 22416 32846
rect 22376 32564 22428 32570
rect 22376 32506 22428 32512
rect 22480 32450 22508 32966
rect 22836 32904 22888 32910
rect 22836 32846 22888 32852
rect 22652 32564 22704 32570
rect 22652 32506 22704 32512
rect 22388 32422 22508 32450
rect 22388 29238 22416 32422
rect 22558 32328 22614 32337
rect 22558 32263 22614 32272
rect 22572 31958 22600 32263
rect 22664 32201 22692 32506
rect 22650 32192 22706 32201
rect 22650 32127 22706 32136
rect 22560 31952 22612 31958
rect 22560 31894 22612 31900
rect 22468 31748 22520 31754
rect 22468 31690 22520 31696
rect 22480 31278 22508 31690
rect 22664 31686 22692 32127
rect 22744 31884 22796 31890
rect 22744 31826 22796 31832
rect 22652 31680 22704 31686
rect 22652 31622 22704 31628
rect 22468 31272 22520 31278
rect 22468 31214 22520 31220
rect 22652 31272 22704 31278
rect 22652 31214 22704 31220
rect 22480 30138 22508 31214
rect 22664 30666 22692 31214
rect 22652 30660 22704 30666
rect 22652 30602 22704 30608
rect 22480 30110 22600 30138
rect 22468 30048 22520 30054
rect 22468 29990 22520 29996
rect 22376 29232 22428 29238
rect 22376 29174 22428 29180
rect 22480 27470 22508 29990
rect 22572 27606 22600 30110
rect 22756 30036 22784 31826
rect 22848 31482 22876 32846
rect 22940 31754 22968 37998
rect 23124 37806 23152 38150
rect 23112 37800 23164 37806
rect 23112 37742 23164 37748
rect 23216 37126 23244 38150
rect 23020 37120 23072 37126
rect 23020 37062 23072 37068
rect 23204 37120 23256 37126
rect 23204 37062 23256 37068
rect 23032 35766 23060 37062
rect 23112 36236 23164 36242
rect 23112 36178 23164 36184
rect 23204 36236 23256 36242
rect 23204 36178 23256 36184
rect 23020 35760 23072 35766
rect 23020 35702 23072 35708
rect 23032 35018 23060 35702
rect 23124 35698 23152 36178
rect 23216 35873 23244 36178
rect 23202 35864 23258 35873
rect 23202 35799 23258 35808
rect 23216 35766 23244 35799
rect 23204 35760 23256 35766
rect 23204 35702 23256 35708
rect 23112 35692 23164 35698
rect 23112 35634 23164 35640
rect 23124 35290 23152 35634
rect 23112 35284 23164 35290
rect 23112 35226 23164 35232
rect 23204 35148 23256 35154
rect 23204 35090 23256 35096
rect 23020 35012 23072 35018
rect 23020 34954 23072 34960
rect 23112 33992 23164 33998
rect 23112 33934 23164 33940
rect 23020 32768 23072 32774
rect 23020 32710 23072 32716
rect 23032 32570 23060 32710
rect 23020 32564 23072 32570
rect 23020 32506 23072 32512
rect 23124 32026 23152 33934
rect 23112 32020 23164 32026
rect 23112 31962 23164 31968
rect 22940 31726 23152 31754
rect 22928 31680 22980 31686
rect 22928 31622 22980 31628
rect 22836 31476 22888 31482
rect 22836 31418 22888 31424
rect 22940 30190 22968 31622
rect 23020 30796 23072 30802
rect 23020 30738 23072 30744
rect 23032 30394 23060 30738
rect 23020 30388 23072 30394
rect 23020 30330 23072 30336
rect 22928 30184 22980 30190
rect 22928 30126 22980 30132
rect 22756 30008 23060 30036
rect 22928 29232 22980 29238
rect 22928 29174 22980 29180
rect 22940 28422 22968 29174
rect 22928 28416 22980 28422
rect 22928 28358 22980 28364
rect 22940 27606 22968 28358
rect 22560 27600 22612 27606
rect 22560 27542 22612 27548
rect 22928 27600 22980 27606
rect 22928 27542 22980 27548
rect 22468 27464 22520 27470
rect 22468 27406 22520 27412
rect 22480 26994 22508 27406
rect 22468 26988 22520 26994
rect 22468 26930 22520 26936
rect 22284 26308 22336 26314
rect 22284 26250 22336 26256
rect 22284 25356 22336 25362
rect 22284 25298 22336 25304
rect 22100 25220 22152 25226
rect 22100 25162 22152 25168
rect 22112 24138 22140 25162
rect 22296 24886 22324 25298
rect 22284 24880 22336 24886
rect 22284 24822 22336 24828
rect 22296 24682 22324 24822
rect 22284 24676 22336 24682
rect 22284 24618 22336 24624
rect 22480 24154 22508 26930
rect 22572 26874 22600 27542
rect 23032 27418 23060 30008
rect 22848 27390 23060 27418
rect 22572 26858 22692 26874
rect 22572 26852 22704 26858
rect 22572 26846 22652 26852
rect 22652 26794 22704 26800
rect 22664 26314 22692 26794
rect 22652 26308 22704 26314
rect 22652 26250 22704 26256
rect 22560 25696 22612 25702
rect 22560 25638 22612 25644
rect 22572 24274 22600 25638
rect 22744 25356 22796 25362
rect 22744 25298 22796 25304
rect 22652 24676 22704 24682
rect 22652 24618 22704 24624
rect 22664 24274 22692 24618
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 22100 24132 22152 24138
rect 22480 24126 22600 24154
rect 22100 24074 22152 24080
rect 22112 20942 22140 24074
rect 22192 22704 22244 22710
rect 22192 22646 22244 22652
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 22100 12912 22152 12918
rect 22100 12854 22152 12860
rect 22112 10674 22140 12854
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 22112 7410 22140 10610
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22008 4752 22060 4758
rect 22008 4694 22060 4700
rect 21916 4480 21968 4486
rect 21916 4422 21968 4428
rect 21928 3670 21956 4422
rect 22204 4146 22232 22646
rect 22468 22160 22520 22166
rect 22468 22102 22520 22108
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 22284 21412 22336 21418
rect 22284 21354 22336 21360
rect 22296 20466 22324 21354
rect 22388 20534 22416 21422
rect 22480 20806 22508 22102
rect 22572 22030 22600 24126
rect 22652 24064 22704 24070
rect 22652 24006 22704 24012
rect 22664 23662 22692 24006
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22756 22710 22784 25298
rect 22744 22704 22796 22710
rect 22744 22646 22796 22652
rect 22744 22160 22796 22166
rect 22744 22102 22796 22108
rect 22560 22024 22612 22030
rect 22612 21984 22692 22012
rect 22560 21966 22612 21972
rect 22560 21412 22612 21418
rect 22560 21354 22612 21360
rect 22572 21146 22600 21354
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22468 20800 22520 20806
rect 22468 20742 22520 20748
rect 22376 20528 22428 20534
rect 22376 20470 22428 20476
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22388 20074 22416 20470
rect 22296 20046 22416 20074
rect 22296 18290 22324 20046
rect 22664 18766 22692 21984
rect 22756 21350 22784 22102
rect 22744 21344 22796 21350
rect 22744 21286 22796 21292
rect 22744 18896 22796 18902
rect 22744 18838 22796 18844
rect 22652 18760 22704 18766
rect 22756 18737 22784 18838
rect 22652 18702 22704 18708
rect 22742 18728 22798 18737
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22388 18222 22416 18566
rect 22376 18216 22428 18222
rect 22376 18158 22428 18164
rect 22664 17354 22692 18702
rect 22742 18663 22798 18672
rect 22572 17326 22692 17354
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22296 16250 22324 16458
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22572 16114 22600 17326
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22560 16108 22612 16114
rect 22560 16050 22612 16056
rect 22284 15904 22336 15910
rect 22284 15846 22336 15852
rect 22296 15502 22324 15846
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22480 13870 22508 14758
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22296 12714 22324 12922
rect 22572 12850 22600 16050
rect 22664 16046 22692 16526
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22744 15972 22796 15978
rect 22744 15914 22796 15920
rect 22756 15570 22784 15914
rect 22744 15564 22796 15570
rect 22744 15506 22796 15512
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22664 14618 22692 14894
rect 22652 14612 22704 14618
rect 22652 14554 22704 14560
rect 22652 14476 22704 14482
rect 22652 14418 22704 14424
rect 22664 14074 22692 14418
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22284 12708 22336 12714
rect 22284 12650 22336 12656
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22572 12442 22600 12582
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22572 11694 22600 12378
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 22560 11688 22612 11694
rect 22560 11630 22612 11636
rect 22756 11558 22784 11766
rect 22744 11552 22796 11558
rect 22744 11494 22796 11500
rect 22560 11008 22612 11014
rect 22560 10950 22612 10956
rect 22284 10600 22336 10606
rect 22284 10542 22336 10548
rect 22296 7342 22324 10542
rect 22572 10470 22600 10950
rect 22652 10532 22704 10538
rect 22652 10474 22704 10480
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22664 9518 22692 10474
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 22664 9110 22692 9454
rect 22652 9104 22704 9110
rect 22652 9046 22704 9052
rect 22756 8974 22784 11494
rect 22744 8968 22796 8974
rect 22744 8910 22796 8916
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22480 7206 22508 7754
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22572 6254 22600 7686
rect 22560 6248 22612 6254
rect 22560 6190 22612 6196
rect 22744 6112 22796 6118
rect 22744 6054 22796 6060
rect 22468 5092 22520 5098
rect 22468 5034 22520 5040
rect 22376 4752 22428 4758
rect 22376 4694 22428 4700
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 21916 3664 21968 3670
rect 21916 3606 21968 3612
rect 22388 3126 22416 4694
rect 22480 3942 22508 5034
rect 22756 4690 22784 6054
rect 22848 5370 22876 27390
rect 23020 26852 23072 26858
rect 23020 26794 23072 26800
rect 23032 26518 23060 26794
rect 23020 26512 23072 26518
rect 23020 26454 23072 26460
rect 23032 25702 23060 26454
rect 23020 25696 23072 25702
rect 23020 25638 23072 25644
rect 23032 25430 23060 25638
rect 23020 25424 23072 25430
rect 23020 25366 23072 25372
rect 22928 25152 22980 25158
rect 22928 25094 22980 25100
rect 23020 25152 23072 25158
rect 23020 25094 23072 25100
rect 22940 24682 22968 25094
rect 22928 24676 22980 24682
rect 22928 24618 22980 24624
rect 23032 24410 23060 25094
rect 23020 24404 23072 24410
rect 23020 24346 23072 24352
rect 23124 22778 23152 31726
rect 23216 30122 23244 35090
rect 23308 33998 23336 38626
rect 23388 36236 23440 36242
rect 23388 36178 23440 36184
rect 23400 36038 23428 36178
rect 23584 36122 23612 39630
rect 23664 39500 23716 39506
rect 23664 39442 23716 39448
rect 23676 39302 23704 39442
rect 23664 39296 23716 39302
rect 23664 39238 23716 39244
rect 23492 36094 23612 36122
rect 23664 36168 23716 36174
rect 23664 36110 23716 36116
rect 23388 36032 23440 36038
rect 23388 35974 23440 35980
rect 23388 35148 23440 35154
rect 23388 35090 23440 35096
rect 23400 34610 23428 35090
rect 23388 34604 23440 34610
rect 23388 34546 23440 34552
rect 23400 34066 23428 34546
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 23296 33992 23348 33998
rect 23296 33934 23348 33940
rect 23294 32464 23350 32473
rect 23492 32450 23520 36094
rect 23572 34400 23624 34406
rect 23572 34342 23624 34348
rect 23294 32399 23350 32408
rect 23400 32422 23520 32450
rect 23308 32298 23336 32399
rect 23296 32292 23348 32298
rect 23296 32234 23348 32240
rect 23296 31816 23348 31822
rect 23296 31758 23348 31764
rect 23400 31770 23428 32422
rect 23584 31890 23612 34342
rect 23676 33454 23704 36110
rect 23664 33448 23716 33454
rect 23664 33390 23716 33396
rect 23768 32570 23796 52906
rect 24492 52488 24544 52494
rect 24492 52430 24544 52436
rect 24116 52252 24412 52272
rect 24172 52250 24196 52252
rect 24252 52250 24276 52252
rect 24332 52250 24356 52252
rect 24194 52198 24196 52250
rect 24258 52198 24270 52250
rect 24332 52198 24334 52250
rect 24172 52196 24196 52198
rect 24252 52196 24276 52198
rect 24332 52196 24356 52198
rect 24116 52176 24412 52196
rect 23848 52080 23900 52086
rect 23848 52022 23900 52028
rect 23860 50454 23888 52022
rect 24504 51950 24532 52430
rect 24596 52057 24624 52974
rect 24688 52958 24900 52986
rect 24688 52902 24716 52958
rect 24676 52896 24728 52902
rect 24676 52838 24728 52844
rect 24768 52896 24820 52902
rect 24768 52838 24820 52844
rect 24858 52864 24914 52873
rect 24676 52556 24728 52562
rect 24676 52498 24728 52504
rect 24688 52465 24716 52498
rect 24674 52456 24730 52465
rect 24674 52391 24730 52400
rect 24582 52048 24638 52057
rect 24582 51983 24638 51992
rect 24492 51944 24544 51950
rect 24492 51886 24544 51892
rect 23940 51876 23992 51882
rect 23940 51818 23992 51824
rect 23952 51474 23980 51818
rect 23940 51468 23992 51474
rect 23940 51410 23992 51416
rect 24032 51468 24084 51474
rect 24032 51410 24084 51416
rect 23940 51264 23992 51270
rect 23940 51206 23992 51212
rect 23952 51066 23980 51206
rect 23940 51060 23992 51066
rect 23940 51002 23992 51008
rect 24044 50522 24072 51410
rect 24116 51164 24412 51184
rect 24172 51162 24196 51164
rect 24252 51162 24276 51164
rect 24332 51162 24356 51164
rect 24194 51110 24196 51162
rect 24258 51110 24270 51162
rect 24332 51110 24334 51162
rect 24172 51108 24196 51110
rect 24252 51108 24276 51110
rect 24332 51108 24356 51110
rect 24116 51088 24412 51108
rect 24124 50720 24176 50726
rect 24124 50662 24176 50668
rect 24032 50516 24084 50522
rect 24032 50458 24084 50464
rect 23848 50448 23900 50454
rect 23848 50390 23900 50396
rect 24136 50386 24164 50662
rect 24676 50448 24728 50454
rect 24780 50436 24808 52838
rect 24858 52799 24914 52808
rect 24872 52630 24900 52799
rect 24860 52624 24912 52630
rect 24860 52566 24912 52572
rect 25044 52556 25096 52562
rect 25044 52498 25096 52504
rect 25056 51649 25084 52498
rect 25042 51640 25098 51649
rect 25042 51575 25098 51584
rect 24728 50408 24808 50436
rect 24950 50416 25006 50425
rect 24676 50390 24728 50396
rect 24124 50380 24176 50386
rect 24950 50351 24952 50360
rect 24124 50322 24176 50328
rect 25004 50351 25006 50360
rect 24952 50322 25004 50328
rect 24768 50312 24820 50318
rect 24768 50254 24820 50260
rect 24116 50076 24412 50096
rect 24172 50074 24196 50076
rect 24252 50074 24276 50076
rect 24332 50074 24356 50076
rect 24194 50022 24196 50074
rect 24258 50022 24270 50074
rect 24332 50022 24334 50074
rect 24172 50020 24196 50022
rect 24252 50020 24276 50022
rect 24332 50020 24356 50022
rect 24116 50000 24412 50020
rect 23848 49768 23900 49774
rect 24032 49768 24084 49774
rect 23848 49710 23900 49716
rect 23952 49716 24032 49722
rect 23952 49710 24084 49716
rect 23860 49298 23888 49710
rect 23952 49694 24072 49710
rect 23848 49292 23900 49298
rect 23848 49234 23900 49240
rect 23860 48006 23888 49234
rect 23952 49230 23980 49694
rect 24032 49632 24084 49638
rect 24032 49574 24084 49580
rect 23940 49224 23992 49230
rect 23940 49166 23992 49172
rect 23952 48618 23980 49166
rect 24044 48754 24072 49574
rect 24676 49292 24728 49298
rect 24676 49234 24728 49240
rect 24116 48988 24412 49008
rect 24172 48986 24196 48988
rect 24252 48986 24276 48988
rect 24332 48986 24356 48988
rect 24194 48934 24196 48986
rect 24258 48934 24270 48986
rect 24332 48934 24334 48986
rect 24172 48932 24196 48934
rect 24252 48932 24276 48934
rect 24332 48932 24356 48934
rect 24116 48912 24412 48932
rect 24032 48748 24084 48754
rect 24032 48690 24084 48696
rect 24688 48686 24716 49234
rect 24780 48822 24808 50254
rect 25148 50250 25176 54839
rect 25136 50244 25188 50250
rect 25136 50186 25188 50192
rect 25136 49904 25188 49910
rect 25136 49846 25188 49852
rect 24860 49292 24912 49298
rect 24860 49234 24912 49240
rect 24768 48816 24820 48822
rect 24768 48758 24820 48764
rect 24676 48680 24728 48686
rect 24872 48634 24900 49234
rect 24676 48622 24728 48628
rect 23940 48612 23992 48618
rect 23940 48554 23992 48560
rect 24032 48612 24084 48618
rect 24032 48554 24084 48560
rect 24780 48606 24900 48634
rect 23952 48278 23980 48554
rect 23940 48272 23992 48278
rect 23940 48214 23992 48220
rect 24044 48210 24072 48554
rect 24780 48550 24808 48606
rect 24584 48544 24636 48550
rect 24584 48486 24636 48492
rect 24768 48544 24820 48550
rect 24768 48486 24820 48492
rect 24596 48346 24624 48486
rect 24584 48340 24636 48346
rect 25148 48314 25176 49846
rect 24584 48282 24636 48288
rect 25056 48286 25176 48314
rect 24032 48204 24084 48210
rect 24032 48146 24084 48152
rect 24492 48204 24544 48210
rect 24492 48146 24544 48152
rect 23848 48000 23900 48006
rect 23848 47942 23900 47948
rect 23940 48000 23992 48006
rect 23940 47942 23992 47948
rect 23860 47598 23888 47942
rect 23952 47802 23980 47942
rect 23940 47796 23992 47802
rect 23940 47738 23992 47744
rect 23848 47592 23900 47598
rect 23848 47534 23900 47540
rect 24044 47258 24072 48146
rect 24116 47900 24412 47920
rect 24172 47898 24196 47900
rect 24252 47898 24276 47900
rect 24332 47898 24356 47900
rect 24194 47846 24196 47898
rect 24258 47846 24270 47898
rect 24332 47846 24334 47898
rect 24172 47844 24196 47846
rect 24252 47844 24276 47846
rect 24332 47844 24356 47846
rect 24116 47824 24412 47844
rect 24504 47802 24532 48146
rect 24492 47796 24544 47802
rect 24492 47738 24544 47744
rect 24032 47252 24084 47258
rect 24032 47194 24084 47200
rect 24308 47116 24360 47122
rect 24360 47076 24532 47104
rect 24308 47058 24360 47064
rect 24116 46812 24412 46832
rect 24172 46810 24196 46812
rect 24252 46810 24276 46812
rect 24332 46810 24356 46812
rect 24194 46758 24196 46810
rect 24258 46758 24270 46810
rect 24332 46758 24334 46810
rect 24172 46756 24196 46758
rect 24252 46756 24276 46758
rect 24332 46756 24356 46758
rect 24116 46736 24412 46756
rect 23848 46504 23900 46510
rect 23848 46446 23900 46452
rect 23860 45286 23888 46446
rect 24504 46374 24532 47076
rect 24492 46368 24544 46374
rect 24492 46310 24544 46316
rect 24032 46028 24084 46034
rect 24032 45970 24084 45976
rect 23940 45348 23992 45354
rect 23940 45290 23992 45296
rect 23848 45280 23900 45286
rect 23848 45222 23900 45228
rect 23952 45014 23980 45290
rect 24044 45014 24072 45970
rect 24116 45724 24412 45744
rect 24172 45722 24196 45724
rect 24252 45722 24276 45724
rect 24332 45722 24356 45724
rect 24194 45670 24196 45722
rect 24258 45670 24270 45722
rect 24332 45670 24334 45722
rect 24172 45668 24196 45670
rect 24252 45668 24276 45670
rect 24332 45668 24356 45670
rect 24116 45648 24412 45668
rect 24504 45490 24532 46310
rect 24596 46170 24624 48282
rect 24676 48136 24728 48142
rect 24676 48078 24728 48084
rect 24584 46164 24636 46170
rect 24584 46106 24636 46112
rect 24584 46028 24636 46034
rect 24584 45970 24636 45976
rect 24596 45558 24624 45970
rect 24584 45552 24636 45558
rect 24584 45494 24636 45500
rect 24492 45484 24544 45490
rect 24492 45426 24544 45432
rect 24124 45416 24176 45422
rect 24124 45358 24176 45364
rect 24136 45082 24164 45358
rect 24308 45280 24360 45286
rect 24308 45222 24360 45228
rect 24124 45076 24176 45082
rect 24124 45018 24176 45024
rect 24320 45014 24348 45222
rect 23940 45008 23992 45014
rect 23940 44950 23992 44956
rect 24032 45008 24084 45014
rect 24032 44950 24084 44956
rect 24308 45008 24360 45014
rect 24308 44950 24360 44956
rect 23940 44804 23992 44810
rect 23940 44746 23992 44752
rect 23952 44538 23980 44746
rect 23940 44532 23992 44538
rect 23940 44474 23992 44480
rect 23848 44396 23900 44402
rect 23848 44338 23900 44344
rect 23860 43926 23888 44338
rect 24044 44282 24072 44950
rect 24320 44724 24348 44950
rect 24320 44696 24532 44724
rect 24116 44636 24412 44656
rect 24172 44634 24196 44636
rect 24252 44634 24276 44636
rect 24332 44634 24356 44636
rect 24194 44582 24196 44634
rect 24258 44582 24270 44634
rect 24332 44582 24334 44634
rect 24172 44580 24196 44582
rect 24252 44580 24276 44582
rect 24332 44580 24356 44582
rect 24116 44560 24412 44580
rect 24504 44402 24532 44696
rect 24492 44396 24544 44402
rect 24492 44338 24544 44344
rect 23952 44254 24072 44282
rect 23952 44198 23980 44254
rect 23940 44192 23992 44198
rect 23940 44134 23992 44140
rect 23848 43920 23900 43926
rect 23848 43862 23900 43868
rect 23860 43654 23888 43862
rect 23848 43648 23900 43654
rect 23848 43590 23900 43596
rect 23848 42764 23900 42770
rect 23848 42706 23900 42712
rect 23860 42226 23888 42706
rect 23848 42220 23900 42226
rect 23848 42162 23900 42168
rect 23952 41546 23980 44134
rect 24116 43548 24412 43568
rect 24172 43546 24196 43548
rect 24252 43546 24276 43548
rect 24332 43546 24356 43548
rect 24194 43494 24196 43546
rect 24258 43494 24270 43546
rect 24332 43494 24334 43546
rect 24172 43492 24196 43494
rect 24252 43492 24276 43494
rect 24332 43492 24356 43494
rect 24116 43472 24412 43492
rect 24032 42764 24084 42770
rect 24032 42706 24084 42712
rect 24044 42362 24072 42706
rect 24492 42696 24544 42702
rect 24492 42638 24544 42644
rect 24116 42460 24412 42480
rect 24172 42458 24196 42460
rect 24252 42458 24276 42460
rect 24332 42458 24356 42460
rect 24194 42406 24196 42458
rect 24258 42406 24270 42458
rect 24332 42406 24334 42458
rect 24172 42404 24196 42406
rect 24252 42404 24276 42406
rect 24332 42404 24356 42406
rect 24116 42384 24412 42404
rect 24032 42356 24084 42362
rect 24032 42298 24084 42304
rect 24504 41682 24532 42638
rect 24124 41676 24176 41682
rect 24124 41618 24176 41624
rect 24492 41676 24544 41682
rect 24492 41618 24544 41624
rect 24136 41562 24164 41618
rect 23940 41540 23992 41546
rect 23940 41482 23992 41488
rect 24044 41534 24164 41562
rect 23848 41064 23900 41070
rect 23848 41006 23900 41012
rect 23860 40594 23888 41006
rect 24044 40662 24072 41534
rect 24116 41372 24412 41392
rect 24172 41370 24196 41372
rect 24252 41370 24276 41372
rect 24332 41370 24356 41372
rect 24194 41318 24196 41370
rect 24258 41318 24270 41370
rect 24332 41318 24334 41370
rect 24172 41316 24196 41318
rect 24252 41316 24276 41318
rect 24332 41316 24356 41318
rect 24116 41296 24412 41316
rect 24032 40656 24084 40662
rect 24032 40598 24084 40604
rect 23848 40588 23900 40594
rect 23848 40530 23900 40536
rect 23860 40050 23888 40530
rect 24044 40066 24072 40598
rect 24492 40520 24544 40526
rect 24492 40462 24544 40468
rect 24116 40284 24412 40304
rect 24172 40282 24196 40284
rect 24252 40282 24276 40284
rect 24332 40282 24356 40284
rect 24194 40230 24196 40282
rect 24258 40230 24270 40282
rect 24332 40230 24334 40282
rect 24172 40228 24196 40230
rect 24252 40228 24276 40230
rect 24332 40228 24356 40230
rect 24116 40208 24412 40228
rect 23848 40044 23900 40050
rect 24044 40038 24256 40066
rect 23848 39986 23900 39992
rect 24228 39982 24256 40038
rect 24216 39976 24268 39982
rect 24216 39918 24268 39924
rect 24228 39506 24256 39918
rect 24504 39914 24532 40462
rect 24492 39908 24544 39914
rect 24492 39850 24544 39856
rect 24400 39840 24452 39846
rect 24400 39782 24452 39788
rect 24216 39500 24268 39506
rect 24216 39442 24268 39448
rect 24412 39438 24440 39782
rect 24400 39432 24452 39438
rect 24400 39374 24452 39380
rect 24504 39302 24532 39850
rect 24492 39296 24544 39302
rect 24492 39238 24544 39244
rect 24116 39196 24412 39216
rect 24172 39194 24196 39196
rect 24252 39194 24276 39196
rect 24332 39194 24356 39196
rect 24194 39142 24196 39194
rect 24258 39142 24270 39194
rect 24332 39142 24334 39194
rect 24172 39140 24196 39142
rect 24252 39140 24276 39142
rect 24332 39140 24356 39142
rect 24116 39120 24412 39140
rect 24116 38108 24412 38128
rect 24172 38106 24196 38108
rect 24252 38106 24276 38108
rect 24332 38106 24356 38108
rect 24194 38054 24196 38106
rect 24258 38054 24270 38106
rect 24332 38054 24334 38106
rect 24172 38052 24196 38054
rect 24252 38052 24276 38054
rect 24332 38052 24356 38054
rect 24116 38032 24412 38052
rect 24032 37800 24084 37806
rect 24032 37742 24084 37748
rect 24044 37126 24072 37742
rect 24032 37120 24084 37126
rect 24032 37062 24084 37068
rect 24044 36174 24072 37062
rect 24116 37020 24412 37040
rect 24172 37018 24196 37020
rect 24252 37018 24276 37020
rect 24332 37018 24356 37020
rect 24194 36966 24196 37018
rect 24258 36966 24270 37018
rect 24332 36966 24334 37018
rect 24172 36964 24196 36966
rect 24252 36964 24276 36966
rect 24332 36964 24356 36966
rect 24116 36944 24412 36964
rect 24032 36168 24084 36174
rect 24032 36110 24084 36116
rect 24116 35932 24412 35952
rect 24172 35930 24196 35932
rect 24252 35930 24276 35932
rect 24332 35930 24356 35932
rect 24194 35878 24196 35930
rect 24258 35878 24270 35930
rect 24332 35878 24334 35930
rect 24172 35876 24196 35878
rect 24252 35876 24276 35878
rect 24332 35876 24356 35878
rect 24116 35856 24412 35876
rect 24400 35692 24452 35698
rect 24400 35634 24452 35640
rect 23848 35624 23900 35630
rect 23848 35566 23900 35572
rect 23860 34610 23888 35566
rect 24412 35154 24440 35634
rect 24216 35148 24268 35154
rect 24216 35090 24268 35096
rect 24400 35148 24452 35154
rect 24400 35090 24452 35096
rect 24228 35018 24256 35090
rect 24216 35012 24268 35018
rect 24216 34954 24268 34960
rect 24116 34844 24412 34864
rect 24172 34842 24196 34844
rect 24252 34842 24276 34844
rect 24332 34842 24356 34844
rect 24194 34790 24196 34842
rect 24258 34790 24270 34842
rect 24332 34790 24334 34842
rect 24172 34788 24196 34790
rect 24252 34788 24276 34790
rect 24332 34788 24356 34790
rect 24116 34768 24412 34788
rect 23848 34604 23900 34610
rect 23848 34546 23900 34552
rect 24504 33998 24532 39238
rect 24584 35624 24636 35630
rect 24584 35566 24636 35572
rect 24596 35290 24624 35566
rect 24584 35284 24636 35290
rect 24584 35226 24636 35232
rect 24584 35148 24636 35154
rect 24584 35090 24636 35096
rect 24596 34746 24624 35090
rect 24584 34740 24636 34746
rect 24584 34682 24636 34688
rect 24688 34626 24716 48078
rect 25056 47054 25084 48286
rect 25044 47048 25096 47054
rect 25044 46990 25096 46996
rect 24860 46028 24912 46034
rect 24860 45970 24912 45976
rect 24768 44736 24820 44742
rect 24872 44724 24900 45970
rect 24820 44696 24900 44724
rect 24768 44678 24820 44684
rect 24872 44402 24900 44696
rect 24952 44736 25004 44742
rect 24952 44678 25004 44684
rect 24860 44396 24912 44402
rect 24860 44338 24912 44344
rect 24860 44260 24912 44266
rect 24860 44202 24912 44208
rect 24872 43994 24900 44202
rect 24860 43988 24912 43994
rect 24860 43930 24912 43936
rect 24964 43926 24992 44678
rect 24952 43920 25004 43926
rect 24952 43862 25004 43868
rect 24858 43480 24914 43489
rect 24858 43415 24914 43424
rect 24872 43246 24900 43415
rect 24860 43240 24912 43246
rect 24860 43182 24912 43188
rect 24952 41064 25004 41070
rect 24952 41006 25004 41012
rect 24860 40588 24912 40594
rect 24860 40530 24912 40536
rect 24872 39438 24900 40530
rect 24860 39432 24912 39438
rect 24860 39374 24912 39380
rect 24860 38208 24912 38214
rect 24860 38150 24912 38156
rect 24872 35698 24900 38150
rect 24860 35692 24912 35698
rect 24860 35634 24912 35640
rect 24872 35442 24900 35634
rect 24780 35414 24900 35442
rect 24780 35154 24808 35414
rect 24860 35284 24912 35290
rect 24860 35226 24912 35232
rect 24768 35148 24820 35154
rect 24768 35090 24820 35096
rect 24872 35018 24900 35226
rect 24860 35012 24912 35018
rect 24860 34954 24912 34960
rect 24596 34598 24716 34626
rect 24492 33992 24544 33998
rect 24492 33934 24544 33940
rect 24492 33856 24544 33862
rect 24492 33798 24544 33804
rect 24116 33756 24412 33776
rect 24172 33754 24196 33756
rect 24252 33754 24276 33756
rect 24332 33754 24356 33756
rect 24194 33702 24196 33754
rect 24258 33702 24270 33754
rect 24332 33702 24334 33754
rect 24172 33700 24196 33702
rect 24252 33700 24276 33702
rect 24332 33700 24356 33702
rect 24116 33680 24412 33700
rect 23848 33584 23900 33590
rect 23846 33552 23848 33561
rect 24400 33584 24452 33590
rect 23900 33552 23902 33561
rect 24400 33526 24452 33532
rect 23846 33487 23902 33496
rect 24308 33448 24360 33454
rect 24308 33390 24360 33396
rect 23848 33380 23900 33386
rect 23848 33322 23900 33328
rect 23940 33380 23992 33386
rect 23940 33322 23992 33328
rect 23860 32910 23888 33322
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 23952 32774 23980 33322
rect 24032 33312 24084 33318
rect 24032 33254 24084 33260
rect 23940 32768 23992 32774
rect 23940 32710 23992 32716
rect 23756 32564 23808 32570
rect 23756 32506 23808 32512
rect 23664 32360 23716 32366
rect 23664 32302 23716 32308
rect 23572 31884 23624 31890
rect 23572 31826 23624 31832
rect 23308 30326 23336 31758
rect 23400 31742 23520 31770
rect 23388 31680 23440 31686
rect 23388 31622 23440 31628
rect 23400 30802 23428 31622
rect 23388 30796 23440 30802
rect 23388 30738 23440 30744
rect 23296 30320 23348 30326
rect 23296 30262 23348 30268
rect 23204 30116 23256 30122
rect 23204 30058 23256 30064
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 22928 22636 22980 22642
rect 22928 22578 22980 22584
rect 22940 21146 22968 22578
rect 23112 22160 23164 22166
rect 23112 22102 23164 22108
rect 22928 21140 22980 21146
rect 22928 21082 22980 21088
rect 22928 21004 22980 21010
rect 22928 20946 22980 20952
rect 22940 20602 22968 20946
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 23032 20482 23060 20878
rect 22940 20454 23060 20482
rect 22940 17762 22968 20454
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 23032 18834 23060 19110
rect 23124 18834 23152 22102
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 23112 18828 23164 18834
rect 23112 18770 23164 18776
rect 22940 17746 23060 17762
rect 22940 17740 23072 17746
rect 22940 17734 23020 17740
rect 23020 17682 23072 17688
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 22940 13258 22968 15982
rect 23032 14482 23060 17682
rect 23124 16590 23152 18770
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 23112 16040 23164 16046
rect 23112 15982 23164 15988
rect 23124 15638 23152 15982
rect 23112 15632 23164 15638
rect 23112 15574 23164 15580
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 22928 13252 22980 13258
rect 22928 13194 22980 13200
rect 22940 10606 22968 13194
rect 23032 12434 23060 14418
rect 23112 13252 23164 13258
rect 23112 13194 23164 13200
rect 23124 12782 23152 13194
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 23032 12406 23152 12434
rect 22928 10600 22980 10606
rect 22928 10542 22980 10548
rect 22928 7948 22980 7954
rect 22928 7890 22980 7896
rect 22940 6730 22968 7890
rect 23124 7886 23152 12406
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 23112 7880 23164 7886
rect 23112 7822 23164 7828
rect 23032 6866 23060 7822
rect 23112 7268 23164 7274
rect 23112 7210 23164 7216
rect 23124 7002 23152 7210
rect 23112 6996 23164 7002
rect 23112 6938 23164 6944
rect 23020 6860 23072 6866
rect 23020 6802 23072 6808
rect 22928 6724 22980 6730
rect 22928 6666 22980 6672
rect 23032 6118 23060 6802
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 22836 5364 22888 5370
rect 22836 5306 22888 5312
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 22468 3936 22520 3942
rect 22652 3936 22704 3942
rect 22468 3878 22520 3884
rect 22572 3884 22652 3890
rect 22572 3878 22704 3884
rect 22480 3534 22508 3878
rect 22572 3862 22692 3878
rect 22572 3602 22600 3862
rect 22756 3618 22784 4626
rect 22848 4282 22876 5306
rect 23112 4752 23164 4758
rect 23112 4694 23164 4700
rect 23020 4548 23072 4554
rect 23020 4490 23072 4496
rect 22836 4276 22888 4282
rect 22836 4218 22888 4224
rect 22560 3596 22612 3602
rect 22756 3590 22876 3618
rect 22560 3538 22612 3544
rect 22848 3534 22876 3590
rect 22928 3596 22980 3602
rect 22928 3538 22980 3544
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 22940 3126 22968 3538
rect 23032 3126 23060 4490
rect 23124 4146 23152 4694
rect 23216 4162 23244 30058
rect 23388 27872 23440 27878
rect 23388 27814 23440 27820
rect 23294 27704 23350 27713
rect 23294 27639 23350 27648
rect 23308 27538 23336 27639
rect 23296 27532 23348 27538
rect 23296 27474 23348 27480
rect 23296 26308 23348 26314
rect 23296 26250 23348 26256
rect 23308 22166 23336 26250
rect 23400 25294 23428 27814
rect 23388 25288 23440 25294
rect 23388 25230 23440 25236
rect 23400 24954 23428 25230
rect 23388 24948 23440 24954
rect 23388 24890 23440 24896
rect 23296 22160 23348 22166
rect 23492 22137 23520 31742
rect 23572 27872 23624 27878
rect 23572 27814 23624 27820
rect 23584 27606 23612 27814
rect 23572 27600 23624 27606
rect 23572 27542 23624 27548
rect 23572 27056 23624 27062
rect 23570 27024 23572 27033
rect 23624 27024 23626 27033
rect 23570 26959 23626 26968
rect 23584 24138 23612 26959
rect 23572 24132 23624 24138
rect 23572 24074 23624 24080
rect 23572 22160 23624 22166
rect 23296 22102 23348 22108
rect 23478 22128 23534 22137
rect 23572 22102 23624 22108
rect 23478 22063 23534 22072
rect 23386 21992 23442 22001
rect 23386 21927 23442 21936
rect 23296 21412 23348 21418
rect 23296 21354 23348 21360
rect 23308 20534 23336 21354
rect 23296 20528 23348 20534
rect 23296 20470 23348 20476
rect 23400 19854 23428 21927
rect 23584 21690 23612 22102
rect 23572 21684 23624 21690
rect 23572 21626 23624 21632
rect 23584 21146 23612 21626
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23572 20936 23624 20942
rect 23572 20878 23624 20884
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 23480 19304 23532 19310
rect 23480 19246 23532 19252
rect 23492 18834 23520 19246
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23492 18358 23520 18770
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23492 17814 23520 18294
rect 23480 17808 23532 17814
rect 23480 17750 23532 17756
rect 23584 16658 23612 20878
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23584 16250 23612 16594
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23480 15428 23532 15434
rect 23480 15370 23532 15376
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 23308 12782 23336 14010
rect 23296 12776 23348 12782
rect 23296 12718 23348 12724
rect 23388 12708 23440 12714
rect 23388 12650 23440 12656
rect 23400 12374 23428 12650
rect 23388 12368 23440 12374
rect 23388 12310 23440 12316
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23296 12164 23348 12170
rect 23296 12106 23348 12112
rect 23308 11762 23336 12106
rect 23400 11898 23428 12174
rect 23388 11892 23440 11898
rect 23388 11834 23440 11840
rect 23296 11756 23348 11762
rect 23296 11698 23348 11704
rect 23388 10192 23440 10198
rect 23388 10134 23440 10140
rect 23400 9586 23428 10134
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 23400 7954 23428 8978
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 23400 7546 23428 7890
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23492 5114 23520 15370
rect 23584 13326 23612 16186
rect 23572 13320 23624 13326
rect 23572 13262 23624 13268
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23584 10674 23612 11086
rect 23572 10668 23624 10674
rect 23572 10610 23624 10616
rect 23584 10130 23612 10610
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23584 6798 23612 9522
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23400 5086 23520 5114
rect 23400 4622 23428 5086
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 23216 4146 23336 4162
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 23216 4140 23348 4146
rect 23216 4134 23296 4140
rect 23216 3942 23244 4134
rect 23296 4082 23348 4088
rect 23492 4078 23520 4966
rect 23676 4758 23704 32302
rect 23848 32224 23900 32230
rect 23848 32166 23900 32172
rect 23756 31884 23808 31890
rect 23756 31826 23808 31832
rect 23768 5166 23796 31826
rect 23860 31686 23888 32166
rect 23952 31754 23980 32710
rect 24044 32298 24072 33254
rect 24320 32842 24348 33390
rect 24308 32836 24360 32842
rect 24308 32778 24360 32784
rect 24412 32756 24440 33526
rect 24504 33522 24532 33798
rect 24492 33516 24544 33522
rect 24492 33458 24544 33464
rect 24492 32972 24544 32978
rect 24492 32914 24544 32920
rect 24504 32881 24532 32914
rect 24490 32872 24546 32881
rect 24490 32807 24546 32816
rect 24412 32728 24532 32756
rect 24116 32668 24412 32688
rect 24172 32666 24196 32668
rect 24252 32666 24276 32668
rect 24332 32666 24356 32668
rect 24194 32614 24196 32666
rect 24258 32614 24270 32666
rect 24332 32614 24334 32666
rect 24172 32612 24196 32614
rect 24252 32612 24276 32614
rect 24332 32612 24356 32614
rect 24116 32592 24412 32612
rect 24124 32496 24176 32502
rect 24124 32438 24176 32444
rect 24136 32337 24164 32438
rect 24400 32428 24452 32434
rect 24400 32370 24452 32376
rect 24122 32328 24178 32337
rect 24032 32292 24084 32298
rect 24122 32263 24178 32272
rect 24032 32234 24084 32240
rect 24032 32020 24084 32026
rect 24032 31962 24084 31968
rect 23940 31748 23992 31754
rect 23940 31690 23992 31696
rect 23848 31680 23900 31686
rect 23848 31622 23900 31628
rect 24044 31498 24072 31962
rect 24412 31890 24440 32370
rect 24400 31884 24452 31890
rect 24400 31826 24452 31832
rect 24412 31793 24440 31826
rect 24398 31784 24454 31793
rect 24398 31719 24454 31728
rect 24116 31580 24412 31600
rect 24172 31578 24196 31580
rect 24252 31578 24276 31580
rect 24332 31578 24356 31580
rect 24194 31526 24196 31578
rect 24258 31526 24270 31578
rect 24332 31526 24334 31578
rect 24172 31524 24196 31526
rect 24252 31524 24276 31526
rect 24332 31524 24356 31526
rect 24116 31504 24412 31524
rect 23860 31470 24072 31498
rect 23860 26042 23888 31470
rect 24124 31408 24176 31414
rect 24124 31350 24176 31356
rect 24136 31278 24164 31350
rect 23940 31272 23992 31278
rect 23938 31240 23940 31249
rect 24124 31272 24176 31278
rect 23992 31240 23994 31249
rect 24124 31214 24176 31220
rect 23938 31175 23994 31184
rect 24032 31136 24084 31142
rect 24032 31078 24084 31084
rect 24044 30394 24072 31078
rect 24116 30492 24412 30512
rect 24172 30490 24196 30492
rect 24252 30490 24276 30492
rect 24332 30490 24356 30492
rect 24194 30438 24196 30490
rect 24258 30438 24270 30490
rect 24332 30438 24334 30490
rect 24172 30436 24196 30438
rect 24252 30436 24276 30438
rect 24332 30436 24356 30438
rect 24116 30416 24412 30436
rect 24032 30388 24084 30394
rect 24032 30330 24084 30336
rect 24116 29404 24412 29424
rect 24172 29402 24196 29404
rect 24252 29402 24276 29404
rect 24332 29402 24356 29404
rect 24194 29350 24196 29402
rect 24258 29350 24270 29402
rect 24332 29350 24334 29402
rect 24172 29348 24196 29350
rect 24252 29348 24276 29350
rect 24332 29348 24356 29350
rect 24116 29328 24412 29348
rect 24116 28316 24412 28336
rect 24172 28314 24196 28316
rect 24252 28314 24276 28316
rect 24332 28314 24356 28316
rect 24194 28262 24196 28314
rect 24258 28262 24270 28314
rect 24332 28262 24334 28314
rect 24172 28260 24196 28262
rect 24252 28260 24276 28262
rect 24332 28260 24356 28262
rect 24116 28240 24412 28260
rect 24032 28008 24084 28014
rect 24030 27976 24032 27985
rect 24124 28008 24176 28014
rect 24084 27976 24086 27985
rect 24124 27950 24176 27956
rect 24030 27911 24086 27920
rect 23940 27668 23992 27674
rect 23940 27610 23992 27616
rect 23952 27577 23980 27610
rect 24032 27600 24084 27606
rect 23938 27568 23994 27577
rect 24032 27542 24084 27548
rect 23938 27503 23994 27512
rect 24044 27452 24072 27542
rect 23952 27424 24072 27452
rect 23952 27130 23980 27424
rect 24136 27316 24164 27950
rect 24044 27288 24164 27316
rect 23940 27124 23992 27130
rect 23940 27066 23992 27072
rect 23848 26036 23900 26042
rect 23848 25978 23900 25984
rect 23848 25900 23900 25906
rect 23848 25842 23900 25848
rect 23860 22710 23888 25842
rect 23848 22704 23900 22710
rect 23848 22646 23900 22652
rect 23952 22574 23980 27066
rect 24044 26858 24072 27288
rect 24116 27228 24412 27248
rect 24172 27226 24196 27228
rect 24252 27226 24276 27228
rect 24332 27226 24356 27228
rect 24194 27174 24196 27226
rect 24258 27174 24270 27226
rect 24332 27174 24334 27226
rect 24172 27172 24196 27174
rect 24252 27172 24276 27174
rect 24332 27172 24356 27174
rect 24116 27152 24412 27172
rect 24032 26852 24084 26858
rect 24032 26794 24084 26800
rect 24116 26140 24412 26160
rect 24172 26138 24196 26140
rect 24252 26138 24276 26140
rect 24332 26138 24356 26140
rect 24194 26086 24196 26138
rect 24258 26086 24270 26138
rect 24332 26086 24334 26138
rect 24172 26084 24196 26086
rect 24252 26084 24276 26086
rect 24332 26084 24356 26086
rect 24116 26064 24412 26084
rect 24504 25838 24532 32728
rect 24032 25832 24084 25838
rect 24032 25774 24084 25780
rect 24492 25832 24544 25838
rect 24492 25774 24544 25780
rect 24044 22692 24072 25774
rect 24492 25356 24544 25362
rect 24492 25298 24544 25304
rect 24116 25052 24412 25072
rect 24172 25050 24196 25052
rect 24252 25050 24276 25052
rect 24332 25050 24356 25052
rect 24194 24998 24196 25050
rect 24258 24998 24270 25050
rect 24332 24998 24334 25050
rect 24172 24996 24196 24998
rect 24252 24996 24276 24998
rect 24332 24996 24356 24998
rect 24116 24976 24412 24996
rect 24504 24206 24532 25298
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 24116 23964 24412 23984
rect 24172 23962 24196 23964
rect 24252 23962 24276 23964
rect 24332 23962 24356 23964
rect 24194 23910 24196 23962
rect 24258 23910 24270 23962
rect 24332 23910 24334 23962
rect 24172 23908 24196 23910
rect 24252 23908 24276 23910
rect 24332 23908 24356 23910
rect 24116 23888 24412 23908
rect 24116 22876 24412 22896
rect 24172 22874 24196 22876
rect 24252 22874 24276 22876
rect 24332 22874 24356 22876
rect 24194 22822 24196 22874
rect 24258 22822 24270 22874
rect 24332 22822 24334 22874
rect 24172 22820 24196 22822
rect 24252 22820 24276 22822
rect 24332 22820 24356 22822
rect 24116 22800 24412 22820
rect 24492 22772 24544 22778
rect 24492 22714 24544 22720
rect 24044 22664 24164 22692
rect 23848 22568 23900 22574
rect 23848 22510 23900 22516
rect 23940 22568 23992 22574
rect 23940 22510 23992 22516
rect 23860 21078 23888 22510
rect 23940 22432 23992 22438
rect 23940 22374 23992 22380
rect 23848 21072 23900 21078
rect 23848 21014 23900 21020
rect 23860 19394 23888 21014
rect 23952 21010 23980 22374
rect 24032 22228 24084 22234
rect 24032 22170 24084 22176
rect 24044 21146 24072 22170
rect 24136 22001 24164 22664
rect 24216 22568 24268 22574
rect 24216 22510 24268 22516
rect 24228 22234 24256 22510
rect 24216 22228 24268 22234
rect 24216 22170 24268 22176
rect 24122 21992 24178 22001
rect 24122 21927 24178 21936
rect 24116 21788 24412 21808
rect 24172 21786 24196 21788
rect 24252 21786 24276 21788
rect 24332 21786 24356 21788
rect 24194 21734 24196 21786
rect 24258 21734 24270 21786
rect 24332 21734 24334 21786
rect 24172 21732 24196 21734
rect 24252 21732 24276 21734
rect 24332 21732 24356 21734
rect 24116 21712 24412 21732
rect 24122 21584 24178 21593
rect 24122 21519 24178 21528
rect 24032 21140 24084 21146
rect 24032 21082 24084 21088
rect 23940 21004 23992 21010
rect 23940 20946 23992 20952
rect 24136 20788 24164 21519
rect 24504 21146 24532 22714
rect 24492 21140 24544 21146
rect 24492 21082 24544 21088
rect 24044 20760 24164 20788
rect 24044 19496 24072 20760
rect 24116 20700 24412 20720
rect 24172 20698 24196 20700
rect 24252 20698 24276 20700
rect 24332 20698 24356 20700
rect 24194 20646 24196 20698
rect 24258 20646 24270 20698
rect 24332 20646 24334 20698
rect 24172 20644 24196 20646
rect 24252 20644 24276 20646
rect 24332 20644 24356 20646
rect 24116 20624 24412 20644
rect 24492 20596 24544 20602
rect 24492 20538 24544 20544
rect 24116 19612 24412 19632
rect 24172 19610 24196 19612
rect 24252 19610 24276 19612
rect 24332 19610 24356 19612
rect 24194 19558 24196 19610
rect 24258 19558 24270 19610
rect 24332 19558 24334 19610
rect 24172 19556 24196 19558
rect 24252 19556 24276 19558
rect 24332 19556 24356 19558
rect 24116 19536 24412 19556
rect 24044 19468 24256 19496
rect 23860 19366 24164 19394
rect 23940 19304 23992 19310
rect 23940 19246 23992 19252
rect 24032 19304 24084 19310
rect 24032 19246 24084 19252
rect 23848 19236 23900 19242
rect 23848 19178 23900 19184
rect 23860 18902 23888 19178
rect 23952 18902 23980 19246
rect 23848 18896 23900 18902
rect 23848 18838 23900 18844
rect 23940 18896 23992 18902
rect 23940 18838 23992 18844
rect 23952 18290 23980 18838
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 24044 18170 24072 19246
rect 24136 18834 24164 19366
rect 24228 19281 24256 19468
rect 24214 19272 24270 19281
rect 24214 19207 24270 19216
rect 24124 18828 24176 18834
rect 24124 18770 24176 18776
rect 24136 18698 24164 18770
rect 24228 18766 24256 19207
rect 24216 18760 24268 18766
rect 24216 18702 24268 18708
rect 24124 18692 24176 18698
rect 24124 18634 24176 18640
rect 24116 18524 24412 18544
rect 24172 18522 24196 18524
rect 24252 18522 24276 18524
rect 24332 18522 24356 18524
rect 24194 18470 24196 18522
rect 24258 18470 24270 18522
rect 24332 18470 24334 18522
rect 24172 18468 24196 18470
rect 24252 18468 24276 18470
rect 24332 18468 24356 18470
rect 24116 18448 24412 18468
rect 23952 18154 24072 18170
rect 23940 18148 24072 18154
rect 23992 18142 24072 18148
rect 23940 18090 23992 18096
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 23860 14006 23888 15438
rect 23848 14000 23900 14006
rect 23848 13942 23900 13948
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 23860 12238 23888 13330
rect 23952 13258 23980 18090
rect 24116 17436 24412 17456
rect 24172 17434 24196 17436
rect 24252 17434 24276 17436
rect 24332 17434 24356 17436
rect 24194 17382 24196 17434
rect 24258 17382 24270 17434
rect 24332 17382 24334 17434
rect 24172 17380 24196 17382
rect 24252 17380 24276 17382
rect 24332 17380 24356 17382
rect 24116 17360 24412 17380
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24032 16652 24084 16658
rect 24032 16594 24084 16600
rect 24044 15144 24072 16594
rect 24216 16584 24268 16590
rect 24214 16552 24216 16561
rect 24268 16552 24270 16561
rect 24412 16522 24440 16934
rect 24214 16487 24270 16496
rect 24400 16516 24452 16522
rect 24400 16458 24452 16464
rect 24116 16348 24412 16368
rect 24172 16346 24196 16348
rect 24252 16346 24276 16348
rect 24332 16346 24356 16348
rect 24194 16294 24196 16346
rect 24258 16294 24270 16346
rect 24332 16294 24334 16346
rect 24172 16292 24196 16294
rect 24252 16292 24276 16294
rect 24332 16292 24356 16294
rect 24116 16272 24412 16292
rect 24504 15434 24532 20538
rect 24492 15428 24544 15434
rect 24492 15370 24544 15376
rect 24116 15260 24412 15280
rect 24172 15258 24196 15260
rect 24252 15258 24276 15260
rect 24332 15258 24356 15260
rect 24194 15206 24196 15258
rect 24258 15206 24270 15258
rect 24332 15206 24334 15258
rect 24172 15204 24196 15206
rect 24252 15204 24276 15206
rect 24332 15204 24356 15206
rect 24116 15184 24412 15204
rect 24044 15116 24532 15144
rect 24116 14172 24412 14192
rect 24172 14170 24196 14172
rect 24252 14170 24276 14172
rect 24332 14170 24356 14172
rect 24194 14118 24196 14170
rect 24258 14118 24270 14170
rect 24332 14118 24334 14170
rect 24172 14116 24196 14118
rect 24252 14116 24276 14118
rect 24332 14116 24356 14118
rect 24116 14096 24412 14116
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 23940 13252 23992 13258
rect 23940 13194 23992 13200
rect 24044 12986 24072 13330
rect 24116 13084 24412 13104
rect 24172 13082 24196 13084
rect 24252 13082 24276 13084
rect 24332 13082 24356 13084
rect 24194 13030 24196 13082
rect 24258 13030 24270 13082
rect 24332 13030 24334 13082
rect 24172 13028 24196 13030
rect 24252 13028 24276 13030
rect 24332 13028 24356 13030
rect 24116 13008 24412 13028
rect 24032 12980 24084 12986
rect 24032 12922 24084 12928
rect 24044 12434 24072 12922
rect 23952 12406 24072 12434
rect 23952 12306 23980 12406
rect 23940 12300 23992 12306
rect 23940 12242 23992 12248
rect 23848 12232 23900 12238
rect 23848 12174 23900 12180
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 23860 10470 23888 11086
rect 23952 10674 23980 12242
rect 24116 11996 24412 12016
rect 24172 11994 24196 11996
rect 24252 11994 24276 11996
rect 24332 11994 24356 11996
rect 24194 11942 24196 11994
rect 24258 11942 24270 11994
rect 24332 11942 24334 11994
rect 24172 11940 24196 11942
rect 24252 11940 24276 11942
rect 24332 11940 24356 11942
rect 24116 11920 24412 11940
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 24044 10810 24072 11086
rect 24116 10908 24412 10928
rect 24172 10906 24196 10908
rect 24252 10906 24276 10908
rect 24332 10906 24356 10908
rect 24194 10854 24196 10906
rect 24258 10854 24270 10906
rect 24332 10854 24334 10906
rect 24172 10852 24196 10854
rect 24252 10852 24276 10854
rect 24332 10852 24356 10854
rect 24116 10832 24412 10852
rect 24504 10810 24532 15116
rect 24032 10804 24084 10810
rect 24032 10746 24084 10752
rect 24492 10804 24544 10810
rect 24492 10746 24544 10752
rect 24596 10690 24624 34598
rect 24872 34218 24900 34954
rect 24780 34190 24900 34218
rect 24676 33992 24728 33998
rect 24676 33934 24728 33940
rect 24688 33590 24716 33934
rect 24676 33584 24728 33590
rect 24676 33526 24728 33532
rect 24674 33416 24730 33425
rect 24674 33351 24730 33360
rect 24688 31906 24716 33351
rect 24780 33130 24808 34190
rect 24860 34060 24912 34066
rect 24860 34002 24912 34008
rect 24872 33289 24900 34002
rect 24858 33280 24914 33289
rect 24858 33215 24914 33224
rect 24780 33102 24900 33130
rect 24768 33040 24820 33046
rect 24768 32982 24820 32988
rect 24780 32842 24808 32982
rect 24872 32978 24900 33102
rect 24860 32972 24912 32978
rect 24860 32914 24912 32920
rect 24768 32836 24820 32842
rect 24768 32778 24820 32784
rect 24860 32836 24912 32842
rect 24860 32778 24912 32784
rect 24780 32026 24808 32778
rect 24872 32298 24900 32778
rect 24860 32292 24912 32298
rect 24860 32234 24912 32240
rect 24768 32020 24820 32026
rect 24768 31962 24820 31968
rect 24964 31929 24992 41006
rect 25056 38654 25084 46990
rect 25136 44736 25188 44742
rect 25136 44678 25188 44684
rect 25148 43790 25176 44678
rect 25136 43784 25188 43790
rect 25136 43726 25188 43732
rect 25136 43240 25188 43246
rect 25136 43182 25188 43188
rect 25148 42838 25176 43182
rect 25136 42832 25188 42838
rect 25136 42774 25188 42780
rect 25240 41698 25268 55655
rect 25502 55200 25558 56800
rect 27250 55200 27306 56800
rect 28998 55200 29054 56800
rect 25516 53582 25544 55200
rect 27068 53780 27120 53786
rect 27068 53722 27120 53728
rect 26700 53712 26752 53718
rect 25686 53680 25742 53689
rect 26700 53654 26752 53660
rect 25686 53615 25688 53624
rect 25740 53615 25742 53624
rect 25688 53586 25740 53592
rect 25504 53576 25556 53582
rect 25504 53518 25556 53524
rect 25780 53032 25832 53038
rect 25780 52974 25832 52980
rect 25504 52896 25556 52902
rect 25504 52838 25556 52844
rect 25516 52562 25544 52838
rect 25412 52556 25464 52562
rect 25412 52498 25464 52504
rect 25504 52556 25556 52562
rect 25504 52498 25556 52504
rect 25320 51060 25372 51066
rect 25320 51002 25372 51008
rect 25332 50674 25360 51002
rect 25424 50833 25452 52498
rect 25688 51264 25740 51270
rect 25792 51241 25820 52974
rect 26240 52964 26292 52970
rect 26240 52906 26292 52912
rect 26608 52964 26660 52970
rect 26608 52906 26660 52912
rect 26252 52562 26280 52906
rect 26424 52896 26476 52902
rect 26424 52838 26476 52844
rect 26240 52556 26292 52562
rect 26240 52498 26292 52504
rect 26332 52488 26384 52494
rect 26332 52430 26384 52436
rect 26056 52352 26108 52358
rect 26056 52294 26108 52300
rect 25872 51808 25924 51814
rect 25872 51750 25924 51756
rect 25884 51377 25912 51750
rect 26068 51610 26096 52294
rect 26056 51604 26108 51610
rect 26056 51546 26108 51552
rect 25870 51368 25926 51377
rect 25870 51303 25926 51312
rect 25688 51206 25740 51212
rect 25778 51232 25834 51241
rect 25700 50862 25728 51206
rect 25778 51167 25834 51176
rect 25688 50856 25740 50862
rect 25410 50824 25466 50833
rect 25688 50798 25740 50804
rect 26056 50856 26108 50862
rect 26056 50798 26108 50804
rect 25410 50759 25466 50768
rect 25332 50646 25452 50674
rect 25424 49774 25452 50646
rect 25596 50380 25648 50386
rect 25596 50322 25648 50328
rect 25412 49768 25464 49774
rect 25412 49710 25464 49716
rect 25320 48680 25372 48686
rect 25320 48622 25372 48628
rect 25332 48550 25360 48622
rect 25320 48544 25372 48550
rect 25320 48486 25372 48492
rect 25424 47598 25452 49710
rect 25608 49609 25636 50322
rect 25594 49600 25650 49609
rect 25594 49535 25650 49544
rect 25596 49224 25648 49230
rect 25596 49166 25648 49172
rect 25504 49088 25556 49094
rect 25504 49030 25556 49036
rect 25516 48686 25544 49030
rect 25504 48680 25556 48686
rect 25504 48622 25556 48628
rect 25608 48498 25636 49166
rect 25516 48470 25636 48498
rect 25412 47592 25464 47598
rect 25412 47534 25464 47540
rect 25320 44940 25372 44946
rect 25320 44882 25372 44888
rect 25332 44538 25360 44882
rect 25320 44532 25372 44538
rect 25320 44474 25372 44480
rect 25424 44470 25452 47534
rect 25412 44464 25464 44470
rect 25412 44406 25464 44412
rect 25412 44328 25464 44334
rect 25412 44270 25464 44276
rect 25320 43920 25372 43926
rect 25320 43862 25372 43868
rect 25332 43450 25360 43862
rect 25320 43444 25372 43450
rect 25320 43386 25372 43392
rect 25424 42294 25452 44270
rect 25516 43994 25544 48470
rect 25596 48204 25648 48210
rect 25596 48146 25648 48152
rect 25608 47569 25636 48146
rect 25700 47818 25728 50798
rect 25872 50720 25924 50726
rect 25872 50662 25924 50668
rect 25884 50454 25912 50662
rect 25872 50448 25924 50454
rect 25872 50390 25924 50396
rect 25872 50176 25924 50182
rect 25872 50118 25924 50124
rect 25884 49774 25912 50118
rect 26068 50017 26096 50798
rect 26344 50794 26372 52430
rect 26436 51882 26464 52838
rect 26516 52692 26568 52698
rect 26516 52634 26568 52640
rect 26528 51950 26556 52634
rect 26516 51944 26568 51950
rect 26516 51886 26568 51892
rect 26424 51876 26476 51882
rect 26424 51818 26476 51824
rect 26620 50930 26648 52906
rect 26712 51474 26740 53654
rect 27080 53038 27108 53722
rect 27264 53446 27292 55200
rect 27252 53440 27304 53446
rect 27252 53382 27304 53388
rect 27896 53236 27948 53242
rect 27896 53178 27948 53184
rect 27252 53100 27304 53106
rect 27252 53042 27304 53048
rect 27068 53032 27120 53038
rect 27068 52974 27120 52980
rect 27158 53000 27214 53009
rect 27158 52935 27214 52944
rect 27172 52902 27200 52935
rect 27160 52896 27212 52902
rect 27160 52838 27212 52844
rect 27264 51950 27292 53042
rect 27908 52630 27936 53178
rect 27988 53168 28040 53174
rect 27988 53110 28040 53116
rect 27528 52624 27580 52630
rect 27528 52566 27580 52572
rect 27896 52624 27948 52630
rect 27896 52566 27948 52572
rect 27540 51950 27568 52566
rect 27620 52488 27672 52494
rect 27620 52430 27672 52436
rect 27252 51944 27304 51950
rect 27252 51886 27304 51892
rect 27528 51944 27580 51950
rect 27528 51886 27580 51892
rect 27632 51513 27660 52430
rect 27618 51504 27674 51513
rect 26700 51468 26752 51474
rect 28000 51474 28028 53110
rect 29012 52086 29040 55200
rect 29000 52080 29052 52086
rect 29000 52022 29052 52028
rect 28078 51912 28134 51921
rect 28078 51847 28134 51856
rect 28092 51814 28120 51847
rect 28080 51808 28132 51814
rect 28080 51750 28132 51756
rect 27618 51439 27674 51448
rect 27988 51468 28040 51474
rect 26700 51410 26752 51416
rect 27988 51410 28040 51416
rect 26792 51264 26844 51270
rect 26792 51206 26844 51212
rect 26608 50924 26660 50930
rect 26608 50866 26660 50872
rect 26700 50856 26752 50862
rect 26700 50798 26752 50804
rect 26332 50788 26384 50794
rect 26332 50730 26384 50736
rect 26240 50380 26292 50386
rect 26240 50322 26292 50328
rect 26054 50008 26110 50017
rect 26054 49943 26110 49952
rect 25780 49768 25832 49774
rect 25780 49710 25832 49716
rect 25872 49768 25924 49774
rect 25872 49710 25924 49716
rect 25792 49434 25820 49710
rect 25872 49632 25924 49638
rect 25872 49574 25924 49580
rect 25780 49428 25832 49434
rect 25780 49370 25832 49376
rect 25780 49292 25832 49298
rect 25780 49234 25832 49240
rect 25792 48890 25820 49234
rect 25884 49230 25912 49574
rect 25872 49224 25924 49230
rect 25872 49166 25924 49172
rect 26148 49224 26200 49230
rect 26148 49166 26200 49172
rect 25780 48884 25832 48890
rect 25780 48826 25832 48832
rect 26160 48550 26188 49166
rect 26252 48793 26280 50322
rect 26424 49836 26476 49842
rect 26424 49778 26476 49784
rect 26238 48784 26294 48793
rect 26238 48719 26294 48728
rect 26148 48544 26200 48550
rect 26148 48486 26200 48492
rect 25964 48000 26016 48006
rect 25964 47942 26016 47948
rect 26056 48000 26108 48006
rect 26056 47942 26108 47948
rect 25700 47790 25820 47818
rect 25594 47560 25650 47569
rect 25594 47495 25650 47504
rect 25596 46028 25648 46034
rect 25596 45970 25648 45976
rect 25608 45529 25636 45970
rect 25688 45552 25740 45558
rect 25594 45520 25650 45529
rect 25688 45494 25740 45500
rect 25594 45455 25650 45464
rect 25596 45416 25648 45422
rect 25700 45404 25728 45494
rect 25648 45376 25728 45404
rect 25596 45358 25648 45364
rect 25596 44328 25648 44334
rect 25596 44270 25648 44276
rect 25504 43988 25556 43994
rect 25504 43930 25556 43936
rect 25504 42628 25556 42634
rect 25504 42570 25556 42576
rect 25412 42288 25464 42294
rect 25412 42230 25464 42236
rect 25412 42152 25464 42158
rect 25412 42094 25464 42100
rect 25516 42106 25544 42570
rect 25608 42226 25636 44270
rect 25688 43988 25740 43994
rect 25688 43930 25740 43936
rect 25596 42220 25648 42226
rect 25596 42162 25648 42168
rect 25240 41670 25360 41698
rect 25228 41608 25280 41614
rect 25228 41550 25280 41556
rect 25240 40050 25268 41550
rect 25332 41070 25360 41670
rect 25424 41206 25452 42094
rect 25516 42078 25636 42106
rect 25608 42022 25636 42078
rect 25596 42016 25648 42022
rect 25596 41958 25648 41964
rect 25502 41440 25558 41449
rect 25502 41375 25558 41384
rect 25412 41200 25464 41206
rect 25412 41142 25464 41148
rect 25516 41070 25544 41375
rect 25320 41064 25372 41070
rect 25320 41006 25372 41012
rect 25504 41064 25556 41070
rect 25504 41006 25556 41012
rect 25228 40044 25280 40050
rect 25228 39986 25280 39992
rect 25320 40044 25372 40050
rect 25320 39986 25372 39992
rect 25228 39840 25280 39846
rect 25228 39782 25280 39788
rect 25240 39574 25268 39782
rect 25228 39568 25280 39574
rect 25228 39510 25280 39516
rect 25056 38626 25176 38654
rect 25044 38412 25096 38418
rect 25044 38354 25096 38360
rect 25056 37398 25084 38354
rect 25044 37392 25096 37398
rect 25044 37334 25096 37340
rect 25148 36564 25176 38626
rect 25332 38214 25360 39986
rect 25412 39976 25464 39982
rect 25412 39918 25464 39924
rect 25424 39817 25452 39918
rect 25410 39808 25466 39817
rect 25410 39743 25466 39752
rect 25504 38752 25556 38758
rect 25504 38694 25556 38700
rect 25320 38208 25372 38214
rect 25320 38150 25372 38156
rect 25320 37732 25372 37738
rect 25320 37674 25372 37680
rect 25332 37330 25360 37674
rect 25412 37664 25464 37670
rect 25412 37606 25464 37612
rect 25424 37330 25452 37606
rect 25320 37324 25372 37330
rect 25320 37266 25372 37272
rect 25412 37324 25464 37330
rect 25412 37266 25464 37272
rect 25056 36536 25176 36564
rect 25228 36576 25280 36582
rect 24950 31920 25006 31929
rect 24688 31878 24900 31906
rect 24872 31754 24900 31878
rect 24950 31855 25006 31864
rect 24872 31726 24992 31754
rect 24768 31408 24820 31414
rect 24768 31350 24820 31356
rect 24674 27840 24730 27849
rect 24674 27775 24730 27784
rect 24688 27674 24716 27775
rect 24676 27668 24728 27674
rect 24676 27610 24728 27616
rect 24688 25974 24716 27610
rect 24676 25968 24728 25974
rect 24676 25910 24728 25916
rect 24780 25242 24808 31350
rect 24860 28960 24912 28966
rect 24860 28902 24912 28908
rect 24872 28558 24900 28902
rect 24860 28552 24912 28558
rect 24860 28494 24912 28500
rect 24860 28416 24912 28422
rect 24860 28358 24912 28364
rect 24872 28014 24900 28358
rect 24860 28008 24912 28014
rect 24860 27950 24912 27956
rect 24858 27432 24914 27441
rect 24858 27367 24860 27376
rect 24912 27367 24914 27376
rect 24860 27338 24912 27344
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 24688 25214 24808 25242
rect 24688 22658 24716 25214
rect 24768 25152 24820 25158
rect 24768 25094 24820 25100
rect 24780 24682 24808 25094
rect 24768 24676 24820 24682
rect 24768 24618 24820 24624
rect 24768 24132 24820 24138
rect 24768 24074 24820 24080
rect 24780 22778 24808 24074
rect 24768 22772 24820 22778
rect 24768 22714 24820 22720
rect 24688 22630 24808 22658
rect 24676 22500 24728 22506
rect 24676 22442 24728 22448
rect 24688 18426 24716 22442
rect 24780 21026 24808 22630
rect 24872 22098 24900 26930
rect 24964 26790 24992 31726
rect 24952 26784 25004 26790
rect 24952 26726 25004 26732
rect 24950 25936 25006 25945
rect 24950 25871 24952 25880
rect 25004 25871 25006 25880
rect 24952 25842 25004 25848
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 24964 22574 24992 25230
rect 24952 22568 25004 22574
rect 24952 22510 25004 22516
rect 24952 22432 25004 22438
rect 24952 22374 25004 22380
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 24872 21486 24900 22034
rect 24964 22030 24992 22374
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 24872 21146 24900 21422
rect 24860 21140 24912 21146
rect 24860 21082 24912 21088
rect 24780 20998 24900 21026
rect 24768 20868 24820 20874
rect 24768 20810 24820 20816
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24780 18306 24808 20810
rect 24688 18278 24808 18306
rect 24688 16726 24716 18278
rect 24872 18170 24900 20998
rect 24964 18873 24992 21966
rect 24950 18864 25006 18873
rect 24950 18799 25006 18808
rect 25056 18630 25084 36536
rect 25228 36518 25280 36524
rect 25240 36310 25268 36518
rect 25228 36304 25280 36310
rect 25228 36246 25280 36252
rect 25228 34604 25280 34610
rect 25228 34546 25280 34552
rect 25136 32836 25188 32842
rect 25136 32778 25188 32784
rect 25148 30580 25176 32778
rect 25240 32366 25268 34546
rect 25332 33425 25360 37266
rect 25516 36786 25544 38694
rect 25504 36780 25556 36786
rect 25504 36722 25556 36728
rect 25412 36712 25464 36718
rect 25412 36654 25464 36660
rect 25424 36553 25452 36654
rect 25504 36644 25556 36650
rect 25504 36586 25556 36592
rect 25410 36544 25466 36553
rect 25410 36479 25466 36488
rect 25516 36378 25544 36586
rect 25504 36372 25556 36378
rect 25504 36314 25556 36320
rect 25412 34536 25464 34542
rect 25412 34478 25464 34484
rect 25318 33416 25374 33425
rect 25318 33351 25374 33360
rect 25318 33144 25374 33153
rect 25318 33079 25374 33088
rect 25228 32360 25280 32366
rect 25228 32302 25280 32308
rect 25228 31884 25280 31890
rect 25228 31826 25280 31832
rect 25240 31657 25268 31826
rect 25226 31648 25282 31657
rect 25226 31583 25282 31592
rect 25228 31272 25280 31278
rect 25228 31214 25280 31220
rect 25240 30734 25268 31214
rect 25228 30728 25280 30734
rect 25228 30670 25280 30676
rect 25228 30592 25280 30598
rect 25148 30552 25228 30580
rect 25228 30534 25280 30540
rect 25240 30326 25268 30534
rect 25228 30320 25280 30326
rect 25228 30262 25280 30268
rect 25240 29073 25268 30262
rect 25226 29064 25282 29073
rect 25226 28999 25282 29008
rect 25136 28960 25188 28966
rect 25136 28902 25188 28908
rect 25148 28762 25176 28902
rect 25136 28756 25188 28762
rect 25136 28698 25188 28704
rect 25136 28620 25188 28626
rect 25136 28562 25188 28568
rect 25148 28218 25176 28562
rect 25228 28552 25280 28558
rect 25228 28494 25280 28500
rect 25136 28212 25188 28218
rect 25136 28154 25188 28160
rect 25240 28082 25268 28494
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 25240 27554 25268 28018
rect 25148 27526 25268 27554
rect 25148 25294 25176 27526
rect 25332 27418 25360 33079
rect 25424 33017 25452 34478
rect 25504 34060 25556 34066
rect 25504 34002 25556 34008
rect 25410 33008 25466 33017
rect 25410 32943 25466 32952
rect 25516 32065 25544 34002
rect 25502 32056 25558 32065
rect 25502 31991 25558 32000
rect 25410 31920 25466 31929
rect 25410 31855 25466 31864
rect 25424 30802 25452 31855
rect 25608 31754 25636 41958
rect 25516 31726 25636 31754
rect 25412 30796 25464 30802
rect 25412 30738 25464 30744
rect 25516 30682 25544 31726
rect 25240 27390 25360 27418
rect 25424 30654 25544 30682
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 25136 25152 25188 25158
rect 25136 25094 25188 25100
rect 25148 24954 25176 25094
rect 25136 24948 25188 24954
rect 25136 24890 25188 24896
rect 25136 23044 25188 23050
rect 25136 22986 25188 22992
rect 25148 22681 25176 22986
rect 25134 22672 25190 22681
rect 25134 22607 25190 22616
rect 25240 22556 25268 27390
rect 25320 27328 25372 27334
rect 25320 27270 25372 27276
rect 25332 26926 25360 27270
rect 25424 26994 25452 30654
rect 25700 30546 25728 43930
rect 25792 37346 25820 47790
rect 25976 47598 26004 47942
rect 25872 47592 25924 47598
rect 25872 47534 25924 47540
rect 25964 47592 26016 47598
rect 25964 47534 26016 47540
rect 25884 47258 25912 47534
rect 25964 47456 26016 47462
rect 25964 47398 26016 47404
rect 25872 47252 25924 47258
rect 25872 47194 25924 47200
rect 25976 47054 26004 47398
rect 25964 47048 26016 47054
rect 25964 46990 26016 46996
rect 25964 46504 26016 46510
rect 25964 46446 26016 46452
rect 25872 46368 25924 46374
rect 25872 46310 25924 46316
rect 25884 38758 25912 46310
rect 25976 45937 26004 46446
rect 26068 46442 26096 47942
rect 26160 47054 26188 48486
rect 26240 48204 26292 48210
rect 26240 48146 26292 48152
rect 26148 47048 26200 47054
rect 26148 46990 26200 46996
rect 26056 46436 26108 46442
rect 26056 46378 26108 46384
rect 25962 45928 26018 45937
rect 25962 45863 26018 45872
rect 26160 45234 26188 46990
rect 26252 46753 26280 48146
rect 26238 46744 26294 46753
rect 26238 46679 26294 46688
rect 26436 46510 26464 49778
rect 26712 49201 26740 50798
rect 26804 50697 26832 51206
rect 27344 51060 27396 51066
rect 27344 51002 27396 51008
rect 27356 50969 27384 51002
rect 27342 50960 27398 50969
rect 27342 50895 27398 50904
rect 27436 50788 27488 50794
rect 27436 50730 27488 50736
rect 27160 50720 27212 50726
rect 26790 50688 26846 50697
rect 27160 50662 27212 50668
rect 26790 50623 26846 50632
rect 26976 50380 27028 50386
rect 26976 50322 27028 50328
rect 26884 49292 26936 49298
rect 26884 49234 26936 49240
rect 26698 49192 26754 49201
rect 26698 49127 26754 49136
rect 26700 48680 26752 48686
rect 26700 48622 26752 48628
rect 26516 48544 26568 48550
rect 26516 48486 26568 48492
rect 26528 47190 26556 48486
rect 26516 47184 26568 47190
rect 26712 47161 26740 48622
rect 26896 47977 26924 49234
rect 26988 48385 27016 50322
rect 27172 48686 27200 50662
rect 27448 50522 27476 50730
rect 28080 50720 28132 50726
rect 28080 50662 28132 50668
rect 27436 50516 27488 50522
rect 27436 50458 27488 50464
rect 28092 50289 28120 50662
rect 28078 50280 28134 50289
rect 27896 50244 27948 50250
rect 28078 50215 28134 50224
rect 27896 50186 27948 50192
rect 27908 49366 27936 50186
rect 27988 50176 28040 50182
rect 27988 50118 28040 50124
rect 27896 49360 27948 49366
rect 27896 49302 27948 49308
rect 27896 49088 27948 49094
rect 27896 49030 27948 49036
rect 27160 48680 27212 48686
rect 27160 48622 27212 48628
rect 26974 48376 27030 48385
rect 26974 48311 27030 48320
rect 27908 48278 27936 49030
rect 28000 48686 28028 50118
rect 28080 49156 28132 49162
rect 28080 49098 28132 49104
rect 28092 48890 28120 49098
rect 28080 48884 28132 48890
rect 28080 48826 28132 48832
rect 27988 48680 28040 48686
rect 27988 48622 28040 48628
rect 27896 48272 27948 48278
rect 27896 48214 27948 48220
rect 26976 48204 27028 48210
rect 26976 48146 27028 48152
rect 26882 47968 26938 47977
rect 26882 47903 26938 47912
rect 26516 47126 26568 47132
rect 26698 47152 26754 47161
rect 26698 47087 26754 47096
rect 26424 46504 26476 46510
rect 26424 46446 26476 46452
rect 26988 46345 27016 48146
rect 27896 48000 27948 48006
rect 27896 47942 27948 47948
rect 27908 47190 27936 47942
rect 27896 47184 27948 47190
rect 27896 47126 27948 47132
rect 26974 46336 27030 46345
rect 26974 46271 27030 46280
rect 26240 46028 26292 46034
rect 26240 45970 26292 45976
rect 26976 46028 27028 46034
rect 26976 45970 27028 45976
rect 25976 45206 26188 45234
rect 25976 43858 26004 45206
rect 26252 45121 26280 45970
rect 26884 45280 26936 45286
rect 26884 45222 26936 45228
rect 26238 45112 26294 45121
rect 26238 45047 26294 45056
rect 26148 44940 26200 44946
rect 26148 44882 26200 44888
rect 26056 44736 26108 44742
rect 26056 44678 26108 44684
rect 26068 43926 26096 44678
rect 26160 44305 26188 44882
rect 26700 44736 26752 44742
rect 26700 44678 26752 44684
rect 26146 44296 26202 44305
rect 26146 44231 26202 44240
rect 26056 43920 26108 43926
rect 26056 43862 26108 43868
rect 25964 43852 26016 43858
rect 25964 43794 26016 43800
rect 26148 43852 26200 43858
rect 26148 43794 26200 43800
rect 26240 43852 26292 43858
rect 26240 43794 26292 43800
rect 25976 41546 26004 43794
rect 26056 43240 26108 43246
rect 26056 43182 26108 43188
rect 26068 42265 26096 43182
rect 26160 42673 26188 43794
rect 26252 43178 26280 43794
rect 26240 43172 26292 43178
rect 26240 43114 26292 43120
rect 26712 42770 26740 44678
rect 26896 44334 26924 45222
rect 26988 44713 27016 45970
rect 27620 45892 27672 45898
rect 27620 45834 27672 45840
rect 27632 45422 27660 45834
rect 27896 45824 27948 45830
rect 27896 45766 27948 45772
rect 27068 45416 27120 45422
rect 27068 45358 27120 45364
rect 27620 45416 27672 45422
rect 27620 45358 27672 45364
rect 26974 44704 27030 44713
rect 26974 44639 27030 44648
rect 26884 44328 26936 44334
rect 26884 44270 26936 44276
rect 27080 43897 27108 45358
rect 27908 45014 27936 45766
rect 27896 45008 27948 45014
rect 27896 44950 27948 44956
rect 27160 44940 27212 44946
rect 27160 44882 27212 44888
rect 27066 43888 27122 43897
rect 27066 43823 27122 43832
rect 26792 43240 26844 43246
rect 26792 43182 26844 43188
rect 26700 42764 26752 42770
rect 26700 42706 26752 42712
rect 26146 42664 26202 42673
rect 26146 42599 26202 42608
rect 26148 42560 26200 42566
rect 26148 42502 26200 42508
rect 26608 42560 26660 42566
rect 26608 42502 26660 42508
rect 26054 42256 26110 42265
rect 26054 42191 26110 42200
rect 26160 41614 26188 42502
rect 26620 42158 26648 42502
rect 26608 42152 26660 42158
rect 26608 42094 26660 42100
rect 26332 42084 26384 42090
rect 26332 42026 26384 42032
rect 26344 41818 26372 42026
rect 26804 41857 26832 43182
rect 27172 43081 27200 44882
rect 28080 44192 28132 44198
rect 28080 44134 28132 44140
rect 28092 43790 28120 44134
rect 28080 43784 28132 43790
rect 28080 43726 28132 43732
rect 27252 43716 27304 43722
rect 27252 43658 27304 43664
rect 27264 43178 27292 43658
rect 28080 43648 28132 43654
rect 28080 43590 28132 43596
rect 27988 43376 28040 43382
rect 27988 43318 28040 43324
rect 27252 43172 27304 43178
rect 27252 43114 27304 43120
rect 27158 43072 27214 43081
rect 27158 43007 27214 43016
rect 28000 42770 28028 43318
rect 28092 42906 28120 43590
rect 28080 42900 28132 42906
rect 28080 42842 28132 42848
rect 27988 42764 28040 42770
rect 27988 42706 28040 42712
rect 28080 42560 28132 42566
rect 28080 42502 28132 42508
rect 28092 42362 28120 42502
rect 28080 42356 28132 42362
rect 28080 42298 28132 42304
rect 27436 42152 27488 42158
rect 27436 42094 27488 42100
rect 26790 41848 26846 41857
rect 26332 41812 26384 41818
rect 26790 41783 26846 41792
rect 26332 41754 26384 41760
rect 27068 41676 27120 41682
rect 27068 41618 27120 41624
rect 26148 41608 26200 41614
rect 26148 41550 26200 41556
rect 25964 41540 26016 41546
rect 25964 41482 26016 41488
rect 25976 40882 26004 41482
rect 27080 41274 27108 41618
rect 27068 41268 27120 41274
rect 27068 41210 27120 41216
rect 26148 41064 26200 41070
rect 26146 41032 26148 41041
rect 26792 41064 26844 41070
rect 26200 41032 26202 41041
rect 26792 41006 26844 41012
rect 26146 40967 26202 40976
rect 26608 40928 26660 40934
rect 25976 40854 26188 40882
rect 26608 40870 26660 40876
rect 26160 40526 26188 40854
rect 26620 40662 26648 40870
rect 26608 40656 26660 40662
rect 26804 40633 26832 41006
rect 27252 40928 27304 40934
rect 27252 40870 27304 40876
rect 26608 40598 26660 40604
rect 26790 40624 26846 40633
rect 26790 40559 26846 40568
rect 26148 40520 26200 40526
rect 26148 40462 26200 40468
rect 25964 40384 26016 40390
rect 25964 40326 26016 40332
rect 25976 39982 26004 40326
rect 25964 39976 26016 39982
rect 25964 39918 26016 39924
rect 26884 39500 26936 39506
rect 26884 39442 26936 39448
rect 26054 38992 26110 39001
rect 26054 38927 26110 38936
rect 26068 38894 26096 38927
rect 26056 38888 26108 38894
rect 26056 38830 26108 38836
rect 26792 38888 26844 38894
rect 26792 38830 26844 38836
rect 25872 38752 25924 38758
rect 25872 38694 25924 38700
rect 26148 38412 26200 38418
rect 26148 38354 26200 38360
rect 25872 38208 25924 38214
rect 25872 38150 25924 38156
rect 26056 38208 26108 38214
rect 26056 38150 26108 38156
rect 25884 37874 25912 38150
rect 25872 37868 25924 37874
rect 25872 37810 25924 37816
rect 25964 37868 26016 37874
rect 25964 37810 26016 37816
rect 25976 37482 26004 37810
rect 26068 37806 26096 38150
rect 26056 37800 26108 37806
rect 26160 37777 26188 38354
rect 26700 38208 26752 38214
rect 26804 38185 26832 38830
rect 26896 38593 26924 39442
rect 27264 38894 27292 40870
rect 27448 40225 27476 42094
rect 27896 42016 27948 42022
rect 27896 41958 27948 41964
rect 27528 41064 27580 41070
rect 27528 41006 27580 41012
rect 27434 40216 27490 40225
rect 27434 40151 27490 40160
rect 27344 39840 27396 39846
rect 27344 39782 27396 39788
rect 27356 39642 27384 39782
rect 27344 39636 27396 39642
rect 27344 39578 27396 39584
rect 27540 39409 27568 41006
rect 27908 39982 27936 41958
rect 27988 40384 28040 40390
rect 27988 40326 28040 40332
rect 28000 40186 28028 40326
rect 27988 40180 28040 40186
rect 27988 40122 28040 40128
rect 27896 39976 27948 39982
rect 27896 39918 27948 39924
rect 27526 39400 27582 39409
rect 27526 39335 27582 39344
rect 28172 39364 28224 39370
rect 28172 39306 28224 39312
rect 27896 39296 27948 39302
rect 27896 39238 27948 39244
rect 28080 39296 28132 39302
rect 28080 39238 28132 39244
rect 27804 39024 27856 39030
rect 27804 38966 27856 38972
rect 27252 38888 27304 38894
rect 27252 38830 27304 38836
rect 26882 38584 26938 38593
rect 26882 38519 26938 38528
rect 27252 38480 27304 38486
rect 27252 38422 27304 38428
rect 26884 38412 26936 38418
rect 26884 38354 26936 38360
rect 26700 38150 26752 38156
rect 26790 38176 26846 38185
rect 26056 37742 26108 37748
rect 26146 37768 26202 37777
rect 26146 37703 26202 37712
rect 25976 37454 26096 37482
rect 25792 37318 26004 37346
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 25792 36922 25820 37198
rect 25870 36952 25926 36961
rect 25780 36916 25832 36922
rect 25870 36887 25926 36896
rect 25780 36858 25832 36864
rect 25780 36712 25832 36718
rect 25780 36654 25832 36660
rect 25792 36582 25820 36654
rect 25780 36576 25832 36582
rect 25780 36518 25832 36524
rect 25792 35290 25820 36518
rect 25884 36242 25912 36887
rect 25872 36236 25924 36242
rect 25872 36178 25924 36184
rect 25976 36122 26004 37318
rect 26068 36582 26096 37454
rect 26712 37398 26740 38150
rect 26790 38111 26846 38120
rect 26700 37392 26752 37398
rect 26896 37369 26924 38354
rect 27264 38010 27292 38422
rect 27252 38004 27304 38010
rect 27252 37946 27304 37952
rect 27816 37806 27844 38966
rect 27908 38486 27936 39238
rect 28092 39098 28120 39238
rect 28080 39092 28132 39098
rect 28080 39034 28132 39040
rect 28184 39030 28212 39306
rect 28172 39024 28224 39030
rect 28172 38966 28224 38972
rect 28080 38548 28132 38554
rect 28080 38490 28132 38496
rect 27896 38480 27948 38486
rect 27896 38422 27948 38428
rect 27988 38208 28040 38214
rect 27988 38150 28040 38156
rect 28000 37942 28028 38150
rect 27988 37936 28040 37942
rect 27988 37878 28040 37884
rect 27804 37800 27856 37806
rect 27804 37742 27856 37748
rect 27344 37664 27396 37670
rect 27344 37606 27396 37612
rect 27356 37466 27384 37606
rect 28092 37466 28120 38490
rect 27344 37460 27396 37466
rect 27344 37402 27396 37408
rect 28080 37460 28132 37466
rect 28080 37402 28132 37408
rect 26700 37334 26752 37340
rect 26882 37360 26938 37369
rect 26882 37295 26938 37304
rect 26976 37324 27028 37330
rect 26976 37266 27028 37272
rect 26608 37256 26660 37262
rect 26608 37198 26660 37204
rect 26056 36576 26108 36582
rect 26056 36518 26108 36524
rect 26148 36236 26200 36242
rect 26148 36178 26200 36184
rect 26160 36145 26188 36178
rect 25884 36094 26004 36122
rect 26146 36136 26202 36145
rect 25780 35284 25832 35290
rect 25780 35226 25832 35232
rect 25780 34196 25832 34202
rect 25780 34138 25832 34144
rect 25792 33590 25820 34138
rect 25780 33584 25832 33590
rect 25780 33526 25832 33532
rect 25884 33130 25912 36094
rect 26146 36071 26202 36080
rect 26056 36032 26108 36038
rect 26056 35974 26108 35980
rect 26068 35630 26096 35974
rect 26056 35624 26108 35630
rect 26056 35566 26108 35572
rect 26620 35494 26648 37198
rect 26792 36712 26844 36718
rect 26792 36654 26844 36660
rect 26804 35737 26832 36654
rect 26884 36236 26936 36242
rect 26884 36178 26936 36184
rect 26790 35728 26846 35737
rect 26790 35663 26846 35672
rect 26608 35488 26660 35494
rect 26608 35430 26660 35436
rect 25964 34740 26016 34746
rect 25964 34682 26016 34688
rect 25976 33538 26004 34682
rect 26620 34610 26648 35430
rect 26896 35329 26924 36178
rect 26882 35320 26938 35329
rect 26882 35255 26938 35264
rect 26608 34604 26660 34610
rect 26608 34546 26660 34552
rect 26056 34536 26108 34542
rect 26054 34504 26056 34513
rect 26700 34536 26752 34542
rect 26108 34504 26110 34513
rect 26700 34478 26752 34484
rect 26054 34439 26110 34448
rect 26516 34400 26568 34406
rect 26516 34342 26568 34348
rect 26528 34134 26556 34342
rect 26516 34128 26568 34134
rect 26146 34096 26202 34105
rect 26516 34070 26568 34076
rect 26146 34031 26148 34040
rect 26200 34031 26202 34040
rect 26148 34002 26200 34008
rect 26516 33856 26568 33862
rect 26516 33798 26568 33804
rect 25976 33510 26280 33538
rect 26252 33454 26280 33510
rect 26332 33516 26384 33522
rect 26332 33458 26384 33464
rect 26056 33448 26108 33454
rect 26056 33390 26108 33396
rect 26240 33448 26292 33454
rect 26240 33390 26292 33396
rect 25884 33102 26004 33130
rect 25780 32768 25832 32774
rect 25778 32736 25780 32745
rect 25832 32736 25834 32745
rect 25778 32671 25834 32680
rect 25780 32360 25832 32366
rect 25780 32302 25832 32308
rect 25792 32201 25820 32302
rect 25872 32292 25924 32298
rect 25872 32234 25924 32240
rect 25778 32192 25834 32201
rect 25778 32127 25834 32136
rect 25792 31278 25820 32127
rect 25780 31272 25832 31278
rect 25884 31249 25912 32234
rect 25780 31214 25832 31220
rect 25870 31240 25926 31249
rect 25870 31175 25926 31184
rect 25884 31142 25912 31175
rect 25872 31136 25924 31142
rect 25872 31078 25924 31084
rect 25780 30796 25832 30802
rect 25780 30738 25832 30744
rect 25516 30518 25728 30546
rect 25412 26988 25464 26994
rect 25412 26930 25464 26936
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 25320 26784 25372 26790
rect 25320 26726 25372 26732
rect 25148 22528 25268 22556
rect 25044 18624 25096 18630
rect 25044 18566 25096 18572
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 24780 18142 24900 18170
rect 24780 16998 24808 18142
rect 25056 17814 25084 18294
rect 25044 17808 25096 17814
rect 25044 17750 25096 17756
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24676 16720 24728 16726
rect 24676 16662 24728 16668
rect 24768 16720 24820 16726
rect 24768 16662 24820 16668
rect 24780 15638 24808 16662
rect 24950 16552 25006 16561
rect 24950 16487 25006 16496
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24768 15632 24820 15638
rect 24768 15574 24820 15580
rect 24872 14890 24900 16390
rect 24964 16046 24992 16487
rect 24952 16040 25004 16046
rect 24952 15982 25004 15988
rect 24860 14884 24912 14890
rect 24860 14826 24912 14832
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24872 13326 24900 13806
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 24860 13184 24912 13190
rect 24860 13126 24912 13132
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24780 11150 24808 12174
rect 24872 11354 24900 13126
rect 25056 12170 25084 13330
rect 25044 12164 25096 12170
rect 25044 12106 25096 12112
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 24044 10662 24624 10690
rect 23940 10532 23992 10538
rect 23940 10474 23992 10480
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23860 10130 23888 10406
rect 23952 10198 23980 10474
rect 23940 10192 23992 10198
rect 23940 10134 23992 10140
rect 23848 10124 23900 10130
rect 23848 10066 23900 10072
rect 23860 8906 23888 10066
rect 23848 8900 23900 8906
rect 23848 8842 23900 8848
rect 23848 7880 23900 7886
rect 23952 7868 23980 10134
rect 23900 7840 23980 7868
rect 23848 7822 23900 7828
rect 23756 5160 23808 5166
rect 23756 5102 23808 5108
rect 23572 4752 23624 4758
rect 23572 4694 23624 4700
rect 23664 4752 23716 4758
rect 23664 4694 23716 4700
rect 23388 4072 23440 4078
rect 23388 4014 23440 4020
rect 23480 4072 23532 4078
rect 23480 4014 23532 4020
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 23204 3732 23256 3738
rect 23204 3674 23256 3680
rect 22376 3120 22428 3126
rect 22376 3062 22428 3068
rect 22928 3120 22980 3126
rect 22928 3062 22980 3068
rect 23020 3120 23072 3126
rect 23020 3062 23072 3068
rect 23112 2984 23164 2990
rect 21914 2952 21970 2961
rect 23216 2972 23244 3674
rect 23164 2944 23244 2972
rect 23112 2926 23164 2932
rect 21914 2887 21916 2896
rect 21968 2887 21970 2896
rect 22008 2916 22060 2922
rect 21916 2858 21968 2864
rect 22008 2858 22060 2864
rect 23020 2916 23072 2922
rect 23020 2858 23072 2864
rect 22020 2825 22048 2858
rect 21362 2751 21418 2760
rect 21652 2746 21772 2774
rect 22006 2816 22062 2825
rect 22006 2751 22062 2760
rect 20350 2544 20406 2553
rect 20350 2479 20406 2488
rect 20444 2508 20496 2514
rect 20444 2450 20496 2456
rect 19720 1414 19840 1442
rect 19720 800 19748 1414
rect 20456 1290 20484 2450
rect 20444 1284 20496 1290
rect 20444 1226 20496 1232
rect 21100 800 21128 2746
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 21376 2446 21404 2586
rect 21652 2582 21680 2746
rect 21640 2576 21692 2582
rect 21640 2518 21692 2524
rect 23032 2514 23060 2858
rect 23400 2514 23428 4014
rect 23584 4010 23612 4694
rect 23768 4282 23796 5102
rect 23860 4554 23888 7822
rect 23940 7200 23992 7206
rect 23940 7142 23992 7148
rect 23952 6866 23980 7142
rect 23940 6860 23992 6866
rect 23940 6802 23992 6808
rect 23952 6458 23980 6802
rect 23940 6452 23992 6458
rect 23940 6394 23992 6400
rect 23940 5568 23992 5574
rect 23940 5510 23992 5516
rect 23952 4826 23980 5510
rect 23940 4820 23992 4826
rect 23940 4762 23992 4768
rect 23940 4616 23992 4622
rect 23940 4558 23992 4564
rect 23848 4548 23900 4554
rect 23848 4490 23900 4496
rect 23756 4276 23808 4282
rect 23756 4218 23808 4224
rect 23664 4208 23716 4214
rect 23664 4150 23716 4156
rect 23572 4004 23624 4010
rect 23572 3946 23624 3952
rect 23676 2990 23704 4150
rect 23664 2984 23716 2990
rect 23664 2926 23716 2932
rect 23952 2922 23980 4558
rect 24044 2961 24072 10662
rect 24688 10198 24716 10950
rect 24676 10192 24728 10198
rect 24676 10134 24728 10140
rect 24780 10062 24808 11086
rect 24768 10056 24820 10062
rect 24768 9998 24820 10004
rect 24116 9820 24412 9840
rect 24172 9818 24196 9820
rect 24252 9818 24276 9820
rect 24332 9818 24356 9820
rect 24194 9766 24196 9818
rect 24258 9766 24270 9818
rect 24332 9766 24334 9818
rect 24172 9764 24196 9766
rect 24252 9764 24276 9766
rect 24332 9764 24356 9766
rect 24116 9744 24412 9764
rect 24858 9616 24914 9625
rect 24858 9551 24914 9560
rect 24872 8974 24900 9551
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 24952 8900 25004 8906
rect 24952 8842 25004 8848
rect 24860 8832 24912 8838
rect 24964 8809 24992 8842
rect 24860 8774 24912 8780
rect 24950 8800 25006 8809
rect 24116 8732 24412 8752
rect 24172 8730 24196 8732
rect 24252 8730 24276 8732
rect 24332 8730 24356 8732
rect 24194 8678 24196 8730
rect 24258 8678 24270 8730
rect 24332 8678 24334 8730
rect 24172 8676 24196 8678
rect 24252 8676 24276 8678
rect 24332 8676 24356 8678
rect 24116 8656 24412 8676
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 24116 7644 24412 7664
rect 24172 7642 24196 7644
rect 24252 7642 24276 7644
rect 24332 7642 24356 7644
rect 24194 7590 24196 7642
rect 24258 7590 24270 7642
rect 24332 7590 24334 7642
rect 24172 7588 24196 7590
rect 24252 7588 24276 7590
rect 24332 7588 24356 7590
rect 24116 7568 24412 7588
rect 24492 7336 24544 7342
rect 24492 7278 24544 7284
rect 24116 6556 24412 6576
rect 24172 6554 24196 6556
rect 24252 6554 24276 6556
rect 24332 6554 24356 6556
rect 24194 6502 24196 6554
rect 24258 6502 24270 6554
rect 24332 6502 24334 6554
rect 24172 6500 24196 6502
rect 24252 6500 24276 6502
rect 24332 6500 24356 6502
rect 24116 6480 24412 6500
rect 24504 5914 24532 7278
rect 24584 6860 24636 6866
rect 24584 6802 24636 6808
rect 24676 6860 24728 6866
rect 24676 6802 24728 6808
rect 24596 6458 24624 6802
rect 24584 6452 24636 6458
rect 24584 6394 24636 6400
rect 24688 6322 24716 6802
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 24780 6254 24808 8366
rect 24872 6934 24900 8774
rect 24950 8735 25006 8744
rect 24860 6928 24912 6934
rect 24860 6870 24912 6876
rect 25056 6730 25084 11834
rect 25148 11778 25176 22528
rect 25332 22094 25360 26726
rect 25412 26308 25464 26314
rect 25412 26250 25464 26256
rect 25424 25537 25452 26250
rect 25410 25528 25466 25537
rect 25410 25463 25466 25472
rect 25516 25412 25544 30518
rect 25686 30424 25742 30433
rect 25686 30359 25742 30368
rect 25700 30190 25728 30359
rect 25688 30184 25740 30190
rect 25688 30126 25740 30132
rect 25596 30048 25648 30054
rect 25596 29990 25648 29996
rect 25608 29306 25636 29990
rect 25596 29300 25648 29306
rect 25596 29242 25648 29248
rect 25686 29200 25742 29209
rect 25686 29135 25688 29144
rect 25740 29135 25742 29144
rect 25688 29106 25740 29112
rect 25686 29064 25742 29073
rect 25596 29028 25648 29034
rect 25686 28999 25742 29008
rect 25596 28970 25648 28976
rect 25608 27878 25636 28970
rect 25700 28014 25728 28999
rect 25688 28008 25740 28014
rect 25688 27950 25740 27956
rect 25596 27872 25648 27878
rect 25596 27814 25648 27820
rect 25700 27690 25728 27950
rect 25240 22066 25360 22094
rect 25424 25384 25544 25412
rect 25608 27662 25728 27690
rect 25240 19922 25268 22066
rect 25424 21162 25452 25384
rect 25504 25288 25556 25294
rect 25608 25242 25636 27662
rect 25792 27554 25820 30738
rect 25700 27526 25820 27554
rect 25884 27928 25912 31078
rect 25976 28098 26004 33102
rect 26068 32570 26096 33390
rect 26240 33312 26292 33318
rect 26240 33254 26292 33260
rect 26252 32910 26280 33254
rect 26344 33153 26372 33458
rect 26424 33380 26476 33386
rect 26424 33322 26476 33328
rect 26330 33144 26386 33153
rect 26330 33079 26386 33088
rect 26240 32904 26292 32910
rect 26240 32846 26292 32852
rect 26332 32904 26384 32910
rect 26436 32892 26464 33322
rect 26384 32864 26464 32892
rect 26332 32846 26384 32852
rect 26056 32564 26108 32570
rect 26056 32506 26108 32512
rect 26252 32230 26280 32846
rect 26344 32502 26372 32846
rect 26332 32496 26384 32502
rect 26332 32438 26384 32444
rect 26240 32224 26292 32230
rect 26240 32166 26292 32172
rect 26528 31890 26556 33798
rect 26712 33697 26740 34478
rect 26792 33856 26844 33862
rect 26792 33798 26844 33804
rect 26698 33688 26754 33697
rect 26804 33658 26832 33798
rect 26698 33623 26754 33632
rect 26792 33652 26844 33658
rect 26792 33594 26844 33600
rect 26608 32020 26660 32026
rect 26608 31962 26660 31968
rect 26148 31884 26200 31890
rect 26148 31826 26200 31832
rect 26516 31884 26568 31890
rect 26516 31826 26568 31832
rect 26054 31240 26110 31249
rect 26054 31175 26110 31184
rect 26068 29714 26096 31175
rect 26160 30841 26188 31826
rect 26332 31204 26384 31210
rect 26332 31146 26384 31152
rect 26146 30832 26202 30841
rect 26146 30767 26202 30776
rect 26148 30184 26200 30190
rect 26148 30126 26200 30132
rect 26160 30025 26188 30126
rect 26146 30016 26202 30025
rect 26146 29951 26202 29960
rect 26344 29850 26372 31146
rect 26620 30870 26648 31962
rect 26608 30864 26660 30870
rect 26608 30806 26660 30812
rect 26332 29844 26384 29850
rect 26332 29786 26384 29792
rect 26056 29708 26108 29714
rect 26056 29650 26108 29656
rect 26700 29708 26752 29714
rect 26700 29650 26752 29656
rect 26240 29572 26292 29578
rect 26240 29514 26292 29520
rect 26148 28620 26200 28626
rect 26148 28562 26200 28568
rect 26056 28416 26108 28422
rect 26056 28358 26108 28364
rect 26068 28098 26096 28358
rect 25976 28070 26096 28098
rect 25964 27940 26016 27946
rect 25884 27900 25964 27928
rect 25700 26314 25728 27526
rect 25780 27396 25832 27402
rect 25780 27338 25832 27344
rect 25792 27130 25820 27338
rect 25780 27124 25832 27130
rect 25780 27066 25832 27072
rect 25688 26308 25740 26314
rect 25688 26250 25740 26256
rect 25688 26036 25740 26042
rect 25688 25978 25740 25984
rect 25700 25362 25728 25978
rect 25884 25430 25912 27900
rect 25964 27882 26016 27888
rect 26068 27878 26096 28070
rect 26056 27872 26108 27878
rect 26056 27814 26108 27820
rect 25964 27668 26016 27674
rect 25964 27610 26016 27616
rect 25976 25786 26004 27610
rect 26068 26450 26096 27814
rect 26160 27674 26188 28562
rect 26252 27878 26280 29514
rect 26516 29232 26568 29238
rect 26516 29174 26568 29180
rect 26528 29102 26556 29174
rect 26516 29096 26568 29102
rect 26516 29038 26568 29044
rect 26424 29028 26476 29034
rect 26424 28970 26476 28976
rect 26436 28393 26464 28970
rect 26712 28966 26740 29650
rect 26884 29572 26936 29578
rect 26884 29514 26936 29520
rect 26700 28960 26752 28966
rect 26700 28902 26752 28908
rect 26712 28762 26740 28902
rect 26896 28801 26924 29514
rect 26882 28792 26938 28801
rect 26700 28756 26752 28762
rect 26882 28727 26938 28736
rect 26700 28698 26752 28704
rect 26422 28384 26478 28393
rect 26422 28319 26478 28328
rect 26712 28014 26740 28698
rect 26700 28008 26752 28014
rect 26422 27976 26478 27985
rect 26700 27950 26752 27956
rect 26422 27911 26478 27920
rect 26240 27872 26292 27878
rect 26240 27814 26292 27820
rect 26330 27840 26386 27849
rect 26330 27775 26386 27784
rect 26148 27668 26200 27674
rect 26148 27610 26200 27616
rect 26344 27606 26372 27775
rect 26332 27600 26384 27606
rect 26146 27568 26202 27577
rect 26332 27542 26384 27548
rect 26146 27503 26202 27512
rect 26240 27532 26292 27538
rect 26160 26518 26188 27503
rect 26240 27474 26292 27480
rect 26252 27441 26280 27474
rect 26238 27432 26294 27441
rect 26436 27402 26464 27911
rect 26698 27704 26754 27713
rect 26698 27639 26754 27648
rect 26712 27606 26740 27639
rect 26700 27600 26752 27606
rect 26700 27542 26752 27548
rect 26238 27367 26294 27376
rect 26424 27396 26476 27402
rect 26424 27338 26476 27344
rect 26240 27328 26292 27334
rect 26240 27270 26292 27276
rect 26792 27328 26844 27334
rect 26792 27270 26844 27276
rect 26252 27033 26280 27270
rect 26804 27169 26832 27270
rect 26790 27160 26846 27169
rect 26790 27095 26846 27104
rect 26332 27056 26384 27062
rect 26238 27024 26294 27033
rect 26332 26998 26384 27004
rect 26238 26959 26294 26968
rect 26148 26512 26200 26518
rect 26148 26454 26200 26460
rect 26056 26444 26108 26450
rect 26056 26386 26108 26392
rect 26240 26376 26292 26382
rect 26240 26318 26292 26324
rect 26148 26308 26200 26314
rect 26148 26250 26200 26256
rect 25976 25770 26096 25786
rect 25976 25764 26108 25770
rect 25976 25758 26056 25764
rect 25872 25424 25924 25430
rect 25792 25372 25872 25378
rect 25792 25366 25924 25372
rect 25688 25356 25740 25362
rect 25688 25298 25740 25304
rect 25792 25350 25912 25366
rect 25556 25236 25636 25242
rect 25504 25230 25636 25236
rect 25516 25214 25636 25230
rect 25516 22574 25544 25214
rect 25596 23180 25648 23186
rect 25596 23122 25648 23128
rect 25504 22568 25556 22574
rect 25504 22510 25556 22516
rect 25504 22432 25556 22438
rect 25504 22374 25556 22380
rect 25516 21486 25544 22374
rect 25608 22234 25636 23122
rect 25596 22228 25648 22234
rect 25596 22170 25648 22176
rect 25688 22092 25740 22098
rect 25608 22052 25688 22080
rect 25504 21480 25556 21486
rect 25504 21422 25556 21428
rect 25424 21134 25544 21162
rect 25412 21004 25464 21010
rect 25412 20946 25464 20952
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 25240 18034 25268 19858
rect 25424 19718 25452 20946
rect 25412 19712 25464 19718
rect 25412 19654 25464 19660
rect 25412 19440 25464 19446
rect 25412 19382 25464 19388
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25332 18222 25360 19110
rect 25424 18902 25452 19382
rect 25412 18896 25464 18902
rect 25412 18838 25464 18844
rect 25412 18624 25464 18630
rect 25412 18566 25464 18572
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 25240 18006 25360 18034
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25240 16250 25268 16594
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 25226 16144 25282 16153
rect 25226 16079 25282 16088
rect 25240 15638 25268 16079
rect 25228 15632 25280 15638
rect 25226 15600 25228 15609
rect 25280 15600 25282 15609
rect 25226 15535 25282 15544
rect 25228 13796 25280 13802
rect 25228 13738 25280 13744
rect 25240 12714 25268 13738
rect 25228 12708 25280 12714
rect 25228 12650 25280 12656
rect 25228 12164 25280 12170
rect 25228 12106 25280 12112
rect 25240 11898 25268 12106
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 25148 11750 25268 11778
rect 25136 11144 25188 11150
rect 25136 11086 25188 11092
rect 25148 10810 25176 11086
rect 25136 10804 25188 10810
rect 25136 10746 25188 10752
rect 25044 6724 25096 6730
rect 25044 6666 25096 6672
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25148 6254 25176 6598
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 24504 5658 24532 5850
rect 24768 5772 24820 5778
rect 24768 5714 24820 5720
rect 24504 5630 24624 5658
rect 24596 5574 24624 5630
rect 24492 5568 24544 5574
rect 24492 5510 24544 5516
rect 24584 5568 24636 5574
rect 24584 5510 24636 5516
rect 24116 5468 24412 5488
rect 24172 5466 24196 5468
rect 24252 5466 24276 5468
rect 24332 5466 24356 5468
rect 24194 5414 24196 5466
rect 24258 5414 24270 5466
rect 24332 5414 24334 5466
rect 24172 5412 24196 5414
rect 24252 5412 24276 5414
rect 24332 5412 24356 5414
rect 24116 5392 24412 5412
rect 24504 4690 24532 5510
rect 24584 4752 24636 4758
rect 24584 4694 24636 4700
rect 24492 4684 24544 4690
rect 24492 4626 24544 4632
rect 24116 4380 24412 4400
rect 24172 4378 24196 4380
rect 24252 4378 24276 4380
rect 24332 4378 24356 4380
rect 24194 4326 24196 4378
rect 24258 4326 24270 4378
rect 24332 4326 24334 4378
rect 24172 4324 24196 4326
rect 24252 4324 24276 4326
rect 24332 4324 24356 4326
rect 24116 4304 24412 4324
rect 24596 3738 24624 4694
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24116 3292 24412 3312
rect 24172 3290 24196 3292
rect 24252 3290 24276 3292
rect 24332 3290 24356 3292
rect 24194 3238 24196 3290
rect 24258 3238 24270 3290
rect 24332 3238 24334 3290
rect 24172 3236 24196 3238
rect 24252 3236 24276 3238
rect 24332 3236 24356 3238
rect 24116 3216 24412 3236
rect 24030 2952 24086 2961
rect 23940 2916 23992 2922
rect 24504 2922 24532 3334
rect 24780 2938 24808 5714
rect 25240 5250 25268 11750
rect 25332 11082 25360 18006
rect 25424 16289 25452 18566
rect 25410 16280 25466 16289
rect 25410 16215 25466 16224
rect 25516 16096 25544 21134
rect 25608 18737 25636 22052
rect 25792 22080 25820 25350
rect 25976 24750 26004 25758
rect 26056 25706 26108 25712
rect 26160 25129 26188 26250
rect 26252 25430 26280 26318
rect 26240 25424 26292 25430
rect 26240 25366 26292 25372
rect 26146 25120 26202 25129
rect 26146 25055 26202 25064
rect 26252 24954 26280 25366
rect 26240 24948 26292 24954
rect 26240 24890 26292 24896
rect 25964 24744 26016 24750
rect 25964 24686 26016 24692
rect 26146 24712 26202 24721
rect 25872 23044 25924 23050
rect 25872 22986 25924 22992
rect 25740 22052 25820 22080
rect 25688 22034 25740 22040
rect 25884 21865 25912 22986
rect 25976 22794 26004 24686
rect 26146 24647 26202 24656
rect 26160 24342 26188 24647
rect 26344 24342 26372 26998
rect 26424 26852 26476 26858
rect 26424 26794 26476 26800
rect 26608 26852 26660 26858
rect 26608 26794 26660 26800
rect 26148 24336 26200 24342
rect 26148 24278 26200 24284
rect 26332 24336 26384 24342
rect 26332 24278 26384 24284
rect 26436 24188 26464 26794
rect 26620 26586 26648 26794
rect 26700 26784 26752 26790
rect 26698 26752 26700 26761
rect 26752 26752 26754 26761
rect 26698 26687 26754 26696
rect 26608 26580 26660 26586
rect 26608 26522 26660 26528
rect 26700 25832 26752 25838
rect 26700 25774 26752 25780
rect 26712 25498 26740 25774
rect 26700 25492 26752 25498
rect 26700 25434 26752 25440
rect 26160 24160 26464 24188
rect 25976 22778 26096 22794
rect 25964 22772 26096 22778
rect 26016 22766 26096 22772
rect 25964 22714 26016 22720
rect 25964 22636 26016 22642
rect 25964 22578 26016 22584
rect 25870 21856 25926 21865
rect 25870 21791 25926 21800
rect 25976 21078 26004 22578
rect 26068 21418 26096 22766
rect 26056 21412 26108 21418
rect 26056 21354 26108 21360
rect 25964 21072 26016 21078
rect 25964 21014 26016 21020
rect 25964 20324 26016 20330
rect 25964 20266 26016 20272
rect 25688 19916 25740 19922
rect 25688 19858 25740 19864
rect 25700 19174 25728 19858
rect 25872 19780 25924 19786
rect 25872 19722 25924 19728
rect 25780 19712 25832 19718
rect 25780 19654 25832 19660
rect 25792 19378 25820 19654
rect 25780 19372 25832 19378
rect 25780 19314 25832 19320
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25688 18896 25740 18902
rect 25688 18838 25740 18844
rect 25594 18728 25650 18737
rect 25594 18663 25650 18672
rect 25424 16068 25544 16096
rect 25424 13530 25452 16068
rect 25504 15972 25556 15978
rect 25504 15914 25556 15920
rect 25516 15502 25544 15914
rect 25608 15638 25636 18663
rect 25700 17678 25728 18838
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 25688 16448 25740 16454
rect 25688 16390 25740 16396
rect 25700 16046 25728 16390
rect 25792 16114 25820 19314
rect 25884 19009 25912 19722
rect 25976 19417 26004 20266
rect 25962 19408 26018 19417
rect 25962 19343 26018 19352
rect 26068 19310 26096 21354
rect 26160 20602 26188 24160
rect 26792 24064 26844 24070
rect 26792 24006 26844 24012
rect 26804 23905 26832 24006
rect 26790 23896 26846 23905
rect 26790 23831 26846 23840
rect 26332 23724 26384 23730
rect 26332 23666 26384 23672
rect 26240 23588 26292 23594
rect 26240 23530 26292 23536
rect 26252 22642 26280 23530
rect 26240 22636 26292 22642
rect 26240 22578 26292 22584
rect 26252 22166 26280 22578
rect 26344 22273 26372 23666
rect 26516 23656 26568 23662
rect 26516 23598 26568 23604
rect 26884 23656 26936 23662
rect 26884 23598 26936 23604
rect 26528 23186 26556 23598
rect 26516 23180 26568 23186
rect 26516 23122 26568 23128
rect 26424 23112 26476 23118
rect 26424 23054 26476 23060
rect 26330 22264 26386 22273
rect 26330 22199 26386 22208
rect 26436 22166 26464 23054
rect 26240 22160 26292 22166
rect 26240 22102 26292 22108
rect 26424 22160 26476 22166
rect 26424 22102 26476 22108
rect 26528 21962 26556 23122
rect 26700 23112 26752 23118
rect 26700 23054 26752 23060
rect 26712 22234 26740 23054
rect 26608 22228 26660 22234
rect 26608 22170 26660 22176
rect 26700 22228 26752 22234
rect 26700 22170 26752 22176
rect 26516 21956 26568 21962
rect 26516 21898 26568 21904
rect 26620 21690 26648 22170
rect 26896 22098 26924 23598
rect 26884 22094 26936 22098
rect 26804 22092 26936 22094
rect 26804 22066 26884 22092
rect 26608 21684 26660 21690
rect 26608 21626 26660 21632
rect 26148 20596 26200 20602
rect 26148 20538 26200 20544
rect 26240 20324 26292 20330
rect 26240 20266 26292 20272
rect 26700 20324 26752 20330
rect 26700 20266 26752 20272
rect 26252 19446 26280 20266
rect 26516 19916 26568 19922
rect 26516 19858 26568 19864
rect 26240 19440 26292 19446
rect 26240 19382 26292 19388
rect 26056 19304 26108 19310
rect 26056 19246 26108 19252
rect 25870 19000 25926 19009
rect 25870 18935 25926 18944
rect 25870 18864 25926 18873
rect 25870 18799 25926 18808
rect 25964 18828 26016 18834
rect 25884 18766 25912 18799
rect 25964 18770 26016 18776
rect 25872 18760 25924 18766
rect 25976 18737 26004 18770
rect 25872 18702 25924 18708
rect 25962 18728 26018 18737
rect 25780 16108 25832 16114
rect 25780 16050 25832 16056
rect 25688 16040 25740 16046
rect 25688 15982 25740 15988
rect 25700 15638 25728 15982
rect 25884 15978 25912 18702
rect 25962 18663 26018 18672
rect 26068 18442 26096 19246
rect 26332 19236 26384 19242
rect 26332 19178 26384 19184
rect 26148 19168 26200 19174
rect 26148 19110 26200 19116
rect 26160 18834 26188 19110
rect 26148 18828 26200 18834
rect 26148 18770 26200 18776
rect 26240 18828 26292 18834
rect 26240 18770 26292 18776
rect 25976 18426 26096 18442
rect 26160 18426 26188 18770
rect 26252 18601 26280 18770
rect 26238 18592 26294 18601
rect 26238 18527 26294 18536
rect 25964 18420 26096 18426
rect 26016 18414 26096 18420
rect 26148 18420 26200 18426
rect 25964 18362 26016 18368
rect 26148 18362 26200 18368
rect 26344 17066 26372 19178
rect 26528 17882 26556 19858
rect 26608 18624 26660 18630
rect 26712 18601 26740 20266
rect 26804 19922 26832 22066
rect 26884 22034 26936 22040
rect 26882 21040 26938 21049
rect 26882 20975 26884 20984
rect 26936 20975 26938 20984
rect 26884 20946 26936 20952
rect 26792 19916 26844 19922
rect 26792 19858 26844 19864
rect 26792 19780 26844 19786
rect 26792 19722 26844 19728
rect 26608 18566 26660 18572
rect 26698 18592 26754 18601
rect 26516 17876 26568 17882
rect 26516 17818 26568 17824
rect 26620 17746 26648 18566
rect 26698 18527 26754 18536
rect 26608 17740 26660 17746
rect 26608 17682 26660 17688
rect 26240 17060 26292 17066
rect 26240 17002 26292 17008
rect 26332 17060 26384 17066
rect 26332 17002 26384 17008
rect 26252 16153 26280 17002
rect 26804 16250 26832 19722
rect 26882 17776 26938 17785
rect 26882 17711 26884 17720
rect 26936 17711 26938 17720
rect 26884 17682 26936 17688
rect 26882 17368 26938 17377
rect 26882 17303 26884 17312
rect 26936 17303 26938 17312
rect 26884 17274 26936 17280
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 26238 16144 26294 16153
rect 26238 16079 26294 16088
rect 26240 16040 26292 16046
rect 26240 15982 26292 15988
rect 26516 16040 26568 16046
rect 26516 15982 26568 15988
rect 25872 15972 25924 15978
rect 25872 15914 25924 15920
rect 25962 15736 26018 15745
rect 25962 15671 26018 15680
rect 25596 15632 25648 15638
rect 25596 15574 25648 15580
rect 25688 15632 25740 15638
rect 25688 15574 25740 15580
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 25412 13524 25464 13530
rect 25412 13466 25464 13472
rect 25516 12782 25544 15438
rect 25608 12782 25636 15574
rect 25700 14550 25728 15574
rect 25872 14884 25924 14890
rect 25872 14826 25924 14832
rect 25688 14544 25740 14550
rect 25688 14486 25740 14492
rect 25688 13524 25740 13530
rect 25688 13466 25740 13472
rect 25504 12776 25556 12782
rect 25504 12718 25556 12724
rect 25596 12776 25648 12782
rect 25596 12718 25648 12724
rect 25412 12436 25464 12442
rect 25412 12378 25464 12384
rect 25424 11694 25452 12378
rect 25412 11688 25464 11694
rect 25516 11676 25544 12718
rect 25700 12714 25728 13466
rect 25884 13190 25912 14826
rect 25976 14550 26004 15671
rect 26056 15020 26108 15026
rect 26056 14962 26108 14968
rect 26068 14618 26096 14962
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 25964 14544 26016 14550
rect 25964 14486 26016 14492
rect 25964 13864 26016 13870
rect 25964 13806 26016 13812
rect 25872 13184 25924 13190
rect 25872 13126 25924 13132
rect 25688 12708 25740 12714
rect 25688 12650 25740 12656
rect 25594 12472 25650 12481
rect 25594 12407 25650 12416
rect 25608 11830 25636 12407
rect 25596 11824 25648 11830
rect 25596 11766 25648 11772
rect 25516 11648 25636 11676
rect 25412 11630 25464 11636
rect 25320 11076 25372 11082
rect 25320 11018 25372 11024
rect 25332 10674 25360 11018
rect 25320 10668 25372 10674
rect 25320 10610 25372 10616
rect 25504 10668 25556 10674
rect 25504 10610 25556 10616
rect 25412 10600 25464 10606
rect 25412 10542 25464 10548
rect 25424 8906 25452 10542
rect 25516 10130 25544 10610
rect 25504 10124 25556 10130
rect 25504 10066 25556 10072
rect 25412 8900 25464 8906
rect 25412 8842 25464 8848
rect 25412 7336 25464 7342
rect 25516 7290 25544 10066
rect 25608 9586 25636 11648
rect 25700 11218 25728 12650
rect 25884 12434 25912 13126
rect 25976 12889 26004 13806
rect 26148 13184 26200 13190
rect 26148 13126 26200 13132
rect 25962 12880 26018 12889
rect 25962 12815 26018 12824
rect 26160 12782 26188 13126
rect 26148 12776 26200 12782
rect 26148 12718 26200 12724
rect 26056 12708 26108 12714
rect 26056 12650 26108 12656
rect 25884 12406 26004 12434
rect 25976 12102 26004 12406
rect 25964 12096 26016 12102
rect 25964 12038 26016 12044
rect 25976 11694 26004 12038
rect 25964 11688 26016 11694
rect 25964 11630 26016 11636
rect 25688 11212 25740 11218
rect 25688 11154 25740 11160
rect 25872 10736 25924 10742
rect 25872 10678 25924 10684
rect 25884 10266 25912 10678
rect 25976 10674 26004 11630
rect 25964 10668 26016 10674
rect 25964 10610 26016 10616
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 25596 9580 25648 9586
rect 25596 9522 25648 9528
rect 25608 8974 25636 9522
rect 25884 9178 25912 10202
rect 26068 9586 26096 12650
rect 26160 12442 26188 12718
rect 26148 12436 26200 12442
rect 26148 12378 26200 12384
rect 26252 12238 26280 15982
rect 26424 15700 26476 15706
rect 26424 15642 26476 15648
rect 26436 14958 26464 15642
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26424 14408 26476 14414
rect 26528 14396 26556 15982
rect 26896 15337 26924 16594
rect 26882 15328 26938 15337
rect 26882 15263 26938 15272
rect 26476 14368 26556 14396
rect 26424 14350 26476 14356
rect 26436 12238 26464 14350
rect 26700 14340 26752 14346
rect 26700 14282 26752 14288
rect 26712 12986 26740 14282
rect 26792 13864 26844 13870
rect 26792 13806 26844 13812
rect 26700 12980 26752 12986
rect 26700 12922 26752 12928
rect 26516 12640 26568 12646
rect 26516 12582 26568 12588
rect 26240 12232 26292 12238
rect 26240 12174 26292 12180
rect 26424 12232 26476 12238
rect 26424 12174 26476 12180
rect 26148 11756 26200 11762
rect 26148 11698 26200 11704
rect 26160 11665 26188 11698
rect 26146 11656 26202 11665
rect 26146 11591 26202 11600
rect 26146 11248 26202 11257
rect 26146 11183 26148 11192
rect 26200 11183 26202 11192
rect 26148 11154 26200 11160
rect 26240 10464 26292 10470
rect 26240 10406 26292 10412
rect 26056 9580 26108 9586
rect 26056 9522 26108 9528
rect 25872 9172 25924 9178
rect 25924 9132 26004 9160
rect 25872 9114 25924 9120
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 25872 8424 25924 8430
rect 25870 8392 25872 8401
rect 25924 8392 25926 8401
rect 25870 8327 25926 8336
rect 25596 8288 25648 8294
rect 25596 8230 25648 8236
rect 25608 7954 25636 8230
rect 25976 8022 26004 9132
rect 26068 8838 26096 9522
rect 26252 9518 26280 10406
rect 26436 9654 26464 12174
rect 26528 11558 26556 12582
rect 26712 12306 26740 12922
rect 26700 12300 26752 12306
rect 26700 12242 26752 12248
rect 26804 12073 26832 13806
rect 26790 12064 26846 12073
rect 26790 11999 26846 12008
rect 26516 11552 26568 11558
rect 26516 11494 26568 11500
rect 26988 11234 27016 37266
rect 27896 36848 27948 36854
rect 27896 36790 27948 36796
rect 27436 36712 27488 36718
rect 27436 36654 27488 36660
rect 27342 35048 27398 35057
rect 27342 34983 27398 34992
rect 27356 34746 27384 34983
rect 27448 34921 27476 36654
rect 27804 36576 27856 36582
rect 27804 36518 27856 36524
rect 27434 34912 27490 34921
rect 27434 34847 27490 34856
rect 27344 34740 27396 34746
rect 27344 34682 27396 34688
rect 27816 34474 27844 36518
rect 27908 35630 27936 36790
rect 27988 36032 28040 36038
rect 27988 35974 28040 35980
rect 27896 35624 27948 35630
rect 27896 35566 27948 35572
rect 28000 35222 28028 35974
rect 27988 35216 28040 35222
rect 27988 35158 28040 35164
rect 27804 34468 27856 34474
rect 27804 34410 27856 34416
rect 27252 33924 27304 33930
rect 27252 33866 27304 33872
rect 27264 33658 27292 33866
rect 27252 33652 27304 33658
rect 27252 33594 27304 33600
rect 27988 33652 28040 33658
rect 27988 33594 28040 33600
rect 28000 33561 28028 33594
rect 27986 33552 28042 33561
rect 27986 33487 28042 33496
rect 27252 32972 27304 32978
rect 27252 32914 27304 32920
rect 27264 31754 27292 32914
rect 27436 32292 27488 32298
rect 27436 32234 27488 32240
rect 27264 31726 27384 31754
rect 27068 30048 27120 30054
rect 27068 29990 27120 29996
rect 27080 29782 27108 29990
rect 27068 29776 27120 29782
rect 27068 29718 27120 29724
rect 27160 29028 27212 29034
rect 27160 28970 27212 28976
rect 27172 27985 27200 28970
rect 27158 27976 27214 27985
rect 27158 27911 27214 27920
rect 27252 27940 27304 27946
rect 27252 27882 27304 27888
rect 27264 27606 27292 27882
rect 27252 27600 27304 27606
rect 27252 27542 27304 27548
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 27172 22030 27200 23598
rect 27264 23118 27292 27542
rect 27252 23112 27304 23118
rect 27252 23054 27304 23060
rect 27160 22024 27212 22030
rect 27160 21966 27212 21972
rect 27172 19786 27200 21966
rect 27160 19780 27212 19786
rect 27160 19722 27212 19728
rect 27252 16040 27304 16046
rect 27252 15982 27304 15988
rect 27264 14346 27292 15982
rect 27252 14340 27304 14346
rect 27252 14282 27304 14288
rect 26804 11206 27016 11234
rect 26424 9648 26476 9654
rect 26424 9590 26476 9596
rect 26240 9512 26292 9518
rect 26240 9454 26292 9460
rect 26146 9208 26202 9217
rect 26146 9143 26202 9152
rect 26056 8832 26108 8838
rect 26056 8774 26108 8780
rect 26160 8022 26188 9143
rect 26436 9110 26464 9590
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26424 9104 26476 9110
rect 26424 9046 26476 9052
rect 26620 8498 26648 9454
rect 26804 9110 26832 11206
rect 26884 11076 26936 11082
rect 26884 11018 26936 11024
rect 26896 10441 26924 11018
rect 26882 10432 26938 10441
rect 26882 10367 26938 10376
rect 27160 9512 27212 9518
rect 27160 9454 27212 9460
rect 26792 9104 26844 9110
rect 26792 9046 26844 9052
rect 26608 8492 26660 8498
rect 26608 8434 26660 8440
rect 26240 8424 26292 8430
rect 26240 8366 26292 8372
rect 25964 8016 26016 8022
rect 25964 7958 26016 7964
rect 26148 8016 26200 8022
rect 26148 7958 26200 7964
rect 25596 7948 25648 7954
rect 25596 7890 25648 7896
rect 25464 7284 25544 7290
rect 25412 7278 25544 7284
rect 25424 7262 25544 7278
rect 25516 6390 25544 7262
rect 25504 6384 25556 6390
rect 25318 6352 25374 6361
rect 25504 6326 25556 6332
rect 25318 6287 25374 6296
rect 25332 5914 25360 6287
rect 25320 5908 25372 5914
rect 25320 5850 25372 5856
rect 25240 5222 25452 5250
rect 25228 5160 25280 5166
rect 25228 5102 25280 5108
rect 25044 5024 25096 5030
rect 25044 4966 25096 4972
rect 25056 4214 25084 4966
rect 25044 4208 25096 4214
rect 25044 4150 25096 4156
rect 25136 3528 25188 3534
rect 25136 3470 25188 3476
rect 25148 3126 25176 3470
rect 25136 3120 25188 3126
rect 25136 3062 25188 3068
rect 24030 2887 24086 2896
rect 24492 2916 24544 2922
rect 23940 2858 23992 2864
rect 24780 2910 25176 2938
rect 24492 2858 24544 2864
rect 24768 2848 24820 2854
rect 24768 2790 24820 2796
rect 24780 2666 24808 2790
rect 24858 2680 24914 2689
rect 24780 2638 24858 2666
rect 24858 2615 24914 2624
rect 24490 2544 24546 2553
rect 23020 2508 23072 2514
rect 23020 2450 23072 2456
rect 23388 2508 23440 2514
rect 24490 2479 24492 2488
rect 23388 2450 23440 2456
rect 24544 2479 24546 2488
rect 24492 2450 24544 2456
rect 21364 2440 21416 2446
rect 21364 2382 21416 2388
rect 22468 2440 22520 2446
rect 22468 2382 22520 2388
rect 22480 800 22508 2382
rect 25044 2372 25096 2378
rect 25044 2314 25096 2320
rect 25056 2281 25084 2314
rect 25042 2272 25098 2281
rect 24116 2204 24412 2224
rect 25042 2207 25098 2216
rect 24172 2202 24196 2204
rect 24252 2202 24276 2204
rect 24332 2202 24356 2204
rect 24194 2150 24196 2202
rect 24258 2150 24270 2202
rect 24332 2150 24334 2202
rect 24172 2148 24196 2150
rect 24252 2148 24276 2150
rect 24332 2148 24356 2150
rect 24116 2128 24412 2148
rect 23756 1284 23808 1290
rect 23756 1226 23808 1232
rect 23768 800 23796 1226
rect 25148 800 25176 2910
rect 25240 2446 25268 5102
rect 25424 4758 25452 5222
rect 25412 4752 25464 4758
rect 25412 4694 25464 4700
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 25332 3738 25360 4626
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 25424 3602 25452 4694
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 25412 3596 25464 3602
rect 25412 3538 25464 3544
rect 25516 3097 25544 3878
rect 25502 3088 25558 3097
rect 25502 3023 25558 3032
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25412 2304 25464 2310
rect 25412 2246 25464 2252
rect 25424 1873 25452 2246
rect 25608 1970 25636 7890
rect 25964 7744 26016 7750
rect 25964 7686 26016 7692
rect 25688 7268 25740 7274
rect 25688 7210 25740 7216
rect 25700 7002 25728 7210
rect 25976 7002 26004 7686
rect 26148 7200 26200 7206
rect 26148 7142 26200 7148
rect 25688 6996 25740 7002
rect 25688 6938 25740 6944
rect 25964 6996 26016 7002
rect 25964 6938 26016 6944
rect 26160 6798 26188 7142
rect 25872 6792 25924 6798
rect 25872 6734 25924 6740
rect 26148 6792 26200 6798
rect 26148 6734 26200 6740
rect 25884 6186 25912 6734
rect 25964 6384 26016 6390
rect 25964 6326 26016 6332
rect 25872 6180 25924 6186
rect 25872 6122 25924 6128
rect 25884 5778 25912 6122
rect 25976 5794 26004 6326
rect 26252 6322 26280 8366
rect 26804 8294 26832 9046
rect 26976 9036 27028 9042
rect 26976 8978 27028 8984
rect 26988 8634 27016 8978
rect 26976 8628 27028 8634
rect 26976 8570 27028 8576
rect 27172 8498 27200 9454
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 26792 8288 26844 8294
rect 26792 8230 26844 8236
rect 26792 7744 26844 7750
rect 26792 7686 26844 7692
rect 26804 7585 26832 7686
rect 26790 7576 26846 7585
rect 26790 7511 26846 7520
rect 26240 6316 26292 6322
rect 26240 6258 26292 6264
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 26148 6112 26200 6118
rect 26148 6054 26200 6060
rect 26054 5944 26110 5953
rect 26054 5879 26056 5888
rect 26108 5879 26110 5888
rect 26056 5850 26108 5856
rect 25780 5772 25832 5778
rect 25780 5714 25832 5720
rect 25872 5772 25924 5778
rect 25976 5766 26096 5794
rect 25872 5714 25924 5720
rect 25792 3602 25820 5714
rect 26068 4486 26096 5766
rect 26160 5710 26188 6054
rect 26424 5772 26476 5778
rect 26424 5714 26476 5720
rect 26148 5704 26200 5710
rect 26148 5646 26200 5652
rect 26056 4480 26108 4486
rect 26056 4422 26108 4428
rect 25964 4208 26016 4214
rect 25964 4150 26016 4156
rect 25872 4004 25924 4010
rect 25872 3946 25924 3952
rect 25780 3596 25832 3602
rect 25780 3538 25832 3544
rect 25792 2990 25820 3538
rect 25884 3126 25912 3946
rect 25872 3120 25924 3126
rect 25872 3062 25924 3068
rect 25976 2990 26004 4150
rect 26068 4078 26096 4422
rect 26056 4072 26108 4078
rect 26056 4014 26108 4020
rect 26146 3632 26202 3641
rect 26146 3567 26202 3576
rect 26160 3534 26188 3567
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 26436 3466 26464 5714
rect 26528 5370 26556 6258
rect 26700 5636 26752 5642
rect 26700 5578 26752 5584
rect 26884 5636 26936 5642
rect 26884 5578 26936 5584
rect 26516 5364 26568 5370
rect 26516 5306 26568 5312
rect 26606 5128 26662 5137
rect 26606 5063 26608 5072
rect 26660 5063 26662 5072
rect 26608 5034 26660 5040
rect 26712 4078 26740 5578
rect 26896 5545 26924 5578
rect 26882 5536 26938 5545
rect 26882 5471 26938 5480
rect 27356 5370 27384 31726
rect 27448 29306 27476 32234
rect 27620 32224 27672 32230
rect 27620 32166 27672 32172
rect 27528 30796 27580 30802
rect 27528 30738 27580 30744
rect 27540 29617 27568 30738
rect 27526 29608 27582 29617
rect 27526 29543 27582 29552
rect 27436 29300 27488 29306
rect 27436 29242 27488 29248
rect 27632 29102 27660 32166
rect 27988 31680 28040 31686
rect 27988 31622 28040 31628
rect 28000 30938 28028 31622
rect 27988 30932 28040 30938
rect 27988 30874 28040 30880
rect 27988 30592 28040 30598
rect 27988 30534 28040 30540
rect 28000 29782 28028 30534
rect 27988 29776 28040 29782
rect 27988 29718 28040 29724
rect 27620 29096 27672 29102
rect 27620 29038 27672 29044
rect 27712 29096 27764 29102
rect 27712 29038 27764 29044
rect 28264 29096 28316 29102
rect 28264 29038 28316 29044
rect 27528 28008 27580 28014
rect 27528 27950 27580 27956
rect 27540 27674 27568 27950
rect 27620 27872 27672 27878
rect 27620 27814 27672 27820
rect 27528 27668 27580 27674
rect 27528 27610 27580 27616
rect 27436 25764 27488 25770
rect 27436 25706 27488 25712
rect 27448 24954 27476 25706
rect 27540 25498 27568 27610
rect 27632 27334 27660 27814
rect 27620 27328 27672 27334
rect 27620 27270 27672 27276
rect 27528 25492 27580 25498
rect 27528 25434 27580 25440
rect 27528 25152 27580 25158
rect 27528 25094 27580 25100
rect 27436 24948 27488 24954
rect 27436 24890 27488 24896
rect 27540 24313 27568 25094
rect 27526 24304 27582 24313
rect 27526 24239 27582 24248
rect 27632 23730 27660 27270
rect 27724 27130 27752 29038
rect 27896 28960 27948 28966
rect 27896 28902 27948 28908
rect 27804 27940 27856 27946
rect 27804 27882 27856 27888
rect 27712 27124 27764 27130
rect 27712 27066 27764 27072
rect 27816 26926 27844 27882
rect 27804 26920 27856 26926
rect 27804 26862 27856 26868
rect 27804 26036 27856 26042
rect 27804 25978 27856 25984
rect 27816 24750 27844 25978
rect 27908 24886 27936 28902
rect 27988 28620 28040 28626
rect 27988 28562 28040 28568
rect 28000 28218 28028 28562
rect 28276 28490 28304 29038
rect 28264 28484 28316 28490
rect 28264 28426 28316 28432
rect 27988 28212 28040 28218
rect 27988 28154 28040 28160
rect 27988 28076 28040 28082
rect 27988 28018 28040 28024
rect 28000 26518 28028 28018
rect 28172 27328 28224 27334
rect 28172 27270 28224 27276
rect 28184 26994 28212 27270
rect 28172 26988 28224 26994
rect 28172 26930 28224 26936
rect 27988 26512 28040 26518
rect 27988 26454 28040 26460
rect 28170 26344 28226 26353
rect 28170 26279 28172 26288
rect 28224 26279 28226 26288
rect 28172 26250 28224 26256
rect 27988 25832 28040 25838
rect 27988 25774 28040 25780
rect 27896 24880 27948 24886
rect 27896 24822 27948 24828
rect 27804 24744 27856 24750
rect 27804 24686 27856 24692
rect 27620 23724 27672 23730
rect 27620 23666 27672 23672
rect 27804 22976 27856 22982
rect 27804 22918 27856 22924
rect 27436 22500 27488 22506
rect 27436 22442 27488 22448
rect 27448 21690 27476 22442
rect 27436 21684 27488 21690
rect 27436 21626 27488 21632
rect 27816 21486 27844 22918
rect 27908 22094 27936 24822
rect 28000 23866 28028 25774
rect 28080 25696 28132 25702
rect 28080 25638 28132 25644
rect 28092 24750 28120 25638
rect 28080 24744 28132 24750
rect 28080 24686 28132 24692
rect 28172 24132 28224 24138
rect 28172 24074 28224 24080
rect 27988 23860 28040 23866
rect 27988 23802 28040 23808
rect 28184 23497 28212 24074
rect 28170 23488 28226 23497
rect 28170 23423 28226 23432
rect 28080 23316 28132 23322
rect 28080 23258 28132 23264
rect 28092 22778 28120 23258
rect 28170 23080 28226 23089
rect 28170 23015 28172 23024
rect 28224 23015 28226 23024
rect 28172 22986 28224 22992
rect 28080 22772 28132 22778
rect 28080 22714 28132 22720
rect 27908 22066 28028 22094
rect 28000 21554 28028 22066
rect 27988 21548 28040 21554
rect 27988 21490 28040 21496
rect 27804 21480 27856 21486
rect 27526 21448 27582 21457
rect 27804 21422 27856 21428
rect 27526 21383 27582 21392
rect 27540 20602 27568 21383
rect 27528 20596 27580 20602
rect 27528 20538 27580 20544
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 27436 19236 27488 19242
rect 27436 19178 27488 19184
rect 27448 18426 27476 19178
rect 27436 18420 27488 18426
rect 27436 18362 27488 18368
rect 27816 18222 27844 19654
rect 28000 18272 28028 21490
rect 28092 21486 28120 22714
rect 28080 21480 28132 21486
rect 28080 21422 28132 21428
rect 28080 20800 28132 20806
rect 28080 20742 28132 20748
rect 28092 20641 28120 20742
rect 28078 20632 28134 20641
rect 28078 20567 28134 20576
rect 28172 20324 28224 20330
rect 28172 20266 28224 20272
rect 28080 20256 28132 20262
rect 28184 20233 28212 20266
rect 28080 20198 28132 20204
rect 28170 20224 28226 20233
rect 28092 19514 28120 20198
rect 28170 20159 28226 20168
rect 28170 19816 28226 19825
rect 28170 19751 28172 19760
rect 28224 19751 28226 19760
rect 28172 19722 28224 19728
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 28092 18426 28120 19450
rect 28172 18692 28224 18698
rect 28172 18634 28224 18640
rect 28080 18420 28132 18426
rect 28080 18362 28132 18368
rect 28080 18284 28132 18290
rect 28000 18244 28080 18272
rect 28080 18226 28132 18232
rect 27804 18216 27856 18222
rect 27804 18158 27856 18164
rect 27712 18080 27764 18086
rect 27712 18022 27764 18028
rect 27436 16992 27488 16998
rect 27436 16934 27488 16940
rect 27448 14958 27476 16934
rect 27724 16726 27752 18022
rect 27804 16992 27856 16998
rect 27804 16934 27856 16940
rect 27896 16992 27948 16998
rect 27896 16934 27948 16940
rect 27712 16720 27764 16726
rect 27712 16662 27764 16668
rect 27528 16040 27580 16046
rect 27528 15982 27580 15988
rect 27540 15706 27568 15982
rect 27528 15700 27580 15706
rect 27528 15642 27580 15648
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 27434 14784 27490 14793
rect 27434 14719 27490 14728
rect 27448 14074 27476 14719
rect 27540 14521 27568 15302
rect 27816 15162 27844 16934
rect 27908 15162 27936 16934
rect 27988 16176 28040 16182
rect 27988 16118 28040 16124
rect 27804 15156 27856 15162
rect 27804 15098 27856 15104
rect 27896 15156 27948 15162
rect 27896 15098 27948 15104
rect 28000 14550 28028 16118
rect 27988 14544 28040 14550
rect 27526 14512 27582 14521
rect 27988 14486 28040 14492
rect 27526 14447 27582 14456
rect 27988 14272 28040 14278
rect 27988 14214 28040 14220
rect 27436 14068 27488 14074
rect 27436 14010 27488 14016
rect 28000 13870 28028 14214
rect 27988 13864 28040 13870
rect 27988 13806 28040 13812
rect 27896 13796 27948 13802
rect 27896 13738 27948 13744
rect 27908 12850 27936 13738
rect 27896 12844 27948 12850
rect 27896 12786 27948 12792
rect 27436 12640 27488 12646
rect 27436 12582 27488 12588
rect 27528 12640 27580 12646
rect 27528 12582 27580 12588
rect 27448 11694 27476 12582
rect 27540 12442 27568 12582
rect 27528 12436 27580 12442
rect 27528 12378 27580 12384
rect 27908 11898 27936 12786
rect 27896 11892 27948 11898
rect 27896 11834 27948 11840
rect 27804 11756 27856 11762
rect 27804 11698 27856 11704
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 27528 11076 27580 11082
rect 27528 11018 27580 11024
rect 27540 10033 27568 11018
rect 27526 10024 27582 10033
rect 27526 9959 27582 9968
rect 27436 9512 27488 9518
rect 27436 9454 27488 9460
rect 27448 8430 27476 9454
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 27540 8498 27568 8774
rect 27528 8492 27580 8498
rect 27528 8434 27580 8440
rect 27436 8424 27488 8430
rect 27436 8366 27488 8372
rect 27436 7200 27488 7206
rect 27436 7142 27488 7148
rect 27528 7200 27580 7206
rect 27528 7142 27580 7148
rect 27448 6254 27476 7142
rect 27540 6458 27568 7142
rect 27816 6914 27844 11698
rect 27988 10532 28040 10538
rect 27988 10474 28040 10480
rect 27896 9920 27948 9926
rect 27896 9862 27948 9868
rect 27908 9110 27936 9862
rect 27896 9104 27948 9110
rect 27896 9046 27948 9052
rect 28000 8634 28028 10474
rect 28092 10266 28120 18226
rect 28184 18193 28212 18634
rect 28170 18184 28226 18193
rect 28170 18119 28226 18128
rect 28172 17604 28224 17610
rect 28172 17546 28224 17552
rect 28184 16969 28212 17546
rect 28170 16960 28226 16969
rect 28170 16895 28226 16904
rect 28172 16652 28224 16658
rect 28172 16594 28224 16600
rect 28184 16561 28212 16594
rect 28170 16552 28226 16561
rect 28170 16487 28226 16496
rect 28172 14340 28224 14346
rect 28172 14282 28224 14288
rect 28184 14113 28212 14282
rect 28170 14104 28226 14113
rect 28170 14039 28226 14048
rect 28172 13864 28224 13870
rect 28172 13806 28224 13812
rect 28184 13705 28212 13806
rect 28170 13696 28226 13705
rect 28170 13631 28226 13640
rect 28170 13288 28226 13297
rect 28170 13223 28172 13232
rect 28224 13223 28226 13232
rect 28172 13194 28224 13200
rect 28276 11762 28304 28426
rect 28356 27056 28408 27062
rect 28356 26998 28408 27004
rect 28368 17202 28396 26998
rect 28356 17196 28408 17202
rect 28356 17138 28408 17144
rect 28368 12850 28396 17138
rect 28356 12844 28408 12850
rect 28356 12786 28408 12792
rect 28264 11756 28316 11762
rect 28264 11698 28316 11704
rect 28264 10464 28316 10470
rect 28264 10406 28316 10412
rect 28080 10260 28132 10266
rect 28132 10220 28212 10248
rect 28080 10202 28132 10208
rect 28080 8832 28132 8838
rect 28080 8774 28132 8780
rect 27988 8628 28040 8634
rect 27988 8570 28040 8576
rect 28092 7993 28120 8774
rect 28184 8498 28212 10220
rect 28276 9178 28304 10406
rect 28368 10130 28396 12786
rect 29000 11076 29052 11082
rect 29000 11018 29052 11024
rect 29012 10849 29040 11018
rect 28998 10840 29054 10849
rect 28998 10775 29054 10784
rect 28356 10124 28408 10130
rect 28356 10066 28408 10072
rect 28264 9172 28316 9178
rect 28264 9114 28316 9120
rect 28172 8492 28224 8498
rect 28172 8434 28224 8440
rect 28276 8430 28304 9114
rect 28264 8424 28316 8430
rect 28264 8366 28316 8372
rect 28078 7984 28134 7993
rect 28078 7919 28134 7928
rect 28368 7886 28396 10066
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 28172 7812 28224 7818
rect 28172 7754 28224 7760
rect 28080 7200 28132 7206
rect 28184 7177 28212 7754
rect 28368 7410 28396 7822
rect 28356 7404 28408 7410
rect 28356 7346 28408 7352
rect 28080 7142 28132 7148
rect 28170 7168 28226 7177
rect 27816 6886 27936 6914
rect 27528 6452 27580 6458
rect 27528 6394 27580 6400
rect 27436 6248 27488 6254
rect 27436 6190 27488 6196
rect 27436 5568 27488 5574
rect 27436 5510 27488 5516
rect 27344 5364 27396 5370
rect 27264 5324 27344 5352
rect 26790 4312 26846 4321
rect 27264 4282 27292 5324
rect 27344 5306 27396 5312
rect 27344 5228 27396 5234
rect 27344 5170 27396 5176
rect 26790 4247 26846 4256
rect 27252 4276 27304 4282
rect 26700 4072 26752 4078
rect 26700 4014 26752 4020
rect 26804 3738 26832 4247
rect 27252 4218 27304 4224
rect 26792 3732 26844 3738
rect 26792 3674 26844 3680
rect 26424 3460 26476 3466
rect 26424 3402 26476 3408
rect 27264 3126 27292 4218
rect 27252 3120 27304 3126
rect 27252 3062 27304 3068
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 25964 2984 26016 2990
rect 25964 2926 26016 2932
rect 26790 2952 26846 2961
rect 26790 2887 26792 2896
rect 26844 2887 26846 2896
rect 26976 2916 27028 2922
rect 26792 2858 26844 2864
rect 26976 2858 27028 2864
rect 25872 2372 25924 2378
rect 25872 2314 25924 2320
rect 26056 2372 26108 2378
rect 26056 2314 26108 2320
rect 25596 1964 25648 1970
rect 25596 1906 25648 1912
rect 25410 1864 25466 1873
rect 25410 1799 25466 1808
rect 25884 1057 25912 2314
rect 25870 1048 25926 1057
rect 25870 983 25926 992
rect 2962 640 3018 649
rect 2962 575 3018 584
rect 3330 -800 3386 800
rect 4710 -800 4766 800
rect 6090 -800 6146 800
rect 7470 -800 7526 800
rect 8758 -800 8814 800
rect 10138 -800 10194 800
rect 11518 -800 11574 800
rect 12898 -800 12954 800
rect 14278 -800 14334 800
rect 15658 -800 15714 800
rect 16946 -800 17002 800
rect 18326 -800 18382 800
rect 19706 -800 19762 800
rect 21086 -800 21142 800
rect 22466 -800 22522 800
rect 23754 -800 23810 800
rect 25134 -800 25190 800
rect 26068 241 26096 2314
rect 26148 2304 26200 2310
rect 26148 2246 26200 2252
rect 26160 649 26188 2246
rect 26516 2100 26568 2106
rect 26516 2042 26568 2048
rect 26528 800 26556 2042
rect 26988 1465 27016 2858
rect 27264 2854 27292 3062
rect 27356 2854 27384 5170
rect 27448 4729 27476 5510
rect 27712 5092 27764 5098
rect 27712 5034 27764 5040
rect 27528 5024 27580 5030
rect 27528 4966 27580 4972
rect 27434 4720 27490 4729
rect 27434 4655 27490 4664
rect 27540 3194 27568 4966
rect 27724 4554 27752 5034
rect 27712 4548 27764 4554
rect 27712 4490 27764 4496
rect 27908 4010 27936 6886
rect 28092 6100 28120 7142
rect 28170 7103 28226 7112
rect 28170 6760 28226 6769
rect 28170 6695 28172 6704
rect 28224 6695 28226 6704
rect 28172 6666 28224 6672
rect 28172 6112 28224 6118
rect 28092 6072 28172 6100
rect 28172 6054 28224 6060
rect 28184 5846 28212 6054
rect 28172 5840 28224 5846
rect 28172 5782 28224 5788
rect 28080 4480 28132 4486
rect 28080 4422 28132 4428
rect 27896 4004 27948 4010
rect 27896 3946 27948 3952
rect 28092 3913 28120 4422
rect 28078 3904 28134 3913
rect 28078 3839 28134 3848
rect 28170 3496 28226 3505
rect 28170 3431 28172 3440
rect 28224 3431 28226 3440
rect 28172 3402 28224 3408
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 29276 3392 29328 3398
rect 29276 3334 29328 3340
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 27908 3058 27936 3334
rect 27896 3052 27948 3058
rect 27896 2994 27948 3000
rect 27252 2848 27304 2854
rect 27252 2790 27304 2796
rect 27344 2848 27396 2854
rect 27344 2790 27396 2796
rect 27896 2848 27948 2854
rect 27896 2790 27948 2796
rect 27160 2508 27212 2514
rect 27160 2450 27212 2456
rect 27172 2038 27200 2450
rect 27160 2032 27212 2038
rect 27160 1974 27212 1980
rect 26974 1456 27030 1465
rect 26974 1391 27030 1400
rect 27908 800 27936 2790
rect 29288 800 29316 3334
rect 26146 640 26202 649
rect 26146 575 26202 584
rect 26054 232 26110 241
rect 26054 167 26110 176
rect 26514 -800 26570 800
rect 27894 -800 27950 800
rect 29274 -800 29330 800
<< via2 >>
rect 2778 55664 2834 55720
rect 3882 55256 3938 55312
rect 3238 54848 3294 54904
rect 3146 54440 3202 54496
rect 2962 54032 3018 54088
rect 1858 51856 1914 51912
rect 1950 51584 2006 51640
rect 1490 50768 1546 50824
rect 1398 50360 1454 50416
rect 1858 50224 1914 50280
rect 1950 49952 2006 50008
rect 1398 49136 1454 49192
rect 1950 47912 2006 47968
rect 1306 42608 1362 42664
rect 1950 45464 2006 45520
rect 1398 42200 1454 42256
rect 1398 38120 1454 38176
rect 1950 43424 2006 43480
rect 1950 40976 2006 41032
rect 2778 52436 2780 52456
rect 2780 52436 2832 52456
rect 2832 52436 2834 52456
rect 2778 52400 2834 52436
rect 2778 52012 2834 52048
rect 2778 51992 2780 52012
rect 2780 51992 2832 52012
rect 2832 51992 2834 52012
rect 2778 51176 2834 51232
rect 2686 50904 2742 50960
rect 2594 50788 2650 50824
rect 2594 50768 2596 50788
rect 2596 50768 2648 50788
rect 2648 50768 2650 50788
rect 23570 55256 23626 55312
rect 4066 53624 4122 53680
rect 3606 53216 3662 53272
rect 3422 52808 3478 52864
rect 5588 53338 5644 53340
rect 5668 53338 5724 53340
rect 5748 53338 5804 53340
rect 5828 53338 5884 53340
rect 5588 53286 5614 53338
rect 5614 53286 5644 53338
rect 5668 53286 5678 53338
rect 5678 53286 5724 53338
rect 5748 53286 5794 53338
rect 5794 53286 5804 53338
rect 5828 53286 5858 53338
rect 5858 53286 5884 53338
rect 5588 53284 5644 53286
rect 5668 53284 5724 53286
rect 5748 53284 5804 53286
rect 5828 53284 5884 53286
rect 3330 51468 3386 51504
rect 3330 51448 3332 51468
rect 3332 51448 3384 51468
rect 3384 51448 3386 51468
rect 2778 49544 2834 49600
rect 2870 48728 2926 48784
rect 2962 48320 3018 48376
rect 2778 47504 2834 47560
rect 1950 38936 2006 38992
rect 1674 36488 1730 36544
rect 1398 33652 1454 33688
rect 1398 33632 1400 33652
rect 1400 33632 1452 33652
rect 1452 33632 1454 33652
rect 1398 30368 1454 30424
rect 1674 34892 1676 34912
rect 1676 34892 1728 34912
rect 1728 34892 1730 34912
rect 1674 34856 1730 34892
rect 1950 35264 2006 35320
rect 2042 34484 2044 34504
rect 2044 34484 2096 34504
rect 2096 34484 2098 34504
rect 2042 34448 2098 34484
rect 2042 34060 2098 34096
rect 2042 34040 2044 34060
rect 2044 34040 2096 34060
rect 2096 34040 2098 34060
rect 2226 38256 2282 38312
rect 1950 29552 2006 29608
rect 1858 29144 1914 29200
rect 1858 28736 1914 28792
rect 2870 46280 2926 46336
rect 2962 45056 3018 45112
rect 2870 44648 2926 44704
rect 3790 47096 3846 47152
rect 2778 44240 2834 44296
rect 2778 43016 2834 43072
rect 2778 41792 2834 41848
rect 3514 46688 3570 46744
rect 3422 45872 3478 45928
rect 3422 43832 3478 43888
rect 2962 41384 3018 41440
rect 3146 40568 3202 40624
rect 2778 39344 2834 39400
rect 2870 38528 2926 38584
rect 2778 37712 2834 37768
rect 2778 36896 2834 36952
rect 2778 36080 2834 36136
rect 2962 37304 3018 37360
rect 2870 35672 2926 35728
rect 2778 32408 2834 32464
rect 1766 28092 1768 28112
rect 1768 28092 1820 28112
rect 1820 28092 1822 28112
rect 1766 28056 1822 28092
rect 1950 27512 2006 27568
rect 1950 26696 2006 26752
rect 1950 26288 2006 26344
rect 1398 22208 1454 22264
rect 1582 22616 1638 22672
rect 1858 25880 1914 25936
rect 1766 25472 1822 25528
rect 2410 28872 2466 28928
rect 3606 39752 3662 39808
rect 2778 29960 2834 30016
rect 1950 23432 2006 23488
rect 1582 20984 1638 21040
rect 1674 20168 1730 20224
rect 1950 19760 2006 19816
rect 1858 19352 1914 19408
rect 1858 18944 1914 19000
rect 1490 10784 1546 10840
rect 1582 9968 1638 10024
rect 1490 6704 1546 6760
rect 1950 16904 2006 16960
rect 1950 16496 2006 16552
rect 1858 16088 1914 16144
rect 1858 15680 1914 15736
rect 1950 15000 2006 15056
rect 1950 13232 2006 13288
rect 1858 12824 1914 12880
rect 1858 12416 1914 12472
rect 1950 10376 2006 10432
rect 1858 9560 1914 9616
rect 2778 27104 2834 27160
rect 3054 32000 3110 32056
rect 3238 30776 3294 30832
rect 3606 33260 3608 33280
rect 3608 33260 3660 33280
rect 3660 33260 3662 33280
rect 3606 33224 3662 33260
rect 3054 27920 3110 27976
rect 3054 24656 3110 24712
rect 2778 23840 2834 23896
rect 2778 23024 2834 23080
rect 3146 21392 3202 21448
rect 2778 20576 2834 20632
rect 3330 24248 3386 24304
rect 3422 18536 3478 18592
rect 2870 18128 2926 18184
rect 3238 17720 3294 17776
rect 2778 17312 2834 17368
rect 2502 15000 2558 15056
rect 2502 14612 2558 14648
rect 2502 14592 2504 14612
rect 2504 14592 2556 14612
rect 2556 14592 2558 14612
rect 2778 14048 2834 14104
rect 2410 11636 2412 11656
rect 2412 11636 2464 11656
rect 2464 11636 2466 11656
rect 2410 11600 2466 11636
rect 1950 7520 2006 7576
rect 2410 8372 2412 8392
rect 2412 8372 2464 8392
rect 2464 8372 2466 8392
rect 2410 8336 2466 8372
rect 3330 15272 3386 15328
rect 3422 14456 3478 14512
rect 3054 13640 3110 13696
rect 2778 12008 2834 12064
rect 2778 11212 2834 11248
rect 3790 40160 3846 40216
rect 4894 38392 4950 38448
rect 5814 52964 5870 53000
rect 5814 52944 5816 52964
rect 5816 52944 5868 52964
rect 5868 52944 5870 52964
rect 5588 52250 5644 52252
rect 5668 52250 5724 52252
rect 5748 52250 5804 52252
rect 5828 52250 5884 52252
rect 5588 52198 5614 52250
rect 5614 52198 5644 52250
rect 5668 52198 5678 52250
rect 5678 52198 5724 52250
rect 5748 52198 5794 52250
rect 5794 52198 5804 52250
rect 5828 52198 5858 52250
rect 5858 52198 5884 52250
rect 5588 52196 5644 52198
rect 5668 52196 5724 52198
rect 5748 52196 5804 52198
rect 5828 52196 5884 52198
rect 14852 53338 14908 53340
rect 14932 53338 14988 53340
rect 15012 53338 15068 53340
rect 15092 53338 15148 53340
rect 14852 53286 14878 53338
rect 14878 53286 14908 53338
rect 14932 53286 14942 53338
rect 14942 53286 14988 53338
rect 15012 53286 15058 53338
rect 15058 53286 15068 53338
rect 15092 53286 15122 53338
rect 15122 53286 15148 53338
rect 14852 53284 14908 53286
rect 14932 53284 14988 53286
rect 15012 53284 15068 53286
rect 15092 53284 15148 53286
rect 20258 54440 20314 54496
rect 5588 51162 5644 51164
rect 5668 51162 5724 51164
rect 5748 51162 5804 51164
rect 5828 51162 5884 51164
rect 5588 51110 5614 51162
rect 5614 51110 5644 51162
rect 5668 51110 5678 51162
rect 5678 51110 5724 51162
rect 5748 51110 5794 51162
rect 5794 51110 5804 51162
rect 5828 51110 5858 51162
rect 5858 51110 5884 51162
rect 5588 51108 5644 51110
rect 5668 51108 5724 51110
rect 5748 51108 5804 51110
rect 5828 51108 5884 51110
rect 5588 50074 5644 50076
rect 5668 50074 5724 50076
rect 5748 50074 5804 50076
rect 5828 50074 5884 50076
rect 5588 50022 5614 50074
rect 5614 50022 5644 50074
rect 5668 50022 5678 50074
rect 5678 50022 5724 50074
rect 5748 50022 5794 50074
rect 5794 50022 5804 50074
rect 5828 50022 5858 50074
rect 5858 50022 5884 50074
rect 5588 50020 5644 50022
rect 5668 50020 5724 50022
rect 5748 50020 5804 50022
rect 5828 50020 5884 50022
rect 5588 48986 5644 48988
rect 5668 48986 5724 48988
rect 5748 48986 5804 48988
rect 5828 48986 5884 48988
rect 5588 48934 5614 48986
rect 5614 48934 5644 48986
rect 5668 48934 5678 48986
rect 5678 48934 5724 48986
rect 5748 48934 5794 48986
rect 5794 48934 5804 48986
rect 5828 48934 5858 48986
rect 5858 48934 5884 48986
rect 5588 48932 5644 48934
rect 5668 48932 5724 48934
rect 5748 48932 5804 48934
rect 5828 48932 5884 48934
rect 5588 47898 5644 47900
rect 5668 47898 5724 47900
rect 5748 47898 5804 47900
rect 5828 47898 5884 47900
rect 5588 47846 5614 47898
rect 5614 47846 5644 47898
rect 5668 47846 5678 47898
rect 5678 47846 5724 47898
rect 5748 47846 5794 47898
rect 5794 47846 5804 47898
rect 5828 47846 5858 47898
rect 5858 47846 5884 47898
rect 5588 47844 5644 47846
rect 5668 47844 5724 47846
rect 5748 47844 5804 47846
rect 5828 47844 5884 47846
rect 5588 46810 5644 46812
rect 5668 46810 5724 46812
rect 5748 46810 5804 46812
rect 5828 46810 5884 46812
rect 5588 46758 5614 46810
rect 5614 46758 5644 46810
rect 5668 46758 5678 46810
rect 5678 46758 5724 46810
rect 5748 46758 5794 46810
rect 5794 46758 5804 46810
rect 5828 46758 5858 46810
rect 5858 46758 5884 46810
rect 5588 46756 5644 46758
rect 5668 46756 5724 46758
rect 5748 46756 5804 46758
rect 5828 46756 5884 46758
rect 5588 45722 5644 45724
rect 5668 45722 5724 45724
rect 5748 45722 5804 45724
rect 5828 45722 5884 45724
rect 5588 45670 5614 45722
rect 5614 45670 5644 45722
rect 5668 45670 5678 45722
rect 5678 45670 5724 45722
rect 5748 45670 5794 45722
rect 5794 45670 5804 45722
rect 5828 45670 5858 45722
rect 5858 45670 5884 45722
rect 5588 45668 5644 45670
rect 5668 45668 5724 45670
rect 5748 45668 5804 45670
rect 5828 45668 5884 45670
rect 5588 44634 5644 44636
rect 5668 44634 5724 44636
rect 5748 44634 5804 44636
rect 5828 44634 5884 44636
rect 5588 44582 5614 44634
rect 5614 44582 5644 44634
rect 5668 44582 5678 44634
rect 5678 44582 5724 44634
rect 5748 44582 5794 44634
rect 5794 44582 5804 44634
rect 5828 44582 5858 44634
rect 5858 44582 5884 44634
rect 5588 44580 5644 44582
rect 5668 44580 5724 44582
rect 5748 44580 5804 44582
rect 5828 44580 5884 44582
rect 5588 43546 5644 43548
rect 5668 43546 5724 43548
rect 5748 43546 5804 43548
rect 5828 43546 5884 43548
rect 5588 43494 5614 43546
rect 5614 43494 5644 43546
rect 5668 43494 5678 43546
rect 5678 43494 5724 43546
rect 5748 43494 5794 43546
rect 5794 43494 5804 43546
rect 5828 43494 5858 43546
rect 5858 43494 5884 43546
rect 5588 43492 5644 43494
rect 5668 43492 5724 43494
rect 5748 43492 5804 43494
rect 5828 43492 5884 43494
rect 5588 42458 5644 42460
rect 5668 42458 5724 42460
rect 5748 42458 5804 42460
rect 5828 42458 5884 42460
rect 5588 42406 5614 42458
rect 5614 42406 5644 42458
rect 5668 42406 5678 42458
rect 5678 42406 5724 42458
rect 5748 42406 5794 42458
rect 5794 42406 5804 42458
rect 5828 42406 5858 42458
rect 5858 42406 5884 42458
rect 5588 42404 5644 42406
rect 5668 42404 5724 42406
rect 5748 42404 5804 42406
rect 5828 42404 5884 42406
rect 5588 41370 5644 41372
rect 5668 41370 5724 41372
rect 5748 41370 5804 41372
rect 5828 41370 5884 41372
rect 5588 41318 5614 41370
rect 5614 41318 5644 41370
rect 5668 41318 5678 41370
rect 5678 41318 5724 41370
rect 5748 41318 5794 41370
rect 5794 41318 5804 41370
rect 5828 41318 5858 41370
rect 5858 41318 5884 41370
rect 5588 41316 5644 41318
rect 5668 41316 5724 41318
rect 5748 41316 5804 41318
rect 5828 41316 5884 41318
rect 5538 41112 5594 41168
rect 4158 32816 4214 32872
rect 3790 31184 3846 31240
rect 3790 28328 3846 28384
rect 4066 31592 4122 31648
rect 4526 34584 4582 34640
rect 3974 28908 3976 28928
rect 3976 28908 4028 28928
rect 4028 28908 4030 28928
rect 3974 28872 4030 28908
rect 4066 25064 4122 25120
rect 4250 22344 4306 22400
rect 4526 21800 4582 21856
rect 4066 14864 4122 14920
rect 2778 11192 2780 11212
rect 2780 11192 2832 11212
rect 2832 11192 2834 11212
rect 2410 7948 2466 7984
rect 2410 7928 2412 7948
rect 2412 7928 2464 7948
rect 2464 7928 2466 7948
rect 2870 9152 2926 9208
rect 3238 8744 3294 8800
rect 3054 7112 3110 7168
rect 2778 3848 2834 3904
rect 1950 3440 2006 3496
rect 1674 3032 1730 3088
rect 2778 1400 2834 1456
rect 1398 176 1454 232
rect 3238 992 3294 1048
rect 3698 5908 3754 5944
rect 3698 5888 3700 5908
rect 3700 5888 3752 5908
rect 3752 5888 3754 5908
rect 4066 6296 4122 6352
rect 3974 5480 4030 5536
rect 4066 5072 4122 5128
rect 4066 4664 4122 4720
rect 3974 4256 4030 4312
rect 3514 2624 3570 2680
rect 5588 40282 5644 40284
rect 5668 40282 5724 40284
rect 5748 40282 5804 40284
rect 5828 40282 5884 40284
rect 5588 40230 5614 40282
rect 5614 40230 5644 40282
rect 5668 40230 5678 40282
rect 5678 40230 5724 40282
rect 5748 40230 5794 40282
rect 5794 40230 5804 40282
rect 5828 40230 5858 40282
rect 5858 40230 5884 40282
rect 5588 40228 5644 40230
rect 5668 40228 5724 40230
rect 5748 40228 5804 40230
rect 5828 40228 5884 40230
rect 5588 39194 5644 39196
rect 5668 39194 5724 39196
rect 5748 39194 5804 39196
rect 5828 39194 5884 39196
rect 5588 39142 5614 39194
rect 5614 39142 5644 39194
rect 5668 39142 5678 39194
rect 5678 39142 5724 39194
rect 5748 39142 5794 39194
rect 5794 39142 5804 39194
rect 5828 39142 5858 39194
rect 5858 39142 5884 39194
rect 5588 39140 5644 39142
rect 5668 39140 5724 39142
rect 5748 39140 5804 39142
rect 5828 39140 5884 39142
rect 5588 38106 5644 38108
rect 5668 38106 5724 38108
rect 5748 38106 5804 38108
rect 5828 38106 5884 38108
rect 5588 38054 5614 38106
rect 5614 38054 5644 38106
rect 5668 38054 5678 38106
rect 5678 38054 5724 38106
rect 5748 38054 5794 38106
rect 5794 38054 5804 38106
rect 5828 38054 5858 38106
rect 5858 38054 5884 38106
rect 5588 38052 5644 38054
rect 5668 38052 5724 38054
rect 5748 38052 5804 38054
rect 5828 38052 5884 38054
rect 5588 37018 5644 37020
rect 5668 37018 5724 37020
rect 5748 37018 5804 37020
rect 5828 37018 5884 37020
rect 5588 36966 5614 37018
rect 5614 36966 5644 37018
rect 5668 36966 5678 37018
rect 5678 36966 5724 37018
rect 5748 36966 5794 37018
rect 5794 36966 5804 37018
rect 5828 36966 5858 37018
rect 5858 36966 5884 37018
rect 5588 36964 5644 36966
rect 5668 36964 5724 36966
rect 5748 36964 5804 36966
rect 5828 36964 5884 36966
rect 5588 35930 5644 35932
rect 5668 35930 5724 35932
rect 5748 35930 5804 35932
rect 5828 35930 5884 35932
rect 5588 35878 5614 35930
rect 5614 35878 5644 35930
rect 5668 35878 5678 35930
rect 5678 35878 5724 35930
rect 5748 35878 5794 35930
rect 5794 35878 5804 35930
rect 5828 35878 5858 35930
rect 5858 35878 5884 35930
rect 5588 35876 5644 35878
rect 5668 35876 5724 35878
rect 5748 35876 5804 35878
rect 5828 35876 5884 35878
rect 5588 34842 5644 34844
rect 5668 34842 5724 34844
rect 5748 34842 5804 34844
rect 5828 34842 5884 34844
rect 5588 34790 5614 34842
rect 5614 34790 5644 34842
rect 5668 34790 5678 34842
rect 5678 34790 5724 34842
rect 5748 34790 5794 34842
rect 5794 34790 5804 34842
rect 5828 34790 5858 34842
rect 5858 34790 5884 34842
rect 5588 34788 5644 34790
rect 5668 34788 5724 34790
rect 5748 34788 5804 34790
rect 5828 34788 5884 34790
rect 5538 34604 5594 34640
rect 5538 34584 5540 34604
rect 5540 34584 5592 34604
rect 5592 34584 5594 34604
rect 5588 33754 5644 33756
rect 5668 33754 5724 33756
rect 5748 33754 5804 33756
rect 5828 33754 5884 33756
rect 5588 33702 5614 33754
rect 5614 33702 5644 33754
rect 5668 33702 5678 33754
rect 5678 33702 5724 33754
rect 5748 33702 5794 33754
rect 5794 33702 5804 33754
rect 5828 33702 5858 33754
rect 5858 33702 5884 33754
rect 5588 33700 5644 33702
rect 5668 33700 5724 33702
rect 5748 33700 5804 33702
rect 5828 33700 5884 33702
rect 5588 32666 5644 32668
rect 5668 32666 5724 32668
rect 5748 32666 5804 32668
rect 5828 32666 5884 32668
rect 5588 32614 5614 32666
rect 5614 32614 5644 32666
rect 5668 32614 5678 32666
rect 5678 32614 5724 32666
rect 5748 32614 5794 32666
rect 5794 32614 5804 32666
rect 5828 32614 5858 32666
rect 5858 32614 5884 32666
rect 5588 32612 5644 32614
rect 5668 32612 5724 32614
rect 5748 32612 5804 32614
rect 5828 32612 5884 32614
rect 5588 31578 5644 31580
rect 5668 31578 5724 31580
rect 5748 31578 5804 31580
rect 5828 31578 5884 31580
rect 5588 31526 5614 31578
rect 5614 31526 5644 31578
rect 5668 31526 5678 31578
rect 5678 31526 5724 31578
rect 5748 31526 5794 31578
rect 5794 31526 5804 31578
rect 5828 31526 5858 31578
rect 5858 31526 5884 31578
rect 5588 31524 5644 31526
rect 5668 31524 5724 31526
rect 5748 31524 5804 31526
rect 5828 31524 5884 31526
rect 5588 30490 5644 30492
rect 5668 30490 5724 30492
rect 5748 30490 5804 30492
rect 5828 30490 5884 30492
rect 5588 30438 5614 30490
rect 5614 30438 5644 30490
rect 5668 30438 5678 30490
rect 5678 30438 5724 30490
rect 5748 30438 5794 30490
rect 5794 30438 5804 30490
rect 5828 30438 5858 30490
rect 5858 30438 5884 30490
rect 5588 30436 5644 30438
rect 5668 30436 5724 30438
rect 5748 30436 5804 30438
rect 5828 30436 5884 30438
rect 5446 29824 5502 29880
rect 6182 38392 6238 38448
rect 5722 29824 5778 29880
rect 5588 29402 5644 29404
rect 5668 29402 5724 29404
rect 5748 29402 5804 29404
rect 5828 29402 5884 29404
rect 5588 29350 5614 29402
rect 5614 29350 5644 29402
rect 5668 29350 5678 29402
rect 5678 29350 5724 29402
rect 5748 29350 5794 29402
rect 5794 29350 5804 29402
rect 5828 29350 5858 29402
rect 5858 29350 5884 29402
rect 5588 29348 5644 29350
rect 5668 29348 5724 29350
rect 5748 29348 5804 29350
rect 5828 29348 5884 29350
rect 5588 28314 5644 28316
rect 5668 28314 5724 28316
rect 5748 28314 5804 28316
rect 5828 28314 5884 28316
rect 5588 28262 5614 28314
rect 5614 28262 5644 28314
rect 5668 28262 5678 28314
rect 5678 28262 5724 28314
rect 5748 28262 5794 28314
rect 5794 28262 5804 28314
rect 5828 28262 5858 28314
rect 5858 28262 5884 28314
rect 5588 28260 5644 28262
rect 5668 28260 5724 28262
rect 5748 28260 5804 28262
rect 5828 28260 5884 28262
rect 5588 27226 5644 27228
rect 5668 27226 5724 27228
rect 5748 27226 5804 27228
rect 5828 27226 5884 27228
rect 5588 27174 5614 27226
rect 5614 27174 5644 27226
rect 5668 27174 5678 27226
rect 5678 27174 5724 27226
rect 5748 27174 5794 27226
rect 5794 27174 5804 27226
rect 5828 27174 5858 27226
rect 5858 27174 5884 27226
rect 5588 27172 5644 27174
rect 5668 27172 5724 27174
rect 5748 27172 5804 27174
rect 5828 27172 5884 27174
rect 5588 26138 5644 26140
rect 5668 26138 5724 26140
rect 5748 26138 5804 26140
rect 5828 26138 5884 26140
rect 5588 26086 5614 26138
rect 5614 26086 5644 26138
rect 5668 26086 5678 26138
rect 5678 26086 5724 26138
rect 5748 26086 5794 26138
rect 5794 26086 5804 26138
rect 5828 26086 5858 26138
rect 5858 26086 5884 26138
rect 5588 26084 5644 26086
rect 5668 26084 5724 26086
rect 5748 26084 5804 26086
rect 5828 26084 5884 26086
rect 5262 22344 5318 22400
rect 5078 21936 5134 21992
rect 4986 18808 5042 18864
rect 5170 15000 5226 15056
rect 5588 25050 5644 25052
rect 5668 25050 5724 25052
rect 5748 25050 5804 25052
rect 5828 25050 5884 25052
rect 5588 24998 5614 25050
rect 5614 24998 5644 25050
rect 5668 24998 5678 25050
rect 5678 24998 5724 25050
rect 5748 24998 5794 25050
rect 5794 24998 5804 25050
rect 5828 24998 5858 25050
rect 5858 24998 5884 25050
rect 5588 24996 5644 24998
rect 5668 24996 5724 24998
rect 5748 24996 5804 24998
rect 5828 24996 5884 24998
rect 5588 23962 5644 23964
rect 5668 23962 5724 23964
rect 5748 23962 5804 23964
rect 5828 23962 5884 23964
rect 5588 23910 5614 23962
rect 5614 23910 5644 23962
rect 5668 23910 5678 23962
rect 5678 23910 5724 23962
rect 5748 23910 5794 23962
rect 5794 23910 5804 23962
rect 5828 23910 5858 23962
rect 5858 23910 5884 23962
rect 5588 23908 5644 23910
rect 5668 23908 5724 23910
rect 5748 23908 5804 23910
rect 5828 23908 5884 23910
rect 5588 22874 5644 22876
rect 5668 22874 5724 22876
rect 5748 22874 5804 22876
rect 5828 22874 5884 22876
rect 5588 22822 5614 22874
rect 5614 22822 5644 22874
rect 5668 22822 5678 22874
rect 5678 22822 5724 22874
rect 5748 22822 5794 22874
rect 5794 22822 5804 22874
rect 5828 22822 5858 22874
rect 5858 22822 5884 22874
rect 5588 22820 5644 22822
rect 5668 22820 5724 22822
rect 5748 22820 5804 22822
rect 5828 22820 5884 22822
rect 5538 21972 5540 21992
rect 5540 21972 5592 21992
rect 5592 21972 5594 21992
rect 5538 21936 5594 21972
rect 5588 21786 5644 21788
rect 5668 21786 5724 21788
rect 5748 21786 5804 21788
rect 5828 21786 5884 21788
rect 5588 21734 5614 21786
rect 5614 21734 5644 21786
rect 5668 21734 5678 21786
rect 5678 21734 5724 21786
rect 5748 21734 5794 21786
rect 5794 21734 5804 21786
rect 5828 21734 5858 21786
rect 5858 21734 5884 21786
rect 5588 21732 5644 21734
rect 5668 21732 5724 21734
rect 5748 21732 5804 21734
rect 5828 21732 5884 21734
rect 5588 20698 5644 20700
rect 5668 20698 5724 20700
rect 5748 20698 5804 20700
rect 5828 20698 5884 20700
rect 5588 20646 5614 20698
rect 5614 20646 5644 20698
rect 5668 20646 5678 20698
rect 5678 20646 5724 20698
rect 5748 20646 5794 20698
rect 5794 20646 5804 20698
rect 5828 20646 5858 20698
rect 5858 20646 5884 20698
rect 5588 20644 5644 20646
rect 5668 20644 5724 20646
rect 5748 20644 5804 20646
rect 5828 20644 5884 20646
rect 5588 19610 5644 19612
rect 5668 19610 5724 19612
rect 5748 19610 5804 19612
rect 5828 19610 5884 19612
rect 5588 19558 5614 19610
rect 5614 19558 5644 19610
rect 5668 19558 5678 19610
rect 5678 19558 5724 19610
rect 5748 19558 5794 19610
rect 5794 19558 5804 19610
rect 5828 19558 5858 19610
rect 5858 19558 5884 19610
rect 5588 19556 5644 19558
rect 5668 19556 5724 19558
rect 5748 19556 5804 19558
rect 5828 19556 5884 19558
rect 5538 18808 5594 18864
rect 5588 18522 5644 18524
rect 5668 18522 5724 18524
rect 5748 18522 5804 18524
rect 5828 18522 5884 18524
rect 5588 18470 5614 18522
rect 5614 18470 5644 18522
rect 5668 18470 5678 18522
rect 5678 18470 5724 18522
rect 5748 18470 5794 18522
rect 5794 18470 5804 18522
rect 5828 18470 5858 18522
rect 5858 18470 5884 18522
rect 5588 18468 5644 18470
rect 5668 18468 5724 18470
rect 5748 18468 5804 18470
rect 5828 18468 5884 18470
rect 5588 17434 5644 17436
rect 5668 17434 5724 17436
rect 5748 17434 5804 17436
rect 5828 17434 5884 17436
rect 5588 17382 5614 17434
rect 5614 17382 5644 17434
rect 5668 17382 5678 17434
rect 5678 17382 5724 17434
rect 5748 17382 5794 17434
rect 5794 17382 5804 17434
rect 5828 17382 5858 17434
rect 5858 17382 5884 17434
rect 5588 17380 5644 17382
rect 5668 17380 5724 17382
rect 5748 17380 5804 17382
rect 5828 17380 5884 17382
rect 5588 16346 5644 16348
rect 5668 16346 5724 16348
rect 5748 16346 5804 16348
rect 5828 16346 5884 16348
rect 5588 16294 5614 16346
rect 5614 16294 5644 16346
rect 5668 16294 5678 16346
rect 5678 16294 5724 16346
rect 5748 16294 5794 16346
rect 5794 16294 5804 16346
rect 5828 16294 5858 16346
rect 5858 16294 5884 16346
rect 5588 16292 5644 16294
rect 5668 16292 5724 16294
rect 5748 16292 5804 16294
rect 5828 16292 5884 16294
rect 5588 15258 5644 15260
rect 5668 15258 5724 15260
rect 5748 15258 5804 15260
rect 5828 15258 5884 15260
rect 5588 15206 5614 15258
rect 5614 15206 5644 15258
rect 5668 15206 5678 15258
rect 5678 15206 5724 15258
rect 5748 15206 5794 15258
rect 5794 15206 5804 15258
rect 5828 15206 5858 15258
rect 5858 15206 5884 15258
rect 5588 15204 5644 15206
rect 5668 15204 5724 15206
rect 5748 15204 5804 15206
rect 5828 15204 5884 15206
rect 5588 14170 5644 14172
rect 5668 14170 5724 14172
rect 5748 14170 5804 14172
rect 5828 14170 5884 14172
rect 5588 14118 5614 14170
rect 5614 14118 5644 14170
rect 5668 14118 5678 14170
rect 5678 14118 5724 14170
rect 5748 14118 5794 14170
rect 5794 14118 5804 14170
rect 5828 14118 5858 14170
rect 5858 14118 5884 14170
rect 5588 14116 5644 14118
rect 5668 14116 5724 14118
rect 5748 14116 5804 14118
rect 5828 14116 5884 14118
rect 5588 13082 5644 13084
rect 5668 13082 5724 13084
rect 5748 13082 5804 13084
rect 5828 13082 5884 13084
rect 5588 13030 5614 13082
rect 5614 13030 5644 13082
rect 5668 13030 5678 13082
rect 5678 13030 5724 13082
rect 5748 13030 5794 13082
rect 5794 13030 5804 13082
rect 5828 13030 5858 13082
rect 5858 13030 5884 13082
rect 5588 13028 5644 13030
rect 5668 13028 5724 13030
rect 5748 13028 5804 13030
rect 5828 13028 5884 13030
rect 5588 11994 5644 11996
rect 5668 11994 5724 11996
rect 5748 11994 5804 11996
rect 5828 11994 5884 11996
rect 5588 11942 5614 11994
rect 5614 11942 5644 11994
rect 5668 11942 5678 11994
rect 5678 11942 5724 11994
rect 5748 11942 5794 11994
rect 5794 11942 5804 11994
rect 5828 11942 5858 11994
rect 5858 11942 5884 11994
rect 5588 11940 5644 11942
rect 5668 11940 5724 11942
rect 5748 11940 5804 11942
rect 5828 11940 5884 11942
rect 5588 10906 5644 10908
rect 5668 10906 5724 10908
rect 5748 10906 5804 10908
rect 5828 10906 5884 10908
rect 5588 10854 5614 10906
rect 5614 10854 5644 10906
rect 5668 10854 5678 10906
rect 5678 10854 5724 10906
rect 5748 10854 5794 10906
rect 5794 10854 5804 10906
rect 5828 10854 5858 10906
rect 5858 10854 5884 10906
rect 5588 10852 5644 10854
rect 5668 10852 5724 10854
rect 5748 10852 5804 10854
rect 5828 10852 5884 10854
rect 5588 9818 5644 9820
rect 5668 9818 5724 9820
rect 5748 9818 5804 9820
rect 5828 9818 5884 9820
rect 5588 9766 5614 9818
rect 5614 9766 5644 9818
rect 5668 9766 5678 9818
rect 5678 9766 5724 9818
rect 5748 9766 5794 9818
rect 5794 9766 5804 9818
rect 5828 9766 5858 9818
rect 5858 9766 5884 9818
rect 5588 9764 5644 9766
rect 5668 9764 5724 9766
rect 5748 9764 5804 9766
rect 5828 9764 5884 9766
rect 5588 8730 5644 8732
rect 5668 8730 5724 8732
rect 5748 8730 5804 8732
rect 5828 8730 5884 8732
rect 5588 8678 5614 8730
rect 5614 8678 5644 8730
rect 5668 8678 5678 8730
rect 5678 8678 5724 8730
rect 5748 8678 5794 8730
rect 5794 8678 5804 8730
rect 5828 8678 5858 8730
rect 5858 8678 5884 8730
rect 5588 8676 5644 8678
rect 5668 8676 5724 8678
rect 5748 8676 5804 8678
rect 5828 8676 5884 8678
rect 3422 2216 3478 2272
rect 3422 1844 3424 1864
rect 3424 1844 3476 1864
rect 3476 1844 3478 1864
rect 3422 1808 3478 1844
rect 5588 7642 5644 7644
rect 5668 7642 5724 7644
rect 5748 7642 5804 7644
rect 5828 7642 5884 7644
rect 5588 7590 5614 7642
rect 5614 7590 5644 7642
rect 5668 7590 5678 7642
rect 5678 7590 5724 7642
rect 5748 7590 5794 7642
rect 5794 7590 5804 7642
rect 5828 7590 5858 7642
rect 5858 7590 5884 7642
rect 5588 7588 5644 7590
rect 5668 7588 5724 7590
rect 5748 7588 5804 7590
rect 5828 7588 5884 7590
rect 5588 6554 5644 6556
rect 5668 6554 5724 6556
rect 5748 6554 5804 6556
rect 5828 6554 5884 6556
rect 5588 6502 5614 6554
rect 5614 6502 5644 6554
rect 5668 6502 5678 6554
rect 5678 6502 5724 6554
rect 5748 6502 5794 6554
rect 5794 6502 5804 6554
rect 5828 6502 5858 6554
rect 5858 6502 5884 6554
rect 5588 6500 5644 6502
rect 5668 6500 5724 6502
rect 5748 6500 5804 6502
rect 5828 6500 5884 6502
rect 5588 5466 5644 5468
rect 5668 5466 5724 5468
rect 5748 5466 5804 5468
rect 5828 5466 5884 5468
rect 5588 5414 5614 5466
rect 5614 5414 5644 5466
rect 5668 5414 5678 5466
rect 5678 5414 5724 5466
rect 5748 5414 5794 5466
rect 5794 5414 5804 5466
rect 5828 5414 5858 5466
rect 5858 5414 5884 5466
rect 5588 5412 5644 5414
rect 5668 5412 5724 5414
rect 5748 5412 5804 5414
rect 5828 5412 5884 5414
rect 5588 4378 5644 4380
rect 5668 4378 5724 4380
rect 5748 4378 5804 4380
rect 5828 4378 5884 4380
rect 5588 4326 5614 4378
rect 5614 4326 5644 4378
rect 5668 4326 5678 4378
rect 5678 4326 5724 4378
rect 5748 4326 5794 4378
rect 5794 4326 5804 4378
rect 5828 4326 5858 4378
rect 5858 4326 5884 4378
rect 5588 4324 5644 4326
rect 5668 4324 5724 4326
rect 5748 4324 5804 4326
rect 5828 4324 5884 4326
rect 5588 3290 5644 3292
rect 5668 3290 5724 3292
rect 5748 3290 5804 3292
rect 5828 3290 5884 3292
rect 5588 3238 5614 3290
rect 5614 3238 5644 3290
rect 5668 3238 5678 3290
rect 5678 3238 5724 3290
rect 5748 3238 5794 3290
rect 5794 3238 5804 3290
rect 5828 3238 5858 3290
rect 5858 3238 5884 3290
rect 5588 3236 5644 3238
rect 5668 3236 5724 3238
rect 5748 3236 5804 3238
rect 5828 3236 5884 3238
rect 5588 2202 5644 2204
rect 5668 2202 5724 2204
rect 5748 2202 5804 2204
rect 5828 2202 5884 2204
rect 5588 2150 5614 2202
rect 5614 2150 5644 2202
rect 5668 2150 5678 2202
rect 5678 2150 5724 2202
rect 5748 2150 5794 2202
rect 5794 2150 5804 2202
rect 5828 2150 5858 2202
rect 5858 2150 5884 2202
rect 5588 2148 5644 2150
rect 5668 2148 5724 2150
rect 5748 2148 5804 2150
rect 5828 2148 5884 2150
rect 7378 28076 7434 28112
rect 7378 28056 7380 28076
rect 7380 28056 7432 28076
rect 7432 28056 7434 28076
rect 7378 14592 7434 14648
rect 9218 41132 9274 41168
rect 9218 41112 9220 41132
rect 9220 41112 9272 41132
rect 9272 41112 9274 41132
rect 9218 38120 9274 38176
rect 10220 52794 10276 52796
rect 10300 52794 10356 52796
rect 10380 52794 10436 52796
rect 10460 52794 10516 52796
rect 10220 52742 10246 52794
rect 10246 52742 10276 52794
rect 10300 52742 10310 52794
rect 10310 52742 10356 52794
rect 10380 52742 10426 52794
rect 10426 52742 10436 52794
rect 10460 52742 10490 52794
rect 10490 52742 10516 52794
rect 10220 52740 10276 52742
rect 10300 52740 10356 52742
rect 10380 52740 10436 52742
rect 10460 52740 10516 52742
rect 10220 51706 10276 51708
rect 10300 51706 10356 51708
rect 10380 51706 10436 51708
rect 10460 51706 10516 51708
rect 10220 51654 10246 51706
rect 10246 51654 10276 51706
rect 10300 51654 10310 51706
rect 10310 51654 10356 51706
rect 10380 51654 10426 51706
rect 10426 51654 10436 51706
rect 10460 51654 10490 51706
rect 10490 51654 10516 51706
rect 10220 51652 10276 51654
rect 10300 51652 10356 51654
rect 10380 51652 10436 51654
rect 10460 51652 10516 51654
rect 10782 51312 10838 51368
rect 10220 50618 10276 50620
rect 10300 50618 10356 50620
rect 10380 50618 10436 50620
rect 10460 50618 10516 50620
rect 10220 50566 10246 50618
rect 10246 50566 10276 50618
rect 10300 50566 10310 50618
rect 10310 50566 10356 50618
rect 10380 50566 10426 50618
rect 10426 50566 10436 50618
rect 10460 50566 10490 50618
rect 10490 50566 10516 50618
rect 10220 50564 10276 50566
rect 10300 50564 10356 50566
rect 10380 50564 10436 50566
rect 10460 50564 10516 50566
rect 10220 49530 10276 49532
rect 10300 49530 10356 49532
rect 10380 49530 10436 49532
rect 10460 49530 10516 49532
rect 10220 49478 10246 49530
rect 10246 49478 10276 49530
rect 10300 49478 10310 49530
rect 10310 49478 10356 49530
rect 10380 49478 10426 49530
rect 10426 49478 10436 49530
rect 10460 49478 10490 49530
rect 10490 49478 10516 49530
rect 10220 49476 10276 49478
rect 10300 49476 10356 49478
rect 10380 49476 10436 49478
rect 10460 49476 10516 49478
rect 10220 48442 10276 48444
rect 10300 48442 10356 48444
rect 10380 48442 10436 48444
rect 10460 48442 10516 48444
rect 10220 48390 10246 48442
rect 10246 48390 10276 48442
rect 10300 48390 10310 48442
rect 10310 48390 10356 48442
rect 10380 48390 10426 48442
rect 10426 48390 10436 48442
rect 10460 48390 10490 48442
rect 10490 48390 10516 48442
rect 10220 48388 10276 48390
rect 10300 48388 10356 48390
rect 10380 48388 10436 48390
rect 10460 48388 10516 48390
rect 10220 47354 10276 47356
rect 10300 47354 10356 47356
rect 10380 47354 10436 47356
rect 10460 47354 10516 47356
rect 10220 47302 10246 47354
rect 10246 47302 10276 47354
rect 10300 47302 10310 47354
rect 10310 47302 10356 47354
rect 10380 47302 10426 47354
rect 10426 47302 10436 47354
rect 10460 47302 10490 47354
rect 10490 47302 10516 47354
rect 10220 47300 10276 47302
rect 10300 47300 10356 47302
rect 10380 47300 10436 47302
rect 10460 47300 10516 47302
rect 10220 46266 10276 46268
rect 10300 46266 10356 46268
rect 10380 46266 10436 46268
rect 10460 46266 10516 46268
rect 10220 46214 10246 46266
rect 10246 46214 10276 46266
rect 10300 46214 10310 46266
rect 10310 46214 10356 46266
rect 10380 46214 10426 46266
rect 10426 46214 10436 46266
rect 10460 46214 10490 46266
rect 10490 46214 10516 46266
rect 10220 46212 10276 46214
rect 10300 46212 10356 46214
rect 10380 46212 10436 46214
rect 10460 46212 10516 46214
rect 10220 45178 10276 45180
rect 10300 45178 10356 45180
rect 10380 45178 10436 45180
rect 10460 45178 10516 45180
rect 10220 45126 10246 45178
rect 10246 45126 10276 45178
rect 10300 45126 10310 45178
rect 10310 45126 10356 45178
rect 10380 45126 10426 45178
rect 10426 45126 10436 45178
rect 10460 45126 10490 45178
rect 10490 45126 10516 45178
rect 10220 45124 10276 45126
rect 10300 45124 10356 45126
rect 10380 45124 10436 45126
rect 10460 45124 10516 45126
rect 10220 44090 10276 44092
rect 10300 44090 10356 44092
rect 10380 44090 10436 44092
rect 10460 44090 10516 44092
rect 10220 44038 10246 44090
rect 10246 44038 10276 44090
rect 10300 44038 10310 44090
rect 10310 44038 10356 44090
rect 10380 44038 10426 44090
rect 10426 44038 10436 44090
rect 10460 44038 10490 44090
rect 10490 44038 10516 44090
rect 10220 44036 10276 44038
rect 10300 44036 10356 44038
rect 10380 44036 10436 44038
rect 10460 44036 10516 44038
rect 9402 38292 9404 38312
rect 9404 38292 9456 38312
rect 9456 38292 9458 38312
rect 9402 38256 9458 38292
rect 10220 43002 10276 43004
rect 10300 43002 10356 43004
rect 10380 43002 10436 43004
rect 10460 43002 10516 43004
rect 10220 42950 10246 43002
rect 10246 42950 10276 43002
rect 10300 42950 10310 43002
rect 10310 42950 10356 43002
rect 10380 42950 10426 43002
rect 10426 42950 10436 43002
rect 10460 42950 10490 43002
rect 10490 42950 10516 43002
rect 10220 42948 10276 42950
rect 10300 42948 10356 42950
rect 10380 42948 10436 42950
rect 10460 42948 10516 42950
rect 10220 41914 10276 41916
rect 10300 41914 10356 41916
rect 10380 41914 10436 41916
rect 10460 41914 10516 41916
rect 10220 41862 10246 41914
rect 10246 41862 10276 41914
rect 10300 41862 10310 41914
rect 10310 41862 10356 41914
rect 10380 41862 10426 41914
rect 10426 41862 10436 41914
rect 10460 41862 10490 41914
rect 10490 41862 10516 41914
rect 10220 41860 10276 41862
rect 10300 41860 10356 41862
rect 10380 41860 10436 41862
rect 10460 41860 10516 41862
rect 9954 26288 10010 26344
rect 10220 40826 10276 40828
rect 10300 40826 10356 40828
rect 10380 40826 10436 40828
rect 10460 40826 10516 40828
rect 10220 40774 10246 40826
rect 10246 40774 10276 40826
rect 10300 40774 10310 40826
rect 10310 40774 10356 40826
rect 10380 40774 10426 40826
rect 10426 40774 10436 40826
rect 10460 40774 10490 40826
rect 10490 40774 10516 40826
rect 10220 40772 10276 40774
rect 10300 40772 10356 40774
rect 10380 40772 10436 40774
rect 10460 40772 10516 40774
rect 10220 39738 10276 39740
rect 10300 39738 10356 39740
rect 10380 39738 10436 39740
rect 10460 39738 10516 39740
rect 10220 39686 10246 39738
rect 10246 39686 10276 39738
rect 10300 39686 10310 39738
rect 10310 39686 10356 39738
rect 10380 39686 10426 39738
rect 10426 39686 10436 39738
rect 10460 39686 10490 39738
rect 10490 39686 10516 39738
rect 10220 39684 10276 39686
rect 10300 39684 10356 39686
rect 10380 39684 10436 39686
rect 10460 39684 10516 39686
rect 10230 39516 10232 39536
rect 10232 39516 10284 39536
rect 10284 39516 10286 39536
rect 10230 39480 10286 39516
rect 10506 39344 10562 39400
rect 10506 38936 10562 38992
rect 10322 38800 10378 38856
rect 10220 38650 10276 38652
rect 10300 38650 10356 38652
rect 10380 38650 10436 38652
rect 10460 38650 10516 38652
rect 10220 38598 10246 38650
rect 10246 38598 10276 38650
rect 10300 38598 10310 38650
rect 10310 38598 10356 38650
rect 10380 38598 10426 38650
rect 10426 38598 10436 38650
rect 10460 38598 10490 38650
rect 10490 38598 10516 38650
rect 10220 38596 10276 38598
rect 10300 38596 10356 38598
rect 10380 38596 10436 38598
rect 10460 38596 10516 38598
rect 10230 38392 10286 38448
rect 10506 38256 10562 38312
rect 10220 37562 10276 37564
rect 10300 37562 10356 37564
rect 10380 37562 10436 37564
rect 10460 37562 10516 37564
rect 10220 37510 10246 37562
rect 10246 37510 10276 37562
rect 10300 37510 10310 37562
rect 10310 37510 10356 37562
rect 10380 37510 10426 37562
rect 10426 37510 10436 37562
rect 10460 37510 10490 37562
rect 10490 37510 10516 37562
rect 10220 37508 10276 37510
rect 10300 37508 10356 37510
rect 10380 37508 10436 37510
rect 10460 37508 10516 37510
rect 10220 36474 10276 36476
rect 10300 36474 10356 36476
rect 10380 36474 10436 36476
rect 10460 36474 10516 36476
rect 10220 36422 10246 36474
rect 10246 36422 10276 36474
rect 10300 36422 10310 36474
rect 10310 36422 10356 36474
rect 10380 36422 10426 36474
rect 10426 36422 10436 36474
rect 10460 36422 10490 36474
rect 10490 36422 10516 36474
rect 10220 36420 10276 36422
rect 10300 36420 10356 36422
rect 10380 36420 10436 36422
rect 10460 36420 10516 36422
rect 10220 35386 10276 35388
rect 10300 35386 10356 35388
rect 10380 35386 10436 35388
rect 10460 35386 10516 35388
rect 10220 35334 10246 35386
rect 10246 35334 10276 35386
rect 10300 35334 10310 35386
rect 10310 35334 10356 35386
rect 10380 35334 10426 35386
rect 10426 35334 10436 35386
rect 10460 35334 10490 35386
rect 10490 35334 10516 35386
rect 10220 35332 10276 35334
rect 10300 35332 10356 35334
rect 10380 35332 10436 35334
rect 10460 35332 10516 35334
rect 10414 35028 10416 35048
rect 10416 35028 10468 35048
rect 10468 35028 10470 35048
rect 10414 34992 10470 35028
rect 10322 34448 10378 34504
rect 10220 34298 10276 34300
rect 10300 34298 10356 34300
rect 10380 34298 10436 34300
rect 10460 34298 10516 34300
rect 10220 34246 10246 34298
rect 10246 34246 10276 34298
rect 10300 34246 10310 34298
rect 10310 34246 10356 34298
rect 10380 34246 10426 34298
rect 10426 34246 10436 34298
rect 10460 34246 10490 34298
rect 10490 34246 10516 34298
rect 10220 34244 10276 34246
rect 10300 34244 10356 34246
rect 10380 34244 10436 34246
rect 10460 34244 10516 34246
rect 10220 33210 10276 33212
rect 10300 33210 10356 33212
rect 10380 33210 10436 33212
rect 10460 33210 10516 33212
rect 10220 33158 10246 33210
rect 10246 33158 10276 33210
rect 10300 33158 10310 33210
rect 10310 33158 10356 33210
rect 10380 33158 10426 33210
rect 10426 33158 10436 33210
rect 10460 33158 10490 33210
rect 10490 33158 10516 33210
rect 10220 33156 10276 33158
rect 10300 33156 10356 33158
rect 10380 33156 10436 33158
rect 10460 33156 10516 33158
rect 10220 32122 10276 32124
rect 10300 32122 10356 32124
rect 10380 32122 10436 32124
rect 10460 32122 10516 32124
rect 10220 32070 10246 32122
rect 10246 32070 10276 32122
rect 10300 32070 10310 32122
rect 10310 32070 10356 32122
rect 10380 32070 10426 32122
rect 10426 32070 10436 32122
rect 10460 32070 10490 32122
rect 10490 32070 10516 32122
rect 10220 32068 10276 32070
rect 10300 32068 10356 32070
rect 10380 32068 10436 32070
rect 10460 32068 10516 32070
rect 10220 31034 10276 31036
rect 10300 31034 10356 31036
rect 10380 31034 10436 31036
rect 10460 31034 10516 31036
rect 10220 30982 10246 31034
rect 10246 30982 10276 31034
rect 10300 30982 10310 31034
rect 10310 30982 10356 31034
rect 10380 30982 10426 31034
rect 10426 30982 10436 31034
rect 10460 30982 10490 31034
rect 10490 30982 10516 31034
rect 10220 30980 10276 30982
rect 10300 30980 10356 30982
rect 10380 30980 10436 30982
rect 10460 30980 10516 30982
rect 10220 29946 10276 29948
rect 10300 29946 10356 29948
rect 10380 29946 10436 29948
rect 10460 29946 10516 29948
rect 10220 29894 10246 29946
rect 10246 29894 10276 29946
rect 10300 29894 10310 29946
rect 10310 29894 10356 29946
rect 10380 29894 10426 29946
rect 10426 29894 10436 29946
rect 10460 29894 10490 29946
rect 10490 29894 10516 29946
rect 10220 29892 10276 29894
rect 10300 29892 10356 29894
rect 10380 29892 10436 29894
rect 10460 29892 10516 29894
rect 10230 29552 10286 29608
rect 10506 29008 10562 29064
rect 10220 28858 10276 28860
rect 10300 28858 10356 28860
rect 10380 28858 10436 28860
rect 10460 28858 10516 28860
rect 10220 28806 10246 28858
rect 10246 28806 10276 28858
rect 10300 28806 10310 28858
rect 10310 28806 10356 28858
rect 10380 28806 10426 28858
rect 10426 28806 10436 28858
rect 10460 28806 10490 28858
rect 10490 28806 10516 28858
rect 10220 28804 10276 28806
rect 10300 28804 10356 28806
rect 10380 28804 10436 28806
rect 10460 28804 10516 28806
rect 10220 27770 10276 27772
rect 10300 27770 10356 27772
rect 10380 27770 10436 27772
rect 10460 27770 10516 27772
rect 10220 27718 10246 27770
rect 10246 27718 10276 27770
rect 10300 27718 10310 27770
rect 10310 27718 10356 27770
rect 10380 27718 10426 27770
rect 10426 27718 10436 27770
rect 10460 27718 10490 27770
rect 10490 27718 10516 27770
rect 10220 27716 10276 27718
rect 10300 27716 10356 27718
rect 10380 27716 10436 27718
rect 10460 27716 10516 27718
rect 10690 38800 10746 38856
rect 10874 38800 10930 38856
rect 10782 38528 10838 38584
rect 11242 39208 11298 39264
rect 12714 51584 12770 51640
rect 13174 51348 13176 51368
rect 13176 51348 13228 51368
rect 13228 51348 13230 51368
rect 12346 51176 12402 51232
rect 11242 38664 11298 38720
rect 10690 28872 10746 28928
rect 10220 26682 10276 26684
rect 10300 26682 10356 26684
rect 10380 26682 10436 26684
rect 10460 26682 10516 26684
rect 10220 26630 10246 26682
rect 10246 26630 10276 26682
rect 10300 26630 10310 26682
rect 10310 26630 10356 26682
rect 10380 26630 10426 26682
rect 10426 26630 10436 26682
rect 10460 26630 10490 26682
rect 10490 26630 10516 26682
rect 10220 26628 10276 26630
rect 10300 26628 10356 26630
rect 10380 26628 10436 26630
rect 10460 26628 10516 26630
rect 10598 26560 10654 26616
rect 10414 26152 10470 26208
rect 10220 25594 10276 25596
rect 10300 25594 10356 25596
rect 10380 25594 10436 25596
rect 10460 25594 10516 25596
rect 10220 25542 10246 25594
rect 10246 25542 10276 25594
rect 10300 25542 10310 25594
rect 10310 25542 10356 25594
rect 10380 25542 10426 25594
rect 10426 25542 10436 25594
rect 10460 25542 10490 25594
rect 10490 25542 10516 25594
rect 10220 25540 10276 25542
rect 10300 25540 10356 25542
rect 10380 25540 10436 25542
rect 10460 25540 10516 25542
rect 10220 24506 10276 24508
rect 10300 24506 10356 24508
rect 10380 24506 10436 24508
rect 10460 24506 10516 24508
rect 10220 24454 10246 24506
rect 10246 24454 10276 24506
rect 10300 24454 10310 24506
rect 10310 24454 10356 24506
rect 10380 24454 10426 24506
rect 10426 24454 10436 24506
rect 10460 24454 10490 24506
rect 10490 24454 10516 24506
rect 10220 24452 10276 24454
rect 10300 24452 10356 24454
rect 10380 24452 10436 24454
rect 10460 24452 10516 24454
rect 10220 23418 10276 23420
rect 10300 23418 10356 23420
rect 10380 23418 10436 23420
rect 10460 23418 10516 23420
rect 10220 23366 10246 23418
rect 10246 23366 10276 23418
rect 10300 23366 10310 23418
rect 10310 23366 10356 23418
rect 10380 23366 10426 23418
rect 10426 23366 10436 23418
rect 10460 23366 10490 23418
rect 10490 23366 10516 23418
rect 10220 23364 10276 23366
rect 10300 23364 10356 23366
rect 10380 23364 10436 23366
rect 10460 23364 10516 23366
rect 10220 22330 10276 22332
rect 10300 22330 10356 22332
rect 10380 22330 10436 22332
rect 10460 22330 10516 22332
rect 10220 22278 10246 22330
rect 10246 22278 10276 22330
rect 10300 22278 10310 22330
rect 10310 22278 10356 22330
rect 10380 22278 10426 22330
rect 10426 22278 10436 22330
rect 10460 22278 10490 22330
rect 10490 22278 10516 22330
rect 10220 22276 10276 22278
rect 10300 22276 10356 22278
rect 10380 22276 10436 22278
rect 10460 22276 10516 22278
rect 10220 21242 10276 21244
rect 10300 21242 10356 21244
rect 10380 21242 10436 21244
rect 10460 21242 10516 21244
rect 10220 21190 10246 21242
rect 10246 21190 10276 21242
rect 10300 21190 10310 21242
rect 10310 21190 10356 21242
rect 10380 21190 10426 21242
rect 10426 21190 10436 21242
rect 10460 21190 10490 21242
rect 10490 21190 10516 21242
rect 10220 21188 10276 21190
rect 10300 21188 10356 21190
rect 10380 21188 10436 21190
rect 10460 21188 10516 21190
rect 10220 20154 10276 20156
rect 10300 20154 10356 20156
rect 10380 20154 10436 20156
rect 10460 20154 10516 20156
rect 10220 20102 10246 20154
rect 10246 20102 10276 20154
rect 10300 20102 10310 20154
rect 10310 20102 10356 20154
rect 10380 20102 10426 20154
rect 10426 20102 10436 20154
rect 10460 20102 10490 20154
rect 10490 20102 10516 20154
rect 10220 20100 10276 20102
rect 10300 20100 10356 20102
rect 10380 20100 10436 20102
rect 10460 20100 10516 20102
rect 10220 19066 10276 19068
rect 10300 19066 10356 19068
rect 10380 19066 10436 19068
rect 10460 19066 10516 19068
rect 10220 19014 10246 19066
rect 10246 19014 10276 19066
rect 10300 19014 10310 19066
rect 10310 19014 10356 19066
rect 10380 19014 10426 19066
rect 10426 19014 10436 19066
rect 10460 19014 10490 19066
rect 10490 19014 10516 19066
rect 10220 19012 10276 19014
rect 10300 19012 10356 19014
rect 10380 19012 10436 19014
rect 10460 19012 10516 19014
rect 10220 17978 10276 17980
rect 10300 17978 10356 17980
rect 10380 17978 10436 17980
rect 10460 17978 10516 17980
rect 10220 17926 10246 17978
rect 10246 17926 10276 17978
rect 10300 17926 10310 17978
rect 10310 17926 10356 17978
rect 10380 17926 10426 17978
rect 10426 17926 10436 17978
rect 10460 17926 10490 17978
rect 10490 17926 10516 17978
rect 10220 17924 10276 17926
rect 10300 17924 10356 17926
rect 10380 17924 10436 17926
rect 10460 17924 10516 17926
rect 10220 16890 10276 16892
rect 10300 16890 10356 16892
rect 10380 16890 10436 16892
rect 10460 16890 10516 16892
rect 10220 16838 10246 16890
rect 10246 16838 10276 16890
rect 10300 16838 10310 16890
rect 10310 16838 10356 16890
rect 10380 16838 10426 16890
rect 10426 16838 10436 16890
rect 10460 16838 10490 16890
rect 10490 16838 10516 16890
rect 10220 16836 10276 16838
rect 10300 16836 10356 16838
rect 10380 16836 10436 16838
rect 10460 16836 10516 16838
rect 10220 15802 10276 15804
rect 10300 15802 10356 15804
rect 10380 15802 10436 15804
rect 10460 15802 10516 15804
rect 10220 15750 10246 15802
rect 10246 15750 10276 15802
rect 10300 15750 10310 15802
rect 10310 15750 10356 15802
rect 10380 15750 10426 15802
rect 10426 15750 10436 15802
rect 10460 15750 10490 15802
rect 10490 15750 10516 15802
rect 10220 15748 10276 15750
rect 10300 15748 10356 15750
rect 10380 15748 10436 15750
rect 10460 15748 10516 15750
rect 10782 26560 10838 26616
rect 11058 27376 11114 27432
rect 11150 26424 11206 26480
rect 10690 17876 10746 17912
rect 10690 17856 10692 17876
rect 10692 17856 10744 17876
rect 10744 17856 10746 17876
rect 10220 14714 10276 14716
rect 10300 14714 10356 14716
rect 10380 14714 10436 14716
rect 10460 14714 10516 14716
rect 10220 14662 10246 14714
rect 10246 14662 10276 14714
rect 10300 14662 10310 14714
rect 10310 14662 10356 14714
rect 10380 14662 10426 14714
rect 10426 14662 10436 14714
rect 10460 14662 10490 14714
rect 10490 14662 10516 14714
rect 10220 14660 10276 14662
rect 10300 14660 10356 14662
rect 10380 14660 10436 14662
rect 10460 14660 10516 14662
rect 10220 13626 10276 13628
rect 10300 13626 10356 13628
rect 10380 13626 10436 13628
rect 10460 13626 10516 13628
rect 10220 13574 10246 13626
rect 10246 13574 10276 13626
rect 10300 13574 10310 13626
rect 10310 13574 10356 13626
rect 10380 13574 10426 13626
rect 10426 13574 10436 13626
rect 10460 13574 10490 13626
rect 10490 13574 10516 13626
rect 10220 13572 10276 13574
rect 10300 13572 10356 13574
rect 10380 13572 10436 13574
rect 10460 13572 10516 13574
rect 10220 12538 10276 12540
rect 10300 12538 10356 12540
rect 10380 12538 10436 12540
rect 10460 12538 10516 12540
rect 10220 12486 10246 12538
rect 10246 12486 10276 12538
rect 10300 12486 10310 12538
rect 10310 12486 10356 12538
rect 10380 12486 10426 12538
rect 10426 12486 10436 12538
rect 10460 12486 10490 12538
rect 10490 12486 10516 12538
rect 10220 12484 10276 12486
rect 10300 12484 10356 12486
rect 10380 12484 10436 12486
rect 10460 12484 10516 12486
rect 10220 11450 10276 11452
rect 10300 11450 10356 11452
rect 10380 11450 10436 11452
rect 10460 11450 10516 11452
rect 10220 11398 10246 11450
rect 10246 11398 10276 11450
rect 10300 11398 10310 11450
rect 10310 11398 10356 11450
rect 10380 11398 10426 11450
rect 10426 11398 10436 11450
rect 10460 11398 10490 11450
rect 10490 11398 10516 11450
rect 10220 11396 10276 11398
rect 10300 11396 10356 11398
rect 10380 11396 10436 11398
rect 10460 11396 10516 11398
rect 8666 7248 8722 7304
rect 10220 10362 10276 10364
rect 10300 10362 10356 10364
rect 10380 10362 10436 10364
rect 10460 10362 10516 10364
rect 10220 10310 10246 10362
rect 10246 10310 10276 10362
rect 10300 10310 10310 10362
rect 10310 10310 10356 10362
rect 10380 10310 10426 10362
rect 10426 10310 10436 10362
rect 10460 10310 10490 10362
rect 10490 10310 10516 10362
rect 10220 10308 10276 10310
rect 10300 10308 10356 10310
rect 10380 10308 10436 10310
rect 10460 10308 10516 10310
rect 10966 19080 11022 19136
rect 11518 38836 11520 38856
rect 11520 38836 11572 38856
rect 11572 38836 11574 38856
rect 11518 38800 11574 38836
rect 11426 38664 11482 38720
rect 11334 38256 11390 38312
rect 11334 28908 11336 28928
rect 11336 28908 11388 28928
rect 11388 28908 11390 28928
rect 11334 28872 11390 28908
rect 11610 38120 11666 38176
rect 11242 20304 11298 20360
rect 10220 9274 10276 9276
rect 10300 9274 10356 9276
rect 10380 9274 10436 9276
rect 10460 9274 10516 9276
rect 10220 9222 10246 9274
rect 10246 9222 10276 9274
rect 10300 9222 10310 9274
rect 10310 9222 10356 9274
rect 10380 9222 10426 9274
rect 10426 9222 10436 9274
rect 10460 9222 10490 9274
rect 10490 9222 10516 9274
rect 10220 9220 10276 9222
rect 10300 9220 10356 9222
rect 10380 9220 10436 9222
rect 10460 9220 10516 9222
rect 10220 8186 10276 8188
rect 10300 8186 10356 8188
rect 10380 8186 10436 8188
rect 10460 8186 10516 8188
rect 10220 8134 10246 8186
rect 10246 8134 10276 8186
rect 10300 8134 10310 8186
rect 10310 8134 10356 8186
rect 10380 8134 10426 8186
rect 10426 8134 10436 8186
rect 10460 8134 10490 8186
rect 10490 8134 10516 8186
rect 10220 8132 10276 8134
rect 10300 8132 10356 8134
rect 10380 8132 10436 8134
rect 10460 8132 10516 8134
rect 10230 7964 10232 7984
rect 10232 7964 10284 7984
rect 10284 7964 10286 7984
rect 10230 7928 10286 7964
rect 10220 7098 10276 7100
rect 10300 7098 10356 7100
rect 10380 7098 10436 7100
rect 10460 7098 10516 7100
rect 10220 7046 10246 7098
rect 10246 7046 10276 7098
rect 10300 7046 10310 7098
rect 10310 7046 10356 7098
rect 10380 7046 10426 7098
rect 10426 7046 10436 7098
rect 10460 7046 10490 7098
rect 10490 7046 10516 7098
rect 10220 7044 10276 7046
rect 10300 7044 10356 7046
rect 10380 7044 10436 7046
rect 10460 7044 10516 7046
rect 10690 7248 10746 7304
rect 10220 6010 10276 6012
rect 10300 6010 10356 6012
rect 10380 6010 10436 6012
rect 10460 6010 10516 6012
rect 10220 5958 10246 6010
rect 10246 5958 10276 6010
rect 10300 5958 10310 6010
rect 10310 5958 10356 6010
rect 10380 5958 10426 6010
rect 10426 5958 10436 6010
rect 10460 5958 10490 6010
rect 10490 5958 10516 6010
rect 10220 5956 10276 5958
rect 10300 5956 10356 5958
rect 10380 5956 10436 5958
rect 10460 5956 10516 5958
rect 9954 5752 10010 5808
rect 11610 26832 11666 26888
rect 13174 51312 13230 51348
rect 11978 38936 12034 38992
rect 12530 39364 12586 39400
rect 12530 39344 12532 39364
rect 12532 39344 12584 39364
rect 12584 39344 12586 39364
rect 12162 37340 12164 37360
rect 12164 37340 12216 37360
rect 12216 37340 12218 37360
rect 12162 37304 12218 37340
rect 12438 37232 12494 37288
rect 12530 35264 12586 35320
rect 12070 35028 12072 35048
rect 12072 35028 12124 35048
rect 12124 35028 12126 35048
rect 12070 34992 12126 35028
rect 11886 29044 11888 29064
rect 11888 29044 11940 29064
rect 11940 29044 11942 29064
rect 11886 29008 11942 29044
rect 11886 26988 11942 27024
rect 11886 26968 11888 26988
rect 11888 26968 11940 26988
rect 11940 26968 11942 26988
rect 11794 20712 11850 20768
rect 11978 24792 12034 24848
rect 12346 30776 12402 30832
rect 12162 26696 12218 26752
rect 11886 18264 11942 18320
rect 11794 17992 11850 18048
rect 12254 24812 12310 24848
rect 12254 24792 12256 24812
rect 12256 24792 12308 24812
rect 12308 24792 12310 24812
rect 12070 18944 12126 19000
rect 10220 4922 10276 4924
rect 10300 4922 10356 4924
rect 10380 4922 10436 4924
rect 10460 4922 10516 4924
rect 10220 4870 10246 4922
rect 10246 4870 10276 4922
rect 10300 4870 10310 4922
rect 10310 4870 10356 4922
rect 10380 4870 10426 4922
rect 10426 4870 10436 4922
rect 10460 4870 10490 4922
rect 10490 4870 10516 4922
rect 10220 4868 10276 4870
rect 10300 4868 10356 4870
rect 10380 4868 10436 4870
rect 10460 4868 10516 4870
rect 11610 13232 11666 13288
rect 11610 12280 11666 12336
rect 11518 9444 11574 9480
rect 11518 9424 11520 9444
rect 11520 9424 11572 9444
rect 11572 9424 11574 9444
rect 11610 8880 11666 8936
rect 11334 3848 11390 3904
rect 10220 3834 10276 3836
rect 10300 3834 10356 3836
rect 10380 3834 10436 3836
rect 10460 3834 10516 3836
rect 10220 3782 10246 3834
rect 10246 3782 10276 3834
rect 10300 3782 10310 3834
rect 10310 3782 10356 3834
rect 10380 3782 10426 3834
rect 10426 3782 10436 3834
rect 10460 3782 10490 3834
rect 10490 3782 10516 3834
rect 10220 3780 10276 3782
rect 10300 3780 10356 3782
rect 10380 3780 10436 3782
rect 10460 3780 10516 3782
rect 10220 2746 10276 2748
rect 10300 2746 10356 2748
rect 10380 2746 10436 2748
rect 10460 2746 10516 2748
rect 10220 2694 10246 2746
rect 10246 2694 10276 2746
rect 10300 2694 10310 2746
rect 10310 2694 10356 2746
rect 10380 2694 10426 2746
rect 10426 2694 10436 2746
rect 10460 2694 10490 2746
rect 10490 2694 10516 2746
rect 10220 2692 10276 2694
rect 10300 2692 10356 2694
rect 10380 2692 10436 2694
rect 10460 2692 10516 2694
rect 12530 26560 12586 26616
rect 12714 37440 12770 37496
rect 12806 31184 12862 31240
rect 12714 27648 12770 27704
rect 12806 26968 12862 27024
rect 12530 21684 12586 21720
rect 12530 21664 12532 21684
rect 12532 21664 12584 21684
rect 12584 21664 12586 21684
rect 12254 4120 12310 4176
rect 12530 7948 12586 7984
rect 12530 7928 12532 7948
rect 12532 7928 12584 7948
rect 12584 7928 12586 7948
rect 13910 51212 13912 51232
rect 13912 51212 13964 51232
rect 13964 51212 13966 51232
rect 13910 51176 13966 51212
rect 13450 39208 13506 39264
rect 13450 37324 13506 37360
rect 13450 37304 13452 37324
rect 13452 37304 13504 37324
rect 13504 37304 13506 37324
rect 13726 37440 13782 37496
rect 13542 31728 13598 31784
rect 13174 26968 13230 27024
rect 13082 26560 13138 26616
rect 13174 26016 13230 26072
rect 12990 21528 13046 21584
rect 12806 10376 12862 10432
rect 13266 11464 13322 11520
rect 13174 10648 13230 10704
rect 14002 37340 14004 37360
rect 14004 37340 14056 37360
rect 14056 37340 14058 37360
rect 14002 37304 14058 37340
rect 14852 52250 14908 52252
rect 14932 52250 14988 52252
rect 15012 52250 15068 52252
rect 15092 52250 15148 52252
rect 14852 52198 14878 52250
rect 14878 52198 14908 52250
rect 14932 52198 14942 52250
rect 14942 52198 14988 52250
rect 15012 52198 15058 52250
rect 15058 52198 15068 52250
rect 15092 52198 15122 52250
rect 15122 52198 15148 52250
rect 14852 52196 14908 52198
rect 14932 52196 14988 52198
rect 15012 52196 15068 52198
rect 15092 52196 15148 52198
rect 14852 51162 14908 51164
rect 14932 51162 14988 51164
rect 15012 51162 15068 51164
rect 15092 51162 15148 51164
rect 14852 51110 14878 51162
rect 14878 51110 14908 51162
rect 14932 51110 14942 51162
rect 14942 51110 14988 51162
rect 15012 51110 15058 51162
rect 15058 51110 15068 51162
rect 15092 51110 15122 51162
rect 15122 51110 15148 51162
rect 14852 51108 14908 51110
rect 14932 51108 14988 51110
rect 15012 51108 15068 51110
rect 15092 51108 15148 51110
rect 14852 50074 14908 50076
rect 14932 50074 14988 50076
rect 15012 50074 15068 50076
rect 15092 50074 15148 50076
rect 14852 50022 14878 50074
rect 14878 50022 14908 50074
rect 14932 50022 14942 50074
rect 14942 50022 14988 50074
rect 15012 50022 15058 50074
rect 15058 50022 15068 50074
rect 15092 50022 15122 50074
rect 15122 50022 15148 50074
rect 14852 50020 14908 50022
rect 14932 50020 14988 50022
rect 15012 50020 15068 50022
rect 15092 50020 15148 50022
rect 14852 48986 14908 48988
rect 14932 48986 14988 48988
rect 15012 48986 15068 48988
rect 15092 48986 15148 48988
rect 14852 48934 14878 48986
rect 14878 48934 14908 48986
rect 14932 48934 14942 48986
rect 14942 48934 14988 48986
rect 15012 48934 15058 48986
rect 15058 48934 15068 48986
rect 15092 48934 15122 48986
rect 15122 48934 15148 48986
rect 14852 48932 14908 48934
rect 14932 48932 14988 48934
rect 15012 48932 15068 48934
rect 15092 48932 15148 48934
rect 15842 51584 15898 51640
rect 14852 47898 14908 47900
rect 14932 47898 14988 47900
rect 15012 47898 15068 47900
rect 15092 47898 15148 47900
rect 14852 47846 14878 47898
rect 14878 47846 14908 47898
rect 14932 47846 14942 47898
rect 14942 47846 14988 47898
rect 15012 47846 15058 47898
rect 15058 47846 15068 47898
rect 15092 47846 15122 47898
rect 15122 47846 15148 47898
rect 14852 47844 14908 47846
rect 14932 47844 14988 47846
rect 15012 47844 15068 47846
rect 15092 47844 15148 47846
rect 14852 46810 14908 46812
rect 14932 46810 14988 46812
rect 15012 46810 15068 46812
rect 15092 46810 15148 46812
rect 14852 46758 14878 46810
rect 14878 46758 14908 46810
rect 14932 46758 14942 46810
rect 14942 46758 14988 46810
rect 15012 46758 15058 46810
rect 15058 46758 15068 46810
rect 15092 46758 15122 46810
rect 15122 46758 15148 46810
rect 14852 46756 14908 46758
rect 14932 46756 14988 46758
rect 15012 46756 15068 46758
rect 15092 46756 15148 46758
rect 13910 34992 13966 35048
rect 13726 34448 13782 34504
rect 13726 32272 13782 32328
rect 13818 29844 13874 29880
rect 13818 29824 13820 29844
rect 13820 29824 13872 29844
rect 13872 29824 13874 29844
rect 13910 26968 13966 27024
rect 13726 21412 13782 21448
rect 13726 21392 13728 21412
rect 13728 21392 13780 21412
rect 13780 21392 13782 21412
rect 13726 20848 13782 20904
rect 13818 18672 13874 18728
rect 13450 11600 13506 11656
rect 14094 26016 14150 26072
rect 14278 26560 14334 26616
rect 14094 25200 14150 25256
rect 14278 25372 14280 25392
rect 14280 25372 14332 25392
rect 14332 25372 14334 25392
rect 14278 25336 14334 25372
rect 14278 24792 14334 24848
rect 14094 20748 14096 20768
rect 14096 20748 14148 20768
rect 14148 20748 14150 20768
rect 14094 20712 14150 20748
rect 14852 45722 14908 45724
rect 14932 45722 14988 45724
rect 15012 45722 15068 45724
rect 15092 45722 15148 45724
rect 14852 45670 14878 45722
rect 14878 45670 14908 45722
rect 14932 45670 14942 45722
rect 14942 45670 14988 45722
rect 15012 45670 15058 45722
rect 15058 45670 15068 45722
rect 15092 45670 15122 45722
rect 15122 45670 15148 45722
rect 14852 45668 14908 45670
rect 14932 45668 14988 45670
rect 15012 45668 15068 45670
rect 15092 45668 15148 45670
rect 14852 44634 14908 44636
rect 14932 44634 14988 44636
rect 15012 44634 15068 44636
rect 15092 44634 15148 44636
rect 14852 44582 14878 44634
rect 14878 44582 14908 44634
rect 14932 44582 14942 44634
rect 14942 44582 14988 44634
rect 15012 44582 15058 44634
rect 15058 44582 15068 44634
rect 15092 44582 15122 44634
rect 15122 44582 15148 44634
rect 14852 44580 14908 44582
rect 14932 44580 14988 44582
rect 15012 44580 15068 44582
rect 15092 44580 15148 44582
rect 14852 43546 14908 43548
rect 14932 43546 14988 43548
rect 15012 43546 15068 43548
rect 15092 43546 15148 43548
rect 14852 43494 14878 43546
rect 14878 43494 14908 43546
rect 14932 43494 14942 43546
rect 14942 43494 14988 43546
rect 15012 43494 15058 43546
rect 15058 43494 15068 43546
rect 15092 43494 15122 43546
rect 15122 43494 15148 43546
rect 14852 43492 14908 43494
rect 14932 43492 14988 43494
rect 15012 43492 15068 43494
rect 15092 43492 15148 43494
rect 14852 42458 14908 42460
rect 14932 42458 14988 42460
rect 15012 42458 15068 42460
rect 15092 42458 15148 42460
rect 14852 42406 14878 42458
rect 14878 42406 14908 42458
rect 14932 42406 14942 42458
rect 14942 42406 14988 42458
rect 15012 42406 15058 42458
rect 15058 42406 15068 42458
rect 15092 42406 15122 42458
rect 15122 42406 15148 42458
rect 14852 42404 14908 42406
rect 14932 42404 14988 42406
rect 15012 42404 15068 42406
rect 15092 42404 15148 42406
rect 14852 41370 14908 41372
rect 14932 41370 14988 41372
rect 15012 41370 15068 41372
rect 15092 41370 15148 41372
rect 14852 41318 14878 41370
rect 14878 41318 14908 41370
rect 14932 41318 14942 41370
rect 14942 41318 14988 41370
rect 15012 41318 15058 41370
rect 15058 41318 15068 41370
rect 15092 41318 15122 41370
rect 15122 41318 15148 41370
rect 14852 41316 14908 41318
rect 14932 41316 14988 41318
rect 15012 41316 15068 41318
rect 15092 41316 15148 41318
rect 14852 40282 14908 40284
rect 14932 40282 14988 40284
rect 15012 40282 15068 40284
rect 15092 40282 15148 40284
rect 14852 40230 14878 40282
rect 14878 40230 14908 40282
rect 14932 40230 14942 40282
rect 14942 40230 14988 40282
rect 15012 40230 15058 40282
rect 15058 40230 15068 40282
rect 15092 40230 15122 40282
rect 15122 40230 15148 40282
rect 14852 40228 14908 40230
rect 14932 40228 14988 40230
rect 15012 40228 15068 40230
rect 15092 40228 15148 40230
rect 14852 39194 14908 39196
rect 14932 39194 14988 39196
rect 15012 39194 15068 39196
rect 15092 39194 15148 39196
rect 14852 39142 14878 39194
rect 14878 39142 14908 39194
rect 14932 39142 14942 39194
rect 14942 39142 14988 39194
rect 15012 39142 15058 39194
rect 15058 39142 15068 39194
rect 15092 39142 15122 39194
rect 15122 39142 15148 39194
rect 14852 39140 14908 39142
rect 14932 39140 14988 39142
rect 15012 39140 15068 39142
rect 15092 39140 15148 39142
rect 15474 38800 15530 38856
rect 14852 38106 14908 38108
rect 14932 38106 14988 38108
rect 15012 38106 15068 38108
rect 15092 38106 15148 38108
rect 14852 38054 14878 38106
rect 14878 38054 14908 38106
rect 14932 38054 14942 38106
rect 14942 38054 14988 38106
rect 15012 38054 15058 38106
rect 15058 38054 15068 38106
rect 15092 38054 15122 38106
rect 15122 38054 15148 38106
rect 14852 38052 14908 38054
rect 14932 38052 14988 38054
rect 15012 38052 15068 38054
rect 15092 38052 15148 38054
rect 14852 37018 14908 37020
rect 14932 37018 14988 37020
rect 15012 37018 15068 37020
rect 15092 37018 15148 37020
rect 14852 36966 14878 37018
rect 14878 36966 14908 37018
rect 14932 36966 14942 37018
rect 14942 36966 14988 37018
rect 15012 36966 15058 37018
rect 15058 36966 15068 37018
rect 15092 36966 15122 37018
rect 15122 36966 15148 37018
rect 14852 36964 14908 36966
rect 14932 36964 14988 36966
rect 15012 36964 15068 36966
rect 15092 36964 15148 36966
rect 14852 35930 14908 35932
rect 14932 35930 14988 35932
rect 15012 35930 15068 35932
rect 15092 35930 15148 35932
rect 14852 35878 14878 35930
rect 14878 35878 14908 35930
rect 14932 35878 14942 35930
rect 14942 35878 14988 35930
rect 15012 35878 15058 35930
rect 15058 35878 15068 35930
rect 15092 35878 15122 35930
rect 15122 35878 15148 35930
rect 14852 35876 14908 35878
rect 14932 35876 14988 35878
rect 15012 35876 15068 35878
rect 15092 35876 15148 35878
rect 14830 34992 14886 35048
rect 14852 34842 14908 34844
rect 14932 34842 14988 34844
rect 15012 34842 15068 34844
rect 15092 34842 15148 34844
rect 14852 34790 14878 34842
rect 14878 34790 14908 34842
rect 14932 34790 14942 34842
rect 14942 34790 14988 34842
rect 15012 34790 15058 34842
rect 15058 34790 15068 34842
rect 15092 34790 15122 34842
rect 15122 34790 15148 34842
rect 14852 34788 14908 34790
rect 14932 34788 14988 34790
rect 15012 34788 15068 34790
rect 15092 34788 15148 34790
rect 14852 33754 14908 33756
rect 14932 33754 14988 33756
rect 15012 33754 15068 33756
rect 15092 33754 15148 33756
rect 14852 33702 14878 33754
rect 14878 33702 14908 33754
rect 14932 33702 14942 33754
rect 14942 33702 14988 33754
rect 15012 33702 15058 33754
rect 15058 33702 15068 33754
rect 15092 33702 15122 33754
rect 15122 33702 15148 33754
rect 14852 33700 14908 33702
rect 14932 33700 14988 33702
rect 15012 33700 15068 33702
rect 15092 33700 15148 33702
rect 14852 32666 14908 32668
rect 14932 32666 14988 32668
rect 15012 32666 15068 32668
rect 15092 32666 15148 32668
rect 14852 32614 14878 32666
rect 14878 32614 14908 32666
rect 14932 32614 14942 32666
rect 14942 32614 14988 32666
rect 15012 32614 15058 32666
rect 15058 32614 15068 32666
rect 15092 32614 15122 32666
rect 15122 32614 15148 32666
rect 14852 32612 14908 32614
rect 14932 32612 14988 32614
rect 15012 32612 15068 32614
rect 15092 32612 15148 32614
rect 14852 31578 14908 31580
rect 14932 31578 14988 31580
rect 15012 31578 15068 31580
rect 15092 31578 15148 31580
rect 14852 31526 14878 31578
rect 14878 31526 14908 31578
rect 14932 31526 14942 31578
rect 14942 31526 14988 31578
rect 15012 31526 15058 31578
rect 15058 31526 15068 31578
rect 15092 31526 15122 31578
rect 15122 31526 15148 31578
rect 14852 31524 14908 31526
rect 14932 31524 14988 31526
rect 15012 31524 15068 31526
rect 15092 31524 15148 31526
rect 15106 31320 15162 31376
rect 14852 30490 14908 30492
rect 14932 30490 14988 30492
rect 15012 30490 15068 30492
rect 15092 30490 15148 30492
rect 14852 30438 14878 30490
rect 14878 30438 14908 30490
rect 14932 30438 14942 30490
rect 14942 30438 14988 30490
rect 15012 30438 15058 30490
rect 15058 30438 15068 30490
rect 15092 30438 15122 30490
rect 15122 30438 15148 30490
rect 14852 30436 14908 30438
rect 14932 30436 14988 30438
rect 15012 30436 15068 30438
rect 15092 30436 15148 30438
rect 15474 36080 15530 36136
rect 15658 36080 15714 36136
rect 15474 31320 15530 31376
rect 15474 30796 15530 30832
rect 15474 30776 15476 30796
rect 15476 30776 15528 30796
rect 15528 30776 15530 30796
rect 15566 29824 15622 29880
rect 14852 29402 14908 29404
rect 14932 29402 14988 29404
rect 15012 29402 15068 29404
rect 15092 29402 15148 29404
rect 14852 29350 14878 29402
rect 14878 29350 14908 29402
rect 14932 29350 14942 29402
rect 14942 29350 14988 29402
rect 15012 29350 15058 29402
rect 15058 29350 15068 29402
rect 15092 29350 15122 29402
rect 15122 29350 15148 29402
rect 14852 29348 14908 29350
rect 14932 29348 14988 29350
rect 15012 29348 15068 29350
rect 15092 29348 15148 29350
rect 14852 28314 14908 28316
rect 14932 28314 14988 28316
rect 15012 28314 15068 28316
rect 15092 28314 15148 28316
rect 14852 28262 14878 28314
rect 14878 28262 14908 28314
rect 14932 28262 14942 28314
rect 14942 28262 14988 28314
rect 15012 28262 15058 28314
rect 15058 28262 15068 28314
rect 15092 28262 15122 28314
rect 15122 28262 15148 28314
rect 14852 28260 14908 28262
rect 14932 28260 14988 28262
rect 15012 28260 15068 28262
rect 15092 28260 15148 28262
rect 14852 27226 14908 27228
rect 14932 27226 14988 27228
rect 15012 27226 15068 27228
rect 15092 27226 15148 27228
rect 14852 27174 14878 27226
rect 14878 27174 14908 27226
rect 14932 27174 14942 27226
rect 14942 27174 14988 27226
rect 15012 27174 15058 27226
rect 15058 27174 15068 27226
rect 15092 27174 15122 27226
rect 15122 27174 15148 27226
rect 14852 27172 14908 27174
rect 14932 27172 14988 27174
rect 15012 27172 15068 27174
rect 15092 27172 15148 27174
rect 14554 26560 14610 26616
rect 14738 26852 14794 26888
rect 14738 26832 14740 26852
rect 14740 26832 14792 26852
rect 14792 26832 14794 26852
rect 14852 26138 14908 26140
rect 14932 26138 14988 26140
rect 15012 26138 15068 26140
rect 15092 26138 15148 26140
rect 14852 26086 14878 26138
rect 14878 26086 14908 26138
rect 14932 26086 14942 26138
rect 14942 26086 14988 26138
rect 15012 26086 15058 26138
rect 15058 26086 15068 26138
rect 15092 26086 15122 26138
rect 15122 26086 15148 26138
rect 14852 26084 14908 26086
rect 14932 26084 14988 26086
rect 15012 26084 15068 26086
rect 15092 26084 15148 26086
rect 15566 29572 15622 29608
rect 15566 29552 15568 29572
rect 15568 29552 15620 29572
rect 15620 29552 15622 29572
rect 15474 29008 15530 29064
rect 14852 25050 14908 25052
rect 14932 25050 14988 25052
rect 15012 25050 15068 25052
rect 15092 25050 15148 25052
rect 14852 24998 14878 25050
rect 14878 24998 14908 25050
rect 14932 24998 14942 25050
rect 14942 24998 14988 25050
rect 15012 24998 15058 25050
rect 15058 24998 15068 25050
rect 15092 24998 15122 25050
rect 15122 24998 15148 25050
rect 14852 24996 14908 24998
rect 14932 24996 14988 24998
rect 15012 24996 15068 24998
rect 15092 24996 15148 24998
rect 14852 23962 14908 23964
rect 14932 23962 14988 23964
rect 15012 23962 15068 23964
rect 15092 23962 15148 23964
rect 14852 23910 14878 23962
rect 14878 23910 14908 23962
rect 14932 23910 14942 23962
rect 14942 23910 14988 23962
rect 15012 23910 15058 23962
rect 15058 23910 15068 23962
rect 15092 23910 15122 23962
rect 15122 23910 15148 23962
rect 14852 23908 14908 23910
rect 14932 23908 14988 23910
rect 15012 23908 15068 23910
rect 15092 23908 15148 23910
rect 14852 22874 14908 22876
rect 14932 22874 14988 22876
rect 15012 22874 15068 22876
rect 15092 22874 15148 22876
rect 14852 22822 14878 22874
rect 14878 22822 14908 22874
rect 14932 22822 14942 22874
rect 14942 22822 14988 22874
rect 15012 22822 15058 22874
rect 15058 22822 15068 22874
rect 15092 22822 15122 22874
rect 15122 22822 15148 22874
rect 14852 22820 14908 22822
rect 14932 22820 14988 22822
rect 15012 22820 15068 22822
rect 15092 22820 15148 22822
rect 14852 21786 14908 21788
rect 14932 21786 14988 21788
rect 15012 21786 15068 21788
rect 15092 21786 15148 21788
rect 14852 21734 14878 21786
rect 14878 21734 14908 21786
rect 14932 21734 14942 21786
rect 14942 21734 14988 21786
rect 15012 21734 15058 21786
rect 15058 21734 15068 21786
rect 15092 21734 15122 21786
rect 15122 21734 15148 21786
rect 14852 21732 14908 21734
rect 14932 21732 14988 21734
rect 15012 21732 15068 21734
rect 15092 21732 15148 21734
rect 14852 20698 14908 20700
rect 14932 20698 14988 20700
rect 15012 20698 15068 20700
rect 15092 20698 15148 20700
rect 14852 20646 14878 20698
rect 14878 20646 14908 20698
rect 14932 20646 14942 20698
rect 14942 20646 14988 20698
rect 15012 20646 15058 20698
rect 15058 20646 15068 20698
rect 15092 20646 15122 20698
rect 15122 20646 15148 20698
rect 14852 20644 14908 20646
rect 14932 20644 14988 20646
rect 15012 20644 15068 20646
rect 15092 20644 15148 20646
rect 14852 19610 14908 19612
rect 14932 19610 14988 19612
rect 15012 19610 15068 19612
rect 15092 19610 15148 19612
rect 14852 19558 14878 19610
rect 14878 19558 14908 19610
rect 14932 19558 14942 19610
rect 14942 19558 14988 19610
rect 15012 19558 15058 19610
rect 15058 19558 15068 19610
rect 15092 19558 15122 19610
rect 15122 19558 15148 19610
rect 14852 19556 14908 19558
rect 14932 19556 14988 19558
rect 15012 19556 15068 19558
rect 15092 19556 15148 19558
rect 14852 18522 14908 18524
rect 14932 18522 14988 18524
rect 15012 18522 15068 18524
rect 15092 18522 15148 18524
rect 14852 18470 14878 18522
rect 14878 18470 14908 18522
rect 14932 18470 14942 18522
rect 14942 18470 14988 18522
rect 15012 18470 15058 18522
rect 15058 18470 15068 18522
rect 15092 18470 15122 18522
rect 15122 18470 15148 18522
rect 14852 18468 14908 18470
rect 14932 18468 14988 18470
rect 15012 18468 15068 18470
rect 15092 18468 15148 18470
rect 14852 17434 14908 17436
rect 14932 17434 14988 17436
rect 15012 17434 15068 17436
rect 15092 17434 15148 17436
rect 14852 17382 14878 17434
rect 14878 17382 14908 17434
rect 14932 17382 14942 17434
rect 14942 17382 14988 17434
rect 15012 17382 15058 17434
rect 15058 17382 15068 17434
rect 15092 17382 15122 17434
rect 15122 17382 15148 17434
rect 14852 17380 14908 17382
rect 14932 17380 14988 17382
rect 15012 17380 15068 17382
rect 15092 17380 15148 17382
rect 14852 16346 14908 16348
rect 14932 16346 14988 16348
rect 15012 16346 15068 16348
rect 15092 16346 15148 16348
rect 14852 16294 14878 16346
rect 14878 16294 14908 16346
rect 14932 16294 14942 16346
rect 14942 16294 14988 16346
rect 15012 16294 15058 16346
rect 15058 16294 15068 16346
rect 15092 16294 15122 16346
rect 15122 16294 15148 16346
rect 14852 16292 14908 16294
rect 14932 16292 14988 16294
rect 15012 16292 15068 16294
rect 15092 16292 15148 16294
rect 14852 15258 14908 15260
rect 14932 15258 14988 15260
rect 15012 15258 15068 15260
rect 15092 15258 15148 15260
rect 14852 15206 14878 15258
rect 14878 15206 14908 15258
rect 14932 15206 14942 15258
rect 14942 15206 14988 15258
rect 15012 15206 15058 15258
rect 15058 15206 15068 15258
rect 15092 15206 15122 15258
rect 15122 15206 15148 15258
rect 14852 15204 14908 15206
rect 14932 15204 14988 15206
rect 15012 15204 15068 15206
rect 15092 15204 15148 15206
rect 14094 3984 14150 4040
rect 14852 14170 14908 14172
rect 14932 14170 14988 14172
rect 15012 14170 15068 14172
rect 15092 14170 15148 14172
rect 14852 14118 14878 14170
rect 14878 14118 14908 14170
rect 14932 14118 14942 14170
rect 14942 14118 14988 14170
rect 15012 14118 15058 14170
rect 15058 14118 15068 14170
rect 15092 14118 15122 14170
rect 15122 14118 15148 14170
rect 14852 14116 14908 14118
rect 14932 14116 14988 14118
rect 15012 14116 15068 14118
rect 15092 14116 15148 14118
rect 14852 13082 14908 13084
rect 14932 13082 14988 13084
rect 15012 13082 15068 13084
rect 15092 13082 15148 13084
rect 14852 13030 14878 13082
rect 14878 13030 14908 13082
rect 14932 13030 14942 13082
rect 14942 13030 14988 13082
rect 15012 13030 15058 13082
rect 15058 13030 15068 13082
rect 15092 13030 15122 13082
rect 15122 13030 15148 13082
rect 14852 13028 14908 13030
rect 14932 13028 14988 13030
rect 15012 13028 15068 13030
rect 15092 13028 15148 13030
rect 14852 11994 14908 11996
rect 14932 11994 14988 11996
rect 15012 11994 15068 11996
rect 15092 11994 15148 11996
rect 14852 11942 14878 11994
rect 14878 11942 14908 11994
rect 14932 11942 14942 11994
rect 14942 11942 14988 11994
rect 15012 11942 15058 11994
rect 15058 11942 15068 11994
rect 15092 11942 15122 11994
rect 15122 11942 15148 11994
rect 14852 11940 14908 11942
rect 14932 11940 14988 11942
rect 15012 11940 15068 11942
rect 15092 11940 15148 11942
rect 14852 10906 14908 10908
rect 14932 10906 14988 10908
rect 15012 10906 15068 10908
rect 15092 10906 15148 10908
rect 14852 10854 14878 10906
rect 14878 10854 14908 10906
rect 14932 10854 14942 10906
rect 14942 10854 14988 10906
rect 15012 10854 15058 10906
rect 15058 10854 15068 10906
rect 15092 10854 15122 10906
rect 15122 10854 15148 10906
rect 14852 10852 14908 10854
rect 14932 10852 14988 10854
rect 15012 10852 15068 10854
rect 15092 10852 15148 10854
rect 14852 9818 14908 9820
rect 14932 9818 14988 9820
rect 15012 9818 15068 9820
rect 15092 9818 15148 9820
rect 14852 9766 14878 9818
rect 14878 9766 14908 9818
rect 14932 9766 14942 9818
rect 14942 9766 14988 9818
rect 15012 9766 15058 9818
rect 15058 9766 15068 9818
rect 15092 9766 15122 9818
rect 15122 9766 15148 9818
rect 14852 9764 14908 9766
rect 14932 9764 14988 9766
rect 15012 9764 15068 9766
rect 15092 9764 15148 9766
rect 15106 8916 15108 8936
rect 15108 8916 15160 8936
rect 15160 8916 15162 8936
rect 15106 8880 15162 8916
rect 14852 8730 14908 8732
rect 14932 8730 14988 8732
rect 15012 8730 15068 8732
rect 15092 8730 15148 8732
rect 14852 8678 14878 8730
rect 14878 8678 14908 8730
rect 14932 8678 14942 8730
rect 14942 8678 14988 8730
rect 15012 8678 15058 8730
rect 15058 8678 15068 8730
rect 15092 8678 15122 8730
rect 15122 8678 15148 8730
rect 14852 8676 14908 8678
rect 14932 8676 14988 8678
rect 15012 8676 15068 8678
rect 15092 8676 15148 8678
rect 14852 7642 14908 7644
rect 14932 7642 14988 7644
rect 15012 7642 15068 7644
rect 15092 7642 15148 7644
rect 14852 7590 14878 7642
rect 14878 7590 14908 7642
rect 14932 7590 14942 7642
rect 14942 7590 14988 7642
rect 15012 7590 15058 7642
rect 15058 7590 15068 7642
rect 15092 7590 15122 7642
rect 15122 7590 15148 7642
rect 14852 7588 14908 7590
rect 14932 7588 14988 7590
rect 15012 7588 15068 7590
rect 15092 7588 15148 7590
rect 15014 7284 15016 7304
rect 15016 7284 15068 7304
rect 15068 7284 15070 7304
rect 15014 7248 15070 7284
rect 14852 6554 14908 6556
rect 14932 6554 14988 6556
rect 15012 6554 15068 6556
rect 15092 6554 15148 6556
rect 14852 6502 14878 6554
rect 14878 6502 14908 6554
rect 14932 6502 14942 6554
rect 14942 6502 14988 6554
rect 15012 6502 15058 6554
rect 15058 6502 15068 6554
rect 15092 6502 15122 6554
rect 15122 6502 15148 6554
rect 14852 6500 14908 6502
rect 14932 6500 14988 6502
rect 15012 6500 15068 6502
rect 15092 6500 15148 6502
rect 14852 5466 14908 5468
rect 14932 5466 14988 5468
rect 15012 5466 15068 5468
rect 15092 5466 15148 5468
rect 14852 5414 14878 5466
rect 14878 5414 14908 5466
rect 14932 5414 14942 5466
rect 14942 5414 14988 5466
rect 15012 5414 15058 5466
rect 15058 5414 15068 5466
rect 15092 5414 15122 5466
rect 15122 5414 15148 5466
rect 14852 5412 14908 5414
rect 14932 5412 14988 5414
rect 15012 5412 15068 5414
rect 15092 5412 15148 5414
rect 15842 39516 15844 39536
rect 15844 39516 15896 39536
rect 15896 39516 15898 39536
rect 15842 39480 15898 39516
rect 15842 39344 15898 39400
rect 16026 35808 16082 35864
rect 19484 52794 19540 52796
rect 19564 52794 19620 52796
rect 19644 52794 19700 52796
rect 19724 52794 19780 52796
rect 19484 52742 19510 52794
rect 19510 52742 19540 52794
rect 19564 52742 19574 52794
rect 19574 52742 19620 52794
rect 19644 52742 19690 52794
rect 19690 52742 19700 52794
rect 19724 52742 19754 52794
rect 19754 52742 19780 52794
rect 19484 52740 19540 52742
rect 19564 52740 19620 52742
rect 19644 52740 19700 52742
rect 19724 52740 19780 52742
rect 19484 51706 19540 51708
rect 19564 51706 19620 51708
rect 19644 51706 19700 51708
rect 19724 51706 19780 51708
rect 19484 51654 19510 51706
rect 19510 51654 19540 51706
rect 19564 51654 19574 51706
rect 19574 51654 19620 51706
rect 19644 51654 19690 51706
rect 19690 51654 19700 51706
rect 19724 51654 19754 51706
rect 19754 51654 19780 51706
rect 19484 51652 19540 51654
rect 19564 51652 19620 51654
rect 19644 51652 19700 51654
rect 19724 51652 19780 51654
rect 16578 38664 16634 38720
rect 16118 32000 16174 32056
rect 16210 31728 16266 31784
rect 15934 26424 15990 26480
rect 16486 31884 16542 31920
rect 16486 31864 16488 31884
rect 16488 31864 16540 31884
rect 16540 31864 16542 31884
rect 15750 21936 15806 21992
rect 15934 20984 15990 21040
rect 15750 17856 15806 17912
rect 16118 20304 16174 20360
rect 14852 4378 14908 4380
rect 14932 4378 14988 4380
rect 15012 4378 15068 4380
rect 15092 4378 15148 4380
rect 14852 4326 14878 4378
rect 14878 4326 14908 4378
rect 14932 4326 14942 4378
rect 14942 4326 14988 4378
rect 15012 4326 15058 4378
rect 15058 4326 15068 4378
rect 15092 4326 15122 4378
rect 15122 4326 15148 4378
rect 14852 4324 14908 4326
rect 14932 4324 14988 4326
rect 15012 4324 15068 4326
rect 15092 4324 15148 4326
rect 14830 3884 14832 3904
rect 14832 3884 14884 3904
rect 14884 3884 14886 3904
rect 14830 3848 14886 3884
rect 14852 3290 14908 3292
rect 14932 3290 14988 3292
rect 15012 3290 15068 3292
rect 15092 3290 15148 3292
rect 14852 3238 14878 3290
rect 14878 3238 14908 3290
rect 14932 3238 14942 3290
rect 14942 3238 14988 3290
rect 15012 3238 15058 3290
rect 15058 3238 15068 3290
rect 15092 3238 15122 3290
rect 15122 3238 15148 3290
rect 14852 3236 14908 3238
rect 14932 3236 14988 3238
rect 15012 3236 15068 3238
rect 15092 3236 15148 3238
rect 15658 7248 15714 7304
rect 15934 10532 15990 10568
rect 15934 10512 15936 10532
rect 15936 10512 15988 10532
rect 15988 10512 15990 10532
rect 16394 19080 16450 19136
rect 16394 18148 16450 18184
rect 16394 18128 16396 18148
rect 16396 18128 16448 18148
rect 16448 18128 16450 18148
rect 15474 4020 15476 4040
rect 15476 4020 15528 4040
rect 15528 4020 15530 4040
rect 15474 3984 15530 4020
rect 16026 5752 16082 5808
rect 16394 12588 16396 12608
rect 16396 12588 16448 12608
rect 16448 12588 16450 12608
rect 16394 12552 16450 12588
rect 16670 17992 16726 18048
rect 16578 12280 16634 12336
rect 17038 30776 17094 30832
rect 17038 26288 17094 26344
rect 16486 4120 16542 4176
rect 17038 18128 17094 18184
rect 17406 35672 17462 35728
rect 17314 26696 17370 26752
rect 17314 24792 17370 24848
rect 17222 18672 17278 18728
rect 16854 3576 16910 3632
rect 17866 38664 17922 38720
rect 18050 34584 18106 34640
rect 17958 34348 17960 34368
rect 17960 34348 18012 34368
rect 18012 34348 18014 34368
rect 17958 34312 18014 34348
rect 17406 12588 17408 12608
rect 17408 12588 17460 12608
rect 17460 12588 17462 12608
rect 17406 12552 17462 12588
rect 17866 27376 17922 27432
rect 17866 26424 17922 26480
rect 18050 27376 18106 27432
rect 18050 18672 18106 18728
rect 19484 50618 19540 50620
rect 19564 50618 19620 50620
rect 19644 50618 19700 50620
rect 19724 50618 19780 50620
rect 19484 50566 19510 50618
rect 19510 50566 19540 50618
rect 19564 50566 19574 50618
rect 19574 50566 19620 50618
rect 19644 50566 19690 50618
rect 19690 50566 19700 50618
rect 19724 50566 19754 50618
rect 19754 50566 19780 50618
rect 19484 50564 19540 50566
rect 19564 50564 19620 50566
rect 19644 50564 19700 50566
rect 19724 50564 19780 50566
rect 19484 49530 19540 49532
rect 19564 49530 19620 49532
rect 19644 49530 19700 49532
rect 19724 49530 19780 49532
rect 19484 49478 19510 49530
rect 19510 49478 19540 49530
rect 19564 49478 19574 49530
rect 19574 49478 19620 49530
rect 19644 49478 19690 49530
rect 19690 49478 19700 49530
rect 19724 49478 19754 49530
rect 19754 49478 19780 49530
rect 19484 49476 19540 49478
rect 19564 49476 19620 49478
rect 19644 49476 19700 49478
rect 19724 49476 19780 49478
rect 19484 48442 19540 48444
rect 19564 48442 19620 48444
rect 19644 48442 19700 48444
rect 19724 48442 19780 48444
rect 19484 48390 19510 48442
rect 19510 48390 19540 48442
rect 19564 48390 19574 48442
rect 19574 48390 19620 48442
rect 19644 48390 19690 48442
rect 19690 48390 19700 48442
rect 19724 48390 19754 48442
rect 19754 48390 19780 48442
rect 19484 48388 19540 48390
rect 19564 48388 19620 48390
rect 19644 48388 19700 48390
rect 19724 48388 19780 48390
rect 18786 35708 18788 35728
rect 18788 35708 18840 35728
rect 18840 35708 18842 35728
rect 18786 35672 18842 35708
rect 18326 27512 18382 27568
rect 18326 27376 18382 27432
rect 18326 20032 18382 20088
rect 18786 32000 18842 32056
rect 18510 27648 18566 27704
rect 18878 31184 18934 31240
rect 18418 10648 18474 10704
rect 18142 10376 18198 10432
rect 18418 9968 18474 10024
rect 18786 27376 18842 27432
rect 19154 34584 19210 34640
rect 19484 47354 19540 47356
rect 19564 47354 19620 47356
rect 19644 47354 19700 47356
rect 19724 47354 19780 47356
rect 19484 47302 19510 47354
rect 19510 47302 19540 47354
rect 19564 47302 19574 47354
rect 19574 47302 19620 47354
rect 19644 47302 19690 47354
rect 19690 47302 19700 47354
rect 19724 47302 19754 47354
rect 19754 47302 19780 47354
rect 19484 47300 19540 47302
rect 19564 47300 19620 47302
rect 19644 47300 19700 47302
rect 19724 47300 19780 47302
rect 19484 46266 19540 46268
rect 19564 46266 19620 46268
rect 19644 46266 19700 46268
rect 19724 46266 19780 46268
rect 19484 46214 19510 46266
rect 19510 46214 19540 46266
rect 19564 46214 19574 46266
rect 19574 46214 19620 46266
rect 19644 46214 19690 46266
rect 19690 46214 19700 46266
rect 19724 46214 19754 46266
rect 19754 46214 19780 46266
rect 19484 46212 19540 46214
rect 19564 46212 19620 46214
rect 19644 46212 19700 46214
rect 19724 46212 19780 46214
rect 19484 45178 19540 45180
rect 19564 45178 19620 45180
rect 19644 45178 19700 45180
rect 19724 45178 19780 45180
rect 19484 45126 19510 45178
rect 19510 45126 19540 45178
rect 19564 45126 19574 45178
rect 19574 45126 19620 45178
rect 19644 45126 19690 45178
rect 19690 45126 19700 45178
rect 19724 45126 19754 45178
rect 19754 45126 19780 45178
rect 19484 45124 19540 45126
rect 19564 45124 19620 45126
rect 19644 45124 19700 45126
rect 19724 45124 19780 45126
rect 19484 44090 19540 44092
rect 19564 44090 19620 44092
rect 19644 44090 19700 44092
rect 19724 44090 19780 44092
rect 19484 44038 19510 44090
rect 19510 44038 19540 44090
rect 19564 44038 19574 44090
rect 19574 44038 19620 44090
rect 19644 44038 19690 44090
rect 19690 44038 19700 44090
rect 19724 44038 19754 44090
rect 19754 44038 19780 44090
rect 19484 44036 19540 44038
rect 19564 44036 19620 44038
rect 19644 44036 19700 44038
rect 19724 44036 19780 44038
rect 19484 43002 19540 43004
rect 19564 43002 19620 43004
rect 19644 43002 19700 43004
rect 19724 43002 19780 43004
rect 19484 42950 19510 43002
rect 19510 42950 19540 43002
rect 19564 42950 19574 43002
rect 19574 42950 19620 43002
rect 19644 42950 19690 43002
rect 19690 42950 19700 43002
rect 19724 42950 19754 43002
rect 19754 42950 19780 43002
rect 19484 42948 19540 42950
rect 19564 42948 19620 42950
rect 19644 42948 19700 42950
rect 19724 42948 19780 42950
rect 19484 41914 19540 41916
rect 19564 41914 19620 41916
rect 19644 41914 19700 41916
rect 19724 41914 19780 41916
rect 19484 41862 19510 41914
rect 19510 41862 19540 41914
rect 19564 41862 19574 41914
rect 19574 41862 19620 41914
rect 19644 41862 19690 41914
rect 19690 41862 19700 41914
rect 19724 41862 19754 41914
rect 19754 41862 19780 41914
rect 19484 41860 19540 41862
rect 19564 41860 19620 41862
rect 19644 41860 19700 41862
rect 19724 41860 19780 41862
rect 19484 40826 19540 40828
rect 19564 40826 19620 40828
rect 19644 40826 19700 40828
rect 19724 40826 19780 40828
rect 19484 40774 19510 40826
rect 19510 40774 19540 40826
rect 19564 40774 19574 40826
rect 19574 40774 19620 40826
rect 19644 40774 19690 40826
rect 19690 40774 19700 40826
rect 19724 40774 19754 40826
rect 19754 40774 19780 40826
rect 19484 40772 19540 40774
rect 19564 40772 19620 40774
rect 19644 40772 19700 40774
rect 19724 40772 19780 40774
rect 19484 39738 19540 39740
rect 19564 39738 19620 39740
rect 19644 39738 19700 39740
rect 19724 39738 19780 39740
rect 19484 39686 19510 39738
rect 19510 39686 19540 39738
rect 19564 39686 19574 39738
rect 19574 39686 19620 39738
rect 19644 39686 19690 39738
rect 19690 39686 19700 39738
rect 19724 39686 19754 39738
rect 19754 39686 19780 39738
rect 19484 39684 19540 39686
rect 19564 39684 19620 39686
rect 19644 39684 19700 39686
rect 19724 39684 19780 39686
rect 19484 38650 19540 38652
rect 19564 38650 19620 38652
rect 19644 38650 19700 38652
rect 19724 38650 19780 38652
rect 19484 38598 19510 38650
rect 19510 38598 19540 38650
rect 19564 38598 19574 38650
rect 19574 38598 19620 38650
rect 19644 38598 19690 38650
rect 19690 38598 19700 38650
rect 19724 38598 19754 38650
rect 19754 38598 19780 38650
rect 19484 38596 19540 38598
rect 19564 38596 19620 38598
rect 19644 38596 19700 38598
rect 19724 38596 19780 38598
rect 19484 37562 19540 37564
rect 19564 37562 19620 37564
rect 19644 37562 19700 37564
rect 19724 37562 19780 37564
rect 19484 37510 19510 37562
rect 19510 37510 19540 37562
rect 19564 37510 19574 37562
rect 19574 37510 19620 37562
rect 19644 37510 19690 37562
rect 19690 37510 19700 37562
rect 19724 37510 19754 37562
rect 19754 37510 19780 37562
rect 19484 37508 19540 37510
rect 19564 37508 19620 37510
rect 19644 37508 19700 37510
rect 19724 37508 19780 37510
rect 19484 36474 19540 36476
rect 19564 36474 19620 36476
rect 19644 36474 19700 36476
rect 19724 36474 19780 36476
rect 19484 36422 19510 36474
rect 19510 36422 19540 36474
rect 19564 36422 19574 36474
rect 19574 36422 19620 36474
rect 19644 36422 19690 36474
rect 19690 36422 19700 36474
rect 19724 36422 19754 36474
rect 19754 36422 19780 36474
rect 19484 36420 19540 36422
rect 19564 36420 19620 36422
rect 19644 36420 19700 36422
rect 19724 36420 19780 36422
rect 19484 35386 19540 35388
rect 19564 35386 19620 35388
rect 19644 35386 19700 35388
rect 19724 35386 19780 35388
rect 19484 35334 19510 35386
rect 19510 35334 19540 35386
rect 19564 35334 19574 35386
rect 19574 35334 19620 35386
rect 19644 35334 19690 35386
rect 19690 35334 19700 35386
rect 19724 35334 19754 35386
rect 19754 35334 19780 35386
rect 19484 35332 19540 35334
rect 19564 35332 19620 35334
rect 19644 35332 19700 35334
rect 19724 35332 19780 35334
rect 19484 34298 19540 34300
rect 19564 34298 19620 34300
rect 19644 34298 19700 34300
rect 19724 34298 19780 34300
rect 19484 34246 19510 34298
rect 19510 34246 19540 34298
rect 19564 34246 19574 34298
rect 19574 34246 19620 34298
rect 19644 34246 19690 34298
rect 19690 34246 19700 34298
rect 19724 34246 19754 34298
rect 19754 34246 19780 34298
rect 19484 34244 19540 34246
rect 19564 34244 19620 34246
rect 19644 34244 19700 34246
rect 19724 34244 19780 34246
rect 19484 33210 19540 33212
rect 19564 33210 19620 33212
rect 19644 33210 19700 33212
rect 19724 33210 19780 33212
rect 19484 33158 19510 33210
rect 19510 33158 19540 33210
rect 19564 33158 19574 33210
rect 19574 33158 19620 33210
rect 19644 33158 19690 33210
rect 19690 33158 19700 33210
rect 19724 33158 19754 33210
rect 19754 33158 19780 33210
rect 19484 33156 19540 33158
rect 19564 33156 19620 33158
rect 19644 33156 19700 33158
rect 19724 33156 19780 33158
rect 19484 32122 19540 32124
rect 19564 32122 19620 32124
rect 19644 32122 19700 32124
rect 19724 32122 19780 32124
rect 19484 32070 19510 32122
rect 19510 32070 19540 32122
rect 19564 32070 19574 32122
rect 19574 32070 19620 32122
rect 19644 32070 19690 32122
rect 19690 32070 19700 32122
rect 19724 32070 19754 32122
rect 19754 32070 19780 32122
rect 19484 32068 19540 32070
rect 19564 32068 19620 32070
rect 19644 32068 19700 32070
rect 19724 32068 19780 32070
rect 18970 15580 18972 15600
rect 18972 15580 19024 15600
rect 19024 15580 19026 15600
rect 18970 15544 19026 15580
rect 18602 12552 18658 12608
rect 18602 12316 18604 12336
rect 18604 12316 18656 12336
rect 18656 12316 18658 12336
rect 18602 12280 18658 12316
rect 18786 12552 18842 12608
rect 19484 31034 19540 31036
rect 19564 31034 19620 31036
rect 19644 31034 19700 31036
rect 19724 31034 19780 31036
rect 19484 30982 19510 31034
rect 19510 30982 19540 31034
rect 19564 30982 19574 31034
rect 19574 30982 19620 31034
rect 19644 30982 19690 31034
rect 19690 30982 19700 31034
rect 19724 30982 19754 31034
rect 19754 30982 19780 31034
rect 19484 30980 19540 30982
rect 19564 30980 19620 30982
rect 19644 30980 19700 30982
rect 19724 30980 19780 30982
rect 19484 29946 19540 29948
rect 19564 29946 19620 29948
rect 19644 29946 19700 29948
rect 19724 29946 19780 29948
rect 19484 29894 19510 29946
rect 19510 29894 19540 29946
rect 19564 29894 19574 29946
rect 19574 29894 19620 29946
rect 19644 29894 19690 29946
rect 19690 29894 19700 29946
rect 19724 29894 19754 29946
rect 19754 29894 19780 29946
rect 19484 29892 19540 29894
rect 19564 29892 19620 29894
rect 19644 29892 19700 29894
rect 19724 29892 19780 29894
rect 19484 28858 19540 28860
rect 19564 28858 19620 28860
rect 19644 28858 19700 28860
rect 19724 28858 19780 28860
rect 19484 28806 19510 28858
rect 19510 28806 19540 28858
rect 19564 28806 19574 28858
rect 19574 28806 19620 28858
rect 19644 28806 19690 28858
rect 19690 28806 19700 28858
rect 19724 28806 19754 28858
rect 19754 28806 19780 28858
rect 19484 28804 19540 28806
rect 19564 28804 19620 28806
rect 19644 28804 19700 28806
rect 19724 28804 19780 28806
rect 19484 27770 19540 27772
rect 19564 27770 19620 27772
rect 19644 27770 19700 27772
rect 19724 27770 19780 27772
rect 19484 27718 19510 27770
rect 19510 27718 19540 27770
rect 19564 27718 19574 27770
rect 19574 27718 19620 27770
rect 19644 27718 19690 27770
rect 19690 27718 19700 27770
rect 19724 27718 19754 27770
rect 19754 27718 19780 27770
rect 19484 27716 19540 27718
rect 19564 27716 19620 27718
rect 19644 27716 19700 27718
rect 19724 27716 19780 27718
rect 19484 26682 19540 26684
rect 19564 26682 19620 26684
rect 19644 26682 19700 26684
rect 19724 26682 19780 26684
rect 19484 26630 19510 26682
rect 19510 26630 19540 26682
rect 19564 26630 19574 26682
rect 19574 26630 19620 26682
rect 19644 26630 19690 26682
rect 19690 26630 19700 26682
rect 19724 26630 19754 26682
rect 19754 26630 19780 26682
rect 19484 26628 19540 26630
rect 19564 26628 19620 26630
rect 19644 26628 19700 26630
rect 19724 26628 19780 26630
rect 19484 25594 19540 25596
rect 19564 25594 19620 25596
rect 19644 25594 19700 25596
rect 19724 25594 19780 25596
rect 19484 25542 19510 25594
rect 19510 25542 19540 25594
rect 19564 25542 19574 25594
rect 19574 25542 19620 25594
rect 19644 25542 19690 25594
rect 19690 25542 19700 25594
rect 19724 25542 19754 25594
rect 19754 25542 19780 25594
rect 19484 25540 19540 25542
rect 19564 25540 19620 25542
rect 19644 25540 19700 25542
rect 19724 25540 19780 25542
rect 19484 24506 19540 24508
rect 19564 24506 19620 24508
rect 19644 24506 19700 24508
rect 19724 24506 19780 24508
rect 19484 24454 19510 24506
rect 19510 24454 19540 24506
rect 19564 24454 19574 24506
rect 19574 24454 19620 24506
rect 19644 24454 19690 24506
rect 19690 24454 19700 24506
rect 19724 24454 19754 24506
rect 19754 24454 19780 24506
rect 19484 24452 19540 24454
rect 19564 24452 19620 24454
rect 19644 24452 19700 24454
rect 19724 24452 19780 24454
rect 19484 23418 19540 23420
rect 19564 23418 19620 23420
rect 19644 23418 19700 23420
rect 19724 23418 19780 23420
rect 19484 23366 19510 23418
rect 19510 23366 19540 23418
rect 19564 23366 19574 23418
rect 19574 23366 19620 23418
rect 19644 23366 19690 23418
rect 19690 23366 19700 23418
rect 19724 23366 19754 23418
rect 19754 23366 19780 23418
rect 19484 23364 19540 23366
rect 19564 23364 19620 23366
rect 19644 23364 19700 23366
rect 19724 23364 19780 23366
rect 19484 22330 19540 22332
rect 19564 22330 19620 22332
rect 19644 22330 19700 22332
rect 19724 22330 19780 22332
rect 19484 22278 19510 22330
rect 19510 22278 19540 22330
rect 19564 22278 19574 22330
rect 19574 22278 19620 22330
rect 19644 22278 19690 22330
rect 19690 22278 19700 22330
rect 19724 22278 19754 22330
rect 19754 22278 19780 22330
rect 19484 22276 19540 22278
rect 19564 22276 19620 22278
rect 19644 22276 19700 22278
rect 19724 22276 19780 22278
rect 19484 21242 19540 21244
rect 19564 21242 19620 21244
rect 19644 21242 19700 21244
rect 19724 21242 19780 21244
rect 19484 21190 19510 21242
rect 19510 21190 19540 21242
rect 19564 21190 19574 21242
rect 19574 21190 19620 21242
rect 19644 21190 19690 21242
rect 19690 21190 19700 21242
rect 19724 21190 19754 21242
rect 19754 21190 19780 21242
rect 19484 21188 19540 21190
rect 19564 21188 19620 21190
rect 19644 21188 19700 21190
rect 19724 21188 19780 21190
rect 19484 20154 19540 20156
rect 19564 20154 19620 20156
rect 19644 20154 19700 20156
rect 19724 20154 19780 20156
rect 19484 20102 19510 20154
rect 19510 20102 19540 20154
rect 19564 20102 19574 20154
rect 19574 20102 19620 20154
rect 19644 20102 19690 20154
rect 19690 20102 19700 20154
rect 19724 20102 19754 20154
rect 19754 20102 19780 20154
rect 19484 20100 19540 20102
rect 19564 20100 19620 20102
rect 19644 20100 19700 20102
rect 19724 20100 19780 20102
rect 19484 19066 19540 19068
rect 19564 19066 19620 19068
rect 19644 19066 19700 19068
rect 19724 19066 19780 19068
rect 19484 19014 19510 19066
rect 19510 19014 19540 19066
rect 19564 19014 19574 19066
rect 19574 19014 19620 19066
rect 19644 19014 19690 19066
rect 19690 19014 19700 19066
rect 19724 19014 19754 19066
rect 19754 19014 19780 19066
rect 19484 19012 19540 19014
rect 19564 19012 19620 19014
rect 19644 19012 19700 19014
rect 19724 19012 19780 19014
rect 19484 17978 19540 17980
rect 19564 17978 19620 17980
rect 19644 17978 19700 17980
rect 19724 17978 19780 17980
rect 19484 17926 19510 17978
rect 19510 17926 19540 17978
rect 19564 17926 19574 17978
rect 19574 17926 19620 17978
rect 19644 17926 19690 17978
rect 19690 17926 19700 17978
rect 19724 17926 19754 17978
rect 19754 17926 19780 17978
rect 19484 17924 19540 17926
rect 19564 17924 19620 17926
rect 19644 17924 19700 17926
rect 19724 17924 19780 17926
rect 19484 16890 19540 16892
rect 19564 16890 19620 16892
rect 19644 16890 19700 16892
rect 19724 16890 19780 16892
rect 19484 16838 19510 16890
rect 19510 16838 19540 16890
rect 19564 16838 19574 16890
rect 19574 16838 19620 16890
rect 19644 16838 19690 16890
rect 19690 16838 19700 16890
rect 19724 16838 19754 16890
rect 19754 16838 19780 16890
rect 19484 16836 19540 16838
rect 19564 16836 19620 16838
rect 19644 16836 19700 16838
rect 19724 16836 19780 16838
rect 19484 15802 19540 15804
rect 19564 15802 19620 15804
rect 19644 15802 19700 15804
rect 19724 15802 19780 15804
rect 19484 15750 19510 15802
rect 19510 15750 19540 15802
rect 19564 15750 19574 15802
rect 19574 15750 19620 15802
rect 19644 15750 19690 15802
rect 19690 15750 19700 15802
rect 19724 15750 19754 15802
rect 19754 15750 19780 15802
rect 19484 15748 19540 15750
rect 19564 15748 19620 15750
rect 19644 15748 19700 15750
rect 19724 15748 19780 15750
rect 19154 13232 19210 13288
rect 19484 14714 19540 14716
rect 19564 14714 19620 14716
rect 19644 14714 19700 14716
rect 19724 14714 19780 14716
rect 19484 14662 19510 14714
rect 19510 14662 19540 14714
rect 19564 14662 19574 14714
rect 19574 14662 19620 14714
rect 19644 14662 19690 14714
rect 19690 14662 19700 14714
rect 19724 14662 19754 14714
rect 19754 14662 19780 14714
rect 19484 14660 19540 14662
rect 19564 14660 19620 14662
rect 19644 14660 19700 14662
rect 19724 14660 19780 14662
rect 19484 13626 19540 13628
rect 19564 13626 19620 13628
rect 19644 13626 19700 13628
rect 19724 13626 19780 13628
rect 19484 13574 19510 13626
rect 19510 13574 19540 13626
rect 19564 13574 19574 13626
rect 19574 13574 19620 13626
rect 19644 13574 19690 13626
rect 19690 13574 19700 13626
rect 19724 13574 19754 13626
rect 19754 13574 19780 13626
rect 19484 13572 19540 13574
rect 19564 13572 19620 13574
rect 19644 13572 19700 13574
rect 19724 13572 19780 13574
rect 19484 12538 19540 12540
rect 19564 12538 19620 12540
rect 19644 12538 19700 12540
rect 19724 12538 19780 12540
rect 19484 12486 19510 12538
rect 19510 12486 19540 12538
rect 19564 12486 19574 12538
rect 19574 12486 19620 12538
rect 19644 12486 19690 12538
rect 19690 12486 19700 12538
rect 19724 12486 19754 12538
rect 19754 12486 19780 12538
rect 19484 12484 19540 12486
rect 19564 12484 19620 12486
rect 19644 12484 19700 12486
rect 19724 12484 19780 12486
rect 18878 9424 18934 9480
rect 20350 30116 20406 30152
rect 20350 30096 20352 30116
rect 20352 30096 20404 30116
rect 20404 30096 20406 30116
rect 20074 28056 20130 28112
rect 20166 27784 20222 27840
rect 19484 11450 19540 11452
rect 19564 11450 19620 11452
rect 19644 11450 19700 11452
rect 19724 11450 19780 11452
rect 19484 11398 19510 11450
rect 19510 11398 19540 11450
rect 19564 11398 19574 11450
rect 19574 11398 19620 11450
rect 19644 11398 19690 11450
rect 19690 11398 19700 11450
rect 19724 11398 19754 11450
rect 19754 11398 19780 11450
rect 19484 11396 19540 11398
rect 19564 11396 19620 11398
rect 19644 11396 19700 11398
rect 19724 11396 19780 11398
rect 19484 10362 19540 10364
rect 19564 10362 19620 10364
rect 19644 10362 19700 10364
rect 19724 10362 19780 10364
rect 19484 10310 19510 10362
rect 19510 10310 19540 10362
rect 19564 10310 19574 10362
rect 19574 10310 19620 10362
rect 19644 10310 19690 10362
rect 19690 10310 19700 10362
rect 19724 10310 19754 10362
rect 19754 10310 19780 10362
rect 19484 10308 19540 10310
rect 19564 10308 19620 10310
rect 19644 10308 19700 10310
rect 19724 10308 19780 10310
rect 18970 8880 19026 8936
rect 19246 9832 19302 9888
rect 14852 2202 14908 2204
rect 14932 2202 14988 2204
rect 15012 2202 15068 2204
rect 15092 2202 15148 2204
rect 14852 2150 14878 2202
rect 14878 2150 14908 2202
rect 14932 2150 14942 2202
rect 14942 2150 14988 2202
rect 15012 2150 15058 2202
rect 15058 2150 15068 2202
rect 15092 2150 15122 2202
rect 15122 2150 15148 2202
rect 14852 2148 14908 2150
rect 14932 2148 14988 2150
rect 15012 2148 15068 2150
rect 15092 2148 15148 2150
rect 19484 9274 19540 9276
rect 19564 9274 19620 9276
rect 19644 9274 19700 9276
rect 19724 9274 19780 9276
rect 19484 9222 19510 9274
rect 19510 9222 19540 9274
rect 19564 9222 19574 9274
rect 19574 9222 19620 9274
rect 19644 9222 19690 9274
rect 19690 9222 19700 9274
rect 19724 9222 19754 9274
rect 19754 9222 19780 9274
rect 19484 9220 19540 9222
rect 19564 9220 19620 9222
rect 19644 9220 19700 9222
rect 19724 9220 19780 9222
rect 19484 8186 19540 8188
rect 19564 8186 19620 8188
rect 19644 8186 19700 8188
rect 19724 8186 19780 8188
rect 19484 8134 19510 8186
rect 19510 8134 19540 8186
rect 19564 8134 19574 8186
rect 19574 8134 19620 8186
rect 19644 8134 19690 8186
rect 19690 8134 19700 8186
rect 19724 8134 19754 8186
rect 19754 8134 19780 8186
rect 19484 8132 19540 8134
rect 19564 8132 19620 8134
rect 19644 8132 19700 8134
rect 19724 8132 19780 8134
rect 19484 7098 19540 7100
rect 19564 7098 19620 7100
rect 19644 7098 19700 7100
rect 19724 7098 19780 7100
rect 19484 7046 19510 7098
rect 19510 7046 19540 7098
rect 19564 7046 19574 7098
rect 19574 7046 19620 7098
rect 19644 7046 19690 7098
rect 19690 7046 19700 7098
rect 19724 7046 19754 7098
rect 19754 7046 19780 7098
rect 19484 7044 19540 7046
rect 19564 7044 19620 7046
rect 19644 7044 19700 7046
rect 19724 7044 19780 7046
rect 19484 6010 19540 6012
rect 19564 6010 19620 6012
rect 19644 6010 19700 6012
rect 19724 6010 19780 6012
rect 19484 5958 19510 6010
rect 19510 5958 19540 6010
rect 19564 5958 19574 6010
rect 19574 5958 19620 6010
rect 19644 5958 19690 6010
rect 19690 5958 19700 6010
rect 19724 5958 19754 6010
rect 19754 5958 19780 6010
rect 19484 5956 19540 5958
rect 19564 5956 19620 5958
rect 19644 5956 19700 5958
rect 19724 5956 19780 5958
rect 19484 4922 19540 4924
rect 19564 4922 19620 4924
rect 19644 4922 19700 4924
rect 19724 4922 19780 4924
rect 19484 4870 19510 4922
rect 19510 4870 19540 4922
rect 19564 4870 19574 4922
rect 19574 4870 19620 4922
rect 19644 4870 19690 4922
rect 19690 4870 19700 4922
rect 19724 4870 19754 4922
rect 19754 4870 19780 4922
rect 19484 4868 19540 4870
rect 19564 4868 19620 4870
rect 19644 4868 19700 4870
rect 19724 4868 19780 4870
rect 19484 3834 19540 3836
rect 19564 3834 19620 3836
rect 19644 3834 19700 3836
rect 19724 3834 19780 3836
rect 19484 3782 19510 3834
rect 19510 3782 19540 3834
rect 19564 3782 19574 3834
rect 19574 3782 19620 3834
rect 19644 3782 19690 3834
rect 19690 3782 19700 3834
rect 19724 3782 19754 3834
rect 19754 3782 19780 3834
rect 19484 3780 19540 3782
rect 19564 3780 19620 3782
rect 19644 3780 19700 3782
rect 19724 3780 19780 3782
rect 19484 2746 19540 2748
rect 19564 2746 19620 2748
rect 19644 2746 19700 2748
rect 19724 2746 19780 2748
rect 19484 2694 19510 2746
rect 19510 2694 19540 2746
rect 19564 2694 19574 2746
rect 19574 2694 19620 2746
rect 19644 2694 19690 2746
rect 19690 2694 19700 2746
rect 19724 2694 19754 2746
rect 19754 2694 19780 2746
rect 19484 2692 19540 2694
rect 19564 2692 19620 2694
rect 19644 2692 19700 2694
rect 19724 2692 19780 2694
rect 20258 12316 20260 12336
rect 20260 12316 20312 12336
rect 20312 12316 20314 12336
rect 20258 12280 20314 12316
rect 20994 35028 20996 35048
rect 20996 35028 21048 35048
rect 21048 35028 21050 35048
rect 20994 34992 21050 35028
rect 21086 31764 21088 31784
rect 21088 31764 21140 31784
rect 21140 31764 21142 31784
rect 21086 31728 21142 31764
rect 22466 51312 22522 51368
rect 25226 55664 25282 55720
rect 25134 54848 25190 54904
rect 25042 54032 25098 54088
rect 24116 53338 24172 53340
rect 24196 53338 24252 53340
rect 24276 53338 24332 53340
rect 24356 53338 24412 53340
rect 24116 53286 24142 53338
rect 24142 53286 24172 53338
rect 24196 53286 24206 53338
rect 24206 53286 24252 53338
rect 24276 53286 24322 53338
rect 24322 53286 24332 53338
rect 24356 53286 24386 53338
rect 24386 53286 24412 53338
rect 24116 53284 24172 53286
rect 24196 53284 24252 53286
rect 24276 53284 24332 53286
rect 24356 53284 24412 53286
rect 24858 53216 24914 53272
rect 20626 19216 20682 19272
rect 20902 18536 20958 18592
rect 21454 27512 21510 27568
rect 21730 30132 21732 30152
rect 21732 30132 21784 30152
rect 21784 30132 21786 30152
rect 21730 30096 21786 30132
rect 21730 18808 21786 18864
rect 21362 2796 21364 2816
rect 21364 2796 21416 2816
rect 21416 2796 21418 2816
rect 21362 2760 21418 2796
rect 22558 32272 22614 32328
rect 22650 32136 22706 32192
rect 23202 35808 23258 35864
rect 22742 18672 22798 18728
rect 23294 32408 23350 32464
rect 24116 52250 24172 52252
rect 24196 52250 24252 52252
rect 24276 52250 24332 52252
rect 24356 52250 24412 52252
rect 24116 52198 24142 52250
rect 24142 52198 24172 52250
rect 24196 52198 24206 52250
rect 24206 52198 24252 52250
rect 24276 52198 24322 52250
rect 24322 52198 24332 52250
rect 24356 52198 24386 52250
rect 24386 52198 24412 52250
rect 24116 52196 24172 52198
rect 24196 52196 24252 52198
rect 24276 52196 24332 52198
rect 24356 52196 24412 52198
rect 24674 52400 24730 52456
rect 24582 51992 24638 52048
rect 24116 51162 24172 51164
rect 24196 51162 24252 51164
rect 24276 51162 24332 51164
rect 24356 51162 24412 51164
rect 24116 51110 24142 51162
rect 24142 51110 24172 51162
rect 24196 51110 24206 51162
rect 24206 51110 24252 51162
rect 24276 51110 24322 51162
rect 24322 51110 24332 51162
rect 24356 51110 24386 51162
rect 24386 51110 24412 51162
rect 24116 51108 24172 51110
rect 24196 51108 24252 51110
rect 24276 51108 24332 51110
rect 24356 51108 24412 51110
rect 24858 52808 24914 52864
rect 25042 51584 25098 51640
rect 24950 50380 25006 50416
rect 24950 50360 24952 50380
rect 24952 50360 25004 50380
rect 25004 50360 25006 50380
rect 24116 50074 24172 50076
rect 24196 50074 24252 50076
rect 24276 50074 24332 50076
rect 24356 50074 24412 50076
rect 24116 50022 24142 50074
rect 24142 50022 24172 50074
rect 24196 50022 24206 50074
rect 24206 50022 24252 50074
rect 24276 50022 24322 50074
rect 24322 50022 24332 50074
rect 24356 50022 24386 50074
rect 24386 50022 24412 50074
rect 24116 50020 24172 50022
rect 24196 50020 24252 50022
rect 24276 50020 24332 50022
rect 24356 50020 24412 50022
rect 24116 48986 24172 48988
rect 24196 48986 24252 48988
rect 24276 48986 24332 48988
rect 24356 48986 24412 48988
rect 24116 48934 24142 48986
rect 24142 48934 24172 48986
rect 24196 48934 24206 48986
rect 24206 48934 24252 48986
rect 24276 48934 24322 48986
rect 24322 48934 24332 48986
rect 24356 48934 24386 48986
rect 24386 48934 24412 48986
rect 24116 48932 24172 48934
rect 24196 48932 24252 48934
rect 24276 48932 24332 48934
rect 24356 48932 24412 48934
rect 24116 47898 24172 47900
rect 24196 47898 24252 47900
rect 24276 47898 24332 47900
rect 24356 47898 24412 47900
rect 24116 47846 24142 47898
rect 24142 47846 24172 47898
rect 24196 47846 24206 47898
rect 24206 47846 24252 47898
rect 24276 47846 24322 47898
rect 24322 47846 24332 47898
rect 24356 47846 24386 47898
rect 24386 47846 24412 47898
rect 24116 47844 24172 47846
rect 24196 47844 24252 47846
rect 24276 47844 24332 47846
rect 24356 47844 24412 47846
rect 24116 46810 24172 46812
rect 24196 46810 24252 46812
rect 24276 46810 24332 46812
rect 24356 46810 24412 46812
rect 24116 46758 24142 46810
rect 24142 46758 24172 46810
rect 24196 46758 24206 46810
rect 24206 46758 24252 46810
rect 24276 46758 24322 46810
rect 24322 46758 24332 46810
rect 24356 46758 24386 46810
rect 24386 46758 24412 46810
rect 24116 46756 24172 46758
rect 24196 46756 24252 46758
rect 24276 46756 24332 46758
rect 24356 46756 24412 46758
rect 24116 45722 24172 45724
rect 24196 45722 24252 45724
rect 24276 45722 24332 45724
rect 24356 45722 24412 45724
rect 24116 45670 24142 45722
rect 24142 45670 24172 45722
rect 24196 45670 24206 45722
rect 24206 45670 24252 45722
rect 24276 45670 24322 45722
rect 24322 45670 24332 45722
rect 24356 45670 24386 45722
rect 24386 45670 24412 45722
rect 24116 45668 24172 45670
rect 24196 45668 24252 45670
rect 24276 45668 24332 45670
rect 24356 45668 24412 45670
rect 24116 44634 24172 44636
rect 24196 44634 24252 44636
rect 24276 44634 24332 44636
rect 24356 44634 24412 44636
rect 24116 44582 24142 44634
rect 24142 44582 24172 44634
rect 24196 44582 24206 44634
rect 24206 44582 24252 44634
rect 24276 44582 24322 44634
rect 24322 44582 24332 44634
rect 24356 44582 24386 44634
rect 24386 44582 24412 44634
rect 24116 44580 24172 44582
rect 24196 44580 24252 44582
rect 24276 44580 24332 44582
rect 24356 44580 24412 44582
rect 24116 43546 24172 43548
rect 24196 43546 24252 43548
rect 24276 43546 24332 43548
rect 24356 43546 24412 43548
rect 24116 43494 24142 43546
rect 24142 43494 24172 43546
rect 24196 43494 24206 43546
rect 24206 43494 24252 43546
rect 24276 43494 24322 43546
rect 24322 43494 24332 43546
rect 24356 43494 24386 43546
rect 24386 43494 24412 43546
rect 24116 43492 24172 43494
rect 24196 43492 24252 43494
rect 24276 43492 24332 43494
rect 24356 43492 24412 43494
rect 24116 42458 24172 42460
rect 24196 42458 24252 42460
rect 24276 42458 24332 42460
rect 24356 42458 24412 42460
rect 24116 42406 24142 42458
rect 24142 42406 24172 42458
rect 24196 42406 24206 42458
rect 24206 42406 24252 42458
rect 24276 42406 24322 42458
rect 24322 42406 24332 42458
rect 24356 42406 24386 42458
rect 24386 42406 24412 42458
rect 24116 42404 24172 42406
rect 24196 42404 24252 42406
rect 24276 42404 24332 42406
rect 24356 42404 24412 42406
rect 24116 41370 24172 41372
rect 24196 41370 24252 41372
rect 24276 41370 24332 41372
rect 24356 41370 24412 41372
rect 24116 41318 24142 41370
rect 24142 41318 24172 41370
rect 24196 41318 24206 41370
rect 24206 41318 24252 41370
rect 24276 41318 24322 41370
rect 24322 41318 24332 41370
rect 24356 41318 24386 41370
rect 24386 41318 24412 41370
rect 24116 41316 24172 41318
rect 24196 41316 24252 41318
rect 24276 41316 24332 41318
rect 24356 41316 24412 41318
rect 24116 40282 24172 40284
rect 24196 40282 24252 40284
rect 24276 40282 24332 40284
rect 24356 40282 24412 40284
rect 24116 40230 24142 40282
rect 24142 40230 24172 40282
rect 24196 40230 24206 40282
rect 24206 40230 24252 40282
rect 24276 40230 24322 40282
rect 24322 40230 24332 40282
rect 24356 40230 24386 40282
rect 24386 40230 24412 40282
rect 24116 40228 24172 40230
rect 24196 40228 24252 40230
rect 24276 40228 24332 40230
rect 24356 40228 24412 40230
rect 24116 39194 24172 39196
rect 24196 39194 24252 39196
rect 24276 39194 24332 39196
rect 24356 39194 24412 39196
rect 24116 39142 24142 39194
rect 24142 39142 24172 39194
rect 24196 39142 24206 39194
rect 24206 39142 24252 39194
rect 24276 39142 24322 39194
rect 24322 39142 24332 39194
rect 24356 39142 24386 39194
rect 24386 39142 24412 39194
rect 24116 39140 24172 39142
rect 24196 39140 24252 39142
rect 24276 39140 24332 39142
rect 24356 39140 24412 39142
rect 24116 38106 24172 38108
rect 24196 38106 24252 38108
rect 24276 38106 24332 38108
rect 24356 38106 24412 38108
rect 24116 38054 24142 38106
rect 24142 38054 24172 38106
rect 24196 38054 24206 38106
rect 24206 38054 24252 38106
rect 24276 38054 24322 38106
rect 24322 38054 24332 38106
rect 24356 38054 24386 38106
rect 24386 38054 24412 38106
rect 24116 38052 24172 38054
rect 24196 38052 24252 38054
rect 24276 38052 24332 38054
rect 24356 38052 24412 38054
rect 24116 37018 24172 37020
rect 24196 37018 24252 37020
rect 24276 37018 24332 37020
rect 24356 37018 24412 37020
rect 24116 36966 24142 37018
rect 24142 36966 24172 37018
rect 24196 36966 24206 37018
rect 24206 36966 24252 37018
rect 24276 36966 24322 37018
rect 24322 36966 24332 37018
rect 24356 36966 24386 37018
rect 24386 36966 24412 37018
rect 24116 36964 24172 36966
rect 24196 36964 24252 36966
rect 24276 36964 24332 36966
rect 24356 36964 24412 36966
rect 24116 35930 24172 35932
rect 24196 35930 24252 35932
rect 24276 35930 24332 35932
rect 24356 35930 24412 35932
rect 24116 35878 24142 35930
rect 24142 35878 24172 35930
rect 24196 35878 24206 35930
rect 24206 35878 24252 35930
rect 24276 35878 24322 35930
rect 24322 35878 24332 35930
rect 24356 35878 24386 35930
rect 24386 35878 24412 35930
rect 24116 35876 24172 35878
rect 24196 35876 24252 35878
rect 24276 35876 24332 35878
rect 24356 35876 24412 35878
rect 24116 34842 24172 34844
rect 24196 34842 24252 34844
rect 24276 34842 24332 34844
rect 24356 34842 24412 34844
rect 24116 34790 24142 34842
rect 24142 34790 24172 34842
rect 24196 34790 24206 34842
rect 24206 34790 24252 34842
rect 24276 34790 24322 34842
rect 24322 34790 24332 34842
rect 24356 34790 24386 34842
rect 24386 34790 24412 34842
rect 24116 34788 24172 34790
rect 24196 34788 24252 34790
rect 24276 34788 24332 34790
rect 24356 34788 24412 34790
rect 24858 43424 24914 43480
rect 24116 33754 24172 33756
rect 24196 33754 24252 33756
rect 24276 33754 24332 33756
rect 24356 33754 24412 33756
rect 24116 33702 24142 33754
rect 24142 33702 24172 33754
rect 24196 33702 24206 33754
rect 24206 33702 24252 33754
rect 24276 33702 24322 33754
rect 24322 33702 24332 33754
rect 24356 33702 24386 33754
rect 24386 33702 24412 33754
rect 24116 33700 24172 33702
rect 24196 33700 24252 33702
rect 24276 33700 24332 33702
rect 24356 33700 24412 33702
rect 23846 33532 23848 33552
rect 23848 33532 23900 33552
rect 23900 33532 23902 33552
rect 23846 33496 23902 33532
rect 23294 27648 23350 27704
rect 23570 27004 23572 27024
rect 23572 27004 23624 27024
rect 23624 27004 23626 27024
rect 23570 26968 23626 27004
rect 23478 22072 23534 22128
rect 23386 21936 23442 21992
rect 24490 32816 24546 32872
rect 24116 32666 24172 32668
rect 24196 32666 24252 32668
rect 24276 32666 24332 32668
rect 24356 32666 24412 32668
rect 24116 32614 24142 32666
rect 24142 32614 24172 32666
rect 24196 32614 24206 32666
rect 24206 32614 24252 32666
rect 24276 32614 24322 32666
rect 24322 32614 24332 32666
rect 24356 32614 24386 32666
rect 24386 32614 24412 32666
rect 24116 32612 24172 32614
rect 24196 32612 24252 32614
rect 24276 32612 24332 32614
rect 24356 32612 24412 32614
rect 24122 32272 24178 32328
rect 24398 31728 24454 31784
rect 24116 31578 24172 31580
rect 24196 31578 24252 31580
rect 24276 31578 24332 31580
rect 24356 31578 24412 31580
rect 24116 31526 24142 31578
rect 24142 31526 24172 31578
rect 24196 31526 24206 31578
rect 24206 31526 24252 31578
rect 24276 31526 24322 31578
rect 24322 31526 24332 31578
rect 24356 31526 24386 31578
rect 24386 31526 24412 31578
rect 24116 31524 24172 31526
rect 24196 31524 24252 31526
rect 24276 31524 24332 31526
rect 24356 31524 24412 31526
rect 23938 31220 23940 31240
rect 23940 31220 23992 31240
rect 23992 31220 23994 31240
rect 23938 31184 23994 31220
rect 24116 30490 24172 30492
rect 24196 30490 24252 30492
rect 24276 30490 24332 30492
rect 24356 30490 24412 30492
rect 24116 30438 24142 30490
rect 24142 30438 24172 30490
rect 24196 30438 24206 30490
rect 24206 30438 24252 30490
rect 24276 30438 24322 30490
rect 24322 30438 24332 30490
rect 24356 30438 24386 30490
rect 24386 30438 24412 30490
rect 24116 30436 24172 30438
rect 24196 30436 24252 30438
rect 24276 30436 24332 30438
rect 24356 30436 24412 30438
rect 24116 29402 24172 29404
rect 24196 29402 24252 29404
rect 24276 29402 24332 29404
rect 24356 29402 24412 29404
rect 24116 29350 24142 29402
rect 24142 29350 24172 29402
rect 24196 29350 24206 29402
rect 24206 29350 24252 29402
rect 24276 29350 24322 29402
rect 24322 29350 24332 29402
rect 24356 29350 24386 29402
rect 24386 29350 24412 29402
rect 24116 29348 24172 29350
rect 24196 29348 24252 29350
rect 24276 29348 24332 29350
rect 24356 29348 24412 29350
rect 24116 28314 24172 28316
rect 24196 28314 24252 28316
rect 24276 28314 24332 28316
rect 24356 28314 24412 28316
rect 24116 28262 24142 28314
rect 24142 28262 24172 28314
rect 24196 28262 24206 28314
rect 24206 28262 24252 28314
rect 24276 28262 24322 28314
rect 24322 28262 24332 28314
rect 24356 28262 24386 28314
rect 24386 28262 24412 28314
rect 24116 28260 24172 28262
rect 24196 28260 24252 28262
rect 24276 28260 24332 28262
rect 24356 28260 24412 28262
rect 24030 27956 24032 27976
rect 24032 27956 24084 27976
rect 24084 27956 24086 27976
rect 24030 27920 24086 27956
rect 23938 27512 23994 27568
rect 24116 27226 24172 27228
rect 24196 27226 24252 27228
rect 24276 27226 24332 27228
rect 24356 27226 24412 27228
rect 24116 27174 24142 27226
rect 24142 27174 24172 27226
rect 24196 27174 24206 27226
rect 24206 27174 24252 27226
rect 24276 27174 24322 27226
rect 24322 27174 24332 27226
rect 24356 27174 24386 27226
rect 24386 27174 24412 27226
rect 24116 27172 24172 27174
rect 24196 27172 24252 27174
rect 24276 27172 24332 27174
rect 24356 27172 24412 27174
rect 24116 26138 24172 26140
rect 24196 26138 24252 26140
rect 24276 26138 24332 26140
rect 24356 26138 24412 26140
rect 24116 26086 24142 26138
rect 24142 26086 24172 26138
rect 24196 26086 24206 26138
rect 24206 26086 24252 26138
rect 24276 26086 24322 26138
rect 24322 26086 24332 26138
rect 24356 26086 24386 26138
rect 24386 26086 24412 26138
rect 24116 26084 24172 26086
rect 24196 26084 24252 26086
rect 24276 26084 24332 26086
rect 24356 26084 24412 26086
rect 24116 25050 24172 25052
rect 24196 25050 24252 25052
rect 24276 25050 24332 25052
rect 24356 25050 24412 25052
rect 24116 24998 24142 25050
rect 24142 24998 24172 25050
rect 24196 24998 24206 25050
rect 24206 24998 24252 25050
rect 24276 24998 24322 25050
rect 24322 24998 24332 25050
rect 24356 24998 24386 25050
rect 24386 24998 24412 25050
rect 24116 24996 24172 24998
rect 24196 24996 24252 24998
rect 24276 24996 24332 24998
rect 24356 24996 24412 24998
rect 24116 23962 24172 23964
rect 24196 23962 24252 23964
rect 24276 23962 24332 23964
rect 24356 23962 24412 23964
rect 24116 23910 24142 23962
rect 24142 23910 24172 23962
rect 24196 23910 24206 23962
rect 24206 23910 24252 23962
rect 24276 23910 24322 23962
rect 24322 23910 24332 23962
rect 24356 23910 24386 23962
rect 24386 23910 24412 23962
rect 24116 23908 24172 23910
rect 24196 23908 24252 23910
rect 24276 23908 24332 23910
rect 24356 23908 24412 23910
rect 24116 22874 24172 22876
rect 24196 22874 24252 22876
rect 24276 22874 24332 22876
rect 24356 22874 24412 22876
rect 24116 22822 24142 22874
rect 24142 22822 24172 22874
rect 24196 22822 24206 22874
rect 24206 22822 24252 22874
rect 24276 22822 24322 22874
rect 24322 22822 24332 22874
rect 24356 22822 24386 22874
rect 24386 22822 24412 22874
rect 24116 22820 24172 22822
rect 24196 22820 24252 22822
rect 24276 22820 24332 22822
rect 24356 22820 24412 22822
rect 24122 21936 24178 21992
rect 24116 21786 24172 21788
rect 24196 21786 24252 21788
rect 24276 21786 24332 21788
rect 24356 21786 24412 21788
rect 24116 21734 24142 21786
rect 24142 21734 24172 21786
rect 24196 21734 24206 21786
rect 24206 21734 24252 21786
rect 24276 21734 24322 21786
rect 24322 21734 24332 21786
rect 24356 21734 24386 21786
rect 24386 21734 24412 21786
rect 24116 21732 24172 21734
rect 24196 21732 24252 21734
rect 24276 21732 24332 21734
rect 24356 21732 24412 21734
rect 24122 21528 24178 21584
rect 24116 20698 24172 20700
rect 24196 20698 24252 20700
rect 24276 20698 24332 20700
rect 24356 20698 24412 20700
rect 24116 20646 24142 20698
rect 24142 20646 24172 20698
rect 24196 20646 24206 20698
rect 24206 20646 24252 20698
rect 24276 20646 24322 20698
rect 24322 20646 24332 20698
rect 24356 20646 24386 20698
rect 24386 20646 24412 20698
rect 24116 20644 24172 20646
rect 24196 20644 24252 20646
rect 24276 20644 24332 20646
rect 24356 20644 24412 20646
rect 24116 19610 24172 19612
rect 24196 19610 24252 19612
rect 24276 19610 24332 19612
rect 24356 19610 24412 19612
rect 24116 19558 24142 19610
rect 24142 19558 24172 19610
rect 24196 19558 24206 19610
rect 24206 19558 24252 19610
rect 24276 19558 24322 19610
rect 24322 19558 24332 19610
rect 24356 19558 24386 19610
rect 24386 19558 24412 19610
rect 24116 19556 24172 19558
rect 24196 19556 24252 19558
rect 24276 19556 24332 19558
rect 24356 19556 24412 19558
rect 24214 19216 24270 19272
rect 24116 18522 24172 18524
rect 24196 18522 24252 18524
rect 24276 18522 24332 18524
rect 24356 18522 24412 18524
rect 24116 18470 24142 18522
rect 24142 18470 24172 18522
rect 24196 18470 24206 18522
rect 24206 18470 24252 18522
rect 24276 18470 24322 18522
rect 24322 18470 24332 18522
rect 24356 18470 24386 18522
rect 24386 18470 24412 18522
rect 24116 18468 24172 18470
rect 24196 18468 24252 18470
rect 24276 18468 24332 18470
rect 24356 18468 24412 18470
rect 24116 17434 24172 17436
rect 24196 17434 24252 17436
rect 24276 17434 24332 17436
rect 24356 17434 24412 17436
rect 24116 17382 24142 17434
rect 24142 17382 24172 17434
rect 24196 17382 24206 17434
rect 24206 17382 24252 17434
rect 24276 17382 24322 17434
rect 24322 17382 24332 17434
rect 24356 17382 24386 17434
rect 24386 17382 24412 17434
rect 24116 17380 24172 17382
rect 24196 17380 24252 17382
rect 24276 17380 24332 17382
rect 24356 17380 24412 17382
rect 24214 16532 24216 16552
rect 24216 16532 24268 16552
rect 24268 16532 24270 16552
rect 24214 16496 24270 16532
rect 24116 16346 24172 16348
rect 24196 16346 24252 16348
rect 24276 16346 24332 16348
rect 24356 16346 24412 16348
rect 24116 16294 24142 16346
rect 24142 16294 24172 16346
rect 24196 16294 24206 16346
rect 24206 16294 24252 16346
rect 24276 16294 24322 16346
rect 24322 16294 24332 16346
rect 24356 16294 24386 16346
rect 24386 16294 24412 16346
rect 24116 16292 24172 16294
rect 24196 16292 24252 16294
rect 24276 16292 24332 16294
rect 24356 16292 24412 16294
rect 24116 15258 24172 15260
rect 24196 15258 24252 15260
rect 24276 15258 24332 15260
rect 24356 15258 24412 15260
rect 24116 15206 24142 15258
rect 24142 15206 24172 15258
rect 24196 15206 24206 15258
rect 24206 15206 24252 15258
rect 24276 15206 24322 15258
rect 24322 15206 24332 15258
rect 24356 15206 24386 15258
rect 24386 15206 24412 15258
rect 24116 15204 24172 15206
rect 24196 15204 24252 15206
rect 24276 15204 24332 15206
rect 24356 15204 24412 15206
rect 24116 14170 24172 14172
rect 24196 14170 24252 14172
rect 24276 14170 24332 14172
rect 24356 14170 24412 14172
rect 24116 14118 24142 14170
rect 24142 14118 24172 14170
rect 24196 14118 24206 14170
rect 24206 14118 24252 14170
rect 24276 14118 24322 14170
rect 24322 14118 24332 14170
rect 24356 14118 24386 14170
rect 24386 14118 24412 14170
rect 24116 14116 24172 14118
rect 24196 14116 24252 14118
rect 24276 14116 24332 14118
rect 24356 14116 24412 14118
rect 24116 13082 24172 13084
rect 24196 13082 24252 13084
rect 24276 13082 24332 13084
rect 24356 13082 24412 13084
rect 24116 13030 24142 13082
rect 24142 13030 24172 13082
rect 24196 13030 24206 13082
rect 24206 13030 24252 13082
rect 24276 13030 24322 13082
rect 24322 13030 24332 13082
rect 24356 13030 24386 13082
rect 24386 13030 24412 13082
rect 24116 13028 24172 13030
rect 24196 13028 24252 13030
rect 24276 13028 24332 13030
rect 24356 13028 24412 13030
rect 24116 11994 24172 11996
rect 24196 11994 24252 11996
rect 24276 11994 24332 11996
rect 24356 11994 24412 11996
rect 24116 11942 24142 11994
rect 24142 11942 24172 11994
rect 24196 11942 24206 11994
rect 24206 11942 24252 11994
rect 24276 11942 24322 11994
rect 24322 11942 24332 11994
rect 24356 11942 24386 11994
rect 24386 11942 24412 11994
rect 24116 11940 24172 11942
rect 24196 11940 24252 11942
rect 24276 11940 24332 11942
rect 24356 11940 24412 11942
rect 24116 10906 24172 10908
rect 24196 10906 24252 10908
rect 24276 10906 24332 10908
rect 24356 10906 24412 10908
rect 24116 10854 24142 10906
rect 24142 10854 24172 10906
rect 24196 10854 24206 10906
rect 24206 10854 24252 10906
rect 24276 10854 24322 10906
rect 24322 10854 24332 10906
rect 24356 10854 24386 10906
rect 24386 10854 24412 10906
rect 24116 10852 24172 10854
rect 24196 10852 24252 10854
rect 24276 10852 24332 10854
rect 24356 10852 24412 10854
rect 24674 33360 24730 33416
rect 24858 33224 24914 33280
rect 25686 53644 25742 53680
rect 25686 53624 25688 53644
rect 25688 53624 25740 53644
rect 25740 53624 25742 53644
rect 25870 51312 25926 51368
rect 25778 51176 25834 51232
rect 25410 50768 25466 50824
rect 25594 49544 25650 49600
rect 27158 52944 27214 53000
rect 27618 51448 27674 51504
rect 28078 51856 28134 51912
rect 26054 49952 26110 50008
rect 26238 48728 26294 48784
rect 25594 47504 25650 47560
rect 25594 45464 25650 45520
rect 25502 41384 25558 41440
rect 25410 39752 25466 39808
rect 24950 31864 25006 31920
rect 24674 27784 24730 27840
rect 24858 27396 24914 27432
rect 24858 27376 24860 27396
rect 24860 27376 24912 27396
rect 24912 27376 24914 27396
rect 24950 25900 25006 25936
rect 24950 25880 24952 25900
rect 24952 25880 25004 25900
rect 25004 25880 25006 25900
rect 24950 18808 25006 18864
rect 25410 36488 25466 36544
rect 25318 33360 25374 33416
rect 25318 33088 25374 33144
rect 25226 31592 25282 31648
rect 25226 29008 25282 29064
rect 25410 32952 25466 33008
rect 25502 32000 25558 32056
rect 25410 31864 25466 31920
rect 25134 22616 25190 22672
rect 25962 45872 26018 45928
rect 26238 46688 26294 46744
rect 27342 50904 27398 50960
rect 26790 50632 26846 50688
rect 26698 49136 26754 49192
rect 28078 50224 28134 50280
rect 26974 48320 27030 48376
rect 26882 47912 26938 47968
rect 26698 47096 26754 47152
rect 26974 46280 27030 46336
rect 26238 45056 26294 45112
rect 26146 44240 26202 44296
rect 26974 44648 27030 44704
rect 27066 43832 27122 43888
rect 26146 42608 26202 42664
rect 26054 42200 26110 42256
rect 27158 43016 27214 43072
rect 26790 41792 26846 41848
rect 26146 41012 26148 41032
rect 26148 41012 26200 41032
rect 26200 41012 26202 41032
rect 26146 40976 26202 41012
rect 26790 40568 26846 40624
rect 26054 38936 26110 38992
rect 27434 40160 27490 40216
rect 27526 39344 27582 39400
rect 26882 38528 26938 38584
rect 26146 37712 26202 37768
rect 25870 36896 25926 36952
rect 26790 38120 26846 38176
rect 26882 37304 26938 37360
rect 26146 36080 26202 36136
rect 26790 35672 26846 35728
rect 26882 35264 26938 35320
rect 26054 34484 26056 34504
rect 26056 34484 26108 34504
rect 26108 34484 26110 34504
rect 26054 34448 26110 34484
rect 26146 34060 26202 34096
rect 26146 34040 26148 34060
rect 26148 34040 26200 34060
rect 26200 34040 26202 34060
rect 25778 32716 25780 32736
rect 25780 32716 25832 32736
rect 25832 32716 25834 32736
rect 25778 32680 25834 32716
rect 25778 32136 25834 32192
rect 25870 31184 25926 31240
rect 24950 16496 25006 16552
rect 21914 2916 21970 2952
rect 21914 2896 21916 2916
rect 21916 2896 21968 2916
rect 21968 2896 21970 2916
rect 22006 2760 22062 2816
rect 20350 2488 20406 2544
rect 24116 9818 24172 9820
rect 24196 9818 24252 9820
rect 24276 9818 24332 9820
rect 24356 9818 24412 9820
rect 24116 9766 24142 9818
rect 24142 9766 24172 9818
rect 24196 9766 24206 9818
rect 24206 9766 24252 9818
rect 24276 9766 24322 9818
rect 24322 9766 24332 9818
rect 24356 9766 24386 9818
rect 24386 9766 24412 9818
rect 24116 9764 24172 9766
rect 24196 9764 24252 9766
rect 24276 9764 24332 9766
rect 24356 9764 24412 9766
rect 24858 9560 24914 9616
rect 24116 8730 24172 8732
rect 24196 8730 24252 8732
rect 24276 8730 24332 8732
rect 24356 8730 24412 8732
rect 24116 8678 24142 8730
rect 24142 8678 24172 8730
rect 24196 8678 24206 8730
rect 24206 8678 24252 8730
rect 24276 8678 24322 8730
rect 24322 8678 24332 8730
rect 24356 8678 24386 8730
rect 24386 8678 24412 8730
rect 24116 8676 24172 8678
rect 24196 8676 24252 8678
rect 24276 8676 24332 8678
rect 24356 8676 24412 8678
rect 24116 7642 24172 7644
rect 24196 7642 24252 7644
rect 24276 7642 24332 7644
rect 24356 7642 24412 7644
rect 24116 7590 24142 7642
rect 24142 7590 24172 7642
rect 24196 7590 24206 7642
rect 24206 7590 24252 7642
rect 24276 7590 24322 7642
rect 24322 7590 24332 7642
rect 24356 7590 24386 7642
rect 24386 7590 24412 7642
rect 24116 7588 24172 7590
rect 24196 7588 24252 7590
rect 24276 7588 24332 7590
rect 24356 7588 24412 7590
rect 24116 6554 24172 6556
rect 24196 6554 24252 6556
rect 24276 6554 24332 6556
rect 24356 6554 24412 6556
rect 24116 6502 24142 6554
rect 24142 6502 24172 6554
rect 24196 6502 24206 6554
rect 24206 6502 24252 6554
rect 24276 6502 24322 6554
rect 24322 6502 24332 6554
rect 24356 6502 24386 6554
rect 24386 6502 24412 6554
rect 24116 6500 24172 6502
rect 24196 6500 24252 6502
rect 24276 6500 24332 6502
rect 24356 6500 24412 6502
rect 24950 8744 25006 8800
rect 25410 25472 25466 25528
rect 25686 30368 25742 30424
rect 25686 29164 25742 29200
rect 25686 29144 25688 29164
rect 25688 29144 25740 29164
rect 25740 29144 25742 29164
rect 25686 29008 25742 29064
rect 26330 33088 26386 33144
rect 26698 33632 26754 33688
rect 26054 31184 26110 31240
rect 26146 30776 26202 30832
rect 26146 29960 26202 30016
rect 26882 28736 26938 28792
rect 26422 28328 26478 28384
rect 26422 27920 26478 27976
rect 26330 27784 26386 27840
rect 26146 27512 26202 27568
rect 26238 27376 26294 27432
rect 26698 27648 26754 27704
rect 26790 27104 26846 27160
rect 26238 26968 26294 27024
rect 25226 16088 25282 16144
rect 25226 15580 25228 15600
rect 25228 15580 25280 15600
rect 25280 15580 25282 15600
rect 25226 15544 25282 15580
rect 24116 5466 24172 5468
rect 24196 5466 24252 5468
rect 24276 5466 24332 5468
rect 24356 5466 24412 5468
rect 24116 5414 24142 5466
rect 24142 5414 24172 5466
rect 24196 5414 24206 5466
rect 24206 5414 24252 5466
rect 24276 5414 24322 5466
rect 24322 5414 24332 5466
rect 24356 5414 24386 5466
rect 24386 5414 24412 5466
rect 24116 5412 24172 5414
rect 24196 5412 24252 5414
rect 24276 5412 24332 5414
rect 24356 5412 24412 5414
rect 24116 4378 24172 4380
rect 24196 4378 24252 4380
rect 24276 4378 24332 4380
rect 24356 4378 24412 4380
rect 24116 4326 24142 4378
rect 24142 4326 24172 4378
rect 24196 4326 24206 4378
rect 24206 4326 24252 4378
rect 24276 4326 24322 4378
rect 24322 4326 24332 4378
rect 24356 4326 24386 4378
rect 24386 4326 24412 4378
rect 24116 4324 24172 4326
rect 24196 4324 24252 4326
rect 24276 4324 24332 4326
rect 24356 4324 24412 4326
rect 24116 3290 24172 3292
rect 24196 3290 24252 3292
rect 24276 3290 24332 3292
rect 24356 3290 24412 3292
rect 24116 3238 24142 3290
rect 24142 3238 24172 3290
rect 24196 3238 24206 3290
rect 24206 3238 24252 3290
rect 24276 3238 24322 3290
rect 24322 3238 24332 3290
rect 24356 3238 24386 3290
rect 24386 3238 24412 3290
rect 24116 3236 24172 3238
rect 24196 3236 24252 3238
rect 24276 3236 24332 3238
rect 24356 3236 24412 3238
rect 24030 2896 24086 2952
rect 25410 16224 25466 16280
rect 26146 25064 26202 25120
rect 26146 24656 26202 24712
rect 26698 26732 26700 26752
rect 26700 26732 26752 26752
rect 26752 26732 26754 26752
rect 26698 26696 26754 26732
rect 25870 21800 25926 21856
rect 25594 18672 25650 18728
rect 25962 19352 26018 19408
rect 26790 23840 26846 23896
rect 26330 22208 26386 22264
rect 25870 18944 25926 19000
rect 25870 18808 25926 18864
rect 25962 18672 26018 18728
rect 26238 18536 26294 18592
rect 26882 21004 26938 21040
rect 26882 20984 26884 21004
rect 26884 20984 26936 21004
rect 26936 20984 26938 21004
rect 26698 18536 26754 18592
rect 26882 17740 26938 17776
rect 26882 17720 26884 17740
rect 26884 17720 26936 17740
rect 26936 17720 26938 17740
rect 26882 17332 26938 17368
rect 26882 17312 26884 17332
rect 26884 17312 26936 17332
rect 26936 17312 26938 17332
rect 26238 16088 26294 16144
rect 25962 15680 26018 15736
rect 25594 12416 25650 12472
rect 25962 12824 26018 12880
rect 26882 15272 26938 15328
rect 26146 11600 26202 11656
rect 26146 11212 26202 11248
rect 26146 11192 26148 11212
rect 26148 11192 26200 11212
rect 26200 11192 26202 11212
rect 25870 8372 25872 8392
rect 25872 8372 25924 8392
rect 25924 8372 25926 8392
rect 25870 8336 25926 8372
rect 26790 12008 26846 12064
rect 27342 34992 27398 35048
rect 27434 34856 27490 34912
rect 27986 33496 28042 33552
rect 27158 27920 27214 27976
rect 26146 9152 26202 9208
rect 26882 10376 26938 10432
rect 25318 6296 25374 6352
rect 24858 2624 24914 2680
rect 24490 2508 24546 2544
rect 24490 2488 24492 2508
rect 24492 2488 24544 2508
rect 24544 2488 24546 2508
rect 25042 2216 25098 2272
rect 24116 2202 24172 2204
rect 24196 2202 24252 2204
rect 24276 2202 24332 2204
rect 24356 2202 24412 2204
rect 24116 2150 24142 2202
rect 24142 2150 24172 2202
rect 24196 2150 24206 2202
rect 24206 2150 24252 2202
rect 24276 2150 24322 2202
rect 24322 2150 24332 2202
rect 24356 2150 24386 2202
rect 24386 2150 24412 2202
rect 24116 2148 24172 2150
rect 24196 2148 24252 2150
rect 24276 2148 24332 2150
rect 24356 2148 24412 2150
rect 25502 3032 25558 3088
rect 26790 7520 26846 7576
rect 26054 5908 26110 5944
rect 26054 5888 26056 5908
rect 26056 5888 26108 5908
rect 26108 5888 26110 5908
rect 26146 3576 26202 3632
rect 26606 5092 26662 5128
rect 26606 5072 26608 5092
rect 26608 5072 26660 5092
rect 26660 5072 26662 5092
rect 26882 5480 26938 5536
rect 27526 29552 27582 29608
rect 27526 24248 27582 24304
rect 28170 26308 28226 26344
rect 28170 26288 28172 26308
rect 28172 26288 28224 26308
rect 28224 26288 28226 26308
rect 28170 23432 28226 23488
rect 28170 23044 28226 23080
rect 28170 23024 28172 23044
rect 28172 23024 28224 23044
rect 28224 23024 28226 23044
rect 27526 21392 27582 21448
rect 28078 20576 28134 20632
rect 28170 20168 28226 20224
rect 28170 19780 28226 19816
rect 28170 19760 28172 19780
rect 28172 19760 28224 19780
rect 28224 19760 28226 19780
rect 27434 14728 27490 14784
rect 27526 14456 27582 14512
rect 27526 9968 27582 10024
rect 28170 18128 28226 18184
rect 28170 16904 28226 16960
rect 28170 16496 28226 16552
rect 28170 14048 28226 14104
rect 28170 13640 28226 13696
rect 28170 13252 28226 13288
rect 28170 13232 28172 13252
rect 28172 13232 28224 13252
rect 28224 13232 28226 13252
rect 28998 10784 29054 10840
rect 28078 7928 28134 7984
rect 26790 4256 26846 4312
rect 26790 2916 26846 2952
rect 26790 2896 26792 2916
rect 26792 2896 26844 2916
rect 26844 2896 26846 2916
rect 25410 1808 25466 1864
rect 25870 992 25926 1048
rect 2962 584 3018 640
rect 27434 4664 27490 4720
rect 28170 7112 28226 7168
rect 28170 6724 28226 6760
rect 28170 6704 28172 6724
rect 28172 6704 28224 6724
rect 28224 6704 28226 6724
rect 28078 3848 28134 3904
rect 28170 3460 28226 3496
rect 28170 3440 28172 3460
rect 28172 3440 28224 3460
rect 28224 3440 28226 3460
rect 26974 1400 27030 1456
rect 26146 584 26202 640
rect 26054 176 26110 232
<< metal3 >>
rect -800 55722 800 55752
rect 2773 55722 2839 55725
rect -800 55720 2839 55722
rect -800 55664 2778 55720
rect 2834 55664 2839 55720
rect -800 55662 2839 55664
rect -800 55632 800 55662
rect 2773 55659 2839 55662
rect 25221 55722 25287 55725
rect 29200 55722 30800 55752
rect 25221 55720 30800 55722
rect 25221 55664 25226 55720
rect 25282 55664 30800 55720
rect 25221 55662 30800 55664
rect 25221 55659 25287 55662
rect 29200 55632 30800 55662
rect -800 55314 800 55344
rect 3877 55314 3943 55317
rect -800 55312 3943 55314
rect -800 55256 3882 55312
rect 3938 55256 3943 55312
rect -800 55254 3943 55256
rect -800 55224 800 55254
rect 3877 55251 3943 55254
rect 23565 55314 23631 55317
rect 29200 55314 30800 55344
rect 23565 55312 30800 55314
rect 23565 55256 23570 55312
rect 23626 55256 30800 55312
rect 23565 55254 30800 55256
rect 23565 55251 23631 55254
rect 29200 55224 30800 55254
rect -800 54906 800 54936
rect 3233 54906 3299 54909
rect -800 54904 3299 54906
rect -800 54848 3238 54904
rect 3294 54848 3299 54904
rect -800 54846 3299 54848
rect -800 54816 800 54846
rect 3233 54843 3299 54846
rect 25129 54906 25195 54909
rect 29200 54906 30800 54936
rect 25129 54904 30800 54906
rect 25129 54848 25134 54904
rect 25190 54848 30800 54904
rect 25129 54846 30800 54848
rect 25129 54843 25195 54846
rect 29200 54816 30800 54846
rect -800 54498 800 54528
rect 3141 54498 3207 54501
rect -800 54496 3207 54498
rect -800 54440 3146 54496
rect 3202 54440 3207 54496
rect -800 54438 3207 54440
rect -800 54408 800 54438
rect 3141 54435 3207 54438
rect 20253 54498 20319 54501
rect 29200 54498 30800 54528
rect 20253 54496 30800 54498
rect 20253 54440 20258 54496
rect 20314 54440 30800 54496
rect 20253 54438 30800 54440
rect 20253 54435 20319 54438
rect 29200 54408 30800 54438
rect -800 54090 800 54120
rect 2957 54090 3023 54093
rect -800 54088 3023 54090
rect -800 54032 2962 54088
rect 3018 54032 3023 54088
rect -800 54030 3023 54032
rect -800 54000 800 54030
rect 2957 54027 3023 54030
rect 25037 54090 25103 54093
rect 29200 54090 30800 54120
rect 25037 54088 30800 54090
rect 25037 54032 25042 54088
rect 25098 54032 30800 54088
rect 25037 54030 30800 54032
rect 25037 54027 25103 54030
rect 29200 54000 30800 54030
rect -800 53682 800 53712
rect 4061 53682 4127 53685
rect -800 53680 4127 53682
rect -800 53624 4066 53680
rect 4122 53624 4127 53680
rect -800 53622 4127 53624
rect -800 53592 800 53622
rect 4061 53619 4127 53622
rect 25681 53682 25747 53685
rect 29200 53682 30800 53712
rect 25681 53680 30800 53682
rect 25681 53624 25686 53680
rect 25742 53624 30800 53680
rect 25681 53622 30800 53624
rect 25681 53619 25747 53622
rect 29200 53592 30800 53622
rect 5576 53344 5896 53345
rect -800 53274 800 53304
rect 5576 53280 5584 53344
rect 5648 53280 5664 53344
rect 5728 53280 5744 53344
rect 5808 53280 5824 53344
rect 5888 53280 5896 53344
rect 5576 53279 5896 53280
rect 14840 53344 15160 53345
rect 14840 53280 14848 53344
rect 14912 53280 14928 53344
rect 14992 53280 15008 53344
rect 15072 53280 15088 53344
rect 15152 53280 15160 53344
rect 14840 53279 15160 53280
rect 24104 53344 24424 53345
rect 24104 53280 24112 53344
rect 24176 53280 24192 53344
rect 24256 53280 24272 53344
rect 24336 53280 24352 53344
rect 24416 53280 24424 53344
rect 24104 53279 24424 53280
rect 3601 53274 3667 53277
rect -800 53272 3667 53274
rect -800 53216 3606 53272
rect 3662 53216 3667 53272
rect -800 53214 3667 53216
rect -800 53184 800 53214
rect 3601 53211 3667 53214
rect 24853 53274 24919 53277
rect 29200 53274 30800 53304
rect 24853 53272 30800 53274
rect 24853 53216 24858 53272
rect 24914 53216 30800 53272
rect 24853 53214 30800 53216
rect 24853 53211 24919 53214
rect 29200 53184 30800 53214
rect 5809 53002 5875 53005
rect 27153 53002 27219 53005
rect 5809 53000 27219 53002
rect 5809 52944 5814 53000
rect 5870 52944 27158 53000
rect 27214 52944 27219 53000
rect 5809 52942 27219 52944
rect 5809 52939 5875 52942
rect 27153 52939 27219 52942
rect -800 52866 800 52896
rect 3417 52866 3483 52869
rect -800 52864 3483 52866
rect -800 52808 3422 52864
rect 3478 52808 3483 52864
rect -800 52806 3483 52808
rect -800 52776 800 52806
rect 3417 52803 3483 52806
rect 24853 52866 24919 52869
rect 29200 52866 30800 52896
rect 24853 52864 30800 52866
rect 24853 52808 24858 52864
rect 24914 52808 30800 52864
rect 24853 52806 30800 52808
rect 24853 52803 24919 52806
rect 10208 52800 10528 52801
rect 10208 52736 10216 52800
rect 10280 52736 10296 52800
rect 10360 52736 10376 52800
rect 10440 52736 10456 52800
rect 10520 52736 10528 52800
rect 10208 52735 10528 52736
rect 19472 52800 19792 52801
rect 19472 52736 19480 52800
rect 19544 52736 19560 52800
rect 19624 52736 19640 52800
rect 19704 52736 19720 52800
rect 19784 52736 19792 52800
rect 29200 52776 30800 52806
rect 19472 52735 19792 52736
rect -800 52458 800 52488
rect 2773 52458 2839 52461
rect -800 52456 2839 52458
rect -800 52400 2778 52456
rect 2834 52400 2839 52456
rect -800 52398 2839 52400
rect -800 52368 800 52398
rect 2773 52395 2839 52398
rect 24669 52458 24735 52461
rect 29200 52458 30800 52488
rect 24669 52456 30800 52458
rect 24669 52400 24674 52456
rect 24730 52400 30800 52456
rect 24669 52398 30800 52400
rect 24669 52395 24735 52398
rect 29200 52368 30800 52398
rect 5576 52256 5896 52257
rect 5576 52192 5584 52256
rect 5648 52192 5664 52256
rect 5728 52192 5744 52256
rect 5808 52192 5824 52256
rect 5888 52192 5896 52256
rect 5576 52191 5896 52192
rect 14840 52256 15160 52257
rect 14840 52192 14848 52256
rect 14912 52192 14928 52256
rect 14992 52192 15008 52256
rect 15072 52192 15088 52256
rect 15152 52192 15160 52256
rect 14840 52191 15160 52192
rect 24104 52256 24424 52257
rect 24104 52192 24112 52256
rect 24176 52192 24192 52256
rect 24256 52192 24272 52256
rect 24336 52192 24352 52256
rect 24416 52192 24424 52256
rect 24104 52191 24424 52192
rect -800 52050 800 52080
rect 2773 52050 2839 52053
rect -800 52048 2839 52050
rect -800 51992 2778 52048
rect 2834 51992 2839 52048
rect -800 51990 2839 51992
rect -800 51960 800 51990
rect 2773 51987 2839 51990
rect 24577 52050 24643 52053
rect 29200 52050 30800 52080
rect 24577 52048 30800 52050
rect 24577 51992 24582 52048
rect 24638 51992 30800 52048
rect 24577 51990 30800 51992
rect 24577 51987 24643 51990
rect 29200 51960 30800 51990
rect 1853 51914 1919 51917
rect 28073 51914 28139 51917
rect 1853 51912 28139 51914
rect 1853 51856 1858 51912
rect 1914 51856 28078 51912
rect 28134 51856 28139 51912
rect 1853 51854 28139 51856
rect 1853 51851 1919 51854
rect 28073 51851 28139 51854
rect 10208 51712 10528 51713
rect -800 51642 800 51672
rect 10208 51648 10216 51712
rect 10280 51648 10296 51712
rect 10360 51648 10376 51712
rect 10440 51648 10456 51712
rect 10520 51648 10528 51712
rect 10208 51647 10528 51648
rect 19472 51712 19792 51713
rect 19472 51648 19480 51712
rect 19544 51648 19560 51712
rect 19624 51648 19640 51712
rect 19704 51648 19720 51712
rect 19784 51648 19792 51712
rect 19472 51647 19792 51648
rect 1945 51642 2011 51645
rect -800 51640 2011 51642
rect -800 51584 1950 51640
rect 2006 51584 2011 51640
rect -800 51582 2011 51584
rect -800 51552 800 51582
rect 1945 51579 2011 51582
rect 12709 51642 12775 51645
rect 15837 51642 15903 51645
rect 12709 51640 15903 51642
rect 12709 51584 12714 51640
rect 12770 51584 15842 51640
rect 15898 51584 15903 51640
rect 12709 51582 15903 51584
rect 12709 51579 12775 51582
rect 15837 51579 15903 51582
rect 25037 51642 25103 51645
rect 29200 51642 30800 51672
rect 25037 51640 30800 51642
rect 25037 51584 25042 51640
rect 25098 51584 30800 51640
rect 25037 51582 30800 51584
rect 25037 51579 25103 51582
rect 29200 51552 30800 51582
rect 3325 51506 3391 51509
rect 27613 51506 27679 51509
rect 3325 51504 27679 51506
rect 3325 51448 3330 51504
rect 3386 51448 27618 51504
rect 27674 51448 27679 51504
rect 3325 51446 27679 51448
rect 3325 51443 3391 51446
rect 27613 51443 27679 51446
rect 10777 51370 10843 51373
rect 13169 51370 13235 51373
rect 10777 51368 13235 51370
rect 10777 51312 10782 51368
rect 10838 51312 13174 51368
rect 13230 51312 13235 51368
rect 10777 51310 13235 51312
rect 10777 51307 10843 51310
rect 13169 51307 13235 51310
rect 22461 51370 22527 51373
rect 25865 51370 25931 51373
rect 22461 51368 25931 51370
rect 22461 51312 22466 51368
rect 22522 51312 25870 51368
rect 25926 51312 25931 51368
rect 22461 51310 25931 51312
rect 22461 51307 22527 51310
rect 25865 51307 25931 51310
rect -800 51234 800 51264
rect 2773 51234 2839 51237
rect -800 51232 2839 51234
rect -800 51176 2778 51232
rect 2834 51176 2839 51232
rect -800 51174 2839 51176
rect -800 51144 800 51174
rect 2773 51171 2839 51174
rect 12341 51234 12407 51237
rect 13905 51234 13971 51237
rect 12341 51232 13971 51234
rect 12341 51176 12346 51232
rect 12402 51176 13910 51232
rect 13966 51176 13971 51232
rect 12341 51174 13971 51176
rect 12341 51171 12407 51174
rect 13905 51171 13971 51174
rect 25773 51234 25839 51237
rect 29200 51234 30800 51264
rect 25773 51232 30800 51234
rect 25773 51176 25778 51232
rect 25834 51176 30800 51232
rect 25773 51174 30800 51176
rect 25773 51171 25839 51174
rect 5576 51168 5896 51169
rect 5576 51104 5584 51168
rect 5648 51104 5664 51168
rect 5728 51104 5744 51168
rect 5808 51104 5824 51168
rect 5888 51104 5896 51168
rect 5576 51103 5896 51104
rect 14840 51168 15160 51169
rect 14840 51104 14848 51168
rect 14912 51104 14928 51168
rect 14992 51104 15008 51168
rect 15072 51104 15088 51168
rect 15152 51104 15160 51168
rect 14840 51103 15160 51104
rect 24104 51168 24424 51169
rect 24104 51104 24112 51168
rect 24176 51104 24192 51168
rect 24256 51104 24272 51168
rect 24336 51104 24352 51168
rect 24416 51104 24424 51168
rect 29200 51144 30800 51174
rect 24104 51103 24424 51104
rect 2681 50962 2747 50965
rect 27337 50962 27403 50965
rect 2681 50960 27403 50962
rect 2681 50904 2686 50960
rect 2742 50904 27342 50960
rect 27398 50904 27403 50960
rect 2681 50902 27403 50904
rect 2681 50899 2747 50902
rect 27337 50899 27403 50902
rect -800 50826 800 50856
rect 1485 50826 1551 50829
rect -800 50824 1551 50826
rect -800 50768 1490 50824
rect 1546 50768 1551 50824
rect -800 50766 1551 50768
rect -800 50736 800 50766
rect 1485 50763 1551 50766
rect 2589 50826 2655 50829
rect 25405 50826 25471 50829
rect 29200 50826 30800 50856
rect 2589 50824 22110 50826
rect 2589 50768 2594 50824
rect 2650 50768 22110 50824
rect 2589 50766 22110 50768
rect 2589 50763 2655 50766
rect 22050 50690 22110 50766
rect 25405 50824 30800 50826
rect 25405 50768 25410 50824
rect 25466 50768 30800 50824
rect 25405 50766 30800 50768
rect 25405 50763 25471 50766
rect 29200 50736 30800 50766
rect 26785 50690 26851 50693
rect 22050 50688 26851 50690
rect 22050 50632 26790 50688
rect 26846 50632 26851 50688
rect 22050 50630 26851 50632
rect 26785 50627 26851 50630
rect 10208 50624 10528 50625
rect 10208 50560 10216 50624
rect 10280 50560 10296 50624
rect 10360 50560 10376 50624
rect 10440 50560 10456 50624
rect 10520 50560 10528 50624
rect 10208 50559 10528 50560
rect 19472 50624 19792 50625
rect 19472 50560 19480 50624
rect 19544 50560 19560 50624
rect 19624 50560 19640 50624
rect 19704 50560 19720 50624
rect 19784 50560 19792 50624
rect 19472 50559 19792 50560
rect -800 50418 800 50448
rect 1393 50418 1459 50421
rect -800 50416 1459 50418
rect -800 50360 1398 50416
rect 1454 50360 1459 50416
rect -800 50358 1459 50360
rect -800 50328 800 50358
rect 1393 50355 1459 50358
rect 24945 50418 25011 50421
rect 29200 50418 30800 50448
rect 24945 50416 30800 50418
rect 24945 50360 24950 50416
rect 25006 50360 30800 50416
rect 24945 50358 30800 50360
rect 24945 50355 25011 50358
rect 29200 50328 30800 50358
rect 1853 50282 1919 50285
rect 28073 50282 28139 50285
rect 1853 50280 28139 50282
rect 1853 50224 1858 50280
rect 1914 50224 28078 50280
rect 28134 50224 28139 50280
rect 1853 50222 28139 50224
rect 1853 50219 1919 50222
rect 28073 50219 28139 50222
rect 5576 50080 5896 50081
rect -800 50010 800 50040
rect 5576 50016 5584 50080
rect 5648 50016 5664 50080
rect 5728 50016 5744 50080
rect 5808 50016 5824 50080
rect 5888 50016 5896 50080
rect 5576 50015 5896 50016
rect 14840 50080 15160 50081
rect 14840 50016 14848 50080
rect 14912 50016 14928 50080
rect 14992 50016 15008 50080
rect 15072 50016 15088 50080
rect 15152 50016 15160 50080
rect 14840 50015 15160 50016
rect 24104 50080 24424 50081
rect 24104 50016 24112 50080
rect 24176 50016 24192 50080
rect 24256 50016 24272 50080
rect 24336 50016 24352 50080
rect 24416 50016 24424 50080
rect 24104 50015 24424 50016
rect 1945 50010 2011 50013
rect -800 50008 2011 50010
rect -800 49952 1950 50008
rect 2006 49952 2011 50008
rect -800 49950 2011 49952
rect -800 49920 800 49950
rect 1945 49947 2011 49950
rect 26049 50010 26115 50013
rect 29200 50010 30800 50040
rect 26049 50008 30800 50010
rect 26049 49952 26054 50008
rect 26110 49952 30800 50008
rect 26049 49950 30800 49952
rect 26049 49947 26115 49950
rect 29200 49920 30800 49950
rect -800 49602 800 49632
rect 2773 49602 2839 49605
rect -800 49600 2839 49602
rect -800 49544 2778 49600
rect 2834 49544 2839 49600
rect -800 49542 2839 49544
rect -800 49512 800 49542
rect 2773 49539 2839 49542
rect 25589 49602 25655 49605
rect 29200 49602 30800 49632
rect 25589 49600 30800 49602
rect 25589 49544 25594 49600
rect 25650 49544 30800 49600
rect 25589 49542 30800 49544
rect 25589 49539 25655 49542
rect 10208 49536 10528 49537
rect 10208 49472 10216 49536
rect 10280 49472 10296 49536
rect 10360 49472 10376 49536
rect 10440 49472 10456 49536
rect 10520 49472 10528 49536
rect 10208 49471 10528 49472
rect 19472 49536 19792 49537
rect 19472 49472 19480 49536
rect 19544 49472 19560 49536
rect 19624 49472 19640 49536
rect 19704 49472 19720 49536
rect 19784 49472 19792 49536
rect 29200 49512 30800 49542
rect 19472 49471 19792 49472
rect -800 49194 800 49224
rect 1393 49194 1459 49197
rect -800 49192 1459 49194
rect -800 49136 1398 49192
rect 1454 49136 1459 49192
rect -800 49134 1459 49136
rect -800 49104 800 49134
rect 1393 49131 1459 49134
rect 26693 49194 26759 49197
rect 29200 49194 30800 49224
rect 26693 49192 30800 49194
rect 26693 49136 26698 49192
rect 26754 49136 30800 49192
rect 26693 49134 30800 49136
rect 26693 49131 26759 49134
rect 29200 49104 30800 49134
rect 5576 48992 5896 48993
rect 5576 48928 5584 48992
rect 5648 48928 5664 48992
rect 5728 48928 5744 48992
rect 5808 48928 5824 48992
rect 5888 48928 5896 48992
rect 5576 48927 5896 48928
rect 14840 48992 15160 48993
rect 14840 48928 14848 48992
rect 14912 48928 14928 48992
rect 14992 48928 15008 48992
rect 15072 48928 15088 48992
rect 15152 48928 15160 48992
rect 14840 48927 15160 48928
rect 24104 48992 24424 48993
rect 24104 48928 24112 48992
rect 24176 48928 24192 48992
rect 24256 48928 24272 48992
rect 24336 48928 24352 48992
rect 24416 48928 24424 48992
rect 24104 48927 24424 48928
rect -800 48786 800 48816
rect 2865 48786 2931 48789
rect -800 48784 2931 48786
rect -800 48728 2870 48784
rect 2926 48728 2931 48784
rect -800 48726 2931 48728
rect -800 48696 800 48726
rect 2865 48723 2931 48726
rect 26233 48786 26299 48789
rect 29200 48786 30800 48816
rect 26233 48784 30800 48786
rect 26233 48728 26238 48784
rect 26294 48728 30800 48784
rect 26233 48726 30800 48728
rect 26233 48723 26299 48726
rect 29200 48696 30800 48726
rect 10208 48448 10528 48449
rect -800 48378 800 48408
rect 10208 48384 10216 48448
rect 10280 48384 10296 48448
rect 10360 48384 10376 48448
rect 10440 48384 10456 48448
rect 10520 48384 10528 48448
rect 10208 48383 10528 48384
rect 19472 48448 19792 48449
rect 19472 48384 19480 48448
rect 19544 48384 19560 48448
rect 19624 48384 19640 48448
rect 19704 48384 19720 48448
rect 19784 48384 19792 48448
rect 19472 48383 19792 48384
rect 2957 48378 3023 48381
rect -800 48376 3023 48378
rect -800 48320 2962 48376
rect 3018 48320 3023 48376
rect -800 48318 3023 48320
rect -800 48288 800 48318
rect 2957 48315 3023 48318
rect 26969 48378 27035 48381
rect 29200 48378 30800 48408
rect 26969 48376 30800 48378
rect 26969 48320 26974 48376
rect 27030 48320 30800 48376
rect 26969 48318 30800 48320
rect 26969 48315 27035 48318
rect 29200 48288 30800 48318
rect -800 47970 800 48000
rect 1945 47970 2011 47973
rect -800 47968 2011 47970
rect -800 47912 1950 47968
rect 2006 47912 2011 47968
rect -800 47910 2011 47912
rect -800 47880 800 47910
rect 1945 47907 2011 47910
rect 26877 47970 26943 47973
rect 29200 47970 30800 48000
rect 26877 47968 30800 47970
rect 26877 47912 26882 47968
rect 26938 47912 30800 47968
rect 26877 47910 30800 47912
rect 26877 47907 26943 47910
rect 5576 47904 5896 47905
rect 5576 47840 5584 47904
rect 5648 47840 5664 47904
rect 5728 47840 5744 47904
rect 5808 47840 5824 47904
rect 5888 47840 5896 47904
rect 5576 47839 5896 47840
rect 14840 47904 15160 47905
rect 14840 47840 14848 47904
rect 14912 47840 14928 47904
rect 14992 47840 15008 47904
rect 15072 47840 15088 47904
rect 15152 47840 15160 47904
rect 14840 47839 15160 47840
rect 24104 47904 24424 47905
rect 24104 47840 24112 47904
rect 24176 47840 24192 47904
rect 24256 47840 24272 47904
rect 24336 47840 24352 47904
rect 24416 47840 24424 47904
rect 29200 47880 30800 47910
rect 24104 47839 24424 47840
rect -800 47562 800 47592
rect 2773 47562 2839 47565
rect -800 47560 2839 47562
rect -800 47504 2778 47560
rect 2834 47504 2839 47560
rect -800 47502 2839 47504
rect -800 47472 800 47502
rect 2773 47499 2839 47502
rect 25589 47562 25655 47565
rect 29200 47562 30800 47592
rect 25589 47560 30800 47562
rect 25589 47504 25594 47560
rect 25650 47504 30800 47560
rect 25589 47502 30800 47504
rect 25589 47499 25655 47502
rect 29200 47472 30800 47502
rect 10208 47360 10528 47361
rect 10208 47296 10216 47360
rect 10280 47296 10296 47360
rect 10360 47296 10376 47360
rect 10440 47296 10456 47360
rect 10520 47296 10528 47360
rect 10208 47295 10528 47296
rect 19472 47360 19792 47361
rect 19472 47296 19480 47360
rect 19544 47296 19560 47360
rect 19624 47296 19640 47360
rect 19704 47296 19720 47360
rect 19784 47296 19792 47360
rect 19472 47295 19792 47296
rect -800 47154 800 47184
rect 3785 47154 3851 47157
rect -800 47152 3851 47154
rect -800 47096 3790 47152
rect 3846 47096 3851 47152
rect -800 47094 3851 47096
rect -800 47064 800 47094
rect 3785 47091 3851 47094
rect 26693 47154 26759 47157
rect 29200 47154 30800 47184
rect 26693 47152 30800 47154
rect 26693 47096 26698 47152
rect 26754 47096 30800 47152
rect 26693 47094 30800 47096
rect 26693 47091 26759 47094
rect 29200 47064 30800 47094
rect 5576 46816 5896 46817
rect -800 46746 800 46776
rect 5576 46752 5584 46816
rect 5648 46752 5664 46816
rect 5728 46752 5744 46816
rect 5808 46752 5824 46816
rect 5888 46752 5896 46816
rect 5576 46751 5896 46752
rect 14840 46816 15160 46817
rect 14840 46752 14848 46816
rect 14912 46752 14928 46816
rect 14992 46752 15008 46816
rect 15072 46752 15088 46816
rect 15152 46752 15160 46816
rect 14840 46751 15160 46752
rect 24104 46816 24424 46817
rect 24104 46752 24112 46816
rect 24176 46752 24192 46816
rect 24256 46752 24272 46816
rect 24336 46752 24352 46816
rect 24416 46752 24424 46816
rect 24104 46751 24424 46752
rect 3509 46746 3575 46749
rect -800 46744 3575 46746
rect -800 46688 3514 46744
rect 3570 46688 3575 46744
rect -800 46686 3575 46688
rect -800 46656 800 46686
rect 3509 46683 3575 46686
rect 26233 46746 26299 46749
rect 29200 46746 30800 46776
rect 26233 46744 30800 46746
rect 26233 46688 26238 46744
rect 26294 46688 30800 46744
rect 26233 46686 30800 46688
rect 26233 46683 26299 46686
rect 29200 46656 30800 46686
rect -800 46338 800 46368
rect 2865 46338 2931 46341
rect -800 46336 2931 46338
rect -800 46280 2870 46336
rect 2926 46280 2931 46336
rect -800 46278 2931 46280
rect -800 46248 800 46278
rect 2865 46275 2931 46278
rect 26969 46338 27035 46341
rect 29200 46338 30800 46368
rect 26969 46336 30800 46338
rect 26969 46280 26974 46336
rect 27030 46280 30800 46336
rect 26969 46278 30800 46280
rect 26969 46275 27035 46278
rect 10208 46272 10528 46273
rect 10208 46208 10216 46272
rect 10280 46208 10296 46272
rect 10360 46208 10376 46272
rect 10440 46208 10456 46272
rect 10520 46208 10528 46272
rect 10208 46207 10528 46208
rect 19472 46272 19792 46273
rect 19472 46208 19480 46272
rect 19544 46208 19560 46272
rect 19624 46208 19640 46272
rect 19704 46208 19720 46272
rect 19784 46208 19792 46272
rect 29200 46248 30800 46278
rect 19472 46207 19792 46208
rect -800 45930 800 45960
rect 3417 45930 3483 45933
rect -800 45928 3483 45930
rect -800 45872 3422 45928
rect 3478 45872 3483 45928
rect -800 45870 3483 45872
rect -800 45840 800 45870
rect 3417 45867 3483 45870
rect 25957 45930 26023 45933
rect 29200 45930 30800 45960
rect 25957 45928 30800 45930
rect 25957 45872 25962 45928
rect 26018 45872 30800 45928
rect 25957 45870 30800 45872
rect 25957 45867 26023 45870
rect 29200 45840 30800 45870
rect 5576 45728 5896 45729
rect 5576 45664 5584 45728
rect 5648 45664 5664 45728
rect 5728 45664 5744 45728
rect 5808 45664 5824 45728
rect 5888 45664 5896 45728
rect 5576 45663 5896 45664
rect 14840 45728 15160 45729
rect 14840 45664 14848 45728
rect 14912 45664 14928 45728
rect 14992 45664 15008 45728
rect 15072 45664 15088 45728
rect 15152 45664 15160 45728
rect 14840 45663 15160 45664
rect 24104 45728 24424 45729
rect 24104 45664 24112 45728
rect 24176 45664 24192 45728
rect 24256 45664 24272 45728
rect 24336 45664 24352 45728
rect 24416 45664 24424 45728
rect 24104 45663 24424 45664
rect -800 45522 800 45552
rect 1945 45522 2011 45525
rect -800 45520 2011 45522
rect -800 45464 1950 45520
rect 2006 45464 2011 45520
rect -800 45462 2011 45464
rect -800 45432 800 45462
rect 1945 45459 2011 45462
rect 25589 45522 25655 45525
rect 29200 45522 30800 45552
rect 25589 45520 30800 45522
rect 25589 45464 25594 45520
rect 25650 45464 30800 45520
rect 25589 45462 30800 45464
rect 25589 45459 25655 45462
rect 29200 45432 30800 45462
rect 10208 45184 10528 45185
rect -800 45114 800 45144
rect 10208 45120 10216 45184
rect 10280 45120 10296 45184
rect 10360 45120 10376 45184
rect 10440 45120 10456 45184
rect 10520 45120 10528 45184
rect 10208 45119 10528 45120
rect 19472 45184 19792 45185
rect 19472 45120 19480 45184
rect 19544 45120 19560 45184
rect 19624 45120 19640 45184
rect 19704 45120 19720 45184
rect 19784 45120 19792 45184
rect 19472 45119 19792 45120
rect 2957 45114 3023 45117
rect -800 45112 3023 45114
rect -800 45056 2962 45112
rect 3018 45056 3023 45112
rect -800 45054 3023 45056
rect -800 45024 800 45054
rect 2957 45051 3023 45054
rect 26233 45114 26299 45117
rect 29200 45114 30800 45144
rect 26233 45112 30800 45114
rect 26233 45056 26238 45112
rect 26294 45056 30800 45112
rect 26233 45054 30800 45056
rect 26233 45051 26299 45054
rect 29200 45024 30800 45054
rect -800 44706 800 44736
rect 2865 44706 2931 44709
rect -800 44704 2931 44706
rect -800 44648 2870 44704
rect 2926 44648 2931 44704
rect -800 44646 2931 44648
rect -800 44616 800 44646
rect 2865 44643 2931 44646
rect 26969 44706 27035 44709
rect 29200 44706 30800 44736
rect 26969 44704 30800 44706
rect 26969 44648 26974 44704
rect 27030 44648 30800 44704
rect 26969 44646 30800 44648
rect 26969 44643 27035 44646
rect 5576 44640 5896 44641
rect 5576 44576 5584 44640
rect 5648 44576 5664 44640
rect 5728 44576 5744 44640
rect 5808 44576 5824 44640
rect 5888 44576 5896 44640
rect 5576 44575 5896 44576
rect 14840 44640 15160 44641
rect 14840 44576 14848 44640
rect 14912 44576 14928 44640
rect 14992 44576 15008 44640
rect 15072 44576 15088 44640
rect 15152 44576 15160 44640
rect 14840 44575 15160 44576
rect 24104 44640 24424 44641
rect 24104 44576 24112 44640
rect 24176 44576 24192 44640
rect 24256 44576 24272 44640
rect 24336 44576 24352 44640
rect 24416 44576 24424 44640
rect 29200 44616 30800 44646
rect 24104 44575 24424 44576
rect -800 44298 800 44328
rect 2773 44298 2839 44301
rect -800 44296 2839 44298
rect -800 44240 2778 44296
rect 2834 44240 2839 44296
rect -800 44238 2839 44240
rect -800 44208 800 44238
rect 2773 44235 2839 44238
rect 26141 44298 26207 44301
rect 29200 44298 30800 44328
rect 26141 44296 30800 44298
rect 26141 44240 26146 44296
rect 26202 44240 30800 44296
rect 26141 44238 30800 44240
rect 26141 44235 26207 44238
rect 29200 44208 30800 44238
rect 10208 44096 10528 44097
rect 10208 44032 10216 44096
rect 10280 44032 10296 44096
rect 10360 44032 10376 44096
rect 10440 44032 10456 44096
rect 10520 44032 10528 44096
rect 10208 44031 10528 44032
rect 19472 44096 19792 44097
rect 19472 44032 19480 44096
rect 19544 44032 19560 44096
rect 19624 44032 19640 44096
rect 19704 44032 19720 44096
rect 19784 44032 19792 44096
rect 19472 44031 19792 44032
rect -800 43890 800 43920
rect 3417 43890 3483 43893
rect -800 43888 3483 43890
rect -800 43832 3422 43888
rect 3478 43832 3483 43888
rect -800 43830 3483 43832
rect -800 43800 800 43830
rect 3417 43827 3483 43830
rect 27061 43890 27127 43893
rect 29200 43890 30800 43920
rect 27061 43888 30800 43890
rect 27061 43832 27066 43888
rect 27122 43832 30800 43888
rect 27061 43830 30800 43832
rect 27061 43827 27127 43830
rect 29200 43800 30800 43830
rect 5576 43552 5896 43553
rect -800 43482 800 43512
rect 5576 43488 5584 43552
rect 5648 43488 5664 43552
rect 5728 43488 5744 43552
rect 5808 43488 5824 43552
rect 5888 43488 5896 43552
rect 5576 43487 5896 43488
rect 14840 43552 15160 43553
rect 14840 43488 14848 43552
rect 14912 43488 14928 43552
rect 14992 43488 15008 43552
rect 15072 43488 15088 43552
rect 15152 43488 15160 43552
rect 14840 43487 15160 43488
rect 24104 43552 24424 43553
rect 24104 43488 24112 43552
rect 24176 43488 24192 43552
rect 24256 43488 24272 43552
rect 24336 43488 24352 43552
rect 24416 43488 24424 43552
rect 24104 43487 24424 43488
rect 1945 43482 2011 43485
rect -800 43480 2011 43482
rect -800 43424 1950 43480
rect 2006 43424 2011 43480
rect -800 43422 2011 43424
rect -800 43392 800 43422
rect 1945 43419 2011 43422
rect 24853 43482 24919 43485
rect 29200 43482 30800 43512
rect 24853 43480 30800 43482
rect 24853 43424 24858 43480
rect 24914 43424 30800 43480
rect 24853 43422 30800 43424
rect 24853 43419 24919 43422
rect 29200 43392 30800 43422
rect -800 43074 800 43104
rect 2773 43074 2839 43077
rect -800 43072 2839 43074
rect -800 43016 2778 43072
rect 2834 43016 2839 43072
rect -800 43014 2839 43016
rect -800 42984 800 43014
rect 2773 43011 2839 43014
rect 27153 43074 27219 43077
rect 29200 43074 30800 43104
rect 27153 43072 30800 43074
rect 27153 43016 27158 43072
rect 27214 43016 30800 43072
rect 27153 43014 30800 43016
rect 27153 43011 27219 43014
rect 10208 43008 10528 43009
rect 10208 42944 10216 43008
rect 10280 42944 10296 43008
rect 10360 42944 10376 43008
rect 10440 42944 10456 43008
rect 10520 42944 10528 43008
rect 10208 42943 10528 42944
rect 19472 43008 19792 43009
rect 19472 42944 19480 43008
rect 19544 42944 19560 43008
rect 19624 42944 19640 43008
rect 19704 42944 19720 43008
rect 19784 42944 19792 43008
rect 29200 42984 30800 43014
rect 19472 42943 19792 42944
rect -800 42666 800 42696
rect 1301 42666 1367 42669
rect -800 42664 1367 42666
rect -800 42608 1306 42664
rect 1362 42608 1367 42664
rect -800 42606 1367 42608
rect -800 42576 800 42606
rect 1301 42603 1367 42606
rect 26141 42666 26207 42669
rect 29200 42666 30800 42696
rect 26141 42664 30800 42666
rect 26141 42608 26146 42664
rect 26202 42608 30800 42664
rect 26141 42606 30800 42608
rect 26141 42603 26207 42606
rect 29200 42576 30800 42606
rect 5576 42464 5896 42465
rect 5576 42400 5584 42464
rect 5648 42400 5664 42464
rect 5728 42400 5744 42464
rect 5808 42400 5824 42464
rect 5888 42400 5896 42464
rect 5576 42399 5896 42400
rect 14840 42464 15160 42465
rect 14840 42400 14848 42464
rect 14912 42400 14928 42464
rect 14992 42400 15008 42464
rect 15072 42400 15088 42464
rect 15152 42400 15160 42464
rect 14840 42399 15160 42400
rect 24104 42464 24424 42465
rect 24104 42400 24112 42464
rect 24176 42400 24192 42464
rect 24256 42400 24272 42464
rect 24336 42400 24352 42464
rect 24416 42400 24424 42464
rect 24104 42399 24424 42400
rect -800 42258 800 42288
rect 1393 42258 1459 42261
rect -800 42256 1459 42258
rect -800 42200 1398 42256
rect 1454 42200 1459 42256
rect -800 42198 1459 42200
rect -800 42168 800 42198
rect 1393 42195 1459 42198
rect 26049 42258 26115 42261
rect 29200 42258 30800 42288
rect 26049 42256 30800 42258
rect 26049 42200 26054 42256
rect 26110 42200 30800 42256
rect 26049 42198 30800 42200
rect 26049 42195 26115 42198
rect 29200 42168 30800 42198
rect 10208 41920 10528 41921
rect -800 41850 800 41880
rect 10208 41856 10216 41920
rect 10280 41856 10296 41920
rect 10360 41856 10376 41920
rect 10440 41856 10456 41920
rect 10520 41856 10528 41920
rect 10208 41855 10528 41856
rect 19472 41920 19792 41921
rect 19472 41856 19480 41920
rect 19544 41856 19560 41920
rect 19624 41856 19640 41920
rect 19704 41856 19720 41920
rect 19784 41856 19792 41920
rect 19472 41855 19792 41856
rect 2773 41850 2839 41853
rect -800 41848 2839 41850
rect -800 41792 2778 41848
rect 2834 41792 2839 41848
rect -800 41790 2839 41792
rect -800 41760 800 41790
rect 2773 41787 2839 41790
rect 26785 41850 26851 41853
rect 29200 41850 30800 41880
rect 26785 41848 30800 41850
rect 26785 41792 26790 41848
rect 26846 41792 30800 41848
rect 26785 41790 30800 41792
rect 26785 41787 26851 41790
rect 29200 41760 30800 41790
rect -800 41442 800 41472
rect 2957 41442 3023 41445
rect -800 41440 3023 41442
rect -800 41384 2962 41440
rect 3018 41384 3023 41440
rect -800 41382 3023 41384
rect -800 41352 800 41382
rect 2957 41379 3023 41382
rect 25497 41442 25563 41445
rect 29200 41442 30800 41472
rect 25497 41440 30800 41442
rect 25497 41384 25502 41440
rect 25558 41384 30800 41440
rect 25497 41382 30800 41384
rect 25497 41379 25563 41382
rect 5576 41376 5896 41377
rect 5576 41312 5584 41376
rect 5648 41312 5664 41376
rect 5728 41312 5744 41376
rect 5808 41312 5824 41376
rect 5888 41312 5896 41376
rect 5576 41311 5896 41312
rect 14840 41376 15160 41377
rect 14840 41312 14848 41376
rect 14912 41312 14928 41376
rect 14992 41312 15008 41376
rect 15072 41312 15088 41376
rect 15152 41312 15160 41376
rect 14840 41311 15160 41312
rect 24104 41376 24424 41377
rect 24104 41312 24112 41376
rect 24176 41312 24192 41376
rect 24256 41312 24272 41376
rect 24336 41312 24352 41376
rect 24416 41312 24424 41376
rect 29200 41352 30800 41382
rect 24104 41311 24424 41312
rect 5533 41170 5599 41173
rect 9213 41170 9279 41173
rect 5533 41168 9279 41170
rect 5533 41112 5538 41168
rect 5594 41112 9218 41168
rect 9274 41112 9279 41168
rect 5533 41110 9279 41112
rect 5533 41107 5599 41110
rect 9213 41107 9279 41110
rect -800 41034 800 41064
rect 1945 41034 2011 41037
rect -800 41032 2011 41034
rect -800 40976 1950 41032
rect 2006 40976 2011 41032
rect -800 40974 2011 40976
rect -800 40944 800 40974
rect 1945 40971 2011 40974
rect 26141 41034 26207 41037
rect 29200 41034 30800 41064
rect 26141 41032 30800 41034
rect 26141 40976 26146 41032
rect 26202 40976 30800 41032
rect 26141 40974 30800 40976
rect 26141 40971 26207 40974
rect 29200 40944 30800 40974
rect 10208 40832 10528 40833
rect 10208 40768 10216 40832
rect 10280 40768 10296 40832
rect 10360 40768 10376 40832
rect 10440 40768 10456 40832
rect 10520 40768 10528 40832
rect 10208 40767 10528 40768
rect 19472 40832 19792 40833
rect 19472 40768 19480 40832
rect 19544 40768 19560 40832
rect 19624 40768 19640 40832
rect 19704 40768 19720 40832
rect 19784 40768 19792 40832
rect 19472 40767 19792 40768
rect -800 40626 800 40656
rect 3141 40626 3207 40629
rect -800 40624 3207 40626
rect -800 40568 3146 40624
rect 3202 40568 3207 40624
rect -800 40566 3207 40568
rect -800 40536 800 40566
rect 3141 40563 3207 40566
rect 26785 40626 26851 40629
rect 29200 40626 30800 40656
rect 26785 40624 30800 40626
rect 26785 40568 26790 40624
rect 26846 40568 30800 40624
rect 26785 40566 30800 40568
rect 26785 40563 26851 40566
rect 29200 40536 30800 40566
rect 5576 40288 5896 40289
rect -800 40218 800 40248
rect 5576 40224 5584 40288
rect 5648 40224 5664 40288
rect 5728 40224 5744 40288
rect 5808 40224 5824 40288
rect 5888 40224 5896 40288
rect 5576 40223 5896 40224
rect 14840 40288 15160 40289
rect 14840 40224 14848 40288
rect 14912 40224 14928 40288
rect 14992 40224 15008 40288
rect 15072 40224 15088 40288
rect 15152 40224 15160 40288
rect 14840 40223 15160 40224
rect 24104 40288 24424 40289
rect 24104 40224 24112 40288
rect 24176 40224 24192 40288
rect 24256 40224 24272 40288
rect 24336 40224 24352 40288
rect 24416 40224 24424 40288
rect 24104 40223 24424 40224
rect 3785 40218 3851 40221
rect -800 40216 3851 40218
rect -800 40160 3790 40216
rect 3846 40160 3851 40216
rect -800 40158 3851 40160
rect -800 40128 800 40158
rect 3785 40155 3851 40158
rect 27429 40218 27495 40221
rect 29200 40218 30800 40248
rect 27429 40216 30800 40218
rect 27429 40160 27434 40216
rect 27490 40160 30800 40216
rect 27429 40158 30800 40160
rect 27429 40155 27495 40158
rect 29200 40128 30800 40158
rect -800 39810 800 39840
rect 3601 39810 3667 39813
rect -800 39808 3667 39810
rect -800 39752 3606 39808
rect 3662 39752 3667 39808
rect -800 39750 3667 39752
rect -800 39720 800 39750
rect 3601 39747 3667 39750
rect 25405 39810 25471 39813
rect 29200 39810 30800 39840
rect 25405 39808 30800 39810
rect 25405 39752 25410 39808
rect 25466 39752 30800 39808
rect 25405 39750 30800 39752
rect 25405 39747 25471 39750
rect 10208 39744 10528 39745
rect 10208 39680 10216 39744
rect 10280 39680 10296 39744
rect 10360 39680 10376 39744
rect 10440 39680 10456 39744
rect 10520 39680 10528 39744
rect 10208 39679 10528 39680
rect 19472 39744 19792 39745
rect 19472 39680 19480 39744
rect 19544 39680 19560 39744
rect 19624 39680 19640 39744
rect 19704 39680 19720 39744
rect 19784 39680 19792 39744
rect 29200 39720 30800 39750
rect 19472 39679 19792 39680
rect 10225 39538 10291 39541
rect 15837 39538 15903 39541
rect 10225 39536 15903 39538
rect 10225 39480 10230 39536
rect 10286 39480 15842 39536
rect 15898 39480 15903 39536
rect 10225 39478 15903 39480
rect 10225 39475 10291 39478
rect 15837 39475 15903 39478
rect -800 39402 800 39432
rect 2773 39402 2839 39405
rect -800 39400 2839 39402
rect -800 39344 2778 39400
rect 2834 39344 2839 39400
rect -800 39342 2839 39344
rect -800 39312 800 39342
rect 2773 39339 2839 39342
rect 10501 39402 10567 39405
rect 12525 39402 12591 39405
rect 15837 39402 15903 39405
rect 10501 39400 11070 39402
rect 10501 39344 10506 39400
rect 10562 39344 11070 39400
rect 10501 39342 11070 39344
rect 10501 39339 10567 39342
rect 11010 39266 11070 39342
rect 12525 39400 15903 39402
rect 12525 39344 12530 39400
rect 12586 39344 15842 39400
rect 15898 39344 15903 39400
rect 12525 39342 15903 39344
rect 12525 39339 12591 39342
rect 15837 39339 15903 39342
rect 27521 39402 27587 39405
rect 29200 39402 30800 39432
rect 27521 39400 30800 39402
rect 27521 39344 27526 39400
rect 27582 39344 30800 39400
rect 27521 39342 30800 39344
rect 27521 39339 27587 39342
rect 29200 39312 30800 39342
rect 11237 39266 11303 39269
rect 13445 39266 13511 39269
rect 11010 39264 13511 39266
rect 11010 39208 11242 39264
rect 11298 39208 13450 39264
rect 13506 39208 13511 39264
rect 11010 39206 13511 39208
rect 11237 39203 11303 39206
rect 13445 39203 13511 39206
rect 5576 39200 5896 39201
rect 5576 39136 5584 39200
rect 5648 39136 5664 39200
rect 5728 39136 5744 39200
rect 5808 39136 5824 39200
rect 5888 39136 5896 39200
rect 5576 39135 5896 39136
rect 14840 39200 15160 39201
rect 14840 39136 14848 39200
rect 14912 39136 14928 39200
rect 14992 39136 15008 39200
rect 15072 39136 15088 39200
rect 15152 39136 15160 39200
rect 14840 39135 15160 39136
rect 24104 39200 24424 39201
rect 24104 39136 24112 39200
rect 24176 39136 24192 39200
rect 24256 39136 24272 39200
rect 24336 39136 24352 39200
rect 24416 39136 24424 39200
rect 24104 39135 24424 39136
rect -800 38994 800 39024
rect 1945 38994 2011 38997
rect -800 38992 2011 38994
rect -800 38936 1950 38992
rect 2006 38936 2011 38992
rect -800 38934 2011 38936
rect -800 38904 800 38934
rect 1945 38931 2011 38934
rect 10501 38994 10567 38997
rect 11973 38994 12039 38997
rect 10501 38992 12039 38994
rect 10501 38936 10506 38992
rect 10562 38936 11978 38992
rect 12034 38936 12039 38992
rect 10501 38934 12039 38936
rect 10501 38931 10567 38934
rect 11973 38931 12039 38934
rect 26049 38994 26115 38997
rect 29200 38994 30800 39024
rect 26049 38992 30800 38994
rect 26049 38936 26054 38992
rect 26110 38936 30800 38992
rect 26049 38934 30800 38936
rect 26049 38931 26115 38934
rect 29200 38904 30800 38934
rect 10317 38858 10383 38861
rect 10685 38858 10751 38861
rect 10317 38856 10751 38858
rect 10317 38800 10322 38856
rect 10378 38800 10690 38856
rect 10746 38800 10751 38856
rect 10317 38798 10751 38800
rect 10317 38795 10383 38798
rect 10685 38795 10751 38798
rect 10869 38858 10935 38861
rect 11513 38858 11579 38861
rect 15469 38858 15535 38861
rect 10869 38856 15535 38858
rect 10869 38800 10874 38856
rect 10930 38800 11518 38856
rect 11574 38800 15474 38856
rect 15530 38800 15535 38856
rect 10869 38798 15535 38800
rect 10869 38795 10935 38798
rect 11513 38795 11579 38798
rect 15469 38795 15535 38798
rect 11237 38722 11303 38725
rect 11421 38722 11487 38725
rect 11237 38720 11487 38722
rect 11237 38664 11242 38720
rect 11298 38664 11426 38720
rect 11482 38664 11487 38720
rect 11237 38662 11487 38664
rect 11237 38659 11303 38662
rect 11421 38659 11487 38662
rect 16573 38722 16639 38725
rect 17861 38722 17927 38725
rect 16573 38720 17927 38722
rect 16573 38664 16578 38720
rect 16634 38664 17866 38720
rect 17922 38664 17927 38720
rect 16573 38662 17927 38664
rect 16573 38659 16639 38662
rect 17861 38659 17927 38662
rect 10208 38656 10528 38657
rect -800 38586 800 38616
rect 10208 38592 10216 38656
rect 10280 38592 10296 38656
rect 10360 38592 10376 38656
rect 10440 38592 10456 38656
rect 10520 38592 10528 38656
rect 10208 38591 10528 38592
rect 19472 38656 19792 38657
rect 19472 38592 19480 38656
rect 19544 38592 19560 38656
rect 19624 38592 19640 38656
rect 19704 38592 19720 38656
rect 19784 38592 19792 38656
rect 19472 38591 19792 38592
rect 2865 38586 2931 38589
rect -800 38584 2931 38586
rect -800 38528 2870 38584
rect 2926 38528 2931 38584
rect -800 38526 2931 38528
rect -800 38496 800 38526
rect 2865 38523 2931 38526
rect 10777 38584 10843 38589
rect 10777 38528 10782 38584
rect 10838 38528 10843 38584
rect 10777 38523 10843 38528
rect 26877 38586 26943 38589
rect 29200 38586 30800 38616
rect 26877 38584 30800 38586
rect 26877 38528 26882 38584
rect 26938 38528 30800 38584
rect 26877 38526 30800 38528
rect 26877 38523 26943 38526
rect 4889 38450 4955 38453
rect 6177 38450 6243 38453
rect 4889 38448 6243 38450
rect 4889 38392 4894 38448
rect 4950 38392 6182 38448
rect 6238 38392 6243 38448
rect 4889 38390 6243 38392
rect 4889 38387 4955 38390
rect 6177 38387 6243 38390
rect 10225 38450 10291 38453
rect 10780 38450 10840 38523
rect 29200 38496 30800 38526
rect 10225 38448 10840 38450
rect 10225 38392 10230 38448
rect 10286 38392 10840 38448
rect 10225 38390 10840 38392
rect 10225 38387 10291 38390
rect 2221 38314 2287 38317
rect 9397 38314 9463 38317
rect 2221 38312 9463 38314
rect 2221 38256 2226 38312
rect 2282 38256 9402 38312
rect 9458 38256 9463 38312
rect 2221 38254 9463 38256
rect 2221 38251 2287 38254
rect 9397 38251 9463 38254
rect 10501 38314 10567 38317
rect 11329 38314 11395 38317
rect 10501 38312 11395 38314
rect 10501 38256 10506 38312
rect 10562 38256 11334 38312
rect 11390 38256 11395 38312
rect 10501 38254 11395 38256
rect 10501 38251 10567 38254
rect 11329 38251 11395 38254
rect -800 38178 800 38208
rect 1393 38178 1459 38181
rect -800 38176 1459 38178
rect -800 38120 1398 38176
rect 1454 38120 1459 38176
rect -800 38118 1459 38120
rect -800 38088 800 38118
rect 1393 38115 1459 38118
rect 9213 38178 9279 38181
rect 11605 38178 11671 38181
rect 9213 38176 11671 38178
rect 9213 38120 9218 38176
rect 9274 38120 11610 38176
rect 11666 38120 11671 38176
rect 9213 38118 11671 38120
rect 9213 38115 9279 38118
rect 11605 38115 11671 38118
rect 26785 38178 26851 38181
rect 29200 38178 30800 38208
rect 26785 38176 30800 38178
rect 26785 38120 26790 38176
rect 26846 38120 30800 38176
rect 26785 38118 30800 38120
rect 26785 38115 26851 38118
rect 5576 38112 5896 38113
rect 5576 38048 5584 38112
rect 5648 38048 5664 38112
rect 5728 38048 5744 38112
rect 5808 38048 5824 38112
rect 5888 38048 5896 38112
rect 5576 38047 5896 38048
rect 14840 38112 15160 38113
rect 14840 38048 14848 38112
rect 14912 38048 14928 38112
rect 14992 38048 15008 38112
rect 15072 38048 15088 38112
rect 15152 38048 15160 38112
rect 14840 38047 15160 38048
rect 24104 38112 24424 38113
rect 24104 38048 24112 38112
rect 24176 38048 24192 38112
rect 24256 38048 24272 38112
rect 24336 38048 24352 38112
rect 24416 38048 24424 38112
rect 29200 38088 30800 38118
rect 24104 38047 24424 38048
rect -800 37770 800 37800
rect 2773 37770 2839 37773
rect -800 37768 2839 37770
rect -800 37712 2778 37768
rect 2834 37712 2839 37768
rect -800 37710 2839 37712
rect -800 37680 800 37710
rect 2773 37707 2839 37710
rect 26141 37770 26207 37773
rect 29200 37770 30800 37800
rect 26141 37768 30800 37770
rect 26141 37712 26146 37768
rect 26202 37712 30800 37768
rect 26141 37710 30800 37712
rect 26141 37707 26207 37710
rect 29200 37680 30800 37710
rect 10208 37568 10528 37569
rect 10208 37504 10216 37568
rect 10280 37504 10296 37568
rect 10360 37504 10376 37568
rect 10440 37504 10456 37568
rect 10520 37504 10528 37568
rect 10208 37503 10528 37504
rect 19472 37568 19792 37569
rect 19472 37504 19480 37568
rect 19544 37504 19560 37568
rect 19624 37504 19640 37568
rect 19704 37504 19720 37568
rect 19784 37504 19792 37568
rect 19472 37503 19792 37504
rect 12709 37498 12775 37501
rect 13721 37498 13787 37501
rect 12709 37496 13787 37498
rect 12709 37440 12714 37496
rect 12770 37440 13726 37496
rect 13782 37440 13787 37496
rect 12709 37438 13787 37440
rect 12709 37435 12775 37438
rect 13721 37435 13787 37438
rect -800 37362 800 37392
rect 2957 37362 3023 37365
rect -800 37360 3023 37362
rect -800 37304 2962 37360
rect 3018 37304 3023 37360
rect -800 37302 3023 37304
rect -800 37272 800 37302
rect 2957 37299 3023 37302
rect 12157 37362 12223 37365
rect 13445 37362 13511 37365
rect 13997 37362 14063 37365
rect 12157 37360 12450 37362
rect 12157 37304 12162 37360
rect 12218 37304 12450 37360
rect 12157 37302 12450 37304
rect 12157 37299 12223 37302
rect 12390 37293 12450 37302
rect 13445 37360 14063 37362
rect 13445 37304 13450 37360
rect 13506 37304 14002 37360
rect 14058 37304 14063 37360
rect 13445 37302 14063 37304
rect 13445 37299 13511 37302
rect 13997 37299 14063 37302
rect 26877 37362 26943 37365
rect 29200 37362 30800 37392
rect 26877 37360 30800 37362
rect 26877 37304 26882 37360
rect 26938 37304 30800 37360
rect 26877 37302 30800 37304
rect 26877 37299 26943 37302
rect 12390 37288 12499 37293
rect 12390 37232 12438 37288
rect 12494 37232 12499 37288
rect 29200 37272 30800 37302
rect 12390 37230 12499 37232
rect 12433 37227 12499 37230
rect 5576 37024 5896 37025
rect -800 36954 800 36984
rect 5576 36960 5584 37024
rect 5648 36960 5664 37024
rect 5728 36960 5744 37024
rect 5808 36960 5824 37024
rect 5888 36960 5896 37024
rect 5576 36959 5896 36960
rect 14840 37024 15160 37025
rect 14840 36960 14848 37024
rect 14912 36960 14928 37024
rect 14992 36960 15008 37024
rect 15072 36960 15088 37024
rect 15152 36960 15160 37024
rect 14840 36959 15160 36960
rect 24104 37024 24424 37025
rect 24104 36960 24112 37024
rect 24176 36960 24192 37024
rect 24256 36960 24272 37024
rect 24336 36960 24352 37024
rect 24416 36960 24424 37024
rect 24104 36959 24424 36960
rect 2773 36954 2839 36957
rect -800 36952 2839 36954
rect -800 36896 2778 36952
rect 2834 36896 2839 36952
rect -800 36894 2839 36896
rect -800 36864 800 36894
rect 2773 36891 2839 36894
rect 25865 36954 25931 36957
rect 29200 36954 30800 36984
rect 25865 36952 30800 36954
rect 25865 36896 25870 36952
rect 25926 36896 30800 36952
rect 25865 36894 30800 36896
rect 25865 36891 25931 36894
rect 29200 36864 30800 36894
rect -800 36546 800 36576
rect 1669 36546 1735 36549
rect -800 36544 1735 36546
rect -800 36488 1674 36544
rect 1730 36488 1735 36544
rect -800 36486 1735 36488
rect -800 36456 800 36486
rect 1669 36483 1735 36486
rect 25405 36546 25471 36549
rect 29200 36546 30800 36576
rect 25405 36544 30800 36546
rect 25405 36488 25410 36544
rect 25466 36488 30800 36544
rect 25405 36486 30800 36488
rect 25405 36483 25471 36486
rect 10208 36480 10528 36481
rect 10208 36416 10216 36480
rect 10280 36416 10296 36480
rect 10360 36416 10376 36480
rect 10440 36416 10456 36480
rect 10520 36416 10528 36480
rect 10208 36415 10528 36416
rect 19472 36480 19792 36481
rect 19472 36416 19480 36480
rect 19544 36416 19560 36480
rect 19624 36416 19640 36480
rect 19704 36416 19720 36480
rect 19784 36416 19792 36480
rect 29200 36456 30800 36486
rect 19472 36415 19792 36416
rect -800 36138 800 36168
rect 2773 36138 2839 36141
rect -800 36136 2839 36138
rect -800 36080 2778 36136
rect 2834 36080 2839 36136
rect -800 36078 2839 36080
rect -800 36048 800 36078
rect 2773 36075 2839 36078
rect 15469 36138 15535 36141
rect 15653 36138 15719 36141
rect 15469 36136 15719 36138
rect 15469 36080 15474 36136
rect 15530 36080 15658 36136
rect 15714 36080 15719 36136
rect 15469 36078 15719 36080
rect 15469 36075 15535 36078
rect 15653 36075 15719 36078
rect 26141 36138 26207 36141
rect 29200 36138 30800 36168
rect 26141 36136 30800 36138
rect 26141 36080 26146 36136
rect 26202 36080 30800 36136
rect 26141 36078 30800 36080
rect 26141 36075 26207 36078
rect 29200 36048 30800 36078
rect 5576 35936 5896 35937
rect 5576 35872 5584 35936
rect 5648 35872 5664 35936
rect 5728 35872 5744 35936
rect 5808 35872 5824 35936
rect 5888 35872 5896 35936
rect 5576 35871 5896 35872
rect 14840 35936 15160 35937
rect 14840 35872 14848 35936
rect 14912 35872 14928 35936
rect 14992 35872 15008 35936
rect 15072 35872 15088 35936
rect 15152 35872 15160 35936
rect 14840 35871 15160 35872
rect 24104 35936 24424 35937
rect 24104 35872 24112 35936
rect 24176 35872 24192 35936
rect 24256 35872 24272 35936
rect 24336 35872 24352 35936
rect 24416 35872 24424 35936
rect 24104 35871 24424 35872
rect 16021 35866 16087 35869
rect 23197 35866 23263 35869
rect 16021 35864 23263 35866
rect 16021 35808 16026 35864
rect 16082 35808 23202 35864
rect 23258 35808 23263 35864
rect 16021 35806 23263 35808
rect 16021 35803 16087 35806
rect 23197 35803 23263 35806
rect -800 35730 800 35760
rect 2865 35730 2931 35733
rect -800 35728 2931 35730
rect -800 35672 2870 35728
rect 2926 35672 2931 35728
rect -800 35670 2931 35672
rect -800 35640 800 35670
rect 2865 35667 2931 35670
rect 17401 35730 17467 35733
rect 18781 35730 18847 35733
rect 17401 35728 18847 35730
rect 17401 35672 17406 35728
rect 17462 35672 18786 35728
rect 18842 35672 18847 35728
rect 17401 35670 18847 35672
rect 17401 35667 17467 35670
rect 18781 35667 18847 35670
rect 26785 35730 26851 35733
rect 29200 35730 30800 35760
rect 26785 35728 30800 35730
rect 26785 35672 26790 35728
rect 26846 35672 30800 35728
rect 26785 35670 30800 35672
rect 26785 35667 26851 35670
rect 29200 35640 30800 35670
rect 10208 35392 10528 35393
rect -800 35322 800 35352
rect 10208 35328 10216 35392
rect 10280 35328 10296 35392
rect 10360 35328 10376 35392
rect 10440 35328 10456 35392
rect 10520 35328 10528 35392
rect 10208 35327 10528 35328
rect 19472 35392 19792 35393
rect 19472 35328 19480 35392
rect 19544 35328 19560 35392
rect 19624 35328 19640 35392
rect 19704 35328 19720 35392
rect 19784 35328 19792 35392
rect 19472 35327 19792 35328
rect 1945 35322 2011 35325
rect -800 35320 2011 35322
rect -800 35264 1950 35320
rect 2006 35264 2011 35320
rect -800 35262 2011 35264
rect -800 35232 800 35262
rect 1945 35259 2011 35262
rect 12525 35322 12591 35325
rect 26877 35322 26943 35325
rect 29200 35322 30800 35352
rect 12525 35320 12818 35322
rect 12525 35264 12530 35320
rect 12586 35264 12818 35320
rect 12525 35262 12818 35264
rect 12525 35259 12591 35262
rect 10409 35050 10475 35053
rect 12065 35050 12131 35053
rect 10409 35048 12131 35050
rect 10409 34992 10414 35048
rect 10470 34992 12070 35048
rect 12126 34992 12131 35048
rect 10409 34990 12131 34992
rect 10409 34987 10475 34990
rect 12065 34987 12131 34990
rect -800 34914 800 34944
rect 1669 34914 1735 34917
rect -800 34912 1735 34914
rect -800 34856 1674 34912
rect 1730 34856 1735 34912
rect -800 34854 1735 34856
rect -800 34824 800 34854
rect 1669 34851 1735 34854
rect 5576 34848 5896 34849
rect 5576 34784 5584 34848
rect 5648 34784 5664 34848
rect 5728 34784 5744 34848
rect 5808 34784 5824 34848
rect 5888 34784 5896 34848
rect 5576 34783 5896 34784
rect 4521 34642 4587 34645
rect 5533 34642 5599 34645
rect 4521 34640 5599 34642
rect 4521 34584 4526 34640
rect 4582 34584 5538 34640
rect 5594 34584 5599 34640
rect 4521 34582 5599 34584
rect 4521 34579 4587 34582
rect 5533 34579 5599 34582
rect -800 34506 800 34536
rect 2037 34506 2103 34509
rect -800 34504 2103 34506
rect -800 34448 2042 34504
rect 2098 34448 2103 34504
rect -800 34446 2103 34448
rect -800 34416 800 34446
rect 2037 34443 2103 34446
rect 10317 34506 10383 34509
rect 12758 34506 12818 35262
rect 26877 35320 30800 35322
rect 26877 35264 26882 35320
rect 26938 35264 30800 35320
rect 26877 35262 30800 35264
rect 26877 35259 26943 35262
rect 29200 35232 30800 35262
rect 13905 35050 13971 35053
rect 14825 35050 14891 35053
rect 13905 35048 14891 35050
rect 13905 34992 13910 35048
rect 13966 34992 14830 35048
rect 14886 34992 14891 35048
rect 13905 34990 14891 34992
rect 13905 34987 13971 34990
rect 14825 34987 14891 34990
rect 20989 35050 21055 35053
rect 27337 35050 27403 35053
rect 20989 35048 27403 35050
rect 20989 34992 20994 35048
rect 21050 34992 27342 35048
rect 27398 34992 27403 35048
rect 20989 34990 27403 34992
rect 20989 34987 21055 34990
rect 27337 34987 27403 34990
rect 27429 34914 27495 34917
rect 29200 34914 30800 34944
rect 27429 34912 30800 34914
rect 27429 34856 27434 34912
rect 27490 34856 30800 34912
rect 27429 34854 30800 34856
rect 27429 34851 27495 34854
rect 14840 34848 15160 34849
rect 14840 34784 14848 34848
rect 14912 34784 14928 34848
rect 14992 34784 15008 34848
rect 15072 34784 15088 34848
rect 15152 34784 15160 34848
rect 14840 34783 15160 34784
rect 24104 34848 24424 34849
rect 24104 34784 24112 34848
rect 24176 34784 24192 34848
rect 24256 34784 24272 34848
rect 24336 34784 24352 34848
rect 24416 34784 24424 34848
rect 29200 34824 30800 34854
rect 24104 34783 24424 34784
rect 18045 34642 18111 34645
rect 19149 34642 19215 34645
rect 18045 34640 19215 34642
rect 18045 34584 18050 34640
rect 18106 34584 19154 34640
rect 19210 34584 19215 34640
rect 18045 34582 19215 34584
rect 18045 34579 18111 34582
rect 19149 34579 19215 34582
rect 13721 34506 13787 34509
rect 10317 34504 10748 34506
rect 10317 34448 10322 34504
rect 10378 34448 10748 34504
rect 10317 34446 10748 34448
rect 12758 34504 13787 34506
rect 12758 34448 13726 34504
rect 13782 34448 13787 34504
rect 12758 34446 13787 34448
rect 10317 34443 10383 34446
rect 10688 34370 10748 34446
rect 13721 34443 13787 34446
rect 26049 34506 26115 34509
rect 29200 34506 30800 34536
rect 26049 34504 30800 34506
rect 26049 34448 26054 34504
rect 26110 34448 30800 34504
rect 26049 34446 30800 34448
rect 26049 34443 26115 34446
rect 29200 34416 30800 34446
rect 17953 34370 18019 34373
rect 10688 34368 18019 34370
rect 10688 34312 17958 34368
rect 18014 34312 18019 34368
rect 10688 34310 18019 34312
rect 17953 34307 18019 34310
rect 10208 34304 10528 34305
rect 10208 34240 10216 34304
rect 10280 34240 10296 34304
rect 10360 34240 10376 34304
rect 10440 34240 10456 34304
rect 10520 34240 10528 34304
rect 10208 34239 10528 34240
rect 19472 34304 19792 34305
rect 19472 34240 19480 34304
rect 19544 34240 19560 34304
rect 19624 34240 19640 34304
rect 19704 34240 19720 34304
rect 19784 34240 19792 34304
rect 19472 34239 19792 34240
rect -800 34098 800 34128
rect 2037 34098 2103 34101
rect -800 34096 2103 34098
rect -800 34040 2042 34096
rect 2098 34040 2103 34096
rect -800 34038 2103 34040
rect -800 34008 800 34038
rect 2037 34035 2103 34038
rect 26141 34098 26207 34101
rect 29200 34098 30800 34128
rect 26141 34096 30800 34098
rect 26141 34040 26146 34096
rect 26202 34040 30800 34096
rect 26141 34038 30800 34040
rect 26141 34035 26207 34038
rect 29200 34008 30800 34038
rect 5576 33760 5896 33761
rect -800 33690 800 33720
rect 5576 33696 5584 33760
rect 5648 33696 5664 33760
rect 5728 33696 5744 33760
rect 5808 33696 5824 33760
rect 5888 33696 5896 33760
rect 5576 33695 5896 33696
rect 14840 33760 15160 33761
rect 14840 33696 14848 33760
rect 14912 33696 14928 33760
rect 14992 33696 15008 33760
rect 15072 33696 15088 33760
rect 15152 33696 15160 33760
rect 14840 33695 15160 33696
rect 24104 33760 24424 33761
rect 24104 33696 24112 33760
rect 24176 33696 24192 33760
rect 24256 33696 24272 33760
rect 24336 33696 24352 33760
rect 24416 33696 24424 33760
rect 24104 33695 24424 33696
rect 1393 33690 1459 33693
rect -800 33688 1459 33690
rect -800 33632 1398 33688
rect 1454 33632 1459 33688
rect -800 33630 1459 33632
rect -800 33600 800 33630
rect 1393 33627 1459 33630
rect 26693 33690 26759 33693
rect 29200 33690 30800 33720
rect 26693 33688 30800 33690
rect 26693 33632 26698 33688
rect 26754 33632 30800 33688
rect 26693 33630 30800 33632
rect 26693 33627 26759 33630
rect 29200 33600 30800 33630
rect 23841 33554 23907 33557
rect 27981 33554 28047 33557
rect 23841 33552 28047 33554
rect 23841 33496 23846 33552
rect 23902 33496 27986 33552
rect 28042 33496 28047 33552
rect 23841 33494 28047 33496
rect 23841 33491 23907 33494
rect 27981 33491 28047 33494
rect 24669 33418 24735 33421
rect 25313 33418 25379 33421
rect 24669 33416 25379 33418
rect 24669 33360 24674 33416
rect 24730 33360 25318 33416
rect 25374 33360 25379 33416
rect 24669 33358 25379 33360
rect 24669 33355 24735 33358
rect 25313 33355 25379 33358
rect -800 33282 800 33312
rect 3601 33282 3667 33285
rect -800 33280 3667 33282
rect -800 33224 3606 33280
rect 3662 33224 3667 33280
rect -800 33222 3667 33224
rect -800 33192 800 33222
rect 3601 33219 3667 33222
rect 24853 33282 24919 33285
rect 29200 33282 30800 33312
rect 24853 33280 30800 33282
rect 24853 33224 24858 33280
rect 24914 33224 30800 33280
rect 24853 33222 30800 33224
rect 24853 33219 24919 33222
rect 10208 33216 10528 33217
rect 10208 33152 10216 33216
rect 10280 33152 10296 33216
rect 10360 33152 10376 33216
rect 10440 33152 10456 33216
rect 10520 33152 10528 33216
rect 10208 33151 10528 33152
rect 19472 33216 19792 33217
rect 19472 33152 19480 33216
rect 19544 33152 19560 33216
rect 19624 33152 19640 33216
rect 19704 33152 19720 33216
rect 19784 33152 19792 33216
rect 29200 33192 30800 33222
rect 19472 33151 19792 33152
rect 25313 33146 25379 33149
rect 26325 33146 26391 33149
rect 25313 33144 26391 33146
rect 25313 33088 25318 33144
rect 25374 33088 26330 33144
rect 26386 33088 26391 33144
rect 25313 33086 26391 33088
rect 25313 33083 25379 33086
rect 26325 33083 26391 33086
rect 25405 33010 25471 33013
rect 25405 33008 25514 33010
rect 25405 32952 25410 33008
rect 25466 32952 25514 33008
rect 25405 32947 25514 32952
rect -800 32874 800 32904
rect 4153 32874 4219 32877
rect -800 32872 4219 32874
rect -800 32816 4158 32872
rect 4214 32816 4219 32872
rect -800 32814 4219 32816
rect -800 32784 800 32814
rect 4153 32811 4219 32814
rect 24485 32874 24551 32877
rect 25454 32874 25514 32947
rect 29200 32874 30800 32904
rect 24485 32872 24778 32874
rect 24485 32816 24490 32872
rect 24546 32816 24778 32872
rect 24485 32814 24778 32816
rect 25454 32814 30800 32874
rect 24485 32811 24551 32814
rect 24718 32738 24778 32814
rect 29200 32784 30800 32814
rect 25773 32738 25839 32741
rect 24718 32736 25839 32738
rect 24718 32680 25778 32736
rect 25834 32680 25839 32736
rect 24718 32678 25839 32680
rect 25773 32675 25839 32678
rect 5576 32672 5896 32673
rect 5576 32608 5584 32672
rect 5648 32608 5664 32672
rect 5728 32608 5744 32672
rect 5808 32608 5824 32672
rect 5888 32608 5896 32672
rect 5576 32607 5896 32608
rect 14840 32672 15160 32673
rect 14840 32608 14848 32672
rect 14912 32608 14928 32672
rect 14992 32608 15008 32672
rect 15072 32608 15088 32672
rect 15152 32608 15160 32672
rect 14840 32607 15160 32608
rect 24104 32672 24424 32673
rect 24104 32608 24112 32672
rect 24176 32608 24192 32672
rect 24256 32608 24272 32672
rect 24336 32608 24352 32672
rect 24416 32608 24424 32672
rect 24104 32607 24424 32608
rect -800 32466 800 32496
rect 2773 32466 2839 32469
rect -800 32464 2839 32466
rect -800 32408 2778 32464
rect 2834 32408 2839 32464
rect -800 32406 2839 32408
rect -800 32376 800 32406
rect 2773 32403 2839 32406
rect 23289 32466 23355 32469
rect 29200 32466 30800 32496
rect 23289 32464 30800 32466
rect 23289 32408 23294 32464
rect 23350 32408 30800 32464
rect 23289 32406 30800 32408
rect 23289 32403 23355 32406
rect 29200 32376 30800 32406
rect 13721 32330 13787 32333
rect 13678 32328 13787 32330
rect 13678 32272 13726 32328
rect 13782 32272 13787 32328
rect 13678 32267 13787 32272
rect 22553 32330 22619 32333
rect 24117 32330 24183 32333
rect 22553 32328 24183 32330
rect 22553 32272 22558 32328
rect 22614 32272 24122 32328
rect 24178 32272 24183 32328
rect 22553 32270 24183 32272
rect 22553 32267 22619 32270
rect 24117 32267 24183 32270
rect 10208 32128 10528 32129
rect -800 32058 800 32088
rect 10208 32064 10216 32128
rect 10280 32064 10296 32128
rect 10360 32064 10376 32128
rect 10440 32064 10456 32128
rect 10520 32064 10528 32128
rect 10208 32063 10528 32064
rect 3049 32058 3115 32061
rect -800 32056 3115 32058
rect -800 32000 3054 32056
rect 3110 32000 3115 32056
rect -800 31998 3115 32000
rect -800 31968 800 31998
rect 3049 31995 3115 31998
rect 13537 31786 13603 31789
rect 13678 31786 13738 32267
rect 22645 32194 22711 32197
rect 25773 32194 25839 32197
rect 22645 32192 25839 32194
rect 22645 32136 22650 32192
rect 22706 32136 25778 32192
rect 25834 32136 25839 32192
rect 22645 32134 25839 32136
rect 22645 32131 22711 32134
rect 25773 32131 25839 32134
rect 19472 32128 19792 32129
rect 19472 32064 19480 32128
rect 19544 32064 19560 32128
rect 19624 32064 19640 32128
rect 19704 32064 19720 32128
rect 19784 32064 19792 32128
rect 19472 32063 19792 32064
rect 16113 32058 16179 32061
rect 18781 32058 18847 32061
rect 16113 32056 18847 32058
rect 16113 32000 16118 32056
rect 16174 32000 18786 32056
rect 18842 32000 18847 32056
rect 16113 31998 18847 32000
rect 16113 31995 16179 31998
rect 18781 31995 18847 31998
rect 25497 32058 25563 32061
rect 29200 32058 30800 32088
rect 25497 32056 30800 32058
rect 25497 32000 25502 32056
rect 25558 32000 30800 32056
rect 25497 31998 30800 32000
rect 25497 31995 25563 31998
rect 29200 31968 30800 31998
rect 16481 31922 16547 31925
rect 16254 31920 16547 31922
rect 16254 31864 16486 31920
rect 16542 31864 16547 31920
rect 16254 31862 16547 31864
rect 16254 31789 16314 31862
rect 16481 31859 16547 31862
rect 24945 31922 25011 31925
rect 25405 31922 25471 31925
rect 24945 31920 25471 31922
rect 24945 31864 24950 31920
rect 25006 31864 25410 31920
rect 25466 31864 25471 31920
rect 24945 31862 25471 31864
rect 24945 31859 25011 31862
rect 25405 31859 25471 31862
rect 13537 31784 13738 31786
rect 13537 31728 13542 31784
rect 13598 31728 13738 31784
rect 13537 31726 13738 31728
rect 16205 31784 16314 31789
rect 16205 31728 16210 31784
rect 16266 31728 16314 31784
rect 16205 31726 16314 31728
rect 21081 31786 21147 31789
rect 24393 31786 24459 31789
rect 21081 31784 24459 31786
rect 21081 31728 21086 31784
rect 21142 31728 24398 31784
rect 24454 31728 24459 31784
rect 21081 31726 24459 31728
rect 13537 31723 13603 31726
rect 16205 31723 16271 31726
rect 21081 31723 21147 31726
rect 24393 31723 24459 31726
rect -800 31650 800 31680
rect 4061 31650 4127 31653
rect -800 31648 4127 31650
rect -800 31592 4066 31648
rect 4122 31592 4127 31648
rect -800 31590 4127 31592
rect -800 31560 800 31590
rect 4061 31587 4127 31590
rect 25221 31650 25287 31653
rect 29200 31650 30800 31680
rect 25221 31648 30800 31650
rect 25221 31592 25226 31648
rect 25282 31592 30800 31648
rect 25221 31590 30800 31592
rect 25221 31587 25287 31590
rect 5576 31584 5896 31585
rect 5576 31520 5584 31584
rect 5648 31520 5664 31584
rect 5728 31520 5744 31584
rect 5808 31520 5824 31584
rect 5888 31520 5896 31584
rect 5576 31519 5896 31520
rect 14840 31584 15160 31585
rect 14840 31520 14848 31584
rect 14912 31520 14928 31584
rect 14992 31520 15008 31584
rect 15072 31520 15088 31584
rect 15152 31520 15160 31584
rect 14840 31519 15160 31520
rect 24104 31584 24424 31585
rect 24104 31520 24112 31584
rect 24176 31520 24192 31584
rect 24256 31520 24272 31584
rect 24336 31520 24352 31584
rect 24416 31520 24424 31584
rect 29200 31560 30800 31590
rect 24104 31519 24424 31520
rect 15101 31378 15167 31381
rect 15469 31378 15535 31381
rect 15101 31376 15535 31378
rect 15101 31320 15106 31376
rect 15162 31320 15474 31376
rect 15530 31320 15535 31376
rect 15101 31318 15535 31320
rect 15101 31315 15167 31318
rect 15469 31315 15535 31318
rect -800 31242 800 31272
rect 3785 31242 3851 31245
rect -800 31240 3851 31242
rect -800 31184 3790 31240
rect 3846 31184 3851 31240
rect -800 31182 3851 31184
rect -800 31152 800 31182
rect 3785 31179 3851 31182
rect 12801 31242 12867 31245
rect 18873 31242 18939 31245
rect 12801 31240 18939 31242
rect 12801 31184 12806 31240
rect 12862 31184 18878 31240
rect 18934 31184 18939 31240
rect 12801 31182 18939 31184
rect 12801 31179 12867 31182
rect 18873 31179 18939 31182
rect 23933 31242 23999 31245
rect 25865 31242 25931 31245
rect 23933 31240 25931 31242
rect 23933 31184 23938 31240
rect 23994 31184 25870 31240
rect 25926 31184 25931 31240
rect 23933 31182 25931 31184
rect 23933 31179 23999 31182
rect 25865 31179 25931 31182
rect 26049 31242 26115 31245
rect 29200 31242 30800 31272
rect 26049 31240 30800 31242
rect 26049 31184 26054 31240
rect 26110 31184 30800 31240
rect 26049 31182 30800 31184
rect 26049 31179 26115 31182
rect 29200 31152 30800 31182
rect 10208 31040 10528 31041
rect 10208 30976 10216 31040
rect 10280 30976 10296 31040
rect 10360 30976 10376 31040
rect 10440 30976 10456 31040
rect 10520 30976 10528 31040
rect 10208 30975 10528 30976
rect 19472 31040 19792 31041
rect 19472 30976 19480 31040
rect 19544 30976 19560 31040
rect 19624 30976 19640 31040
rect 19704 30976 19720 31040
rect 19784 30976 19792 31040
rect 19472 30975 19792 30976
rect -800 30834 800 30864
rect 3233 30834 3299 30837
rect -800 30832 3299 30834
rect -800 30776 3238 30832
rect 3294 30776 3299 30832
rect -800 30774 3299 30776
rect -800 30744 800 30774
rect 3233 30771 3299 30774
rect 12341 30834 12407 30837
rect 15469 30834 15535 30837
rect 17033 30834 17099 30837
rect 12341 30832 17099 30834
rect 12341 30776 12346 30832
rect 12402 30776 15474 30832
rect 15530 30776 17038 30832
rect 17094 30776 17099 30832
rect 12341 30774 17099 30776
rect 12341 30771 12407 30774
rect 15469 30771 15535 30774
rect 17033 30771 17099 30774
rect 26141 30834 26207 30837
rect 29200 30834 30800 30864
rect 26141 30832 30800 30834
rect 26141 30776 26146 30832
rect 26202 30776 30800 30832
rect 26141 30774 30800 30776
rect 26141 30771 26207 30774
rect 29200 30744 30800 30774
rect 5576 30496 5896 30497
rect -800 30426 800 30456
rect 5576 30432 5584 30496
rect 5648 30432 5664 30496
rect 5728 30432 5744 30496
rect 5808 30432 5824 30496
rect 5888 30432 5896 30496
rect 5576 30431 5896 30432
rect 14840 30496 15160 30497
rect 14840 30432 14848 30496
rect 14912 30432 14928 30496
rect 14992 30432 15008 30496
rect 15072 30432 15088 30496
rect 15152 30432 15160 30496
rect 14840 30431 15160 30432
rect 24104 30496 24424 30497
rect 24104 30432 24112 30496
rect 24176 30432 24192 30496
rect 24256 30432 24272 30496
rect 24336 30432 24352 30496
rect 24416 30432 24424 30496
rect 24104 30431 24424 30432
rect 1393 30426 1459 30429
rect -800 30424 1459 30426
rect -800 30368 1398 30424
rect 1454 30368 1459 30424
rect -800 30366 1459 30368
rect -800 30336 800 30366
rect 1393 30363 1459 30366
rect 25681 30426 25747 30429
rect 29200 30426 30800 30456
rect 25681 30424 30800 30426
rect 25681 30368 25686 30424
rect 25742 30368 30800 30424
rect 25681 30366 30800 30368
rect 25681 30363 25747 30366
rect 29200 30336 30800 30366
rect 20345 30154 20411 30157
rect 21725 30154 21791 30157
rect 20345 30152 21791 30154
rect 20345 30096 20350 30152
rect 20406 30096 21730 30152
rect 21786 30096 21791 30152
rect 20345 30094 21791 30096
rect 20345 30091 20411 30094
rect 21725 30091 21791 30094
rect -800 30018 800 30048
rect 2773 30018 2839 30021
rect -800 30016 2839 30018
rect -800 29960 2778 30016
rect 2834 29960 2839 30016
rect -800 29958 2839 29960
rect -800 29928 800 29958
rect 2773 29955 2839 29958
rect 26141 30018 26207 30021
rect 29200 30018 30800 30048
rect 26141 30016 30800 30018
rect 26141 29960 26146 30016
rect 26202 29960 30800 30016
rect 26141 29958 30800 29960
rect 26141 29955 26207 29958
rect 10208 29952 10528 29953
rect 10208 29888 10216 29952
rect 10280 29888 10296 29952
rect 10360 29888 10376 29952
rect 10440 29888 10456 29952
rect 10520 29888 10528 29952
rect 10208 29887 10528 29888
rect 19472 29952 19792 29953
rect 19472 29888 19480 29952
rect 19544 29888 19560 29952
rect 19624 29888 19640 29952
rect 19704 29888 19720 29952
rect 19784 29888 19792 29952
rect 29200 29928 30800 29958
rect 19472 29887 19792 29888
rect 5441 29882 5507 29885
rect 5717 29882 5783 29885
rect 5441 29880 5783 29882
rect 5441 29824 5446 29880
rect 5502 29824 5722 29880
rect 5778 29824 5783 29880
rect 5441 29822 5783 29824
rect 5441 29819 5507 29822
rect 5717 29819 5783 29822
rect 13813 29882 13879 29885
rect 15561 29882 15627 29885
rect 13813 29880 15627 29882
rect 13813 29824 13818 29880
rect 13874 29824 15566 29880
rect 15622 29824 15627 29880
rect 13813 29822 15627 29824
rect 13813 29819 13879 29822
rect 15561 29819 15627 29822
rect -800 29610 800 29640
rect 1945 29610 2011 29613
rect -800 29608 2011 29610
rect -800 29552 1950 29608
rect 2006 29552 2011 29608
rect -800 29550 2011 29552
rect -800 29520 800 29550
rect 1945 29547 2011 29550
rect 10225 29610 10291 29613
rect 15561 29610 15627 29613
rect 10225 29608 15627 29610
rect 10225 29552 10230 29608
rect 10286 29552 15566 29608
rect 15622 29552 15627 29608
rect 10225 29550 15627 29552
rect 10225 29547 10291 29550
rect 15561 29547 15627 29550
rect 27521 29610 27587 29613
rect 29200 29610 30800 29640
rect 27521 29608 30800 29610
rect 27521 29552 27526 29608
rect 27582 29552 30800 29608
rect 27521 29550 30800 29552
rect 27521 29547 27587 29550
rect 29200 29520 30800 29550
rect 5576 29408 5896 29409
rect 5576 29344 5584 29408
rect 5648 29344 5664 29408
rect 5728 29344 5744 29408
rect 5808 29344 5824 29408
rect 5888 29344 5896 29408
rect 5576 29343 5896 29344
rect 14840 29408 15160 29409
rect 14840 29344 14848 29408
rect 14912 29344 14928 29408
rect 14992 29344 15008 29408
rect 15072 29344 15088 29408
rect 15152 29344 15160 29408
rect 14840 29343 15160 29344
rect 24104 29408 24424 29409
rect 24104 29344 24112 29408
rect 24176 29344 24192 29408
rect 24256 29344 24272 29408
rect 24336 29344 24352 29408
rect 24416 29344 24424 29408
rect 24104 29343 24424 29344
rect -800 29202 800 29232
rect 1853 29202 1919 29205
rect -800 29200 1919 29202
rect -800 29144 1858 29200
rect 1914 29144 1919 29200
rect -800 29142 1919 29144
rect -800 29112 800 29142
rect 1853 29139 1919 29142
rect 25681 29202 25747 29205
rect 29200 29202 30800 29232
rect 25681 29200 30800 29202
rect 25681 29144 25686 29200
rect 25742 29144 30800 29200
rect 25681 29142 30800 29144
rect 25681 29139 25747 29142
rect 29200 29112 30800 29142
rect 10501 29066 10567 29069
rect 11881 29066 11947 29069
rect 15469 29066 15535 29069
rect 10501 29064 15535 29066
rect 10501 29008 10506 29064
rect 10562 29008 11886 29064
rect 11942 29008 15474 29064
rect 15530 29008 15535 29064
rect 10501 29006 15535 29008
rect 10501 29003 10567 29006
rect 11881 29003 11947 29006
rect 15469 29003 15535 29006
rect 25221 29066 25287 29069
rect 25681 29066 25747 29069
rect 25221 29064 25747 29066
rect 25221 29008 25226 29064
rect 25282 29008 25686 29064
rect 25742 29008 25747 29064
rect 25221 29006 25747 29008
rect 25221 29003 25287 29006
rect 25681 29003 25747 29006
rect 2405 28930 2471 28933
rect 3969 28930 4035 28933
rect 2405 28928 4035 28930
rect 2405 28872 2410 28928
rect 2466 28872 3974 28928
rect 4030 28872 4035 28928
rect 2405 28870 4035 28872
rect 2405 28867 2471 28870
rect 3969 28867 4035 28870
rect 10685 28930 10751 28933
rect 11329 28930 11395 28933
rect 10685 28928 11395 28930
rect 10685 28872 10690 28928
rect 10746 28872 11334 28928
rect 11390 28872 11395 28928
rect 10685 28870 11395 28872
rect 10685 28867 10751 28870
rect 11329 28867 11395 28870
rect 10208 28864 10528 28865
rect -800 28794 800 28824
rect 10208 28800 10216 28864
rect 10280 28800 10296 28864
rect 10360 28800 10376 28864
rect 10440 28800 10456 28864
rect 10520 28800 10528 28864
rect 10208 28799 10528 28800
rect 19472 28864 19792 28865
rect 19472 28800 19480 28864
rect 19544 28800 19560 28864
rect 19624 28800 19640 28864
rect 19704 28800 19720 28864
rect 19784 28800 19792 28864
rect 19472 28799 19792 28800
rect 1853 28794 1919 28797
rect -800 28792 1919 28794
rect -800 28736 1858 28792
rect 1914 28736 1919 28792
rect -800 28734 1919 28736
rect -800 28704 800 28734
rect 1853 28731 1919 28734
rect 26877 28794 26943 28797
rect 29200 28794 30800 28824
rect 26877 28792 30800 28794
rect 26877 28736 26882 28792
rect 26938 28736 30800 28792
rect 26877 28734 30800 28736
rect 26877 28731 26943 28734
rect 29200 28704 30800 28734
rect -800 28386 800 28416
rect 3785 28386 3851 28389
rect -800 28384 3851 28386
rect -800 28328 3790 28384
rect 3846 28328 3851 28384
rect -800 28326 3851 28328
rect -800 28296 800 28326
rect 3785 28323 3851 28326
rect 26417 28386 26483 28389
rect 29200 28386 30800 28416
rect 26417 28384 30800 28386
rect 26417 28328 26422 28384
rect 26478 28328 30800 28384
rect 26417 28326 30800 28328
rect 26417 28323 26483 28326
rect 5576 28320 5896 28321
rect 5576 28256 5584 28320
rect 5648 28256 5664 28320
rect 5728 28256 5744 28320
rect 5808 28256 5824 28320
rect 5888 28256 5896 28320
rect 5576 28255 5896 28256
rect 14840 28320 15160 28321
rect 14840 28256 14848 28320
rect 14912 28256 14928 28320
rect 14992 28256 15008 28320
rect 15072 28256 15088 28320
rect 15152 28256 15160 28320
rect 14840 28255 15160 28256
rect 24104 28320 24424 28321
rect 24104 28256 24112 28320
rect 24176 28256 24192 28320
rect 24256 28256 24272 28320
rect 24336 28256 24352 28320
rect 24416 28256 24424 28320
rect 29200 28296 30800 28326
rect 24104 28255 24424 28256
rect 1761 28114 1827 28117
rect 7373 28114 7439 28117
rect 1761 28112 7439 28114
rect 1761 28056 1766 28112
rect 1822 28056 7378 28112
rect 7434 28056 7439 28112
rect 1761 28054 7439 28056
rect 1761 28051 1827 28054
rect 7373 28051 7439 28054
rect 20069 28114 20135 28117
rect 20069 28112 20178 28114
rect 20069 28056 20074 28112
rect 20130 28056 20178 28112
rect 20069 28051 20178 28056
rect -800 27978 800 28008
rect 3049 27978 3115 27981
rect -800 27976 3115 27978
rect -800 27920 3054 27976
rect 3110 27920 3115 27976
rect -800 27918 3115 27920
rect -800 27888 800 27918
rect 3049 27915 3115 27918
rect 20118 27845 20178 28051
rect 24025 27978 24091 27981
rect 26417 27978 26483 27981
rect 24025 27976 26483 27978
rect 24025 27920 24030 27976
rect 24086 27920 26422 27976
rect 26478 27920 26483 27976
rect 24025 27918 26483 27920
rect 24025 27915 24091 27918
rect 26417 27915 26483 27918
rect 27153 27978 27219 27981
rect 29200 27978 30800 28008
rect 27153 27976 30800 27978
rect 27153 27920 27158 27976
rect 27214 27920 30800 27976
rect 27153 27918 30800 27920
rect 27153 27915 27219 27918
rect 29200 27888 30800 27918
rect 20118 27840 20227 27845
rect 20118 27784 20166 27840
rect 20222 27784 20227 27840
rect 20118 27782 20227 27784
rect 20161 27779 20227 27782
rect 24669 27842 24735 27845
rect 26325 27842 26391 27845
rect 24669 27840 26391 27842
rect 24669 27784 24674 27840
rect 24730 27784 26330 27840
rect 26386 27784 26391 27840
rect 24669 27782 26391 27784
rect 24669 27779 24735 27782
rect 26325 27779 26391 27782
rect 10208 27776 10528 27777
rect 10208 27712 10216 27776
rect 10280 27712 10296 27776
rect 10360 27712 10376 27776
rect 10440 27712 10456 27776
rect 10520 27712 10528 27776
rect 10208 27711 10528 27712
rect 19472 27776 19792 27777
rect 19472 27712 19480 27776
rect 19544 27712 19560 27776
rect 19624 27712 19640 27776
rect 19704 27712 19720 27776
rect 19784 27712 19792 27776
rect 19472 27711 19792 27712
rect 12709 27706 12775 27709
rect 18505 27706 18571 27709
rect 12709 27704 18571 27706
rect 12709 27648 12714 27704
rect 12770 27648 18510 27704
rect 18566 27648 18571 27704
rect 12709 27646 18571 27648
rect 12709 27643 12775 27646
rect 18505 27643 18571 27646
rect 23289 27706 23355 27709
rect 26693 27706 26759 27709
rect 23289 27704 26759 27706
rect 23289 27648 23294 27704
rect 23350 27648 26698 27704
rect 26754 27648 26759 27704
rect 23289 27646 26759 27648
rect 23289 27643 23355 27646
rect 26693 27643 26759 27646
rect -800 27570 800 27600
rect 1945 27570 2011 27573
rect 18321 27570 18387 27573
rect -800 27568 2011 27570
rect -800 27512 1950 27568
rect 2006 27512 2011 27568
rect -800 27510 2011 27512
rect -800 27480 800 27510
rect 1945 27507 2011 27510
rect 18094 27568 18387 27570
rect 18094 27512 18326 27568
rect 18382 27512 18387 27568
rect 18094 27510 18387 27512
rect 18094 27437 18154 27510
rect 18321 27507 18387 27510
rect 21449 27570 21515 27573
rect 23933 27570 23999 27573
rect 21449 27568 23999 27570
rect 21449 27512 21454 27568
rect 21510 27512 23938 27568
rect 23994 27512 23999 27568
rect 21449 27510 23999 27512
rect 21449 27507 21515 27510
rect 23933 27507 23999 27510
rect 26141 27570 26207 27573
rect 29200 27570 30800 27600
rect 26141 27568 30800 27570
rect 26141 27512 26146 27568
rect 26202 27512 30800 27568
rect 26141 27510 30800 27512
rect 26141 27507 26207 27510
rect 29200 27480 30800 27510
rect 11053 27434 11119 27437
rect 17861 27434 17927 27437
rect 11053 27432 17927 27434
rect 11053 27376 11058 27432
rect 11114 27376 17866 27432
rect 17922 27376 17927 27432
rect 11053 27374 17927 27376
rect 11053 27371 11119 27374
rect 17861 27371 17927 27374
rect 18045 27432 18154 27437
rect 18045 27376 18050 27432
rect 18106 27376 18154 27432
rect 18045 27374 18154 27376
rect 18321 27434 18387 27437
rect 18781 27434 18847 27437
rect 18321 27432 18847 27434
rect 18321 27376 18326 27432
rect 18382 27376 18786 27432
rect 18842 27376 18847 27432
rect 18321 27374 18847 27376
rect 18045 27371 18111 27374
rect 18321 27371 18387 27374
rect 18781 27371 18847 27374
rect 24853 27434 24919 27437
rect 26233 27434 26299 27437
rect 24853 27432 26299 27434
rect 24853 27376 24858 27432
rect 24914 27376 26238 27432
rect 26294 27376 26299 27432
rect 24853 27374 26299 27376
rect 24853 27371 24919 27374
rect 26233 27371 26299 27374
rect 5576 27232 5896 27233
rect -800 27162 800 27192
rect 5576 27168 5584 27232
rect 5648 27168 5664 27232
rect 5728 27168 5744 27232
rect 5808 27168 5824 27232
rect 5888 27168 5896 27232
rect 5576 27167 5896 27168
rect 14840 27232 15160 27233
rect 14840 27168 14848 27232
rect 14912 27168 14928 27232
rect 14992 27168 15008 27232
rect 15072 27168 15088 27232
rect 15152 27168 15160 27232
rect 14840 27167 15160 27168
rect 24104 27232 24424 27233
rect 24104 27168 24112 27232
rect 24176 27168 24192 27232
rect 24256 27168 24272 27232
rect 24336 27168 24352 27232
rect 24416 27168 24424 27232
rect 24104 27167 24424 27168
rect 2773 27162 2839 27165
rect -800 27160 2839 27162
rect -800 27104 2778 27160
rect 2834 27104 2839 27160
rect -800 27102 2839 27104
rect -800 27072 800 27102
rect 2773 27099 2839 27102
rect 26785 27162 26851 27165
rect 29200 27162 30800 27192
rect 26785 27160 30800 27162
rect 26785 27104 26790 27160
rect 26846 27104 30800 27160
rect 26785 27102 30800 27104
rect 26785 27099 26851 27102
rect 29200 27072 30800 27102
rect 11881 27026 11947 27029
rect 12801 27026 12867 27029
rect 11881 27024 12867 27026
rect 11881 26968 11886 27024
rect 11942 26968 12806 27024
rect 12862 26968 12867 27024
rect 11881 26966 12867 26968
rect 11881 26963 11947 26966
rect 12801 26963 12867 26966
rect 13169 27026 13235 27029
rect 13905 27026 13971 27029
rect 13169 27024 13971 27026
rect 13169 26968 13174 27024
rect 13230 26968 13910 27024
rect 13966 26968 13971 27024
rect 13169 26966 13971 26968
rect 13169 26963 13235 26966
rect 13905 26963 13971 26966
rect 23565 27026 23631 27029
rect 26233 27026 26299 27029
rect 23565 27024 26299 27026
rect 23565 26968 23570 27024
rect 23626 26968 26238 27024
rect 26294 26968 26299 27024
rect 23565 26966 26299 26968
rect 23565 26963 23631 26966
rect 26233 26963 26299 26966
rect 11605 26890 11671 26893
rect 14733 26890 14799 26893
rect 11605 26888 14799 26890
rect 11605 26832 11610 26888
rect 11666 26832 14738 26888
rect 14794 26832 14799 26888
rect 11605 26830 14799 26832
rect 11605 26827 11671 26830
rect -800 26754 800 26784
rect 12206 26757 12266 26830
rect 14733 26827 14799 26830
rect 1945 26754 2011 26757
rect -800 26752 2011 26754
rect -800 26696 1950 26752
rect 2006 26696 2011 26752
rect -800 26694 2011 26696
rect -800 26664 800 26694
rect 1945 26691 2011 26694
rect 12157 26752 12266 26757
rect 17309 26754 17375 26757
rect 12157 26696 12162 26752
rect 12218 26696 12266 26752
rect 12157 26694 12266 26696
rect 12344 26752 17375 26754
rect 12344 26696 17314 26752
rect 17370 26696 17375 26752
rect 12344 26694 17375 26696
rect 12157 26691 12223 26694
rect 10208 26688 10528 26689
rect 10208 26624 10216 26688
rect 10280 26624 10296 26688
rect 10360 26624 10376 26688
rect 10440 26624 10456 26688
rect 10520 26624 10528 26688
rect 10208 26623 10528 26624
rect 10593 26618 10659 26621
rect 10777 26618 10843 26621
rect 12344 26618 12404 26694
rect 17309 26691 17375 26694
rect 26693 26754 26759 26757
rect 29200 26754 30800 26784
rect 26693 26752 30800 26754
rect 26693 26696 26698 26752
rect 26754 26696 30800 26752
rect 26693 26694 30800 26696
rect 26693 26691 26759 26694
rect 19472 26688 19792 26689
rect 19472 26624 19480 26688
rect 19544 26624 19560 26688
rect 19624 26624 19640 26688
rect 19704 26624 19720 26688
rect 19784 26624 19792 26688
rect 29200 26664 30800 26694
rect 19472 26623 19792 26624
rect 10593 26616 12404 26618
rect 10593 26560 10598 26616
rect 10654 26560 10782 26616
rect 10838 26560 12404 26616
rect 10593 26558 12404 26560
rect 12525 26618 12591 26621
rect 13077 26618 13143 26621
rect 12525 26616 13143 26618
rect 12525 26560 12530 26616
rect 12586 26560 13082 26616
rect 13138 26560 13143 26616
rect 12525 26558 13143 26560
rect 10593 26555 10659 26558
rect 10777 26555 10843 26558
rect 12525 26555 12591 26558
rect 13077 26555 13143 26558
rect 14273 26618 14339 26621
rect 14549 26618 14615 26621
rect 14273 26616 14615 26618
rect 14273 26560 14278 26616
rect 14334 26560 14554 26616
rect 14610 26560 14615 26616
rect 14273 26558 14615 26560
rect 14273 26555 14339 26558
rect 14549 26555 14615 26558
rect 11145 26482 11211 26485
rect 15929 26482 15995 26485
rect 17861 26482 17927 26485
rect 11145 26480 17927 26482
rect 11145 26424 11150 26480
rect 11206 26424 15934 26480
rect 15990 26424 17866 26480
rect 17922 26424 17927 26480
rect 11145 26422 17927 26424
rect 11145 26419 11211 26422
rect 15929 26419 15995 26422
rect 17861 26419 17927 26422
rect -800 26346 800 26376
rect 1945 26346 2011 26349
rect -800 26344 2011 26346
rect -800 26288 1950 26344
rect 2006 26288 2011 26344
rect -800 26286 2011 26288
rect -800 26256 800 26286
rect 1945 26283 2011 26286
rect 9949 26346 10015 26349
rect 11148 26346 11208 26419
rect 17033 26346 17099 26349
rect 9949 26344 11208 26346
rect 9949 26288 9954 26344
rect 10010 26288 11208 26344
rect 9949 26286 11208 26288
rect 14230 26344 17099 26346
rect 14230 26288 17038 26344
rect 17094 26288 17099 26344
rect 14230 26286 17099 26288
rect 9949 26283 10015 26286
rect 10409 26210 10475 26213
rect 14230 26210 14290 26286
rect 17033 26283 17099 26286
rect 28165 26346 28231 26349
rect 29200 26346 30800 26376
rect 28165 26344 30800 26346
rect 28165 26288 28170 26344
rect 28226 26288 30800 26344
rect 28165 26286 30800 26288
rect 28165 26283 28231 26286
rect 29200 26256 30800 26286
rect 10409 26208 14290 26210
rect 10409 26152 10414 26208
rect 10470 26152 14290 26208
rect 10409 26150 14290 26152
rect 10409 26147 10475 26150
rect 5576 26144 5896 26145
rect 5576 26080 5584 26144
rect 5648 26080 5664 26144
rect 5728 26080 5744 26144
rect 5808 26080 5824 26144
rect 5888 26080 5896 26144
rect 5576 26079 5896 26080
rect 14840 26144 15160 26145
rect 14840 26080 14848 26144
rect 14912 26080 14928 26144
rect 14992 26080 15008 26144
rect 15072 26080 15088 26144
rect 15152 26080 15160 26144
rect 14840 26079 15160 26080
rect 24104 26144 24424 26145
rect 24104 26080 24112 26144
rect 24176 26080 24192 26144
rect 24256 26080 24272 26144
rect 24336 26080 24352 26144
rect 24416 26080 24424 26144
rect 24104 26079 24424 26080
rect 13169 26074 13235 26077
rect 14089 26074 14155 26077
rect 13169 26072 14155 26074
rect 13169 26016 13174 26072
rect 13230 26016 14094 26072
rect 14150 26016 14155 26072
rect 13169 26014 14155 26016
rect 13169 26011 13235 26014
rect 14089 26011 14155 26014
rect -800 25938 800 25968
rect 1853 25938 1919 25941
rect -800 25936 1919 25938
rect -800 25880 1858 25936
rect 1914 25880 1919 25936
rect -800 25878 1919 25880
rect -800 25848 800 25878
rect 1853 25875 1919 25878
rect 24945 25938 25011 25941
rect 29200 25938 30800 25968
rect 24945 25936 30800 25938
rect 24945 25880 24950 25936
rect 25006 25880 30800 25936
rect 24945 25878 30800 25880
rect 24945 25875 25011 25878
rect 29200 25848 30800 25878
rect 10208 25600 10528 25601
rect -800 25530 800 25560
rect 10208 25536 10216 25600
rect 10280 25536 10296 25600
rect 10360 25536 10376 25600
rect 10440 25536 10456 25600
rect 10520 25536 10528 25600
rect 10208 25535 10528 25536
rect 19472 25600 19792 25601
rect 19472 25536 19480 25600
rect 19544 25536 19560 25600
rect 19624 25536 19640 25600
rect 19704 25536 19720 25600
rect 19784 25536 19792 25600
rect 19472 25535 19792 25536
rect 1761 25530 1827 25533
rect -800 25528 1827 25530
rect -800 25472 1766 25528
rect 1822 25472 1827 25528
rect -800 25470 1827 25472
rect -800 25440 800 25470
rect 1761 25467 1827 25470
rect 25405 25530 25471 25533
rect 29200 25530 30800 25560
rect 25405 25528 30800 25530
rect 25405 25472 25410 25528
rect 25466 25472 30800 25528
rect 25405 25470 30800 25472
rect 25405 25467 25471 25470
rect 29200 25440 30800 25470
rect 14273 25394 14339 25397
rect 14092 25392 14339 25394
rect 14092 25336 14278 25392
rect 14334 25336 14339 25392
rect 14092 25334 14339 25336
rect 14092 25261 14152 25334
rect 14273 25331 14339 25334
rect 14089 25256 14155 25261
rect 14089 25200 14094 25256
rect 14150 25200 14155 25256
rect 14089 25195 14155 25200
rect -800 25122 800 25152
rect 4061 25122 4127 25125
rect -800 25120 4127 25122
rect -800 25064 4066 25120
rect 4122 25064 4127 25120
rect -800 25062 4127 25064
rect -800 25032 800 25062
rect 4061 25059 4127 25062
rect 5576 25056 5896 25057
rect 5576 24992 5584 25056
rect 5648 24992 5664 25056
rect 5728 24992 5744 25056
rect 5808 24992 5824 25056
rect 5888 24992 5896 25056
rect 5576 24991 5896 24992
rect 14092 24986 14152 25195
rect 26141 25122 26207 25125
rect 29200 25122 30800 25152
rect 26141 25120 30800 25122
rect 26141 25064 26146 25120
rect 26202 25064 30800 25120
rect 26141 25062 30800 25064
rect 26141 25059 26207 25062
rect 14840 25056 15160 25057
rect 14840 24992 14848 25056
rect 14912 24992 14928 25056
rect 14992 24992 15008 25056
rect 15072 24992 15088 25056
rect 15152 24992 15160 25056
rect 14840 24991 15160 24992
rect 24104 25056 24424 25057
rect 24104 24992 24112 25056
rect 24176 24992 24192 25056
rect 24256 24992 24272 25056
rect 24336 24992 24352 25056
rect 24416 24992 24424 25056
rect 29200 25032 30800 25062
rect 24104 24991 24424 24992
rect 14092 24926 14336 24986
rect 14276 24853 14336 24926
rect 11973 24850 12039 24853
rect 12249 24850 12315 24853
rect 11973 24848 12315 24850
rect 11973 24792 11978 24848
rect 12034 24792 12254 24848
rect 12310 24792 12315 24848
rect 11973 24790 12315 24792
rect 11973 24787 12039 24790
rect 12249 24787 12315 24790
rect 14273 24850 14339 24853
rect 17309 24850 17375 24853
rect 14273 24848 17375 24850
rect 14273 24792 14278 24848
rect 14334 24792 17314 24848
rect 17370 24792 17375 24848
rect 14273 24790 17375 24792
rect 14273 24787 14339 24790
rect 17309 24787 17375 24790
rect -800 24714 800 24744
rect 3049 24714 3115 24717
rect -800 24712 3115 24714
rect -800 24656 3054 24712
rect 3110 24656 3115 24712
rect -800 24654 3115 24656
rect -800 24624 800 24654
rect 3049 24651 3115 24654
rect 26141 24714 26207 24717
rect 29200 24714 30800 24744
rect 26141 24712 30800 24714
rect 26141 24656 26146 24712
rect 26202 24656 30800 24712
rect 26141 24654 30800 24656
rect 26141 24651 26207 24654
rect 29200 24624 30800 24654
rect 10208 24512 10528 24513
rect 10208 24448 10216 24512
rect 10280 24448 10296 24512
rect 10360 24448 10376 24512
rect 10440 24448 10456 24512
rect 10520 24448 10528 24512
rect 10208 24447 10528 24448
rect 19472 24512 19792 24513
rect 19472 24448 19480 24512
rect 19544 24448 19560 24512
rect 19624 24448 19640 24512
rect 19704 24448 19720 24512
rect 19784 24448 19792 24512
rect 19472 24447 19792 24448
rect -800 24306 800 24336
rect 3325 24306 3391 24309
rect -800 24304 3391 24306
rect -800 24248 3330 24304
rect 3386 24248 3391 24304
rect -800 24246 3391 24248
rect -800 24216 800 24246
rect 3325 24243 3391 24246
rect 27521 24306 27587 24309
rect 29200 24306 30800 24336
rect 27521 24304 30800 24306
rect 27521 24248 27526 24304
rect 27582 24248 30800 24304
rect 27521 24246 30800 24248
rect 27521 24243 27587 24246
rect 29200 24216 30800 24246
rect 5576 23968 5896 23969
rect -800 23898 800 23928
rect 5576 23904 5584 23968
rect 5648 23904 5664 23968
rect 5728 23904 5744 23968
rect 5808 23904 5824 23968
rect 5888 23904 5896 23968
rect 5576 23903 5896 23904
rect 14840 23968 15160 23969
rect 14840 23904 14848 23968
rect 14912 23904 14928 23968
rect 14992 23904 15008 23968
rect 15072 23904 15088 23968
rect 15152 23904 15160 23968
rect 14840 23903 15160 23904
rect 24104 23968 24424 23969
rect 24104 23904 24112 23968
rect 24176 23904 24192 23968
rect 24256 23904 24272 23968
rect 24336 23904 24352 23968
rect 24416 23904 24424 23968
rect 24104 23903 24424 23904
rect 2773 23898 2839 23901
rect -800 23896 2839 23898
rect -800 23840 2778 23896
rect 2834 23840 2839 23896
rect -800 23838 2839 23840
rect -800 23808 800 23838
rect 2773 23835 2839 23838
rect 26785 23898 26851 23901
rect 29200 23898 30800 23928
rect 26785 23896 30800 23898
rect 26785 23840 26790 23896
rect 26846 23840 30800 23896
rect 26785 23838 30800 23840
rect 26785 23835 26851 23838
rect 29200 23808 30800 23838
rect -800 23490 800 23520
rect 1945 23490 2011 23493
rect -800 23488 2011 23490
rect -800 23432 1950 23488
rect 2006 23432 2011 23488
rect -800 23430 2011 23432
rect -800 23400 800 23430
rect 1945 23427 2011 23430
rect 28165 23490 28231 23493
rect 29200 23490 30800 23520
rect 28165 23488 30800 23490
rect 28165 23432 28170 23488
rect 28226 23432 30800 23488
rect 28165 23430 30800 23432
rect 28165 23427 28231 23430
rect 10208 23424 10528 23425
rect 10208 23360 10216 23424
rect 10280 23360 10296 23424
rect 10360 23360 10376 23424
rect 10440 23360 10456 23424
rect 10520 23360 10528 23424
rect 10208 23359 10528 23360
rect 19472 23424 19792 23425
rect 19472 23360 19480 23424
rect 19544 23360 19560 23424
rect 19624 23360 19640 23424
rect 19704 23360 19720 23424
rect 19784 23360 19792 23424
rect 29200 23400 30800 23430
rect 19472 23359 19792 23360
rect -800 23082 800 23112
rect 2773 23082 2839 23085
rect -800 23080 2839 23082
rect -800 23024 2778 23080
rect 2834 23024 2839 23080
rect -800 23022 2839 23024
rect -800 22992 800 23022
rect 2773 23019 2839 23022
rect 28165 23082 28231 23085
rect 29200 23082 30800 23112
rect 28165 23080 30800 23082
rect 28165 23024 28170 23080
rect 28226 23024 30800 23080
rect 28165 23022 30800 23024
rect 28165 23019 28231 23022
rect 29200 22992 30800 23022
rect 5576 22880 5896 22881
rect 5576 22816 5584 22880
rect 5648 22816 5664 22880
rect 5728 22816 5744 22880
rect 5808 22816 5824 22880
rect 5888 22816 5896 22880
rect 5576 22815 5896 22816
rect 14840 22880 15160 22881
rect 14840 22816 14848 22880
rect 14912 22816 14928 22880
rect 14992 22816 15008 22880
rect 15072 22816 15088 22880
rect 15152 22816 15160 22880
rect 14840 22815 15160 22816
rect 24104 22880 24424 22881
rect 24104 22816 24112 22880
rect 24176 22816 24192 22880
rect 24256 22816 24272 22880
rect 24336 22816 24352 22880
rect 24416 22816 24424 22880
rect 24104 22815 24424 22816
rect -800 22674 800 22704
rect 1577 22674 1643 22677
rect -800 22672 1643 22674
rect -800 22616 1582 22672
rect 1638 22616 1643 22672
rect -800 22614 1643 22616
rect -800 22584 800 22614
rect 1577 22611 1643 22614
rect 25129 22674 25195 22677
rect 29200 22674 30800 22704
rect 25129 22672 30800 22674
rect 25129 22616 25134 22672
rect 25190 22616 30800 22672
rect 25129 22614 30800 22616
rect 25129 22611 25195 22614
rect 29200 22584 30800 22614
rect 4245 22402 4311 22405
rect 5257 22402 5323 22405
rect 4245 22400 5323 22402
rect 4245 22344 4250 22400
rect 4306 22344 5262 22400
rect 5318 22344 5323 22400
rect 4245 22342 5323 22344
rect 4245 22339 4311 22342
rect 5257 22339 5323 22342
rect 10208 22336 10528 22337
rect -800 22266 800 22296
rect 10208 22272 10216 22336
rect 10280 22272 10296 22336
rect 10360 22272 10376 22336
rect 10440 22272 10456 22336
rect 10520 22272 10528 22336
rect 10208 22271 10528 22272
rect 19472 22336 19792 22337
rect 19472 22272 19480 22336
rect 19544 22272 19560 22336
rect 19624 22272 19640 22336
rect 19704 22272 19720 22336
rect 19784 22272 19792 22336
rect 19472 22271 19792 22272
rect 1393 22266 1459 22269
rect -800 22264 1459 22266
rect -800 22208 1398 22264
rect 1454 22208 1459 22264
rect -800 22206 1459 22208
rect -800 22176 800 22206
rect 1393 22203 1459 22206
rect 26325 22266 26391 22269
rect 29200 22266 30800 22296
rect 26325 22264 30800 22266
rect 26325 22208 26330 22264
rect 26386 22208 30800 22264
rect 26325 22206 30800 22208
rect 26325 22203 26391 22206
rect 29200 22176 30800 22206
rect 23473 22130 23539 22133
rect 23430 22128 23539 22130
rect 23430 22072 23478 22128
rect 23534 22072 23539 22128
rect 23430 22067 23539 22072
rect 23430 21997 23490 22067
rect 5073 21994 5139 21997
rect 5533 21994 5599 21997
rect 5073 21992 5599 21994
rect 5073 21936 5078 21992
rect 5134 21936 5538 21992
rect 5594 21936 5599 21992
rect 5073 21934 5599 21936
rect 5073 21931 5139 21934
rect 5533 21931 5599 21934
rect 15745 21994 15811 21997
rect 15745 21992 15946 21994
rect 15745 21936 15750 21992
rect 15806 21936 15946 21992
rect 15745 21934 15946 21936
rect 15745 21931 15811 21934
rect -800 21858 800 21888
rect 4521 21858 4587 21861
rect -800 21856 4587 21858
rect -800 21800 4526 21856
rect 4582 21800 4587 21856
rect -800 21798 4587 21800
rect -800 21768 800 21798
rect 4521 21795 4587 21798
rect 5576 21792 5896 21793
rect 5576 21728 5584 21792
rect 5648 21728 5664 21792
rect 5728 21728 5744 21792
rect 5808 21728 5824 21792
rect 5888 21728 5896 21792
rect 5576 21727 5896 21728
rect 14840 21792 15160 21793
rect 14840 21728 14848 21792
rect 14912 21728 14928 21792
rect 14992 21728 15008 21792
rect 15072 21728 15088 21792
rect 15152 21728 15160 21792
rect 14840 21727 15160 21728
rect 12525 21722 12591 21725
rect 12525 21720 13784 21722
rect 12525 21664 12530 21720
rect 12586 21664 13784 21720
rect 12525 21662 13784 21664
rect 12525 21659 12591 21662
rect 12985 21586 13051 21589
rect 12985 21584 13554 21586
rect 12985 21528 12990 21584
rect 13046 21528 13554 21584
rect 12985 21526 13554 21528
rect 12985 21523 13051 21526
rect -800 21450 800 21480
rect 3141 21450 3207 21453
rect -800 21448 3207 21450
rect -800 21392 3146 21448
rect 3202 21392 3207 21448
rect -800 21390 3207 21392
rect -800 21360 800 21390
rect 3141 21387 3207 21390
rect 10208 21248 10528 21249
rect 10208 21184 10216 21248
rect 10280 21184 10296 21248
rect 10360 21184 10376 21248
rect 10440 21184 10456 21248
rect 10520 21184 10528 21248
rect 10208 21183 10528 21184
rect -800 21042 800 21072
rect 1577 21042 1643 21045
rect -800 21040 1643 21042
rect -800 20984 1582 21040
rect 1638 20984 1643 21040
rect -800 20982 1643 20984
rect -800 20952 800 20982
rect 1577 20979 1643 20982
rect 13494 20906 13554 21526
rect 13724 21453 13784 21662
rect 13721 21448 13787 21453
rect 13721 21392 13726 21448
rect 13782 21392 13787 21448
rect 13721 21387 13787 21392
rect 15886 21045 15946 21934
rect 23381 21992 23490 21997
rect 24117 21994 24183 21997
rect 23381 21936 23386 21992
rect 23442 21936 23490 21992
rect 23381 21934 23490 21936
rect 23982 21992 24183 21994
rect 23982 21936 24122 21992
rect 24178 21936 24183 21992
rect 23982 21934 24183 21936
rect 23381 21931 23447 21934
rect 23982 21586 24042 21934
rect 24117 21931 24183 21934
rect 25865 21858 25931 21861
rect 29200 21858 30800 21888
rect 25865 21856 30800 21858
rect 25865 21800 25870 21856
rect 25926 21800 30800 21856
rect 25865 21798 30800 21800
rect 25865 21795 25931 21798
rect 24104 21792 24424 21793
rect 24104 21728 24112 21792
rect 24176 21728 24192 21792
rect 24256 21728 24272 21792
rect 24336 21728 24352 21792
rect 24416 21728 24424 21792
rect 29200 21768 30800 21798
rect 24104 21727 24424 21728
rect 24117 21586 24183 21589
rect 23982 21584 24183 21586
rect 23982 21528 24122 21584
rect 24178 21528 24183 21584
rect 23982 21526 24183 21528
rect 24117 21523 24183 21526
rect 27521 21450 27587 21453
rect 29200 21450 30800 21480
rect 27521 21448 30800 21450
rect 27521 21392 27526 21448
rect 27582 21392 30800 21448
rect 27521 21390 30800 21392
rect 27521 21387 27587 21390
rect 29200 21360 30800 21390
rect 19472 21248 19792 21249
rect 19472 21184 19480 21248
rect 19544 21184 19560 21248
rect 19624 21184 19640 21248
rect 19704 21184 19720 21248
rect 19784 21184 19792 21248
rect 19472 21183 19792 21184
rect 15886 21040 15995 21045
rect 15886 20984 15934 21040
rect 15990 20984 15995 21040
rect 15886 20982 15995 20984
rect 15929 20979 15995 20982
rect 26877 21042 26943 21045
rect 29200 21042 30800 21072
rect 26877 21040 30800 21042
rect 26877 20984 26882 21040
rect 26938 20984 30800 21040
rect 26877 20982 30800 20984
rect 26877 20979 26943 20982
rect 29200 20952 30800 20982
rect 13721 20906 13787 20909
rect 13494 20904 13787 20906
rect 13494 20848 13726 20904
rect 13782 20848 13787 20904
rect 13494 20846 13787 20848
rect 13721 20843 13787 20846
rect 11789 20770 11855 20773
rect 14089 20770 14155 20773
rect 11789 20768 14155 20770
rect 11789 20712 11794 20768
rect 11850 20712 14094 20768
rect 14150 20712 14155 20768
rect 11789 20710 14155 20712
rect 11789 20707 11855 20710
rect 14089 20707 14155 20710
rect 5576 20704 5896 20705
rect -800 20634 800 20664
rect 5576 20640 5584 20704
rect 5648 20640 5664 20704
rect 5728 20640 5744 20704
rect 5808 20640 5824 20704
rect 5888 20640 5896 20704
rect 5576 20639 5896 20640
rect 14840 20704 15160 20705
rect 14840 20640 14848 20704
rect 14912 20640 14928 20704
rect 14992 20640 15008 20704
rect 15072 20640 15088 20704
rect 15152 20640 15160 20704
rect 14840 20639 15160 20640
rect 24104 20704 24424 20705
rect 24104 20640 24112 20704
rect 24176 20640 24192 20704
rect 24256 20640 24272 20704
rect 24336 20640 24352 20704
rect 24416 20640 24424 20704
rect 24104 20639 24424 20640
rect 2773 20634 2839 20637
rect -800 20632 2839 20634
rect -800 20576 2778 20632
rect 2834 20576 2839 20632
rect -800 20574 2839 20576
rect -800 20544 800 20574
rect 2773 20571 2839 20574
rect 28073 20634 28139 20637
rect 29200 20634 30800 20664
rect 28073 20632 30800 20634
rect 28073 20576 28078 20632
rect 28134 20576 30800 20632
rect 28073 20574 30800 20576
rect 28073 20571 28139 20574
rect 29200 20544 30800 20574
rect 11237 20362 11303 20365
rect 16113 20362 16179 20365
rect 11237 20360 16179 20362
rect 11237 20304 11242 20360
rect 11298 20304 16118 20360
rect 16174 20304 16179 20360
rect 11237 20302 16179 20304
rect 11237 20299 11303 20302
rect 16113 20299 16179 20302
rect -800 20226 800 20256
rect 1669 20226 1735 20229
rect -800 20224 1735 20226
rect -800 20168 1674 20224
rect 1730 20168 1735 20224
rect -800 20166 1735 20168
rect -800 20136 800 20166
rect 1669 20163 1735 20166
rect 28165 20226 28231 20229
rect 29200 20226 30800 20256
rect 28165 20224 30800 20226
rect 28165 20168 28170 20224
rect 28226 20168 30800 20224
rect 28165 20166 30800 20168
rect 28165 20163 28231 20166
rect 10208 20160 10528 20161
rect 10208 20096 10216 20160
rect 10280 20096 10296 20160
rect 10360 20096 10376 20160
rect 10440 20096 10456 20160
rect 10520 20096 10528 20160
rect 10208 20095 10528 20096
rect 19472 20160 19792 20161
rect 19472 20096 19480 20160
rect 19544 20096 19560 20160
rect 19624 20096 19640 20160
rect 19704 20096 19720 20160
rect 19784 20096 19792 20160
rect 29200 20136 30800 20166
rect 19472 20095 19792 20096
rect 18321 20090 18387 20093
rect 18278 20088 18387 20090
rect 18278 20032 18326 20088
rect 18382 20032 18387 20088
rect 18278 20027 18387 20032
rect -800 19818 800 19848
rect 1945 19818 2011 19821
rect -800 19816 2011 19818
rect -800 19760 1950 19816
rect 2006 19760 2011 19816
rect -800 19758 2011 19760
rect -800 19728 800 19758
rect 1945 19755 2011 19758
rect 5576 19616 5896 19617
rect 5576 19552 5584 19616
rect 5648 19552 5664 19616
rect 5728 19552 5744 19616
rect 5808 19552 5824 19616
rect 5888 19552 5896 19616
rect 5576 19551 5896 19552
rect 14840 19616 15160 19617
rect 14840 19552 14848 19616
rect 14912 19552 14928 19616
rect 14992 19552 15008 19616
rect 15072 19552 15088 19616
rect 15152 19552 15160 19616
rect 14840 19551 15160 19552
rect -800 19410 800 19440
rect 1853 19410 1919 19413
rect -800 19408 1919 19410
rect -800 19352 1858 19408
rect 1914 19352 1919 19408
rect -800 19350 1919 19352
rect -800 19320 800 19350
rect 1853 19347 1919 19350
rect 10961 19138 11027 19141
rect 16389 19138 16455 19141
rect 10961 19136 16455 19138
rect 10961 19080 10966 19136
rect 11022 19080 16394 19136
rect 16450 19080 16455 19136
rect 10961 19078 16455 19080
rect 10961 19075 11027 19078
rect 16389 19075 16455 19078
rect 10208 19072 10528 19073
rect -800 19002 800 19032
rect 10208 19008 10216 19072
rect 10280 19008 10296 19072
rect 10360 19008 10376 19072
rect 10440 19008 10456 19072
rect 10520 19008 10528 19072
rect 10208 19007 10528 19008
rect 1853 19002 1919 19005
rect 12065 19002 12131 19005
rect -800 19000 1919 19002
rect -800 18944 1858 19000
rect 1914 18944 1919 19000
rect -800 18942 1919 18944
rect -800 18912 800 18942
rect 1853 18939 1919 18942
rect 12022 19000 12131 19002
rect 12022 18944 12070 19000
rect 12126 18944 12131 19000
rect 12022 18939 12131 18944
rect 4981 18866 5047 18869
rect 5533 18866 5599 18869
rect 4981 18864 5599 18866
rect 4981 18808 4986 18864
rect 5042 18808 5538 18864
rect 5594 18808 5599 18864
rect 4981 18806 5599 18808
rect 4981 18803 5047 18806
rect 5533 18803 5599 18806
rect -800 18594 800 18624
rect 3417 18594 3483 18597
rect -800 18592 3483 18594
rect -800 18536 3422 18592
rect 3478 18536 3483 18592
rect -800 18534 3483 18536
rect -800 18504 800 18534
rect 3417 18531 3483 18534
rect 5576 18528 5896 18529
rect 5576 18464 5584 18528
rect 5648 18464 5664 18528
rect 5728 18464 5744 18528
rect 5808 18464 5824 18528
rect 5888 18464 5896 18528
rect 5576 18463 5896 18464
rect 11881 18322 11947 18325
rect 12022 18322 12082 18939
rect 13813 18730 13879 18733
rect 17217 18730 17283 18733
rect 13813 18728 17283 18730
rect 13813 18672 13818 18728
rect 13874 18672 17222 18728
rect 17278 18672 17283 18728
rect 13813 18670 17283 18672
rect 13813 18667 13879 18670
rect 17217 18667 17283 18670
rect 18045 18730 18111 18733
rect 18278 18730 18338 20027
rect 28165 19818 28231 19821
rect 29200 19818 30800 19848
rect 28165 19816 30800 19818
rect 28165 19760 28170 19816
rect 28226 19760 30800 19816
rect 28165 19758 30800 19760
rect 28165 19755 28231 19758
rect 29200 19728 30800 19758
rect 24104 19616 24424 19617
rect 24104 19552 24112 19616
rect 24176 19552 24192 19616
rect 24256 19552 24272 19616
rect 24336 19552 24352 19616
rect 24416 19552 24424 19616
rect 24104 19551 24424 19552
rect 25957 19410 26023 19413
rect 29200 19410 30800 19440
rect 25957 19408 30800 19410
rect 25957 19352 25962 19408
rect 26018 19352 30800 19408
rect 25957 19350 30800 19352
rect 25957 19347 26023 19350
rect 29200 19320 30800 19350
rect 20621 19274 20687 19277
rect 24209 19274 24275 19277
rect 20621 19272 24275 19274
rect 20621 19216 20626 19272
rect 20682 19216 24214 19272
rect 24270 19216 24275 19272
rect 20621 19214 24275 19216
rect 20621 19211 20687 19214
rect 24209 19211 24275 19214
rect 19472 19072 19792 19073
rect 19472 19008 19480 19072
rect 19544 19008 19560 19072
rect 19624 19008 19640 19072
rect 19704 19008 19720 19072
rect 19784 19008 19792 19072
rect 19472 19007 19792 19008
rect 25865 19002 25931 19005
rect 29200 19002 30800 19032
rect 25865 19000 30800 19002
rect 25865 18944 25870 19000
rect 25926 18944 30800 19000
rect 25865 18942 30800 18944
rect 25865 18939 25931 18942
rect 29200 18912 30800 18942
rect 21725 18864 21791 18869
rect 21725 18808 21730 18864
rect 21786 18808 21791 18864
rect 21725 18803 21791 18808
rect 24945 18866 25011 18869
rect 25865 18866 25931 18869
rect 24945 18864 25931 18866
rect 24945 18808 24950 18864
rect 25006 18808 25870 18864
rect 25926 18808 25931 18864
rect 24945 18806 25931 18808
rect 24945 18803 25011 18806
rect 25865 18803 25931 18806
rect 18045 18728 18338 18730
rect 18045 18672 18050 18728
rect 18106 18672 18338 18728
rect 18045 18670 18338 18672
rect 18045 18667 18111 18670
rect 20897 18594 20963 18597
rect 21728 18594 21788 18803
rect 22737 18730 22803 18733
rect 25589 18730 25655 18733
rect 25957 18730 26023 18733
rect 22737 18728 24594 18730
rect 22737 18672 22742 18728
rect 22798 18672 24594 18728
rect 22737 18670 24594 18672
rect 22737 18667 22803 18670
rect 20897 18592 21788 18594
rect 20897 18536 20902 18592
rect 20958 18536 21788 18592
rect 20897 18534 21788 18536
rect 24534 18594 24594 18670
rect 25589 18728 26023 18730
rect 25589 18672 25594 18728
rect 25650 18672 25962 18728
rect 26018 18672 26023 18728
rect 25589 18670 26023 18672
rect 25589 18667 25655 18670
rect 25957 18667 26023 18670
rect 26233 18594 26299 18597
rect 24534 18592 26299 18594
rect 24534 18536 26238 18592
rect 26294 18536 26299 18592
rect 24534 18534 26299 18536
rect 20897 18531 20963 18534
rect 26233 18531 26299 18534
rect 26693 18594 26759 18597
rect 29200 18594 30800 18624
rect 26693 18592 30800 18594
rect 26693 18536 26698 18592
rect 26754 18536 30800 18592
rect 26693 18534 30800 18536
rect 26693 18531 26759 18534
rect 14840 18528 15160 18529
rect 14840 18464 14848 18528
rect 14912 18464 14928 18528
rect 14992 18464 15008 18528
rect 15072 18464 15088 18528
rect 15152 18464 15160 18528
rect 14840 18463 15160 18464
rect 24104 18528 24424 18529
rect 24104 18464 24112 18528
rect 24176 18464 24192 18528
rect 24256 18464 24272 18528
rect 24336 18464 24352 18528
rect 24416 18464 24424 18528
rect 29200 18504 30800 18534
rect 24104 18463 24424 18464
rect 11881 18320 12082 18322
rect 11881 18264 11886 18320
rect 11942 18264 12082 18320
rect 11881 18262 12082 18264
rect 11881 18259 11947 18262
rect -800 18186 800 18216
rect 2865 18186 2931 18189
rect -800 18184 2931 18186
rect -800 18128 2870 18184
rect 2926 18128 2931 18184
rect -800 18126 2931 18128
rect -800 18096 800 18126
rect 2865 18123 2931 18126
rect 16389 18186 16455 18189
rect 17033 18186 17099 18189
rect 16389 18184 17099 18186
rect 16389 18128 16394 18184
rect 16450 18128 17038 18184
rect 17094 18128 17099 18184
rect 16389 18126 17099 18128
rect 16389 18123 16455 18126
rect 17033 18123 17099 18126
rect 28165 18186 28231 18189
rect 29200 18186 30800 18216
rect 28165 18184 30800 18186
rect 28165 18128 28170 18184
rect 28226 18128 30800 18184
rect 28165 18126 30800 18128
rect 28165 18123 28231 18126
rect 29200 18096 30800 18126
rect 11789 18050 11855 18053
rect 16665 18050 16731 18053
rect 11789 18048 16731 18050
rect 11789 17992 11794 18048
rect 11850 17992 16670 18048
rect 16726 17992 16731 18048
rect 11789 17990 16731 17992
rect 11789 17987 11855 17990
rect 16665 17987 16731 17990
rect 10208 17984 10528 17985
rect 10208 17920 10216 17984
rect 10280 17920 10296 17984
rect 10360 17920 10376 17984
rect 10440 17920 10456 17984
rect 10520 17920 10528 17984
rect 10208 17919 10528 17920
rect 19472 17984 19792 17985
rect 19472 17920 19480 17984
rect 19544 17920 19560 17984
rect 19624 17920 19640 17984
rect 19704 17920 19720 17984
rect 19784 17920 19792 17984
rect 19472 17919 19792 17920
rect 10685 17914 10751 17917
rect 15745 17914 15811 17917
rect 10685 17912 15811 17914
rect 10685 17856 10690 17912
rect 10746 17856 15750 17912
rect 15806 17856 15811 17912
rect 10685 17854 15811 17856
rect 10685 17851 10751 17854
rect 15745 17851 15811 17854
rect -800 17778 800 17808
rect 3233 17778 3299 17781
rect -800 17776 3299 17778
rect -800 17720 3238 17776
rect 3294 17720 3299 17776
rect -800 17718 3299 17720
rect -800 17688 800 17718
rect 3233 17715 3299 17718
rect 26877 17778 26943 17781
rect 29200 17778 30800 17808
rect 26877 17776 30800 17778
rect 26877 17720 26882 17776
rect 26938 17720 30800 17776
rect 26877 17718 30800 17720
rect 26877 17715 26943 17718
rect 29200 17688 30800 17718
rect 5576 17440 5896 17441
rect -800 17370 800 17400
rect 5576 17376 5584 17440
rect 5648 17376 5664 17440
rect 5728 17376 5744 17440
rect 5808 17376 5824 17440
rect 5888 17376 5896 17440
rect 5576 17375 5896 17376
rect 14840 17440 15160 17441
rect 14840 17376 14848 17440
rect 14912 17376 14928 17440
rect 14992 17376 15008 17440
rect 15072 17376 15088 17440
rect 15152 17376 15160 17440
rect 14840 17375 15160 17376
rect 24104 17440 24424 17441
rect 24104 17376 24112 17440
rect 24176 17376 24192 17440
rect 24256 17376 24272 17440
rect 24336 17376 24352 17440
rect 24416 17376 24424 17440
rect 24104 17375 24424 17376
rect 2773 17370 2839 17373
rect -800 17368 2839 17370
rect -800 17312 2778 17368
rect 2834 17312 2839 17368
rect -800 17310 2839 17312
rect -800 17280 800 17310
rect 2773 17307 2839 17310
rect 26877 17370 26943 17373
rect 29200 17370 30800 17400
rect 26877 17368 30800 17370
rect 26877 17312 26882 17368
rect 26938 17312 30800 17368
rect 26877 17310 30800 17312
rect 26877 17307 26943 17310
rect 29200 17280 30800 17310
rect -800 16962 800 16992
rect 1945 16962 2011 16965
rect -800 16960 2011 16962
rect -800 16904 1950 16960
rect 2006 16904 2011 16960
rect -800 16902 2011 16904
rect -800 16872 800 16902
rect 1945 16899 2011 16902
rect 28165 16962 28231 16965
rect 29200 16962 30800 16992
rect 28165 16960 30800 16962
rect 28165 16904 28170 16960
rect 28226 16904 30800 16960
rect 28165 16902 30800 16904
rect 28165 16899 28231 16902
rect 10208 16896 10528 16897
rect 10208 16832 10216 16896
rect 10280 16832 10296 16896
rect 10360 16832 10376 16896
rect 10440 16832 10456 16896
rect 10520 16832 10528 16896
rect 10208 16831 10528 16832
rect 19472 16896 19792 16897
rect 19472 16832 19480 16896
rect 19544 16832 19560 16896
rect 19624 16832 19640 16896
rect 19704 16832 19720 16896
rect 19784 16832 19792 16896
rect 29200 16872 30800 16902
rect 19472 16831 19792 16832
rect -800 16554 800 16584
rect 1945 16554 2011 16557
rect -800 16552 2011 16554
rect -800 16496 1950 16552
rect 2006 16496 2011 16552
rect -800 16494 2011 16496
rect -800 16464 800 16494
rect 1945 16491 2011 16494
rect 24209 16554 24275 16557
rect 24945 16554 25011 16557
rect 24209 16552 25011 16554
rect 24209 16496 24214 16552
rect 24270 16496 24950 16552
rect 25006 16496 25011 16552
rect 24209 16494 25011 16496
rect 24209 16491 24275 16494
rect 24945 16491 25011 16494
rect 28165 16554 28231 16557
rect 29200 16554 30800 16584
rect 28165 16552 30800 16554
rect 28165 16496 28170 16552
rect 28226 16496 30800 16552
rect 28165 16494 30800 16496
rect 28165 16491 28231 16494
rect 29200 16464 30800 16494
rect 5576 16352 5896 16353
rect 5576 16288 5584 16352
rect 5648 16288 5664 16352
rect 5728 16288 5744 16352
rect 5808 16288 5824 16352
rect 5888 16288 5896 16352
rect 5576 16287 5896 16288
rect 14840 16352 15160 16353
rect 14840 16288 14848 16352
rect 14912 16288 14928 16352
rect 14992 16288 15008 16352
rect 15072 16288 15088 16352
rect 15152 16288 15160 16352
rect 14840 16287 15160 16288
rect 24104 16352 24424 16353
rect 24104 16288 24112 16352
rect 24176 16288 24192 16352
rect 24256 16288 24272 16352
rect 24336 16288 24352 16352
rect 24416 16288 24424 16352
rect 24104 16287 24424 16288
rect 25405 16282 25471 16285
rect 25270 16280 25471 16282
rect 25270 16224 25410 16280
rect 25466 16224 25471 16280
rect 25270 16222 25471 16224
rect -800 16146 800 16176
rect 25270 16149 25330 16222
rect 25405 16219 25471 16222
rect 1853 16146 1919 16149
rect -800 16144 1919 16146
rect -800 16088 1858 16144
rect 1914 16088 1919 16144
rect -800 16086 1919 16088
rect -800 16056 800 16086
rect 1853 16083 1919 16086
rect 25221 16144 25330 16149
rect 25221 16088 25226 16144
rect 25282 16088 25330 16144
rect 25221 16086 25330 16088
rect 26233 16146 26299 16149
rect 29200 16146 30800 16176
rect 26233 16144 30800 16146
rect 26233 16088 26238 16144
rect 26294 16088 30800 16144
rect 26233 16086 30800 16088
rect 25221 16083 25287 16086
rect 26233 16083 26299 16086
rect 29200 16056 30800 16086
rect 10208 15808 10528 15809
rect -800 15738 800 15768
rect 10208 15744 10216 15808
rect 10280 15744 10296 15808
rect 10360 15744 10376 15808
rect 10440 15744 10456 15808
rect 10520 15744 10528 15808
rect 10208 15743 10528 15744
rect 19472 15808 19792 15809
rect 19472 15744 19480 15808
rect 19544 15744 19560 15808
rect 19624 15744 19640 15808
rect 19704 15744 19720 15808
rect 19784 15744 19792 15808
rect 19472 15743 19792 15744
rect 1853 15738 1919 15741
rect -800 15736 1919 15738
rect -800 15680 1858 15736
rect 1914 15680 1919 15736
rect -800 15678 1919 15680
rect -800 15648 800 15678
rect 1853 15675 1919 15678
rect 25957 15738 26023 15741
rect 29200 15738 30800 15768
rect 25957 15736 30800 15738
rect 25957 15680 25962 15736
rect 26018 15680 30800 15736
rect 25957 15678 30800 15680
rect 25957 15675 26023 15678
rect 29200 15648 30800 15678
rect 18965 15602 19031 15605
rect 25221 15602 25287 15605
rect 18965 15600 25287 15602
rect 18965 15544 18970 15600
rect 19026 15544 25226 15600
rect 25282 15544 25287 15600
rect 18965 15542 25287 15544
rect 18965 15539 19031 15542
rect 25221 15539 25287 15542
rect -800 15330 800 15360
rect 3325 15330 3391 15333
rect -800 15328 3391 15330
rect -800 15272 3330 15328
rect 3386 15272 3391 15328
rect -800 15270 3391 15272
rect -800 15240 800 15270
rect 3325 15267 3391 15270
rect 26877 15330 26943 15333
rect 29200 15330 30800 15360
rect 26877 15328 30800 15330
rect 26877 15272 26882 15328
rect 26938 15272 30800 15328
rect 26877 15270 30800 15272
rect 26877 15267 26943 15270
rect 5576 15264 5896 15265
rect 5576 15200 5584 15264
rect 5648 15200 5664 15264
rect 5728 15200 5744 15264
rect 5808 15200 5824 15264
rect 5888 15200 5896 15264
rect 5576 15199 5896 15200
rect 14840 15264 15160 15265
rect 14840 15200 14848 15264
rect 14912 15200 14928 15264
rect 14992 15200 15008 15264
rect 15072 15200 15088 15264
rect 15152 15200 15160 15264
rect 14840 15199 15160 15200
rect 24104 15264 24424 15265
rect 24104 15200 24112 15264
rect 24176 15200 24192 15264
rect 24256 15200 24272 15264
rect 24336 15200 24352 15264
rect 24416 15200 24424 15264
rect 29200 15240 30800 15270
rect 24104 15199 24424 15200
rect 1945 15058 2011 15061
rect 2497 15058 2563 15061
rect 5165 15058 5231 15061
rect 1945 15056 5231 15058
rect 1945 15000 1950 15056
rect 2006 15000 2502 15056
rect 2558 15000 5170 15056
rect 5226 15000 5231 15056
rect 1945 14998 5231 15000
rect 1945 14995 2011 14998
rect 2497 14995 2563 14998
rect 5165 14995 5231 14998
rect -800 14922 800 14952
rect 4061 14922 4127 14925
rect 29200 14922 30800 14952
rect -800 14920 4127 14922
rect -800 14864 4066 14920
rect 4122 14864 4127 14920
rect -800 14862 4127 14864
rect -800 14832 800 14862
rect 4061 14859 4127 14862
rect 27478 14862 30800 14922
rect 27478 14789 27538 14862
rect 29200 14832 30800 14862
rect 27429 14784 27538 14789
rect 27429 14728 27434 14784
rect 27490 14728 27538 14784
rect 27429 14726 27538 14728
rect 27429 14723 27495 14726
rect 10208 14720 10528 14721
rect 10208 14656 10216 14720
rect 10280 14656 10296 14720
rect 10360 14656 10376 14720
rect 10440 14656 10456 14720
rect 10520 14656 10528 14720
rect 10208 14655 10528 14656
rect 19472 14720 19792 14721
rect 19472 14656 19480 14720
rect 19544 14656 19560 14720
rect 19624 14656 19640 14720
rect 19704 14656 19720 14720
rect 19784 14656 19792 14720
rect 19472 14655 19792 14656
rect 2497 14650 2563 14653
rect 7373 14650 7439 14653
rect 2497 14648 7439 14650
rect 2497 14592 2502 14648
rect 2558 14592 7378 14648
rect 7434 14592 7439 14648
rect 2497 14590 7439 14592
rect 2497 14587 2563 14590
rect 7373 14587 7439 14590
rect -800 14514 800 14544
rect 3417 14514 3483 14517
rect -800 14512 3483 14514
rect -800 14456 3422 14512
rect 3478 14456 3483 14512
rect -800 14454 3483 14456
rect -800 14424 800 14454
rect 3417 14451 3483 14454
rect 27521 14514 27587 14517
rect 29200 14514 30800 14544
rect 27521 14512 30800 14514
rect 27521 14456 27526 14512
rect 27582 14456 30800 14512
rect 27521 14454 30800 14456
rect 27521 14451 27587 14454
rect 29200 14424 30800 14454
rect 5576 14176 5896 14177
rect -800 14106 800 14136
rect 5576 14112 5584 14176
rect 5648 14112 5664 14176
rect 5728 14112 5744 14176
rect 5808 14112 5824 14176
rect 5888 14112 5896 14176
rect 5576 14111 5896 14112
rect 14840 14176 15160 14177
rect 14840 14112 14848 14176
rect 14912 14112 14928 14176
rect 14992 14112 15008 14176
rect 15072 14112 15088 14176
rect 15152 14112 15160 14176
rect 14840 14111 15160 14112
rect 24104 14176 24424 14177
rect 24104 14112 24112 14176
rect 24176 14112 24192 14176
rect 24256 14112 24272 14176
rect 24336 14112 24352 14176
rect 24416 14112 24424 14176
rect 24104 14111 24424 14112
rect 2773 14106 2839 14109
rect -800 14104 2839 14106
rect -800 14048 2778 14104
rect 2834 14048 2839 14104
rect -800 14046 2839 14048
rect -800 14016 800 14046
rect 2773 14043 2839 14046
rect 28165 14106 28231 14109
rect 29200 14106 30800 14136
rect 28165 14104 30800 14106
rect 28165 14048 28170 14104
rect 28226 14048 30800 14104
rect 28165 14046 30800 14048
rect 28165 14043 28231 14046
rect 29200 14016 30800 14046
rect -800 13698 800 13728
rect 3049 13698 3115 13701
rect -800 13696 3115 13698
rect -800 13640 3054 13696
rect 3110 13640 3115 13696
rect -800 13638 3115 13640
rect -800 13608 800 13638
rect 3049 13635 3115 13638
rect 28165 13698 28231 13701
rect 29200 13698 30800 13728
rect 28165 13696 30800 13698
rect 28165 13640 28170 13696
rect 28226 13640 30800 13696
rect 28165 13638 30800 13640
rect 28165 13635 28231 13638
rect 10208 13632 10528 13633
rect 10208 13568 10216 13632
rect 10280 13568 10296 13632
rect 10360 13568 10376 13632
rect 10440 13568 10456 13632
rect 10520 13568 10528 13632
rect 10208 13567 10528 13568
rect 19472 13632 19792 13633
rect 19472 13568 19480 13632
rect 19544 13568 19560 13632
rect 19624 13568 19640 13632
rect 19704 13568 19720 13632
rect 19784 13568 19792 13632
rect 29200 13608 30800 13638
rect 19472 13567 19792 13568
rect -800 13290 800 13320
rect 1945 13290 2011 13293
rect -800 13288 2011 13290
rect -800 13232 1950 13288
rect 2006 13232 2011 13288
rect -800 13230 2011 13232
rect -800 13200 800 13230
rect 1945 13227 2011 13230
rect 11605 13290 11671 13293
rect 19149 13290 19215 13293
rect 11605 13288 19215 13290
rect 11605 13232 11610 13288
rect 11666 13232 19154 13288
rect 19210 13232 19215 13288
rect 11605 13230 19215 13232
rect 11605 13227 11671 13230
rect 19149 13227 19215 13230
rect 28165 13290 28231 13293
rect 29200 13290 30800 13320
rect 28165 13288 30800 13290
rect 28165 13232 28170 13288
rect 28226 13232 30800 13288
rect 28165 13230 30800 13232
rect 28165 13227 28231 13230
rect 29200 13200 30800 13230
rect 5576 13088 5896 13089
rect 5576 13024 5584 13088
rect 5648 13024 5664 13088
rect 5728 13024 5744 13088
rect 5808 13024 5824 13088
rect 5888 13024 5896 13088
rect 5576 13023 5896 13024
rect 14840 13088 15160 13089
rect 14840 13024 14848 13088
rect 14912 13024 14928 13088
rect 14992 13024 15008 13088
rect 15072 13024 15088 13088
rect 15152 13024 15160 13088
rect 14840 13023 15160 13024
rect 24104 13088 24424 13089
rect 24104 13024 24112 13088
rect 24176 13024 24192 13088
rect 24256 13024 24272 13088
rect 24336 13024 24352 13088
rect 24416 13024 24424 13088
rect 24104 13023 24424 13024
rect -800 12882 800 12912
rect 1853 12882 1919 12885
rect -800 12880 1919 12882
rect -800 12824 1858 12880
rect 1914 12824 1919 12880
rect -800 12822 1919 12824
rect -800 12792 800 12822
rect 1853 12819 1919 12822
rect 25957 12882 26023 12885
rect 29200 12882 30800 12912
rect 25957 12880 30800 12882
rect 25957 12824 25962 12880
rect 26018 12824 30800 12880
rect 25957 12822 30800 12824
rect 25957 12819 26023 12822
rect 29200 12792 30800 12822
rect 16389 12610 16455 12613
rect 17401 12610 17467 12613
rect 16389 12608 17467 12610
rect 16389 12552 16394 12608
rect 16450 12552 17406 12608
rect 17462 12552 17467 12608
rect 16389 12550 17467 12552
rect 16389 12547 16455 12550
rect 17401 12547 17467 12550
rect 18597 12610 18663 12613
rect 18781 12610 18847 12613
rect 18597 12608 18847 12610
rect 18597 12552 18602 12608
rect 18658 12552 18786 12608
rect 18842 12552 18847 12608
rect 18597 12550 18847 12552
rect 18597 12547 18663 12550
rect 18781 12547 18847 12550
rect 10208 12544 10528 12545
rect -800 12474 800 12504
rect 10208 12480 10216 12544
rect 10280 12480 10296 12544
rect 10360 12480 10376 12544
rect 10440 12480 10456 12544
rect 10520 12480 10528 12544
rect 10208 12479 10528 12480
rect 19472 12544 19792 12545
rect 19472 12480 19480 12544
rect 19544 12480 19560 12544
rect 19624 12480 19640 12544
rect 19704 12480 19720 12544
rect 19784 12480 19792 12544
rect 19472 12479 19792 12480
rect 1853 12474 1919 12477
rect -800 12472 1919 12474
rect -800 12416 1858 12472
rect 1914 12416 1919 12472
rect -800 12414 1919 12416
rect -800 12384 800 12414
rect 1853 12411 1919 12414
rect 25589 12474 25655 12477
rect 29200 12474 30800 12504
rect 25589 12472 30800 12474
rect 25589 12416 25594 12472
rect 25650 12416 30800 12472
rect 25589 12414 30800 12416
rect 25589 12411 25655 12414
rect 29200 12384 30800 12414
rect 11605 12338 11671 12341
rect 16573 12338 16639 12341
rect 11605 12336 16639 12338
rect 11605 12280 11610 12336
rect 11666 12280 16578 12336
rect 16634 12280 16639 12336
rect 11605 12278 16639 12280
rect 11605 12275 11671 12278
rect 16573 12275 16639 12278
rect 18597 12338 18663 12341
rect 20253 12338 20319 12341
rect 18597 12336 20319 12338
rect 18597 12280 18602 12336
rect 18658 12280 20258 12336
rect 20314 12280 20319 12336
rect 18597 12278 20319 12280
rect 18597 12275 18663 12278
rect 20253 12275 20319 12278
rect -800 12066 800 12096
rect 2773 12066 2839 12069
rect -800 12064 2839 12066
rect -800 12008 2778 12064
rect 2834 12008 2839 12064
rect -800 12006 2839 12008
rect -800 11976 800 12006
rect 2773 12003 2839 12006
rect 26785 12066 26851 12069
rect 29200 12066 30800 12096
rect 26785 12064 30800 12066
rect 26785 12008 26790 12064
rect 26846 12008 30800 12064
rect 26785 12006 30800 12008
rect 26785 12003 26851 12006
rect 5576 12000 5896 12001
rect 5576 11936 5584 12000
rect 5648 11936 5664 12000
rect 5728 11936 5744 12000
rect 5808 11936 5824 12000
rect 5888 11936 5896 12000
rect 5576 11935 5896 11936
rect 14840 12000 15160 12001
rect 14840 11936 14848 12000
rect 14912 11936 14928 12000
rect 14992 11936 15008 12000
rect 15072 11936 15088 12000
rect 15152 11936 15160 12000
rect 14840 11935 15160 11936
rect 24104 12000 24424 12001
rect 24104 11936 24112 12000
rect 24176 11936 24192 12000
rect 24256 11936 24272 12000
rect 24336 11936 24352 12000
rect 24416 11936 24424 12000
rect 29200 11976 30800 12006
rect 24104 11935 24424 11936
rect -800 11658 800 11688
rect 2405 11658 2471 11661
rect 13445 11658 13511 11661
rect -800 11656 2471 11658
rect -800 11600 2410 11656
rect 2466 11600 2471 11656
rect -800 11598 2471 11600
rect -800 11568 800 11598
rect 2405 11595 2471 11598
rect 13310 11656 13511 11658
rect 13310 11600 13450 11656
rect 13506 11600 13511 11656
rect 13310 11598 13511 11600
rect 13310 11525 13370 11598
rect 13445 11595 13511 11598
rect 26141 11658 26207 11661
rect 29200 11658 30800 11688
rect 26141 11656 30800 11658
rect 26141 11600 26146 11656
rect 26202 11600 30800 11656
rect 26141 11598 30800 11600
rect 26141 11595 26207 11598
rect 29200 11568 30800 11598
rect 13261 11520 13370 11525
rect 13261 11464 13266 11520
rect 13322 11464 13370 11520
rect 13261 11462 13370 11464
rect 13261 11459 13327 11462
rect 10208 11456 10528 11457
rect 10208 11392 10216 11456
rect 10280 11392 10296 11456
rect 10360 11392 10376 11456
rect 10440 11392 10456 11456
rect 10520 11392 10528 11456
rect 10208 11391 10528 11392
rect 19472 11456 19792 11457
rect 19472 11392 19480 11456
rect 19544 11392 19560 11456
rect 19624 11392 19640 11456
rect 19704 11392 19720 11456
rect 19784 11392 19792 11456
rect 19472 11391 19792 11392
rect -800 11250 800 11280
rect 2773 11250 2839 11253
rect -800 11248 2839 11250
rect -800 11192 2778 11248
rect 2834 11192 2839 11248
rect -800 11190 2839 11192
rect -800 11160 800 11190
rect 2773 11187 2839 11190
rect 26141 11250 26207 11253
rect 29200 11250 30800 11280
rect 26141 11248 30800 11250
rect 26141 11192 26146 11248
rect 26202 11192 30800 11248
rect 26141 11190 30800 11192
rect 26141 11187 26207 11190
rect 29200 11160 30800 11190
rect 5576 10912 5896 10913
rect -800 10842 800 10872
rect 5576 10848 5584 10912
rect 5648 10848 5664 10912
rect 5728 10848 5744 10912
rect 5808 10848 5824 10912
rect 5888 10848 5896 10912
rect 5576 10847 5896 10848
rect 14840 10912 15160 10913
rect 14840 10848 14848 10912
rect 14912 10848 14928 10912
rect 14992 10848 15008 10912
rect 15072 10848 15088 10912
rect 15152 10848 15160 10912
rect 14840 10847 15160 10848
rect 24104 10912 24424 10913
rect 24104 10848 24112 10912
rect 24176 10848 24192 10912
rect 24256 10848 24272 10912
rect 24336 10848 24352 10912
rect 24416 10848 24424 10912
rect 24104 10847 24424 10848
rect 1485 10842 1551 10845
rect -800 10840 1551 10842
rect -800 10784 1490 10840
rect 1546 10784 1551 10840
rect -800 10782 1551 10784
rect -800 10752 800 10782
rect 1485 10779 1551 10782
rect 28993 10842 29059 10845
rect 29200 10842 30800 10872
rect 28993 10840 30800 10842
rect 28993 10784 28998 10840
rect 29054 10784 30800 10840
rect 28993 10782 30800 10784
rect 28993 10779 29059 10782
rect 29200 10752 30800 10782
rect 13169 10706 13235 10709
rect 13126 10704 13235 10706
rect 13126 10648 13174 10704
rect 13230 10648 13235 10704
rect 13126 10643 13235 10648
rect 18413 10704 18479 10709
rect 18413 10648 18418 10704
rect 18474 10648 18479 10704
rect 18413 10643 18479 10648
rect -800 10434 800 10464
rect 1945 10434 2011 10437
rect -800 10432 2011 10434
rect -800 10376 1950 10432
rect 2006 10376 2011 10432
rect -800 10374 2011 10376
rect -800 10344 800 10374
rect 1945 10371 2011 10374
rect 12801 10434 12867 10437
rect 13126 10434 13186 10643
rect 15929 10570 15995 10573
rect 18416 10570 18476 10643
rect 15929 10568 18476 10570
rect 15929 10512 15934 10568
rect 15990 10512 18476 10568
rect 15929 10510 18476 10512
rect 15929 10507 15995 10510
rect 12801 10432 13186 10434
rect 12801 10376 12806 10432
rect 12862 10376 13186 10432
rect 12801 10374 13186 10376
rect 18137 10434 18203 10437
rect 18137 10432 18338 10434
rect 18137 10376 18142 10432
rect 18198 10376 18338 10432
rect 18137 10374 18338 10376
rect 12801 10371 12867 10374
rect 18137 10371 18203 10374
rect 10208 10368 10528 10369
rect 10208 10304 10216 10368
rect 10280 10304 10296 10368
rect 10360 10304 10376 10368
rect 10440 10304 10456 10368
rect 10520 10304 10528 10368
rect 10208 10303 10528 10304
rect -800 10026 800 10056
rect 1577 10026 1643 10029
rect -800 10024 1643 10026
rect -800 9968 1582 10024
rect 1638 9968 1643 10024
rect -800 9966 1643 9968
rect -800 9936 800 9966
rect 1577 9963 1643 9966
rect 18278 9890 18338 10374
rect 18416 10029 18476 10510
rect 26877 10434 26943 10437
rect 29200 10434 30800 10464
rect 26877 10432 30800 10434
rect 26877 10376 26882 10432
rect 26938 10376 30800 10432
rect 26877 10374 30800 10376
rect 26877 10371 26943 10374
rect 19472 10368 19792 10369
rect 19472 10304 19480 10368
rect 19544 10304 19560 10368
rect 19624 10304 19640 10368
rect 19704 10304 19720 10368
rect 19784 10304 19792 10368
rect 29200 10344 30800 10374
rect 19472 10303 19792 10304
rect 18413 10024 18479 10029
rect 18413 9968 18418 10024
rect 18474 9968 18479 10024
rect 18413 9963 18479 9968
rect 27521 10026 27587 10029
rect 29200 10026 30800 10056
rect 27521 10024 30800 10026
rect 27521 9968 27526 10024
rect 27582 9968 30800 10024
rect 27521 9966 30800 9968
rect 27521 9963 27587 9966
rect 29200 9936 30800 9966
rect 19241 9890 19307 9893
rect 18278 9888 19307 9890
rect 18278 9832 19246 9888
rect 19302 9832 19307 9888
rect 18278 9830 19307 9832
rect 19241 9827 19307 9830
rect 5576 9824 5896 9825
rect 5576 9760 5584 9824
rect 5648 9760 5664 9824
rect 5728 9760 5744 9824
rect 5808 9760 5824 9824
rect 5888 9760 5896 9824
rect 5576 9759 5896 9760
rect 14840 9824 15160 9825
rect 14840 9760 14848 9824
rect 14912 9760 14928 9824
rect 14992 9760 15008 9824
rect 15072 9760 15088 9824
rect 15152 9760 15160 9824
rect 14840 9759 15160 9760
rect 24104 9824 24424 9825
rect 24104 9760 24112 9824
rect 24176 9760 24192 9824
rect 24256 9760 24272 9824
rect 24336 9760 24352 9824
rect 24416 9760 24424 9824
rect 24104 9759 24424 9760
rect -800 9618 800 9648
rect 1853 9618 1919 9621
rect -800 9616 1919 9618
rect -800 9560 1858 9616
rect 1914 9560 1919 9616
rect -800 9558 1919 9560
rect -800 9528 800 9558
rect 1853 9555 1919 9558
rect 24853 9618 24919 9621
rect 29200 9618 30800 9648
rect 24853 9616 30800 9618
rect 24853 9560 24858 9616
rect 24914 9560 30800 9616
rect 24853 9558 30800 9560
rect 24853 9555 24919 9558
rect 29200 9528 30800 9558
rect 11513 9482 11579 9485
rect 18873 9482 18939 9485
rect 11513 9480 18939 9482
rect 11513 9424 11518 9480
rect 11574 9424 18878 9480
rect 18934 9424 18939 9480
rect 11513 9422 18939 9424
rect 11513 9419 11579 9422
rect 18873 9419 18939 9422
rect 10208 9280 10528 9281
rect -800 9210 800 9240
rect 10208 9216 10216 9280
rect 10280 9216 10296 9280
rect 10360 9216 10376 9280
rect 10440 9216 10456 9280
rect 10520 9216 10528 9280
rect 10208 9215 10528 9216
rect 19472 9280 19792 9281
rect 19472 9216 19480 9280
rect 19544 9216 19560 9280
rect 19624 9216 19640 9280
rect 19704 9216 19720 9280
rect 19784 9216 19792 9280
rect 19472 9215 19792 9216
rect 2865 9210 2931 9213
rect -800 9208 2931 9210
rect -800 9152 2870 9208
rect 2926 9152 2931 9208
rect -800 9150 2931 9152
rect -800 9120 800 9150
rect 2865 9147 2931 9150
rect 26141 9210 26207 9213
rect 29200 9210 30800 9240
rect 26141 9208 30800 9210
rect 26141 9152 26146 9208
rect 26202 9152 30800 9208
rect 26141 9150 30800 9152
rect 26141 9147 26207 9150
rect 29200 9120 30800 9150
rect 11605 8938 11671 8941
rect 15101 8938 15167 8941
rect 18965 8938 19031 8941
rect 11605 8936 19031 8938
rect 11605 8880 11610 8936
rect 11666 8880 15106 8936
rect 15162 8880 18970 8936
rect 19026 8880 19031 8936
rect 11605 8878 19031 8880
rect 11605 8875 11671 8878
rect 15101 8875 15167 8878
rect 18965 8875 19031 8878
rect -800 8802 800 8832
rect 3233 8802 3299 8805
rect -800 8800 3299 8802
rect -800 8744 3238 8800
rect 3294 8744 3299 8800
rect -800 8742 3299 8744
rect -800 8712 800 8742
rect 3233 8739 3299 8742
rect 24945 8802 25011 8805
rect 29200 8802 30800 8832
rect 24945 8800 30800 8802
rect 24945 8744 24950 8800
rect 25006 8744 30800 8800
rect 24945 8742 30800 8744
rect 24945 8739 25011 8742
rect 5576 8736 5896 8737
rect 5576 8672 5584 8736
rect 5648 8672 5664 8736
rect 5728 8672 5744 8736
rect 5808 8672 5824 8736
rect 5888 8672 5896 8736
rect 5576 8671 5896 8672
rect 14840 8736 15160 8737
rect 14840 8672 14848 8736
rect 14912 8672 14928 8736
rect 14992 8672 15008 8736
rect 15072 8672 15088 8736
rect 15152 8672 15160 8736
rect 14840 8671 15160 8672
rect 24104 8736 24424 8737
rect 24104 8672 24112 8736
rect 24176 8672 24192 8736
rect 24256 8672 24272 8736
rect 24336 8672 24352 8736
rect 24416 8672 24424 8736
rect 29200 8712 30800 8742
rect 24104 8671 24424 8672
rect -800 8394 800 8424
rect 2405 8394 2471 8397
rect -800 8392 2471 8394
rect -800 8336 2410 8392
rect 2466 8336 2471 8392
rect -800 8334 2471 8336
rect -800 8304 800 8334
rect 2405 8331 2471 8334
rect 25865 8394 25931 8397
rect 29200 8394 30800 8424
rect 25865 8392 30800 8394
rect 25865 8336 25870 8392
rect 25926 8336 30800 8392
rect 25865 8334 30800 8336
rect 25865 8331 25931 8334
rect 29200 8304 30800 8334
rect 10208 8192 10528 8193
rect 10208 8128 10216 8192
rect 10280 8128 10296 8192
rect 10360 8128 10376 8192
rect 10440 8128 10456 8192
rect 10520 8128 10528 8192
rect 10208 8127 10528 8128
rect 19472 8192 19792 8193
rect 19472 8128 19480 8192
rect 19544 8128 19560 8192
rect 19624 8128 19640 8192
rect 19704 8128 19720 8192
rect 19784 8128 19792 8192
rect 19472 8127 19792 8128
rect -800 7986 800 8016
rect 2405 7986 2471 7989
rect -800 7984 2471 7986
rect -800 7928 2410 7984
rect 2466 7928 2471 7984
rect -800 7926 2471 7928
rect -800 7896 800 7926
rect 2405 7923 2471 7926
rect 10225 7986 10291 7989
rect 12525 7986 12591 7989
rect 10225 7984 12591 7986
rect 10225 7928 10230 7984
rect 10286 7928 12530 7984
rect 12586 7928 12591 7984
rect 10225 7926 12591 7928
rect 10225 7923 10291 7926
rect 12525 7923 12591 7926
rect 28073 7986 28139 7989
rect 29200 7986 30800 8016
rect 28073 7984 30800 7986
rect 28073 7928 28078 7984
rect 28134 7928 30800 7984
rect 28073 7926 30800 7928
rect 28073 7923 28139 7926
rect 29200 7896 30800 7926
rect 5576 7648 5896 7649
rect -800 7578 800 7608
rect 5576 7584 5584 7648
rect 5648 7584 5664 7648
rect 5728 7584 5744 7648
rect 5808 7584 5824 7648
rect 5888 7584 5896 7648
rect 5576 7583 5896 7584
rect 14840 7648 15160 7649
rect 14840 7584 14848 7648
rect 14912 7584 14928 7648
rect 14992 7584 15008 7648
rect 15072 7584 15088 7648
rect 15152 7584 15160 7648
rect 14840 7583 15160 7584
rect 24104 7648 24424 7649
rect 24104 7584 24112 7648
rect 24176 7584 24192 7648
rect 24256 7584 24272 7648
rect 24336 7584 24352 7648
rect 24416 7584 24424 7648
rect 24104 7583 24424 7584
rect 1945 7578 2011 7581
rect -800 7576 2011 7578
rect -800 7520 1950 7576
rect 2006 7520 2011 7576
rect -800 7518 2011 7520
rect -800 7488 800 7518
rect 1945 7515 2011 7518
rect 26785 7578 26851 7581
rect 29200 7578 30800 7608
rect 26785 7576 30800 7578
rect 26785 7520 26790 7576
rect 26846 7520 30800 7576
rect 26785 7518 30800 7520
rect 26785 7515 26851 7518
rect 29200 7488 30800 7518
rect 8661 7306 8727 7309
rect 10685 7306 10751 7309
rect 8661 7304 10751 7306
rect 8661 7248 8666 7304
rect 8722 7248 10690 7304
rect 10746 7248 10751 7304
rect 8661 7246 10751 7248
rect 8661 7243 8727 7246
rect 10685 7243 10751 7246
rect 15009 7306 15075 7309
rect 15653 7306 15719 7309
rect 15009 7304 15719 7306
rect 15009 7248 15014 7304
rect 15070 7248 15658 7304
rect 15714 7248 15719 7304
rect 15009 7246 15719 7248
rect 15009 7243 15075 7246
rect 15653 7243 15719 7246
rect -800 7170 800 7200
rect 3049 7170 3115 7173
rect -800 7168 3115 7170
rect -800 7112 3054 7168
rect 3110 7112 3115 7168
rect -800 7110 3115 7112
rect -800 7080 800 7110
rect 3049 7107 3115 7110
rect 28165 7170 28231 7173
rect 29200 7170 30800 7200
rect 28165 7168 30800 7170
rect 28165 7112 28170 7168
rect 28226 7112 30800 7168
rect 28165 7110 30800 7112
rect 28165 7107 28231 7110
rect 10208 7104 10528 7105
rect 10208 7040 10216 7104
rect 10280 7040 10296 7104
rect 10360 7040 10376 7104
rect 10440 7040 10456 7104
rect 10520 7040 10528 7104
rect 10208 7039 10528 7040
rect 19472 7104 19792 7105
rect 19472 7040 19480 7104
rect 19544 7040 19560 7104
rect 19624 7040 19640 7104
rect 19704 7040 19720 7104
rect 19784 7040 19792 7104
rect 29200 7080 30800 7110
rect 19472 7039 19792 7040
rect -800 6762 800 6792
rect 1485 6762 1551 6765
rect -800 6760 1551 6762
rect -800 6704 1490 6760
rect 1546 6704 1551 6760
rect -800 6702 1551 6704
rect -800 6672 800 6702
rect 1485 6699 1551 6702
rect 28165 6762 28231 6765
rect 29200 6762 30800 6792
rect 28165 6760 30800 6762
rect 28165 6704 28170 6760
rect 28226 6704 30800 6760
rect 28165 6702 30800 6704
rect 28165 6699 28231 6702
rect 29200 6672 30800 6702
rect 5576 6560 5896 6561
rect 5576 6496 5584 6560
rect 5648 6496 5664 6560
rect 5728 6496 5744 6560
rect 5808 6496 5824 6560
rect 5888 6496 5896 6560
rect 5576 6495 5896 6496
rect 14840 6560 15160 6561
rect 14840 6496 14848 6560
rect 14912 6496 14928 6560
rect 14992 6496 15008 6560
rect 15072 6496 15088 6560
rect 15152 6496 15160 6560
rect 14840 6495 15160 6496
rect 24104 6560 24424 6561
rect 24104 6496 24112 6560
rect 24176 6496 24192 6560
rect 24256 6496 24272 6560
rect 24336 6496 24352 6560
rect 24416 6496 24424 6560
rect 24104 6495 24424 6496
rect -800 6354 800 6384
rect 4061 6354 4127 6357
rect -800 6352 4127 6354
rect -800 6296 4066 6352
rect 4122 6296 4127 6352
rect -800 6294 4127 6296
rect -800 6264 800 6294
rect 4061 6291 4127 6294
rect 25313 6354 25379 6357
rect 29200 6354 30800 6384
rect 25313 6352 30800 6354
rect 25313 6296 25318 6352
rect 25374 6296 30800 6352
rect 25313 6294 30800 6296
rect 25313 6291 25379 6294
rect 29200 6264 30800 6294
rect 10208 6016 10528 6017
rect -800 5946 800 5976
rect 10208 5952 10216 6016
rect 10280 5952 10296 6016
rect 10360 5952 10376 6016
rect 10440 5952 10456 6016
rect 10520 5952 10528 6016
rect 10208 5951 10528 5952
rect 19472 6016 19792 6017
rect 19472 5952 19480 6016
rect 19544 5952 19560 6016
rect 19624 5952 19640 6016
rect 19704 5952 19720 6016
rect 19784 5952 19792 6016
rect 19472 5951 19792 5952
rect 3693 5946 3759 5949
rect -800 5944 3759 5946
rect -800 5888 3698 5944
rect 3754 5888 3759 5944
rect -800 5886 3759 5888
rect -800 5856 800 5886
rect 3693 5883 3759 5886
rect 26049 5946 26115 5949
rect 29200 5946 30800 5976
rect 26049 5944 30800 5946
rect 26049 5888 26054 5944
rect 26110 5888 30800 5944
rect 26049 5886 30800 5888
rect 26049 5883 26115 5886
rect 29200 5856 30800 5886
rect 9949 5810 10015 5813
rect 16021 5810 16087 5813
rect 9949 5808 16087 5810
rect 9949 5752 9954 5808
rect 10010 5752 16026 5808
rect 16082 5752 16087 5808
rect 9949 5750 16087 5752
rect 9949 5747 10015 5750
rect 16021 5747 16087 5750
rect -800 5538 800 5568
rect 3969 5538 4035 5541
rect -800 5536 4035 5538
rect -800 5480 3974 5536
rect 4030 5480 4035 5536
rect -800 5478 4035 5480
rect -800 5448 800 5478
rect 3969 5475 4035 5478
rect 26877 5538 26943 5541
rect 29200 5538 30800 5568
rect 26877 5536 30800 5538
rect 26877 5480 26882 5536
rect 26938 5480 30800 5536
rect 26877 5478 30800 5480
rect 26877 5475 26943 5478
rect 5576 5472 5896 5473
rect 5576 5408 5584 5472
rect 5648 5408 5664 5472
rect 5728 5408 5744 5472
rect 5808 5408 5824 5472
rect 5888 5408 5896 5472
rect 5576 5407 5896 5408
rect 14840 5472 15160 5473
rect 14840 5408 14848 5472
rect 14912 5408 14928 5472
rect 14992 5408 15008 5472
rect 15072 5408 15088 5472
rect 15152 5408 15160 5472
rect 14840 5407 15160 5408
rect 24104 5472 24424 5473
rect 24104 5408 24112 5472
rect 24176 5408 24192 5472
rect 24256 5408 24272 5472
rect 24336 5408 24352 5472
rect 24416 5408 24424 5472
rect 29200 5448 30800 5478
rect 24104 5407 24424 5408
rect -800 5130 800 5160
rect 4061 5130 4127 5133
rect -800 5128 4127 5130
rect -800 5072 4066 5128
rect 4122 5072 4127 5128
rect -800 5070 4127 5072
rect -800 5040 800 5070
rect 4061 5067 4127 5070
rect 26601 5130 26667 5133
rect 29200 5130 30800 5160
rect 26601 5128 30800 5130
rect 26601 5072 26606 5128
rect 26662 5072 30800 5128
rect 26601 5070 30800 5072
rect 26601 5067 26667 5070
rect 29200 5040 30800 5070
rect 10208 4928 10528 4929
rect 10208 4864 10216 4928
rect 10280 4864 10296 4928
rect 10360 4864 10376 4928
rect 10440 4864 10456 4928
rect 10520 4864 10528 4928
rect 10208 4863 10528 4864
rect 19472 4928 19792 4929
rect 19472 4864 19480 4928
rect 19544 4864 19560 4928
rect 19624 4864 19640 4928
rect 19704 4864 19720 4928
rect 19784 4864 19792 4928
rect 19472 4863 19792 4864
rect -800 4722 800 4752
rect 4061 4722 4127 4725
rect -800 4720 4127 4722
rect -800 4664 4066 4720
rect 4122 4664 4127 4720
rect -800 4662 4127 4664
rect -800 4632 800 4662
rect 4061 4659 4127 4662
rect 27429 4722 27495 4725
rect 29200 4722 30800 4752
rect 27429 4720 30800 4722
rect 27429 4664 27434 4720
rect 27490 4664 30800 4720
rect 27429 4662 30800 4664
rect 27429 4659 27495 4662
rect 29200 4632 30800 4662
rect 5576 4384 5896 4385
rect -800 4314 800 4344
rect 5576 4320 5584 4384
rect 5648 4320 5664 4384
rect 5728 4320 5744 4384
rect 5808 4320 5824 4384
rect 5888 4320 5896 4384
rect 5576 4319 5896 4320
rect 14840 4384 15160 4385
rect 14840 4320 14848 4384
rect 14912 4320 14928 4384
rect 14992 4320 15008 4384
rect 15072 4320 15088 4384
rect 15152 4320 15160 4384
rect 14840 4319 15160 4320
rect 24104 4384 24424 4385
rect 24104 4320 24112 4384
rect 24176 4320 24192 4384
rect 24256 4320 24272 4384
rect 24336 4320 24352 4384
rect 24416 4320 24424 4384
rect 24104 4319 24424 4320
rect 3969 4314 4035 4317
rect -800 4312 4035 4314
rect -800 4256 3974 4312
rect 4030 4256 4035 4312
rect -800 4254 4035 4256
rect -800 4224 800 4254
rect 3969 4251 4035 4254
rect 26785 4314 26851 4317
rect 29200 4314 30800 4344
rect 26785 4312 30800 4314
rect 26785 4256 26790 4312
rect 26846 4256 30800 4312
rect 26785 4254 30800 4256
rect 26785 4251 26851 4254
rect 29200 4224 30800 4254
rect 12249 4178 12315 4181
rect 16481 4178 16547 4181
rect 12249 4176 16547 4178
rect 12249 4120 12254 4176
rect 12310 4120 16486 4176
rect 16542 4120 16547 4176
rect 12249 4118 16547 4120
rect 12249 4115 12315 4118
rect 16481 4115 16547 4118
rect 14089 4042 14155 4045
rect 15469 4042 15535 4045
rect 14089 4040 15535 4042
rect 14089 3984 14094 4040
rect 14150 3984 15474 4040
rect 15530 3984 15535 4040
rect 14089 3982 15535 3984
rect 14089 3979 14155 3982
rect 15469 3979 15535 3982
rect -800 3906 800 3936
rect 2773 3906 2839 3909
rect -800 3904 2839 3906
rect -800 3848 2778 3904
rect 2834 3848 2839 3904
rect -800 3846 2839 3848
rect -800 3816 800 3846
rect 2773 3843 2839 3846
rect 11329 3906 11395 3909
rect 14825 3906 14891 3909
rect 11329 3904 14891 3906
rect 11329 3848 11334 3904
rect 11390 3848 14830 3904
rect 14886 3848 14891 3904
rect 11329 3846 14891 3848
rect 11329 3843 11395 3846
rect 14825 3843 14891 3846
rect 28073 3906 28139 3909
rect 29200 3906 30800 3936
rect 28073 3904 30800 3906
rect 28073 3848 28078 3904
rect 28134 3848 30800 3904
rect 28073 3846 30800 3848
rect 28073 3843 28139 3846
rect 10208 3840 10528 3841
rect 10208 3776 10216 3840
rect 10280 3776 10296 3840
rect 10360 3776 10376 3840
rect 10440 3776 10456 3840
rect 10520 3776 10528 3840
rect 10208 3775 10528 3776
rect 19472 3840 19792 3841
rect 19472 3776 19480 3840
rect 19544 3776 19560 3840
rect 19624 3776 19640 3840
rect 19704 3776 19720 3840
rect 19784 3776 19792 3840
rect 29200 3816 30800 3846
rect 19472 3775 19792 3776
rect 16849 3634 16915 3637
rect 26141 3634 26207 3637
rect 16849 3632 26207 3634
rect 16849 3576 16854 3632
rect 16910 3576 26146 3632
rect 26202 3576 26207 3632
rect 16849 3574 26207 3576
rect 16849 3571 16915 3574
rect 26141 3571 26207 3574
rect -800 3498 800 3528
rect 1945 3498 2011 3501
rect -800 3496 2011 3498
rect -800 3440 1950 3496
rect 2006 3440 2011 3496
rect -800 3438 2011 3440
rect -800 3408 800 3438
rect 1945 3435 2011 3438
rect 28165 3498 28231 3501
rect 29200 3498 30800 3528
rect 28165 3496 30800 3498
rect 28165 3440 28170 3496
rect 28226 3440 30800 3496
rect 28165 3438 30800 3440
rect 28165 3435 28231 3438
rect 29200 3408 30800 3438
rect 5576 3296 5896 3297
rect 5576 3232 5584 3296
rect 5648 3232 5664 3296
rect 5728 3232 5744 3296
rect 5808 3232 5824 3296
rect 5888 3232 5896 3296
rect 5576 3231 5896 3232
rect 14840 3296 15160 3297
rect 14840 3232 14848 3296
rect 14912 3232 14928 3296
rect 14992 3232 15008 3296
rect 15072 3232 15088 3296
rect 15152 3232 15160 3296
rect 14840 3231 15160 3232
rect 24104 3296 24424 3297
rect 24104 3232 24112 3296
rect 24176 3232 24192 3296
rect 24256 3232 24272 3296
rect 24336 3232 24352 3296
rect 24416 3232 24424 3296
rect 24104 3231 24424 3232
rect -800 3090 800 3120
rect 1669 3090 1735 3093
rect -800 3088 1735 3090
rect -800 3032 1674 3088
rect 1730 3032 1735 3088
rect -800 3030 1735 3032
rect -800 3000 800 3030
rect 1669 3027 1735 3030
rect 25497 3090 25563 3093
rect 29200 3090 30800 3120
rect 25497 3088 30800 3090
rect 25497 3032 25502 3088
rect 25558 3032 30800 3088
rect 25497 3030 30800 3032
rect 25497 3027 25563 3030
rect 29200 3000 30800 3030
rect 21909 2954 21975 2957
rect 24025 2954 24091 2957
rect 26785 2954 26851 2957
rect 21909 2952 26851 2954
rect 21909 2896 21914 2952
rect 21970 2896 24030 2952
rect 24086 2896 26790 2952
rect 26846 2896 26851 2952
rect 21909 2894 26851 2896
rect 21909 2891 21975 2894
rect 24025 2891 24091 2894
rect 26785 2891 26851 2894
rect 21357 2818 21423 2821
rect 22001 2818 22067 2821
rect 21357 2816 22067 2818
rect 21357 2760 21362 2816
rect 21418 2760 22006 2816
rect 22062 2760 22067 2816
rect 21357 2758 22067 2760
rect 21357 2755 21423 2758
rect 22001 2755 22067 2758
rect 10208 2752 10528 2753
rect -800 2682 800 2712
rect 10208 2688 10216 2752
rect 10280 2688 10296 2752
rect 10360 2688 10376 2752
rect 10440 2688 10456 2752
rect 10520 2688 10528 2752
rect 10208 2687 10528 2688
rect 19472 2752 19792 2753
rect 19472 2688 19480 2752
rect 19544 2688 19560 2752
rect 19624 2688 19640 2752
rect 19704 2688 19720 2752
rect 19784 2688 19792 2752
rect 19472 2687 19792 2688
rect 3509 2682 3575 2685
rect -800 2680 3575 2682
rect -800 2624 3514 2680
rect 3570 2624 3575 2680
rect -800 2622 3575 2624
rect -800 2592 800 2622
rect 3509 2619 3575 2622
rect 24853 2682 24919 2685
rect 29200 2682 30800 2712
rect 24853 2680 30800 2682
rect 24853 2624 24858 2680
rect 24914 2624 30800 2680
rect 24853 2622 30800 2624
rect 24853 2619 24919 2622
rect 29200 2592 30800 2622
rect 20345 2546 20411 2549
rect 24485 2546 24551 2549
rect 20345 2544 24551 2546
rect 20345 2488 20350 2544
rect 20406 2488 24490 2544
rect 24546 2488 24551 2544
rect 20345 2486 24551 2488
rect 20345 2483 20411 2486
rect 24485 2483 24551 2486
rect -800 2274 800 2304
rect 3417 2274 3483 2277
rect -800 2272 3483 2274
rect -800 2216 3422 2272
rect 3478 2216 3483 2272
rect -800 2214 3483 2216
rect -800 2184 800 2214
rect 3417 2211 3483 2214
rect 25037 2274 25103 2277
rect 29200 2274 30800 2304
rect 25037 2272 30800 2274
rect 25037 2216 25042 2272
rect 25098 2216 30800 2272
rect 25037 2214 30800 2216
rect 25037 2211 25103 2214
rect 5576 2208 5896 2209
rect 5576 2144 5584 2208
rect 5648 2144 5664 2208
rect 5728 2144 5744 2208
rect 5808 2144 5824 2208
rect 5888 2144 5896 2208
rect 5576 2143 5896 2144
rect 14840 2208 15160 2209
rect 14840 2144 14848 2208
rect 14912 2144 14928 2208
rect 14992 2144 15008 2208
rect 15072 2144 15088 2208
rect 15152 2144 15160 2208
rect 14840 2143 15160 2144
rect 24104 2208 24424 2209
rect 24104 2144 24112 2208
rect 24176 2144 24192 2208
rect 24256 2144 24272 2208
rect 24336 2144 24352 2208
rect 24416 2144 24424 2208
rect 29200 2184 30800 2214
rect 24104 2143 24424 2144
rect -800 1866 800 1896
rect 3417 1866 3483 1869
rect -800 1864 3483 1866
rect -800 1808 3422 1864
rect 3478 1808 3483 1864
rect -800 1806 3483 1808
rect -800 1776 800 1806
rect 3417 1803 3483 1806
rect 25405 1866 25471 1869
rect 29200 1866 30800 1896
rect 25405 1864 30800 1866
rect 25405 1808 25410 1864
rect 25466 1808 30800 1864
rect 25405 1806 30800 1808
rect 25405 1803 25471 1806
rect 29200 1776 30800 1806
rect -800 1458 800 1488
rect 2773 1458 2839 1461
rect -800 1456 2839 1458
rect -800 1400 2778 1456
rect 2834 1400 2839 1456
rect -800 1398 2839 1400
rect -800 1368 800 1398
rect 2773 1395 2839 1398
rect 26969 1458 27035 1461
rect 29200 1458 30800 1488
rect 26969 1456 30800 1458
rect 26969 1400 26974 1456
rect 27030 1400 30800 1456
rect 26969 1398 30800 1400
rect 26969 1395 27035 1398
rect 29200 1368 30800 1398
rect -800 1050 800 1080
rect 3233 1050 3299 1053
rect -800 1048 3299 1050
rect -800 992 3238 1048
rect 3294 992 3299 1048
rect -800 990 3299 992
rect -800 960 800 990
rect 3233 987 3299 990
rect 25865 1050 25931 1053
rect 29200 1050 30800 1080
rect 25865 1048 30800 1050
rect 25865 992 25870 1048
rect 25926 992 30800 1048
rect 25865 990 30800 992
rect 25865 987 25931 990
rect 29200 960 30800 990
rect -800 642 800 672
rect 2957 642 3023 645
rect -800 640 3023 642
rect -800 584 2962 640
rect 3018 584 3023 640
rect -800 582 3023 584
rect -800 552 800 582
rect 2957 579 3023 582
rect 26141 642 26207 645
rect 29200 642 30800 672
rect 26141 640 30800 642
rect 26141 584 26146 640
rect 26202 584 30800 640
rect 26141 582 30800 584
rect 26141 579 26207 582
rect 29200 552 30800 582
rect -800 234 800 264
rect 1393 234 1459 237
rect -800 232 1459 234
rect -800 176 1398 232
rect 1454 176 1459 232
rect -800 174 1459 176
rect -800 144 800 174
rect 1393 171 1459 174
rect 26049 234 26115 237
rect 29200 234 30800 264
rect 26049 232 30800 234
rect 26049 176 26054 232
rect 26110 176 30800 232
rect 26049 174 30800 176
rect 26049 171 26115 174
rect 29200 144 30800 174
<< via3 >>
rect 5584 53340 5648 53344
rect 5584 53284 5588 53340
rect 5588 53284 5644 53340
rect 5644 53284 5648 53340
rect 5584 53280 5648 53284
rect 5664 53340 5728 53344
rect 5664 53284 5668 53340
rect 5668 53284 5724 53340
rect 5724 53284 5728 53340
rect 5664 53280 5728 53284
rect 5744 53340 5808 53344
rect 5744 53284 5748 53340
rect 5748 53284 5804 53340
rect 5804 53284 5808 53340
rect 5744 53280 5808 53284
rect 5824 53340 5888 53344
rect 5824 53284 5828 53340
rect 5828 53284 5884 53340
rect 5884 53284 5888 53340
rect 5824 53280 5888 53284
rect 14848 53340 14912 53344
rect 14848 53284 14852 53340
rect 14852 53284 14908 53340
rect 14908 53284 14912 53340
rect 14848 53280 14912 53284
rect 14928 53340 14992 53344
rect 14928 53284 14932 53340
rect 14932 53284 14988 53340
rect 14988 53284 14992 53340
rect 14928 53280 14992 53284
rect 15008 53340 15072 53344
rect 15008 53284 15012 53340
rect 15012 53284 15068 53340
rect 15068 53284 15072 53340
rect 15008 53280 15072 53284
rect 15088 53340 15152 53344
rect 15088 53284 15092 53340
rect 15092 53284 15148 53340
rect 15148 53284 15152 53340
rect 15088 53280 15152 53284
rect 24112 53340 24176 53344
rect 24112 53284 24116 53340
rect 24116 53284 24172 53340
rect 24172 53284 24176 53340
rect 24112 53280 24176 53284
rect 24192 53340 24256 53344
rect 24192 53284 24196 53340
rect 24196 53284 24252 53340
rect 24252 53284 24256 53340
rect 24192 53280 24256 53284
rect 24272 53340 24336 53344
rect 24272 53284 24276 53340
rect 24276 53284 24332 53340
rect 24332 53284 24336 53340
rect 24272 53280 24336 53284
rect 24352 53340 24416 53344
rect 24352 53284 24356 53340
rect 24356 53284 24412 53340
rect 24412 53284 24416 53340
rect 24352 53280 24416 53284
rect 10216 52796 10280 52800
rect 10216 52740 10220 52796
rect 10220 52740 10276 52796
rect 10276 52740 10280 52796
rect 10216 52736 10280 52740
rect 10296 52796 10360 52800
rect 10296 52740 10300 52796
rect 10300 52740 10356 52796
rect 10356 52740 10360 52796
rect 10296 52736 10360 52740
rect 10376 52796 10440 52800
rect 10376 52740 10380 52796
rect 10380 52740 10436 52796
rect 10436 52740 10440 52796
rect 10376 52736 10440 52740
rect 10456 52796 10520 52800
rect 10456 52740 10460 52796
rect 10460 52740 10516 52796
rect 10516 52740 10520 52796
rect 10456 52736 10520 52740
rect 19480 52796 19544 52800
rect 19480 52740 19484 52796
rect 19484 52740 19540 52796
rect 19540 52740 19544 52796
rect 19480 52736 19544 52740
rect 19560 52796 19624 52800
rect 19560 52740 19564 52796
rect 19564 52740 19620 52796
rect 19620 52740 19624 52796
rect 19560 52736 19624 52740
rect 19640 52796 19704 52800
rect 19640 52740 19644 52796
rect 19644 52740 19700 52796
rect 19700 52740 19704 52796
rect 19640 52736 19704 52740
rect 19720 52796 19784 52800
rect 19720 52740 19724 52796
rect 19724 52740 19780 52796
rect 19780 52740 19784 52796
rect 19720 52736 19784 52740
rect 5584 52252 5648 52256
rect 5584 52196 5588 52252
rect 5588 52196 5644 52252
rect 5644 52196 5648 52252
rect 5584 52192 5648 52196
rect 5664 52252 5728 52256
rect 5664 52196 5668 52252
rect 5668 52196 5724 52252
rect 5724 52196 5728 52252
rect 5664 52192 5728 52196
rect 5744 52252 5808 52256
rect 5744 52196 5748 52252
rect 5748 52196 5804 52252
rect 5804 52196 5808 52252
rect 5744 52192 5808 52196
rect 5824 52252 5888 52256
rect 5824 52196 5828 52252
rect 5828 52196 5884 52252
rect 5884 52196 5888 52252
rect 5824 52192 5888 52196
rect 14848 52252 14912 52256
rect 14848 52196 14852 52252
rect 14852 52196 14908 52252
rect 14908 52196 14912 52252
rect 14848 52192 14912 52196
rect 14928 52252 14992 52256
rect 14928 52196 14932 52252
rect 14932 52196 14988 52252
rect 14988 52196 14992 52252
rect 14928 52192 14992 52196
rect 15008 52252 15072 52256
rect 15008 52196 15012 52252
rect 15012 52196 15068 52252
rect 15068 52196 15072 52252
rect 15008 52192 15072 52196
rect 15088 52252 15152 52256
rect 15088 52196 15092 52252
rect 15092 52196 15148 52252
rect 15148 52196 15152 52252
rect 15088 52192 15152 52196
rect 24112 52252 24176 52256
rect 24112 52196 24116 52252
rect 24116 52196 24172 52252
rect 24172 52196 24176 52252
rect 24112 52192 24176 52196
rect 24192 52252 24256 52256
rect 24192 52196 24196 52252
rect 24196 52196 24252 52252
rect 24252 52196 24256 52252
rect 24192 52192 24256 52196
rect 24272 52252 24336 52256
rect 24272 52196 24276 52252
rect 24276 52196 24332 52252
rect 24332 52196 24336 52252
rect 24272 52192 24336 52196
rect 24352 52252 24416 52256
rect 24352 52196 24356 52252
rect 24356 52196 24412 52252
rect 24412 52196 24416 52252
rect 24352 52192 24416 52196
rect 10216 51708 10280 51712
rect 10216 51652 10220 51708
rect 10220 51652 10276 51708
rect 10276 51652 10280 51708
rect 10216 51648 10280 51652
rect 10296 51708 10360 51712
rect 10296 51652 10300 51708
rect 10300 51652 10356 51708
rect 10356 51652 10360 51708
rect 10296 51648 10360 51652
rect 10376 51708 10440 51712
rect 10376 51652 10380 51708
rect 10380 51652 10436 51708
rect 10436 51652 10440 51708
rect 10376 51648 10440 51652
rect 10456 51708 10520 51712
rect 10456 51652 10460 51708
rect 10460 51652 10516 51708
rect 10516 51652 10520 51708
rect 10456 51648 10520 51652
rect 19480 51708 19544 51712
rect 19480 51652 19484 51708
rect 19484 51652 19540 51708
rect 19540 51652 19544 51708
rect 19480 51648 19544 51652
rect 19560 51708 19624 51712
rect 19560 51652 19564 51708
rect 19564 51652 19620 51708
rect 19620 51652 19624 51708
rect 19560 51648 19624 51652
rect 19640 51708 19704 51712
rect 19640 51652 19644 51708
rect 19644 51652 19700 51708
rect 19700 51652 19704 51708
rect 19640 51648 19704 51652
rect 19720 51708 19784 51712
rect 19720 51652 19724 51708
rect 19724 51652 19780 51708
rect 19780 51652 19784 51708
rect 19720 51648 19784 51652
rect 5584 51164 5648 51168
rect 5584 51108 5588 51164
rect 5588 51108 5644 51164
rect 5644 51108 5648 51164
rect 5584 51104 5648 51108
rect 5664 51164 5728 51168
rect 5664 51108 5668 51164
rect 5668 51108 5724 51164
rect 5724 51108 5728 51164
rect 5664 51104 5728 51108
rect 5744 51164 5808 51168
rect 5744 51108 5748 51164
rect 5748 51108 5804 51164
rect 5804 51108 5808 51164
rect 5744 51104 5808 51108
rect 5824 51164 5888 51168
rect 5824 51108 5828 51164
rect 5828 51108 5884 51164
rect 5884 51108 5888 51164
rect 5824 51104 5888 51108
rect 14848 51164 14912 51168
rect 14848 51108 14852 51164
rect 14852 51108 14908 51164
rect 14908 51108 14912 51164
rect 14848 51104 14912 51108
rect 14928 51164 14992 51168
rect 14928 51108 14932 51164
rect 14932 51108 14988 51164
rect 14988 51108 14992 51164
rect 14928 51104 14992 51108
rect 15008 51164 15072 51168
rect 15008 51108 15012 51164
rect 15012 51108 15068 51164
rect 15068 51108 15072 51164
rect 15008 51104 15072 51108
rect 15088 51164 15152 51168
rect 15088 51108 15092 51164
rect 15092 51108 15148 51164
rect 15148 51108 15152 51164
rect 15088 51104 15152 51108
rect 24112 51164 24176 51168
rect 24112 51108 24116 51164
rect 24116 51108 24172 51164
rect 24172 51108 24176 51164
rect 24112 51104 24176 51108
rect 24192 51164 24256 51168
rect 24192 51108 24196 51164
rect 24196 51108 24252 51164
rect 24252 51108 24256 51164
rect 24192 51104 24256 51108
rect 24272 51164 24336 51168
rect 24272 51108 24276 51164
rect 24276 51108 24332 51164
rect 24332 51108 24336 51164
rect 24272 51104 24336 51108
rect 24352 51164 24416 51168
rect 24352 51108 24356 51164
rect 24356 51108 24412 51164
rect 24412 51108 24416 51164
rect 24352 51104 24416 51108
rect 10216 50620 10280 50624
rect 10216 50564 10220 50620
rect 10220 50564 10276 50620
rect 10276 50564 10280 50620
rect 10216 50560 10280 50564
rect 10296 50620 10360 50624
rect 10296 50564 10300 50620
rect 10300 50564 10356 50620
rect 10356 50564 10360 50620
rect 10296 50560 10360 50564
rect 10376 50620 10440 50624
rect 10376 50564 10380 50620
rect 10380 50564 10436 50620
rect 10436 50564 10440 50620
rect 10376 50560 10440 50564
rect 10456 50620 10520 50624
rect 10456 50564 10460 50620
rect 10460 50564 10516 50620
rect 10516 50564 10520 50620
rect 10456 50560 10520 50564
rect 19480 50620 19544 50624
rect 19480 50564 19484 50620
rect 19484 50564 19540 50620
rect 19540 50564 19544 50620
rect 19480 50560 19544 50564
rect 19560 50620 19624 50624
rect 19560 50564 19564 50620
rect 19564 50564 19620 50620
rect 19620 50564 19624 50620
rect 19560 50560 19624 50564
rect 19640 50620 19704 50624
rect 19640 50564 19644 50620
rect 19644 50564 19700 50620
rect 19700 50564 19704 50620
rect 19640 50560 19704 50564
rect 19720 50620 19784 50624
rect 19720 50564 19724 50620
rect 19724 50564 19780 50620
rect 19780 50564 19784 50620
rect 19720 50560 19784 50564
rect 5584 50076 5648 50080
rect 5584 50020 5588 50076
rect 5588 50020 5644 50076
rect 5644 50020 5648 50076
rect 5584 50016 5648 50020
rect 5664 50076 5728 50080
rect 5664 50020 5668 50076
rect 5668 50020 5724 50076
rect 5724 50020 5728 50076
rect 5664 50016 5728 50020
rect 5744 50076 5808 50080
rect 5744 50020 5748 50076
rect 5748 50020 5804 50076
rect 5804 50020 5808 50076
rect 5744 50016 5808 50020
rect 5824 50076 5888 50080
rect 5824 50020 5828 50076
rect 5828 50020 5884 50076
rect 5884 50020 5888 50076
rect 5824 50016 5888 50020
rect 14848 50076 14912 50080
rect 14848 50020 14852 50076
rect 14852 50020 14908 50076
rect 14908 50020 14912 50076
rect 14848 50016 14912 50020
rect 14928 50076 14992 50080
rect 14928 50020 14932 50076
rect 14932 50020 14988 50076
rect 14988 50020 14992 50076
rect 14928 50016 14992 50020
rect 15008 50076 15072 50080
rect 15008 50020 15012 50076
rect 15012 50020 15068 50076
rect 15068 50020 15072 50076
rect 15008 50016 15072 50020
rect 15088 50076 15152 50080
rect 15088 50020 15092 50076
rect 15092 50020 15148 50076
rect 15148 50020 15152 50076
rect 15088 50016 15152 50020
rect 24112 50076 24176 50080
rect 24112 50020 24116 50076
rect 24116 50020 24172 50076
rect 24172 50020 24176 50076
rect 24112 50016 24176 50020
rect 24192 50076 24256 50080
rect 24192 50020 24196 50076
rect 24196 50020 24252 50076
rect 24252 50020 24256 50076
rect 24192 50016 24256 50020
rect 24272 50076 24336 50080
rect 24272 50020 24276 50076
rect 24276 50020 24332 50076
rect 24332 50020 24336 50076
rect 24272 50016 24336 50020
rect 24352 50076 24416 50080
rect 24352 50020 24356 50076
rect 24356 50020 24412 50076
rect 24412 50020 24416 50076
rect 24352 50016 24416 50020
rect 10216 49532 10280 49536
rect 10216 49476 10220 49532
rect 10220 49476 10276 49532
rect 10276 49476 10280 49532
rect 10216 49472 10280 49476
rect 10296 49532 10360 49536
rect 10296 49476 10300 49532
rect 10300 49476 10356 49532
rect 10356 49476 10360 49532
rect 10296 49472 10360 49476
rect 10376 49532 10440 49536
rect 10376 49476 10380 49532
rect 10380 49476 10436 49532
rect 10436 49476 10440 49532
rect 10376 49472 10440 49476
rect 10456 49532 10520 49536
rect 10456 49476 10460 49532
rect 10460 49476 10516 49532
rect 10516 49476 10520 49532
rect 10456 49472 10520 49476
rect 19480 49532 19544 49536
rect 19480 49476 19484 49532
rect 19484 49476 19540 49532
rect 19540 49476 19544 49532
rect 19480 49472 19544 49476
rect 19560 49532 19624 49536
rect 19560 49476 19564 49532
rect 19564 49476 19620 49532
rect 19620 49476 19624 49532
rect 19560 49472 19624 49476
rect 19640 49532 19704 49536
rect 19640 49476 19644 49532
rect 19644 49476 19700 49532
rect 19700 49476 19704 49532
rect 19640 49472 19704 49476
rect 19720 49532 19784 49536
rect 19720 49476 19724 49532
rect 19724 49476 19780 49532
rect 19780 49476 19784 49532
rect 19720 49472 19784 49476
rect 5584 48988 5648 48992
rect 5584 48932 5588 48988
rect 5588 48932 5644 48988
rect 5644 48932 5648 48988
rect 5584 48928 5648 48932
rect 5664 48988 5728 48992
rect 5664 48932 5668 48988
rect 5668 48932 5724 48988
rect 5724 48932 5728 48988
rect 5664 48928 5728 48932
rect 5744 48988 5808 48992
rect 5744 48932 5748 48988
rect 5748 48932 5804 48988
rect 5804 48932 5808 48988
rect 5744 48928 5808 48932
rect 5824 48988 5888 48992
rect 5824 48932 5828 48988
rect 5828 48932 5884 48988
rect 5884 48932 5888 48988
rect 5824 48928 5888 48932
rect 14848 48988 14912 48992
rect 14848 48932 14852 48988
rect 14852 48932 14908 48988
rect 14908 48932 14912 48988
rect 14848 48928 14912 48932
rect 14928 48988 14992 48992
rect 14928 48932 14932 48988
rect 14932 48932 14988 48988
rect 14988 48932 14992 48988
rect 14928 48928 14992 48932
rect 15008 48988 15072 48992
rect 15008 48932 15012 48988
rect 15012 48932 15068 48988
rect 15068 48932 15072 48988
rect 15008 48928 15072 48932
rect 15088 48988 15152 48992
rect 15088 48932 15092 48988
rect 15092 48932 15148 48988
rect 15148 48932 15152 48988
rect 15088 48928 15152 48932
rect 24112 48988 24176 48992
rect 24112 48932 24116 48988
rect 24116 48932 24172 48988
rect 24172 48932 24176 48988
rect 24112 48928 24176 48932
rect 24192 48988 24256 48992
rect 24192 48932 24196 48988
rect 24196 48932 24252 48988
rect 24252 48932 24256 48988
rect 24192 48928 24256 48932
rect 24272 48988 24336 48992
rect 24272 48932 24276 48988
rect 24276 48932 24332 48988
rect 24332 48932 24336 48988
rect 24272 48928 24336 48932
rect 24352 48988 24416 48992
rect 24352 48932 24356 48988
rect 24356 48932 24412 48988
rect 24412 48932 24416 48988
rect 24352 48928 24416 48932
rect 10216 48444 10280 48448
rect 10216 48388 10220 48444
rect 10220 48388 10276 48444
rect 10276 48388 10280 48444
rect 10216 48384 10280 48388
rect 10296 48444 10360 48448
rect 10296 48388 10300 48444
rect 10300 48388 10356 48444
rect 10356 48388 10360 48444
rect 10296 48384 10360 48388
rect 10376 48444 10440 48448
rect 10376 48388 10380 48444
rect 10380 48388 10436 48444
rect 10436 48388 10440 48444
rect 10376 48384 10440 48388
rect 10456 48444 10520 48448
rect 10456 48388 10460 48444
rect 10460 48388 10516 48444
rect 10516 48388 10520 48444
rect 10456 48384 10520 48388
rect 19480 48444 19544 48448
rect 19480 48388 19484 48444
rect 19484 48388 19540 48444
rect 19540 48388 19544 48444
rect 19480 48384 19544 48388
rect 19560 48444 19624 48448
rect 19560 48388 19564 48444
rect 19564 48388 19620 48444
rect 19620 48388 19624 48444
rect 19560 48384 19624 48388
rect 19640 48444 19704 48448
rect 19640 48388 19644 48444
rect 19644 48388 19700 48444
rect 19700 48388 19704 48444
rect 19640 48384 19704 48388
rect 19720 48444 19784 48448
rect 19720 48388 19724 48444
rect 19724 48388 19780 48444
rect 19780 48388 19784 48444
rect 19720 48384 19784 48388
rect 5584 47900 5648 47904
rect 5584 47844 5588 47900
rect 5588 47844 5644 47900
rect 5644 47844 5648 47900
rect 5584 47840 5648 47844
rect 5664 47900 5728 47904
rect 5664 47844 5668 47900
rect 5668 47844 5724 47900
rect 5724 47844 5728 47900
rect 5664 47840 5728 47844
rect 5744 47900 5808 47904
rect 5744 47844 5748 47900
rect 5748 47844 5804 47900
rect 5804 47844 5808 47900
rect 5744 47840 5808 47844
rect 5824 47900 5888 47904
rect 5824 47844 5828 47900
rect 5828 47844 5884 47900
rect 5884 47844 5888 47900
rect 5824 47840 5888 47844
rect 14848 47900 14912 47904
rect 14848 47844 14852 47900
rect 14852 47844 14908 47900
rect 14908 47844 14912 47900
rect 14848 47840 14912 47844
rect 14928 47900 14992 47904
rect 14928 47844 14932 47900
rect 14932 47844 14988 47900
rect 14988 47844 14992 47900
rect 14928 47840 14992 47844
rect 15008 47900 15072 47904
rect 15008 47844 15012 47900
rect 15012 47844 15068 47900
rect 15068 47844 15072 47900
rect 15008 47840 15072 47844
rect 15088 47900 15152 47904
rect 15088 47844 15092 47900
rect 15092 47844 15148 47900
rect 15148 47844 15152 47900
rect 15088 47840 15152 47844
rect 24112 47900 24176 47904
rect 24112 47844 24116 47900
rect 24116 47844 24172 47900
rect 24172 47844 24176 47900
rect 24112 47840 24176 47844
rect 24192 47900 24256 47904
rect 24192 47844 24196 47900
rect 24196 47844 24252 47900
rect 24252 47844 24256 47900
rect 24192 47840 24256 47844
rect 24272 47900 24336 47904
rect 24272 47844 24276 47900
rect 24276 47844 24332 47900
rect 24332 47844 24336 47900
rect 24272 47840 24336 47844
rect 24352 47900 24416 47904
rect 24352 47844 24356 47900
rect 24356 47844 24412 47900
rect 24412 47844 24416 47900
rect 24352 47840 24416 47844
rect 10216 47356 10280 47360
rect 10216 47300 10220 47356
rect 10220 47300 10276 47356
rect 10276 47300 10280 47356
rect 10216 47296 10280 47300
rect 10296 47356 10360 47360
rect 10296 47300 10300 47356
rect 10300 47300 10356 47356
rect 10356 47300 10360 47356
rect 10296 47296 10360 47300
rect 10376 47356 10440 47360
rect 10376 47300 10380 47356
rect 10380 47300 10436 47356
rect 10436 47300 10440 47356
rect 10376 47296 10440 47300
rect 10456 47356 10520 47360
rect 10456 47300 10460 47356
rect 10460 47300 10516 47356
rect 10516 47300 10520 47356
rect 10456 47296 10520 47300
rect 19480 47356 19544 47360
rect 19480 47300 19484 47356
rect 19484 47300 19540 47356
rect 19540 47300 19544 47356
rect 19480 47296 19544 47300
rect 19560 47356 19624 47360
rect 19560 47300 19564 47356
rect 19564 47300 19620 47356
rect 19620 47300 19624 47356
rect 19560 47296 19624 47300
rect 19640 47356 19704 47360
rect 19640 47300 19644 47356
rect 19644 47300 19700 47356
rect 19700 47300 19704 47356
rect 19640 47296 19704 47300
rect 19720 47356 19784 47360
rect 19720 47300 19724 47356
rect 19724 47300 19780 47356
rect 19780 47300 19784 47356
rect 19720 47296 19784 47300
rect 5584 46812 5648 46816
rect 5584 46756 5588 46812
rect 5588 46756 5644 46812
rect 5644 46756 5648 46812
rect 5584 46752 5648 46756
rect 5664 46812 5728 46816
rect 5664 46756 5668 46812
rect 5668 46756 5724 46812
rect 5724 46756 5728 46812
rect 5664 46752 5728 46756
rect 5744 46812 5808 46816
rect 5744 46756 5748 46812
rect 5748 46756 5804 46812
rect 5804 46756 5808 46812
rect 5744 46752 5808 46756
rect 5824 46812 5888 46816
rect 5824 46756 5828 46812
rect 5828 46756 5884 46812
rect 5884 46756 5888 46812
rect 5824 46752 5888 46756
rect 14848 46812 14912 46816
rect 14848 46756 14852 46812
rect 14852 46756 14908 46812
rect 14908 46756 14912 46812
rect 14848 46752 14912 46756
rect 14928 46812 14992 46816
rect 14928 46756 14932 46812
rect 14932 46756 14988 46812
rect 14988 46756 14992 46812
rect 14928 46752 14992 46756
rect 15008 46812 15072 46816
rect 15008 46756 15012 46812
rect 15012 46756 15068 46812
rect 15068 46756 15072 46812
rect 15008 46752 15072 46756
rect 15088 46812 15152 46816
rect 15088 46756 15092 46812
rect 15092 46756 15148 46812
rect 15148 46756 15152 46812
rect 15088 46752 15152 46756
rect 24112 46812 24176 46816
rect 24112 46756 24116 46812
rect 24116 46756 24172 46812
rect 24172 46756 24176 46812
rect 24112 46752 24176 46756
rect 24192 46812 24256 46816
rect 24192 46756 24196 46812
rect 24196 46756 24252 46812
rect 24252 46756 24256 46812
rect 24192 46752 24256 46756
rect 24272 46812 24336 46816
rect 24272 46756 24276 46812
rect 24276 46756 24332 46812
rect 24332 46756 24336 46812
rect 24272 46752 24336 46756
rect 24352 46812 24416 46816
rect 24352 46756 24356 46812
rect 24356 46756 24412 46812
rect 24412 46756 24416 46812
rect 24352 46752 24416 46756
rect 10216 46268 10280 46272
rect 10216 46212 10220 46268
rect 10220 46212 10276 46268
rect 10276 46212 10280 46268
rect 10216 46208 10280 46212
rect 10296 46268 10360 46272
rect 10296 46212 10300 46268
rect 10300 46212 10356 46268
rect 10356 46212 10360 46268
rect 10296 46208 10360 46212
rect 10376 46268 10440 46272
rect 10376 46212 10380 46268
rect 10380 46212 10436 46268
rect 10436 46212 10440 46268
rect 10376 46208 10440 46212
rect 10456 46268 10520 46272
rect 10456 46212 10460 46268
rect 10460 46212 10516 46268
rect 10516 46212 10520 46268
rect 10456 46208 10520 46212
rect 19480 46268 19544 46272
rect 19480 46212 19484 46268
rect 19484 46212 19540 46268
rect 19540 46212 19544 46268
rect 19480 46208 19544 46212
rect 19560 46268 19624 46272
rect 19560 46212 19564 46268
rect 19564 46212 19620 46268
rect 19620 46212 19624 46268
rect 19560 46208 19624 46212
rect 19640 46268 19704 46272
rect 19640 46212 19644 46268
rect 19644 46212 19700 46268
rect 19700 46212 19704 46268
rect 19640 46208 19704 46212
rect 19720 46268 19784 46272
rect 19720 46212 19724 46268
rect 19724 46212 19780 46268
rect 19780 46212 19784 46268
rect 19720 46208 19784 46212
rect 5584 45724 5648 45728
rect 5584 45668 5588 45724
rect 5588 45668 5644 45724
rect 5644 45668 5648 45724
rect 5584 45664 5648 45668
rect 5664 45724 5728 45728
rect 5664 45668 5668 45724
rect 5668 45668 5724 45724
rect 5724 45668 5728 45724
rect 5664 45664 5728 45668
rect 5744 45724 5808 45728
rect 5744 45668 5748 45724
rect 5748 45668 5804 45724
rect 5804 45668 5808 45724
rect 5744 45664 5808 45668
rect 5824 45724 5888 45728
rect 5824 45668 5828 45724
rect 5828 45668 5884 45724
rect 5884 45668 5888 45724
rect 5824 45664 5888 45668
rect 14848 45724 14912 45728
rect 14848 45668 14852 45724
rect 14852 45668 14908 45724
rect 14908 45668 14912 45724
rect 14848 45664 14912 45668
rect 14928 45724 14992 45728
rect 14928 45668 14932 45724
rect 14932 45668 14988 45724
rect 14988 45668 14992 45724
rect 14928 45664 14992 45668
rect 15008 45724 15072 45728
rect 15008 45668 15012 45724
rect 15012 45668 15068 45724
rect 15068 45668 15072 45724
rect 15008 45664 15072 45668
rect 15088 45724 15152 45728
rect 15088 45668 15092 45724
rect 15092 45668 15148 45724
rect 15148 45668 15152 45724
rect 15088 45664 15152 45668
rect 24112 45724 24176 45728
rect 24112 45668 24116 45724
rect 24116 45668 24172 45724
rect 24172 45668 24176 45724
rect 24112 45664 24176 45668
rect 24192 45724 24256 45728
rect 24192 45668 24196 45724
rect 24196 45668 24252 45724
rect 24252 45668 24256 45724
rect 24192 45664 24256 45668
rect 24272 45724 24336 45728
rect 24272 45668 24276 45724
rect 24276 45668 24332 45724
rect 24332 45668 24336 45724
rect 24272 45664 24336 45668
rect 24352 45724 24416 45728
rect 24352 45668 24356 45724
rect 24356 45668 24412 45724
rect 24412 45668 24416 45724
rect 24352 45664 24416 45668
rect 10216 45180 10280 45184
rect 10216 45124 10220 45180
rect 10220 45124 10276 45180
rect 10276 45124 10280 45180
rect 10216 45120 10280 45124
rect 10296 45180 10360 45184
rect 10296 45124 10300 45180
rect 10300 45124 10356 45180
rect 10356 45124 10360 45180
rect 10296 45120 10360 45124
rect 10376 45180 10440 45184
rect 10376 45124 10380 45180
rect 10380 45124 10436 45180
rect 10436 45124 10440 45180
rect 10376 45120 10440 45124
rect 10456 45180 10520 45184
rect 10456 45124 10460 45180
rect 10460 45124 10516 45180
rect 10516 45124 10520 45180
rect 10456 45120 10520 45124
rect 19480 45180 19544 45184
rect 19480 45124 19484 45180
rect 19484 45124 19540 45180
rect 19540 45124 19544 45180
rect 19480 45120 19544 45124
rect 19560 45180 19624 45184
rect 19560 45124 19564 45180
rect 19564 45124 19620 45180
rect 19620 45124 19624 45180
rect 19560 45120 19624 45124
rect 19640 45180 19704 45184
rect 19640 45124 19644 45180
rect 19644 45124 19700 45180
rect 19700 45124 19704 45180
rect 19640 45120 19704 45124
rect 19720 45180 19784 45184
rect 19720 45124 19724 45180
rect 19724 45124 19780 45180
rect 19780 45124 19784 45180
rect 19720 45120 19784 45124
rect 5584 44636 5648 44640
rect 5584 44580 5588 44636
rect 5588 44580 5644 44636
rect 5644 44580 5648 44636
rect 5584 44576 5648 44580
rect 5664 44636 5728 44640
rect 5664 44580 5668 44636
rect 5668 44580 5724 44636
rect 5724 44580 5728 44636
rect 5664 44576 5728 44580
rect 5744 44636 5808 44640
rect 5744 44580 5748 44636
rect 5748 44580 5804 44636
rect 5804 44580 5808 44636
rect 5744 44576 5808 44580
rect 5824 44636 5888 44640
rect 5824 44580 5828 44636
rect 5828 44580 5884 44636
rect 5884 44580 5888 44636
rect 5824 44576 5888 44580
rect 14848 44636 14912 44640
rect 14848 44580 14852 44636
rect 14852 44580 14908 44636
rect 14908 44580 14912 44636
rect 14848 44576 14912 44580
rect 14928 44636 14992 44640
rect 14928 44580 14932 44636
rect 14932 44580 14988 44636
rect 14988 44580 14992 44636
rect 14928 44576 14992 44580
rect 15008 44636 15072 44640
rect 15008 44580 15012 44636
rect 15012 44580 15068 44636
rect 15068 44580 15072 44636
rect 15008 44576 15072 44580
rect 15088 44636 15152 44640
rect 15088 44580 15092 44636
rect 15092 44580 15148 44636
rect 15148 44580 15152 44636
rect 15088 44576 15152 44580
rect 24112 44636 24176 44640
rect 24112 44580 24116 44636
rect 24116 44580 24172 44636
rect 24172 44580 24176 44636
rect 24112 44576 24176 44580
rect 24192 44636 24256 44640
rect 24192 44580 24196 44636
rect 24196 44580 24252 44636
rect 24252 44580 24256 44636
rect 24192 44576 24256 44580
rect 24272 44636 24336 44640
rect 24272 44580 24276 44636
rect 24276 44580 24332 44636
rect 24332 44580 24336 44636
rect 24272 44576 24336 44580
rect 24352 44636 24416 44640
rect 24352 44580 24356 44636
rect 24356 44580 24412 44636
rect 24412 44580 24416 44636
rect 24352 44576 24416 44580
rect 10216 44092 10280 44096
rect 10216 44036 10220 44092
rect 10220 44036 10276 44092
rect 10276 44036 10280 44092
rect 10216 44032 10280 44036
rect 10296 44092 10360 44096
rect 10296 44036 10300 44092
rect 10300 44036 10356 44092
rect 10356 44036 10360 44092
rect 10296 44032 10360 44036
rect 10376 44092 10440 44096
rect 10376 44036 10380 44092
rect 10380 44036 10436 44092
rect 10436 44036 10440 44092
rect 10376 44032 10440 44036
rect 10456 44092 10520 44096
rect 10456 44036 10460 44092
rect 10460 44036 10516 44092
rect 10516 44036 10520 44092
rect 10456 44032 10520 44036
rect 19480 44092 19544 44096
rect 19480 44036 19484 44092
rect 19484 44036 19540 44092
rect 19540 44036 19544 44092
rect 19480 44032 19544 44036
rect 19560 44092 19624 44096
rect 19560 44036 19564 44092
rect 19564 44036 19620 44092
rect 19620 44036 19624 44092
rect 19560 44032 19624 44036
rect 19640 44092 19704 44096
rect 19640 44036 19644 44092
rect 19644 44036 19700 44092
rect 19700 44036 19704 44092
rect 19640 44032 19704 44036
rect 19720 44092 19784 44096
rect 19720 44036 19724 44092
rect 19724 44036 19780 44092
rect 19780 44036 19784 44092
rect 19720 44032 19784 44036
rect 5584 43548 5648 43552
rect 5584 43492 5588 43548
rect 5588 43492 5644 43548
rect 5644 43492 5648 43548
rect 5584 43488 5648 43492
rect 5664 43548 5728 43552
rect 5664 43492 5668 43548
rect 5668 43492 5724 43548
rect 5724 43492 5728 43548
rect 5664 43488 5728 43492
rect 5744 43548 5808 43552
rect 5744 43492 5748 43548
rect 5748 43492 5804 43548
rect 5804 43492 5808 43548
rect 5744 43488 5808 43492
rect 5824 43548 5888 43552
rect 5824 43492 5828 43548
rect 5828 43492 5884 43548
rect 5884 43492 5888 43548
rect 5824 43488 5888 43492
rect 14848 43548 14912 43552
rect 14848 43492 14852 43548
rect 14852 43492 14908 43548
rect 14908 43492 14912 43548
rect 14848 43488 14912 43492
rect 14928 43548 14992 43552
rect 14928 43492 14932 43548
rect 14932 43492 14988 43548
rect 14988 43492 14992 43548
rect 14928 43488 14992 43492
rect 15008 43548 15072 43552
rect 15008 43492 15012 43548
rect 15012 43492 15068 43548
rect 15068 43492 15072 43548
rect 15008 43488 15072 43492
rect 15088 43548 15152 43552
rect 15088 43492 15092 43548
rect 15092 43492 15148 43548
rect 15148 43492 15152 43548
rect 15088 43488 15152 43492
rect 24112 43548 24176 43552
rect 24112 43492 24116 43548
rect 24116 43492 24172 43548
rect 24172 43492 24176 43548
rect 24112 43488 24176 43492
rect 24192 43548 24256 43552
rect 24192 43492 24196 43548
rect 24196 43492 24252 43548
rect 24252 43492 24256 43548
rect 24192 43488 24256 43492
rect 24272 43548 24336 43552
rect 24272 43492 24276 43548
rect 24276 43492 24332 43548
rect 24332 43492 24336 43548
rect 24272 43488 24336 43492
rect 24352 43548 24416 43552
rect 24352 43492 24356 43548
rect 24356 43492 24412 43548
rect 24412 43492 24416 43548
rect 24352 43488 24416 43492
rect 10216 43004 10280 43008
rect 10216 42948 10220 43004
rect 10220 42948 10276 43004
rect 10276 42948 10280 43004
rect 10216 42944 10280 42948
rect 10296 43004 10360 43008
rect 10296 42948 10300 43004
rect 10300 42948 10356 43004
rect 10356 42948 10360 43004
rect 10296 42944 10360 42948
rect 10376 43004 10440 43008
rect 10376 42948 10380 43004
rect 10380 42948 10436 43004
rect 10436 42948 10440 43004
rect 10376 42944 10440 42948
rect 10456 43004 10520 43008
rect 10456 42948 10460 43004
rect 10460 42948 10516 43004
rect 10516 42948 10520 43004
rect 10456 42944 10520 42948
rect 19480 43004 19544 43008
rect 19480 42948 19484 43004
rect 19484 42948 19540 43004
rect 19540 42948 19544 43004
rect 19480 42944 19544 42948
rect 19560 43004 19624 43008
rect 19560 42948 19564 43004
rect 19564 42948 19620 43004
rect 19620 42948 19624 43004
rect 19560 42944 19624 42948
rect 19640 43004 19704 43008
rect 19640 42948 19644 43004
rect 19644 42948 19700 43004
rect 19700 42948 19704 43004
rect 19640 42944 19704 42948
rect 19720 43004 19784 43008
rect 19720 42948 19724 43004
rect 19724 42948 19780 43004
rect 19780 42948 19784 43004
rect 19720 42944 19784 42948
rect 5584 42460 5648 42464
rect 5584 42404 5588 42460
rect 5588 42404 5644 42460
rect 5644 42404 5648 42460
rect 5584 42400 5648 42404
rect 5664 42460 5728 42464
rect 5664 42404 5668 42460
rect 5668 42404 5724 42460
rect 5724 42404 5728 42460
rect 5664 42400 5728 42404
rect 5744 42460 5808 42464
rect 5744 42404 5748 42460
rect 5748 42404 5804 42460
rect 5804 42404 5808 42460
rect 5744 42400 5808 42404
rect 5824 42460 5888 42464
rect 5824 42404 5828 42460
rect 5828 42404 5884 42460
rect 5884 42404 5888 42460
rect 5824 42400 5888 42404
rect 14848 42460 14912 42464
rect 14848 42404 14852 42460
rect 14852 42404 14908 42460
rect 14908 42404 14912 42460
rect 14848 42400 14912 42404
rect 14928 42460 14992 42464
rect 14928 42404 14932 42460
rect 14932 42404 14988 42460
rect 14988 42404 14992 42460
rect 14928 42400 14992 42404
rect 15008 42460 15072 42464
rect 15008 42404 15012 42460
rect 15012 42404 15068 42460
rect 15068 42404 15072 42460
rect 15008 42400 15072 42404
rect 15088 42460 15152 42464
rect 15088 42404 15092 42460
rect 15092 42404 15148 42460
rect 15148 42404 15152 42460
rect 15088 42400 15152 42404
rect 24112 42460 24176 42464
rect 24112 42404 24116 42460
rect 24116 42404 24172 42460
rect 24172 42404 24176 42460
rect 24112 42400 24176 42404
rect 24192 42460 24256 42464
rect 24192 42404 24196 42460
rect 24196 42404 24252 42460
rect 24252 42404 24256 42460
rect 24192 42400 24256 42404
rect 24272 42460 24336 42464
rect 24272 42404 24276 42460
rect 24276 42404 24332 42460
rect 24332 42404 24336 42460
rect 24272 42400 24336 42404
rect 24352 42460 24416 42464
rect 24352 42404 24356 42460
rect 24356 42404 24412 42460
rect 24412 42404 24416 42460
rect 24352 42400 24416 42404
rect 10216 41916 10280 41920
rect 10216 41860 10220 41916
rect 10220 41860 10276 41916
rect 10276 41860 10280 41916
rect 10216 41856 10280 41860
rect 10296 41916 10360 41920
rect 10296 41860 10300 41916
rect 10300 41860 10356 41916
rect 10356 41860 10360 41916
rect 10296 41856 10360 41860
rect 10376 41916 10440 41920
rect 10376 41860 10380 41916
rect 10380 41860 10436 41916
rect 10436 41860 10440 41916
rect 10376 41856 10440 41860
rect 10456 41916 10520 41920
rect 10456 41860 10460 41916
rect 10460 41860 10516 41916
rect 10516 41860 10520 41916
rect 10456 41856 10520 41860
rect 19480 41916 19544 41920
rect 19480 41860 19484 41916
rect 19484 41860 19540 41916
rect 19540 41860 19544 41916
rect 19480 41856 19544 41860
rect 19560 41916 19624 41920
rect 19560 41860 19564 41916
rect 19564 41860 19620 41916
rect 19620 41860 19624 41916
rect 19560 41856 19624 41860
rect 19640 41916 19704 41920
rect 19640 41860 19644 41916
rect 19644 41860 19700 41916
rect 19700 41860 19704 41916
rect 19640 41856 19704 41860
rect 19720 41916 19784 41920
rect 19720 41860 19724 41916
rect 19724 41860 19780 41916
rect 19780 41860 19784 41916
rect 19720 41856 19784 41860
rect 5584 41372 5648 41376
rect 5584 41316 5588 41372
rect 5588 41316 5644 41372
rect 5644 41316 5648 41372
rect 5584 41312 5648 41316
rect 5664 41372 5728 41376
rect 5664 41316 5668 41372
rect 5668 41316 5724 41372
rect 5724 41316 5728 41372
rect 5664 41312 5728 41316
rect 5744 41372 5808 41376
rect 5744 41316 5748 41372
rect 5748 41316 5804 41372
rect 5804 41316 5808 41372
rect 5744 41312 5808 41316
rect 5824 41372 5888 41376
rect 5824 41316 5828 41372
rect 5828 41316 5884 41372
rect 5884 41316 5888 41372
rect 5824 41312 5888 41316
rect 14848 41372 14912 41376
rect 14848 41316 14852 41372
rect 14852 41316 14908 41372
rect 14908 41316 14912 41372
rect 14848 41312 14912 41316
rect 14928 41372 14992 41376
rect 14928 41316 14932 41372
rect 14932 41316 14988 41372
rect 14988 41316 14992 41372
rect 14928 41312 14992 41316
rect 15008 41372 15072 41376
rect 15008 41316 15012 41372
rect 15012 41316 15068 41372
rect 15068 41316 15072 41372
rect 15008 41312 15072 41316
rect 15088 41372 15152 41376
rect 15088 41316 15092 41372
rect 15092 41316 15148 41372
rect 15148 41316 15152 41372
rect 15088 41312 15152 41316
rect 24112 41372 24176 41376
rect 24112 41316 24116 41372
rect 24116 41316 24172 41372
rect 24172 41316 24176 41372
rect 24112 41312 24176 41316
rect 24192 41372 24256 41376
rect 24192 41316 24196 41372
rect 24196 41316 24252 41372
rect 24252 41316 24256 41372
rect 24192 41312 24256 41316
rect 24272 41372 24336 41376
rect 24272 41316 24276 41372
rect 24276 41316 24332 41372
rect 24332 41316 24336 41372
rect 24272 41312 24336 41316
rect 24352 41372 24416 41376
rect 24352 41316 24356 41372
rect 24356 41316 24412 41372
rect 24412 41316 24416 41372
rect 24352 41312 24416 41316
rect 10216 40828 10280 40832
rect 10216 40772 10220 40828
rect 10220 40772 10276 40828
rect 10276 40772 10280 40828
rect 10216 40768 10280 40772
rect 10296 40828 10360 40832
rect 10296 40772 10300 40828
rect 10300 40772 10356 40828
rect 10356 40772 10360 40828
rect 10296 40768 10360 40772
rect 10376 40828 10440 40832
rect 10376 40772 10380 40828
rect 10380 40772 10436 40828
rect 10436 40772 10440 40828
rect 10376 40768 10440 40772
rect 10456 40828 10520 40832
rect 10456 40772 10460 40828
rect 10460 40772 10516 40828
rect 10516 40772 10520 40828
rect 10456 40768 10520 40772
rect 19480 40828 19544 40832
rect 19480 40772 19484 40828
rect 19484 40772 19540 40828
rect 19540 40772 19544 40828
rect 19480 40768 19544 40772
rect 19560 40828 19624 40832
rect 19560 40772 19564 40828
rect 19564 40772 19620 40828
rect 19620 40772 19624 40828
rect 19560 40768 19624 40772
rect 19640 40828 19704 40832
rect 19640 40772 19644 40828
rect 19644 40772 19700 40828
rect 19700 40772 19704 40828
rect 19640 40768 19704 40772
rect 19720 40828 19784 40832
rect 19720 40772 19724 40828
rect 19724 40772 19780 40828
rect 19780 40772 19784 40828
rect 19720 40768 19784 40772
rect 5584 40284 5648 40288
rect 5584 40228 5588 40284
rect 5588 40228 5644 40284
rect 5644 40228 5648 40284
rect 5584 40224 5648 40228
rect 5664 40284 5728 40288
rect 5664 40228 5668 40284
rect 5668 40228 5724 40284
rect 5724 40228 5728 40284
rect 5664 40224 5728 40228
rect 5744 40284 5808 40288
rect 5744 40228 5748 40284
rect 5748 40228 5804 40284
rect 5804 40228 5808 40284
rect 5744 40224 5808 40228
rect 5824 40284 5888 40288
rect 5824 40228 5828 40284
rect 5828 40228 5884 40284
rect 5884 40228 5888 40284
rect 5824 40224 5888 40228
rect 14848 40284 14912 40288
rect 14848 40228 14852 40284
rect 14852 40228 14908 40284
rect 14908 40228 14912 40284
rect 14848 40224 14912 40228
rect 14928 40284 14992 40288
rect 14928 40228 14932 40284
rect 14932 40228 14988 40284
rect 14988 40228 14992 40284
rect 14928 40224 14992 40228
rect 15008 40284 15072 40288
rect 15008 40228 15012 40284
rect 15012 40228 15068 40284
rect 15068 40228 15072 40284
rect 15008 40224 15072 40228
rect 15088 40284 15152 40288
rect 15088 40228 15092 40284
rect 15092 40228 15148 40284
rect 15148 40228 15152 40284
rect 15088 40224 15152 40228
rect 24112 40284 24176 40288
rect 24112 40228 24116 40284
rect 24116 40228 24172 40284
rect 24172 40228 24176 40284
rect 24112 40224 24176 40228
rect 24192 40284 24256 40288
rect 24192 40228 24196 40284
rect 24196 40228 24252 40284
rect 24252 40228 24256 40284
rect 24192 40224 24256 40228
rect 24272 40284 24336 40288
rect 24272 40228 24276 40284
rect 24276 40228 24332 40284
rect 24332 40228 24336 40284
rect 24272 40224 24336 40228
rect 24352 40284 24416 40288
rect 24352 40228 24356 40284
rect 24356 40228 24412 40284
rect 24412 40228 24416 40284
rect 24352 40224 24416 40228
rect 10216 39740 10280 39744
rect 10216 39684 10220 39740
rect 10220 39684 10276 39740
rect 10276 39684 10280 39740
rect 10216 39680 10280 39684
rect 10296 39740 10360 39744
rect 10296 39684 10300 39740
rect 10300 39684 10356 39740
rect 10356 39684 10360 39740
rect 10296 39680 10360 39684
rect 10376 39740 10440 39744
rect 10376 39684 10380 39740
rect 10380 39684 10436 39740
rect 10436 39684 10440 39740
rect 10376 39680 10440 39684
rect 10456 39740 10520 39744
rect 10456 39684 10460 39740
rect 10460 39684 10516 39740
rect 10516 39684 10520 39740
rect 10456 39680 10520 39684
rect 19480 39740 19544 39744
rect 19480 39684 19484 39740
rect 19484 39684 19540 39740
rect 19540 39684 19544 39740
rect 19480 39680 19544 39684
rect 19560 39740 19624 39744
rect 19560 39684 19564 39740
rect 19564 39684 19620 39740
rect 19620 39684 19624 39740
rect 19560 39680 19624 39684
rect 19640 39740 19704 39744
rect 19640 39684 19644 39740
rect 19644 39684 19700 39740
rect 19700 39684 19704 39740
rect 19640 39680 19704 39684
rect 19720 39740 19784 39744
rect 19720 39684 19724 39740
rect 19724 39684 19780 39740
rect 19780 39684 19784 39740
rect 19720 39680 19784 39684
rect 5584 39196 5648 39200
rect 5584 39140 5588 39196
rect 5588 39140 5644 39196
rect 5644 39140 5648 39196
rect 5584 39136 5648 39140
rect 5664 39196 5728 39200
rect 5664 39140 5668 39196
rect 5668 39140 5724 39196
rect 5724 39140 5728 39196
rect 5664 39136 5728 39140
rect 5744 39196 5808 39200
rect 5744 39140 5748 39196
rect 5748 39140 5804 39196
rect 5804 39140 5808 39196
rect 5744 39136 5808 39140
rect 5824 39196 5888 39200
rect 5824 39140 5828 39196
rect 5828 39140 5884 39196
rect 5884 39140 5888 39196
rect 5824 39136 5888 39140
rect 14848 39196 14912 39200
rect 14848 39140 14852 39196
rect 14852 39140 14908 39196
rect 14908 39140 14912 39196
rect 14848 39136 14912 39140
rect 14928 39196 14992 39200
rect 14928 39140 14932 39196
rect 14932 39140 14988 39196
rect 14988 39140 14992 39196
rect 14928 39136 14992 39140
rect 15008 39196 15072 39200
rect 15008 39140 15012 39196
rect 15012 39140 15068 39196
rect 15068 39140 15072 39196
rect 15008 39136 15072 39140
rect 15088 39196 15152 39200
rect 15088 39140 15092 39196
rect 15092 39140 15148 39196
rect 15148 39140 15152 39196
rect 15088 39136 15152 39140
rect 24112 39196 24176 39200
rect 24112 39140 24116 39196
rect 24116 39140 24172 39196
rect 24172 39140 24176 39196
rect 24112 39136 24176 39140
rect 24192 39196 24256 39200
rect 24192 39140 24196 39196
rect 24196 39140 24252 39196
rect 24252 39140 24256 39196
rect 24192 39136 24256 39140
rect 24272 39196 24336 39200
rect 24272 39140 24276 39196
rect 24276 39140 24332 39196
rect 24332 39140 24336 39196
rect 24272 39136 24336 39140
rect 24352 39196 24416 39200
rect 24352 39140 24356 39196
rect 24356 39140 24412 39196
rect 24412 39140 24416 39196
rect 24352 39136 24416 39140
rect 10216 38652 10280 38656
rect 10216 38596 10220 38652
rect 10220 38596 10276 38652
rect 10276 38596 10280 38652
rect 10216 38592 10280 38596
rect 10296 38652 10360 38656
rect 10296 38596 10300 38652
rect 10300 38596 10356 38652
rect 10356 38596 10360 38652
rect 10296 38592 10360 38596
rect 10376 38652 10440 38656
rect 10376 38596 10380 38652
rect 10380 38596 10436 38652
rect 10436 38596 10440 38652
rect 10376 38592 10440 38596
rect 10456 38652 10520 38656
rect 10456 38596 10460 38652
rect 10460 38596 10516 38652
rect 10516 38596 10520 38652
rect 10456 38592 10520 38596
rect 19480 38652 19544 38656
rect 19480 38596 19484 38652
rect 19484 38596 19540 38652
rect 19540 38596 19544 38652
rect 19480 38592 19544 38596
rect 19560 38652 19624 38656
rect 19560 38596 19564 38652
rect 19564 38596 19620 38652
rect 19620 38596 19624 38652
rect 19560 38592 19624 38596
rect 19640 38652 19704 38656
rect 19640 38596 19644 38652
rect 19644 38596 19700 38652
rect 19700 38596 19704 38652
rect 19640 38592 19704 38596
rect 19720 38652 19784 38656
rect 19720 38596 19724 38652
rect 19724 38596 19780 38652
rect 19780 38596 19784 38652
rect 19720 38592 19784 38596
rect 5584 38108 5648 38112
rect 5584 38052 5588 38108
rect 5588 38052 5644 38108
rect 5644 38052 5648 38108
rect 5584 38048 5648 38052
rect 5664 38108 5728 38112
rect 5664 38052 5668 38108
rect 5668 38052 5724 38108
rect 5724 38052 5728 38108
rect 5664 38048 5728 38052
rect 5744 38108 5808 38112
rect 5744 38052 5748 38108
rect 5748 38052 5804 38108
rect 5804 38052 5808 38108
rect 5744 38048 5808 38052
rect 5824 38108 5888 38112
rect 5824 38052 5828 38108
rect 5828 38052 5884 38108
rect 5884 38052 5888 38108
rect 5824 38048 5888 38052
rect 14848 38108 14912 38112
rect 14848 38052 14852 38108
rect 14852 38052 14908 38108
rect 14908 38052 14912 38108
rect 14848 38048 14912 38052
rect 14928 38108 14992 38112
rect 14928 38052 14932 38108
rect 14932 38052 14988 38108
rect 14988 38052 14992 38108
rect 14928 38048 14992 38052
rect 15008 38108 15072 38112
rect 15008 38052 15012 38108
rect 15012 38052 15068 38108
rect 15068 38052 15072 38108
rect 15008 38048 15072 38052
rect 15088 38108 15152 38112
rect 15088 38052 15092 38108
rect 15092 38052 15148 38108
rect 15148 38052 15152 38108
rect 15088 38048 15152 38052
rect 24112 38108 24176 38112
rect 24112 38052 24116 38108
rect 24116 38052 24172 38108
rect 24172 38052 24176 38108
rect 24112 38048 24176 38052
rect 24192 38108 24256 38112
rect 24192 38052 24196 38108
rect 24196 38052 24252 38108
rect 24252 38052 24256 38108
rect 24192 38048 24256 38052
rect 24272 38108 24336 38112
rect 24272 38052 24276 38108
rect 24276 38052 24332 38108
rect 24332 38052 24336 38108
rect 24272 38048 24336 38052
rect 24352 38108 24416 38112
rect 24352 38052 24356 38108
rect 24356 38052 24412 38108
rect 24412 38052 24416 38108
rect 24352 38048 24416 38052
rect 10216 37564 10280 37568
rect 10216 37508 10220 37564
rect 10220 37508 10276 37564
rect 10276 37508 10280 37564
rect 10216 37504 10280 37508
rect 10296 37564 10360 37568
rect 10296 37508 10300 37564
rect 10300 37508 10356 37564
rect 10356 37508 10360 37564
rect 10296 37504 10360 37508
rect 10376 37564 10440 37568
rect 10376 37508 10380 37564
rect 10380 37508 10436 37564
rect 10436 37508 10440 37564
rect 10376 37504 10440 37508
rect 10456 37564 10520 37568
rect 10456 37508 10460 37564
rect 10460 37508 10516 37564
rect 10516 37508 10520 37564
rect 10456 37504 10520 37508
rect 19480 37564 19544 37568
rect 19480 37508 19484 37564
rect 19484 37508 19540 37564
rect 19540 37508 19544 37564
rect 19480 37504 19544 37508
rect 19560 37564 19624 37568
rect 19560 37508 19564 37564
rect 19564 37508 19620 37564
rect 19620 37508 19624 37564
rect 19560 37504 19624 37508
rect 19640 37564 19704 37568
rect 19640 37508 19644 37564
rect 19644 37508 19700 37564
rect 19700 37508 19704 37564
rect 19640 37504 19704 37508
rect 19720 37564 19784 37568
rect 19720 37508 19724 37564
rect 19724 37508 19780 37564
rect 19780 37508 19784 37564
rect 19720 37504 19784 37508
rect 5584 37020 5648 37024
rect 5584 36964 5588 37020
rect 5588 36964 5644 37020
rect 5644 36964 5648 37020
rect 5584 36960 5648 36964
rect 5664 37020 5728 37024
rect 5664 36964 5668 37020
rect 5668 36964 5724 37020
rect 5724 36964 5728 37020
rect 5664 36960 5728 36964
rect 5744 37020 5808 37024
rect 5744 36964 5748 37020
rect 5748 36964 5804 37020
rect 5804 36964 5808 37020
rect 5744 36960 5808 36964
rect 5824 37020 5888 37024
rect 5824 36964 5828 37020
rect 5828 36964 5884 37020
rect 5884 36964 5888 37020
rect 5824 36960 5888 36964
rect 14848 37020 14912 37024
rect 14848 36964 14852 37020
rect 14852 36964 14908 37020
rect 14908 36964 14912 37020
rect 14848 36960 14912 36964
rect 14928 37020 14992 37024
rect 14928 36964 14932 37020
rect 14932 36964 14988 37020
rect 14988 36964 14992 37020
rect 14928 36960 14992 36964
rect 15008 37020 15072 37024
rect 15008 36964 15012 37020
rect 15012 36964 15068 37020
rect 15068 36964 15072 37020
rect 15008 36960 15072 36964
rect 15088 37020 15152 37024
rect 15088 36964 15092 37020
rect 15092 36964 15148 37020
rect 15148 36964 15152 37020
rect 15088 36960 15152 36964
rect 24112 37020 24176 37024
rect 24112 36964 24116 37020
rect 24116 36964 24172 37020
rect 24172 36964 24176 37020
rect 24112 36960 24176 36964
rect 24192 37020 24256 37024
rect 24192 36964 24196 37020
rect 24196 36964 24252 37020
rect 24252 36964 24256 37020
rect 24192 36960 24256 36964
rect 24272 37020 24336 37024
rect 24272 36964 24276 37020
rect 24276 36964 24332 37020
rect 24332 36964 24336 37020
rect 24272 36960 24336 36964
rect 24352 37020 24416 37024
rect 24352 36964 24356 37020
rect 24356 36964 24412 37020
rect 24412 36964 24416 37020
rect 24352 36960 24416 36964
rect 10216 36476 10280 36480
rect 10216 36420 10220 36476
rect 10220 36420 10276 36476
rect 10276 36420 10280 36476
rect 10216 36416 10280 36420
rect 10296 36476 10360 36480
rect 10296 36420 10300 36476
rect 10300 36420 10356 36476
rect 10356 36420 10360 36476
rect 10296 36416 10360 36420
rect 10376 36476 10440 36480
rect 10376 36420 10380 36476
rect 10380 36420 10436 36476
rect 10436 36420 10440 36476
rect 10376 36416 10440 36420
rect 10456 36476 10520 36480
rect 10456 36420 10460 36476
rect 10460 36420 10516 36476
rect 10516 36420 10520 36476
rect 10456 36416 10520 36420
rect 19480 36476 19544 36480
rect 19480 36420 19484 36476
rect 19484 36420 19540 36476
rect 19540 36420 19544 36476
rect 19480 36416 19544 36420
rect 19560 36476 19624 36480
rect 19560 36420 19564 36476
rect 19564 36420 19620 36476
rect 19620 36420 19624 36476
rect 19560 36416 19624 36420
rect 19640 36476 19704 36480
rect 19640 36420 19644 36476
rect 19644 36420 19700 36476
rect 19700 36420 19704 36476
rect 19640 36416 19704 36420
rect 19720 36476 19784 36480
rect 19720 36420 19724 36476
rect 19724 36420 19780 36476
rect 19780 36420 19784 36476
rect 19720 36416 19784 36420
rect 5584 35932 5648 35936
rect 5584 35876 5588 35932
rect 5588 35876 5644 35932
rect 5644 35876 5648 35932
rect 5584 35872 5648 35876
rect 5664 35932 5728 35936
rect 5664 35876 5668 35932
rect 5668 35876 5724 35932
rect 5724 35876 5728 35932
rect 5664 35872 5728 35876
rect 5744 35932 5808 35936
rect 5744 35876 5748 35932
rect 5748 35876 5804 35932
rect 5804 35876 5808 35932
rect 5744 35872 5808 35876
rect 5824 35932 5888 35936
rect 5824 35876 5828 35932
rect 5828 35876 5884 35932
rect 5884 35876 5888 35932
rect 5824 35872 5888 35876
rect 14848 35932 14912 35936
rect 14848 35876 14852 35932
rect 14852 35876 14908 35932
rect 14908 35876 14912 35932
rect 14848 35872 14912 35876
rect 14928 35932 14992 35936
rect 14928 35876 14932 35932
rect 14932 35876 14988 35932
rect 14988 35876 14992 35932
rect 14928 35872 14992 35876
rect 15008 35932 15072 35936
rect 15008 35876 15012 35932
rect 15012 35876 15068 35932
rect 15068 35876 15072 35932
rect 15008 35872 15072 35876
rect 15088 35932 15152 35936
rect 15088 35876 15092 35932
rect 15092 35876 15148 35932
rect 15148 35876 15152 35932
rect 15088 35872 15152 35876
rect 24112 35932 24176 35936
rect 24112 35876 24116 35932
rect 24116 35876 24172 35932
rect 24172 35876 24176 35932
rect 24112 35872 24176 35876
rect 24192 35932 24256 35936
rect 24192 35876 24196 35932
rect 24196 35876 24252 35932
rect 24252 35876 24256 35932
rect 24192 35872 24256 35876
rect 24272 35932 24336 35936
rect 24272 35876 24276 35932
rect 24276 35876 24332 35932
rect 24332 35876 24336 35932
rect 24272 35872 24336 35876
rect 24352 35932 24416 35936
rect 24352 35876 24356 35932
rect 24356 35876 24412 35932
rect 24412 35876 24416 35932
rect 24352 35872 24416 35876
rect 10216 35388 10280 35392
rect 10216 35332 10220 35388
rect 10220 35332 10276 35388
rect 10276 35332 10280 35388
rect 10216 35328 10280 35332
rect 10296 35388 10360 35392
rect 10296 35332 10300 35388
rect 10300 35332 10356 35388
rect 10356 35332 10360 35388
rect 10296 35328 10360 35332
rect 10376 35388 10440 35392
rect 10376 35332 10380 35388
rect 10380 35332 10436 35388
rect 10436 35332 10440 35388
rect 10376 35328 10440 35332
rect 10456 35388 10520 35392
rect 10456 35332 10460 35388
rect 10460 35332 10516 35388
rect 10516 35332 10520 35388
rect 10456 35328 10520 35332
rect 19480 35388 19544 35392
rect 19480 35332 19484 35388
rect 19484 35332 19540 35388
rect 19540 35332 19544 35388
rect 19480 35328 19544 35332
rect 19560 35388 19624 35392
rect 19560 35332 19564 35388
rect 19564 35332 19620 35388
rect 19620 35332 19624 35388
rect 19560 35328 19624 35332
rect 19640 35388 19704 35392
rect 19640 35332 19644 35388
rect 19644 35332 19700 35388
rect 19700 35332 19704 35388
rect 19640 35328 19704 35332
rect 19720 35388 19784 35392
rect 19720 35332 19724 35388
rect 19724 35332 19780 35388
rect 19780 35332 19784 35388
rect 19720 35328 19784 35332
rect 5584 34844 5648 34848
rect 5584 34788 5588 34844
rect 5588 34788 5644 34844
rect 5644 34788 5648 34844
rect 5584 34784 5648 34788
rect 5664 34844 5728 34848
rect 5664 34788 5668 34844
rect 5668 34788 5724 34844
rect 5724 34788 5728 34844
rect 5664 34784 5728 34788
rect 5744 34844 5808 34848
rect 5744 34788 5748 34844
rect 5748 34788 5804 34844
rect 5804 34788 5808 34844
rect 5744 34784 5808 34788
rect 5824 34844 5888 34848
rect 5824 34788 5828 34844
rect 5828 34788 5884 34844
rect 5884 34788 5888 34844
rect 5824 34784 5888 34788
rect 14848 34844 14912 34848
rect 14848 34788 14852 34844
rect 14852 34788 14908 34844
rect 14908 34788 14912 34844
rect 14848 34784 14912 34788
rect 14928 34844 14992 34848
rect 14928 34788 14932 34844
rect 14932 34788 14988 34844
rect 14988 34788 14992 34844
rect 14928 34784 14992 34788
rect 15008 34844 15072 34848
rect 15008 34788 15012 34844
rect 15012 34788 15068 34844
rect 15068 34788 15072 34844
rect 15008 34784 15072 34788
rect 15088 34844 15152 34848
rect 15088 34788 15092 34844
rect 15092 34788 15148 34844
rect 15148 34788 15152 34844
rect 15088 34784 15152 34788
rect 24112 34844 24176 34848
rect 24112 34788 24116 34844
rect 24116 34788 24172 34844
rect 24172 34788 24176 34844
rect 24112 34784 24176 34788
rect 24192 34844 24256 34848
rect 24192 34788 24196 34844
rect 24196 34788 24252 34844
rect 24252 34788 24256 34844
rect 24192 34784 24256 34788
rect 24272 34844 24336 34848
rect 24272 34788 24276 34844
rect 24276 34788 24332 34844
rect 24332 34788 24336 34844
rect 24272 34784 24336 34788
rect 24352 34844 24416 34848
rect 24352 34788 24356 34844
rect 24356 34788 24412 34844
rect 24412 34788 24416 34844
rect 24352 34784 24416 34788
rect 10216 34300 10280 34304
rect 10216 34244 10220 34300
rect 10220 34244 10276 34300
rect 10276 34244 10280 34300
rect 10216 34240 10280 34244
rect 10296 34300 10360 34304
rect 10296 34244 10300 34300
rect 10300 34244 10356 34300
rect 10356 34244 10360 34300
rect 10296 34240 10360 34244
rect 10376 34300 10440 34304
rect 10376 34244 10380 34300
rect 10380 34244 10436 34300
rect 10436 34244 10440 34300
rect 10376 34240 10440 34244
rect 10456 34300 10520 34304
rect 10456 34244 10460 34300
rect 10460 34244 10516 34300
rect 10516 34244 10520 34300
rect 10456 34240 10520 34244
rect 19480 34300 19544 34304
rect 19480 34244 19484 34300
rect 19484 34244 19540 34300
rect 19540 34244 19544 34300
rect 19480 34240 19544 34244
rect 19560 34300 19624 34304
rect 19560 34244 19564 34300
rect 19564 34244 19620 34300
rect 19620 34244 19624 34300
rect 19560 34240 19624 34244
rect 19640 34300 19704 34304
rect 19640 34244 19644 34300
rect 19644 34244 19700 34300
rect 19700 34244 19704 34300
rect 19640 34240 19704 34244
rect 19720 34300 19784 34304
rect 19720 34244 19724 34300
rect 19724 34244 19780 34300
rect 19780 34244 19784 34300
rect 19720 34240 19784 34244
rect 5584 33756 5648 33760
rect 5584 33700 5588 33756
rect 5588 33700 5644 33756
rect 5644 33700 5648 33756
rect 5584 33696 5648 33700
rect 5664 33756 5728 33760
rect 5664 33700 5668 33756
rect 5668 33700 5724 33756
rect 5724 33700 5728 33756
rect 5664 33696 5728 33700
rect 5744 33756 5808 33760
rect 5744 33700 5748 33756
rect 5748 33700 5804 33756
rect 5804 33700 5808 33756
rect 5744 33696 5808 33700
rect 5824 33756 5888 33760
rect 5824 33700 5828 33756
rect 5828 33700 5884 33756
rect 5884 33700 5888 33756
rect 5824 33696 5888 33700
rect 14848 33756 14912 33760
rect 14848 33700 14852 33756
rect 14852 33700 14908 33756
rect 14908 33700 14912 33756
rect 14848 33696 14912 33700
rect 14928 33756 14992 33760
rect 14928 33700 14932 33756
rect 14932 33700 14988 33756
rect 14988 33700 14992 33756
rect 14928 33696 14992 33700
rect 15008 33756 15072 33760
rect 15008 33700 15012 33756
rect 15012 33700 15068 33756
rect 15068 33700 15072 33756
rect 15008 33696 15072 33700
rect 15088 33756 15152 33760
rect 15088 33700 15092 33756
rect 15092 33700 15148 33756
rect 15148 33700 15152 33756
rect 15088 33696 15152 33700
rect 24112 33756 24176 33760
rect 24112 33700 24116 33756
rect 24116 33700 24172 33756
rect 24172 33700 24176 33756
rect 24112 33696 24176 33700
rect 24192 33756 24256 33760
rect 24192 33700 24196 33756
rect 24196 33700 24252 33756
rect 24252 33700 24256 33756
rect 24192 33696 24256 33700
rect 24272 33756 24336 33760
rect 24272 33700 24276 33756
rect 24276 33700 24332 33756
rect 24332 33700 24336 33756
rect 24272 33696 24336 33700
rect 24352 33756 24416 33760
rect 24352 33700 24356 33756
rect 24356 33700 24412 33756
rect 24412 33700 24416 33756
rect 24352 33696 24416 33700
rect 10216 33212 10280 33216
rect 10216 33156 10220 33212
rect 10220 33156 10276 33212
rect 10276 33156 10280 33212
rect 10216 33152 10280 33156
rect 10296 33212 10360 33216
rect 10296 33156 10300 33212
rect 10300 33156 10356 33212
rect 10356 33156 10360 33212
rect 10296 33152 10360 33156
rect 10376 33212 10440 33216
rect 10376 33156 10380 33212
rect 10380 33156 10436 33212
rect 10436 33156 10440 33212
rect 10376 33152 10440 33156
rect 10456 33212 10520 33216
rect 10456 33156 10460 33212
rect 10460 33156 10516 33212
rect 10516 33156 10520 33212
rect 10456 33152 10520 33156
rect 19480 33212 19544 33216
rect 19480 33156 19484 33212
rect 19484 33156 19540 33212
rect 19540 33156 19544 33212
rect 19480 33152 19544 33156
rect 19560 33212 19624 33216
rect 19560 33156 19564 33212
rect 19564 33156 19620 33212
rect 19620 33156 19624 33212
rect 19560 33152 19624 33156
rect 19640 33212 19704 33216
rect 19640 33156 19644 33212
rect 19644 33156 19700 33212
rect 19700 33156 19704 33212
rect 19640 33152 19704 33156
rect 19720 33212 19784 33216
rect 19720 33156 19724 33212
rect 19724 33156 19780 33212
rect 19780 33156 19784 33212
rect 19720 33152 19784 33156
rect 5584 32668 5648 32672
rect 5584 32612 5588 32668
rect 5588 32612 5644 32668
rect 5644 32612 5648 32668
rect 5584 32608 5648 32612
rect 5664 32668 5728 32672
rect 5664 32612 5668 32668
rect 5668 32612 5724 32668
rect 5724 32612 5728 32668
rect 5664 32608 5728 32612
rect 5744 32668 5808 32672
rect 5744 32612 5748 32668
rect 5748 32612 5804 32668
rect 5804 32612 5808 32668
rect 5744 32608 5808 32612
rect 5824 32668 5888 32672
rect 5824 32612 5828 32668
rect 5828 32612 5884 32668
rect 5884 32612 5888 32668
rect 5824 32608 5888 32612
rect 14848 32668 14912 32672
rect 14848 32612 14852 32668
rect 14852 32612 14908 32668
rect 14908 32612 14912 32668
rect 14848 32608 14912 32612
rect 14928 32668 14992 32672
rect 14928 32612 14932 32668
rect 14932 32612 14988 32668
rect 14988 32612 14992 32668
rect 14928 32608 14992 32612
rect 15008 32668 15072 32672
rect 15008 32612 15012 32668
rect 15012 32612 15068 32668
rect 15068 32612 15072 32668
rect 15008 32608 15072 32612
rect 15088 32668 15152 32672
rect 15088 32612 15092 32668
rect 15092 32612 15148 32668
rect 15148 32612 15152 32668
rect 15088 32608 15152 32612
rect 24112 32668 24176 32672
rect 24112 32612 24116 32668
rect 24116 32612 24172 32668
rect 24172 32612 24176 32668
rect 24112 32608 24176 32612
rect 24192 32668 24256 32672
rect 24192 32612 24196 32668
rect 24196 32612 24252 32668
rect 24252 32612 24256 32668
rect 24192 32608 24256 32612
rect 24272 32668 24336 32672
rect 24272 32612 24276 32668
rect 24276 32612 24332 32668
rect 24332 32612 24336 32668
rect 24272 32608 24336 32612
rect 24352 32668 24416 32672
rect 24352 32612 24356 32668
rect 24356 32612 24412 32668
rect 24412 32612 24416 32668
rect 24352 32608 24416 32612
rect 10216 32124 10280 32128
rect 10216 32068 10220 32124
rect 10220 32068 10276 32124
rect 10276 32068 10280 32124
rect 10216 32064 10280 32068
rect 10296 32124 10360 32128
rect 10296 32068 10300 32124
rect 10300 32068 10356 32124
rect 10356 32068 10360 32124
rect 10296 32064 10360 32068
rect 10376 32124 10440 32128
rect 10376 32068 10380 32124
rect 10380 32068 10436 32124
rect 10436 32068 10440 32124
rect 10376 32064 10440 32068
rect 10456 32124 10520 32128
rect 10456 32068 10460 32124
rect 10460 32068 10516 32124
rect 10516 32068 10520 32124
rect 10456 32064 10520 32068
rect 19480 32124 19544 32128
rect 19480 32068 19484 32124
rect 19484 32068 19540 32124
rect 19540 32068 19544 32124
rect 19480 32064 19544 32068
rect 19560 32124 19624 32128
rect 19560 32068 19564 32124
rect 19564 32068 19620 32124
rect 19620 32068 19624 32124
rect 19560 32064 19624 32068
rect 19640 32124 19704 32128
rect 19640 32068 19644 32124
rect 19644 32068 19700 32124
rect 19700 32068 19704 32124
rect 19640 32064 19704 32068
rect 19720 32124 19784 32128
rect 19720 32068 19724 32124
rect 19724 32068 19780 32124
rect 19780 32068 19784 32124
rect 19720 32064 19784 32068
rect 5584 31580 5648 31584
rect 5584 31524 5588 31580
rect 5588 31524 5644 31580
rect 5644 31524 5648 31580
rect 5584 31520 5648 31524
rect 5664 31580 5728 31584
rect 5664 31524 5668 31580
rect 5668 31524 5724 31580
rect 5724 31524 5728 31580
rect 5664 31520 5728 31524
rect 5744 31580 5808 31584
rect 5744 31524 5748 31580
rect 5748 31524 5804 31580
rect 5804 31524 5808 31580
rect 5744 31520 5808 31524
rect 5824 31580 5888 31584
rect 5824 31524 5828 31580
rect 5828 31524 5884 31580
rect 5884 31524 5888 31580
rect 5824 31520 5888 31524
rect 14848 31580 14912 31584
rect 14848 31524 14852 31580
rect 14852 31524 14908 31580
rect 14908 31524 14912 31580
rect 14848 31520 14912 31524
rect 14928 31580 14992 31584
rect 14928 31524 14932 31580
rect 14932 31524 14988 31580
rect 14988 31524 14992 31580
rect 14928 31520 14992 31524
rect 15008 31580 15072 31584
rect 15008 31524 15012 31580
rect 15012 31524 15068 31580
rect 15068 31524 15072 31580
rect 15008 31520 15072 31524
rect 15088 31580 15152 31584
rect 15088 31524 15092 31580
rect 15092 31524 15148 31580
rect 15148 31524 15152 31580
rect 15088 31520 15152 31524
rect 24112 31580 24176 31584
rect 24112 31524 24116 31580
rect 24116 31524 24172 31580
rect 24172 31524 24176 31580
rect 24112 31520 24176 31524
rect 24192 31580 24256 31584
rect 24192 31524 24196 31580
rect 24196 31524 24252 31580
rect 24252 31524 24256 31580
rect 24192 31520 24256 31524
rect 24272 31580 24336 31584
rect 24272 31524 24276 31580
rect 24276 31524 24332 31580
rect 24332 31524 24336 31580
rect 24272 31520 24336 31524
rect 24352 31580 24416 31584
rect 24352 31524 24356 31580
rect 24356 31524 24412 31580
rect 24412 31524 24416 31580
rect 24352 31520 24416 31524
rect 10216 31036 10280 31040
rect 10216 30980 10220 31036
rect 10220 30980 10276 31036
rect 10276 30980 10280 31036
rect 10216 30976 10280 30980
rect 10296 31036 10360 31040
rect 10296 30980 10300 31036
rect 10300 30980 10356 31036
rect 10356 30980 10360 31036
rect 10296 30976 10360 30980
rect 10376 31036 10440 31040
rect 10376 30980 10380 31036
rect 10380 30980 10436 31036
rect 10436 30980 10440 31036
rect 10376 30976 10440 30980
rect 10456 31036 10520 31040
rect 10456 30980 10460 31036
rect 10460 30980 10516 31036
rect 10516 30980 10520 31036
rect 10456 30976 10520 30980
rect 19480 31036 19544 31040
rect 19480 30980 19484 31036
rect 19484 30980 19540 31036
rect 19540 30980 19544 31036
rect 19480 30976 19544 30980
rect 19560 31036 19624 31040
rect 19560 30980 19564 31036
rect 19564 30980 19620 31036
rect 19620 30980 19624 31036
rect 19560 30976 19624 30980
rect 19640 31036 19704 31040
rect 19640 30980 19644 31036
rect 19644 30980 19700 31036
rect 19700 30980 19704 31036
rect 19640 30976 19704 30980
rect 19720 31036 19784 31040
rect 19720 30980 19724 31036
rect 19724 30980 19780 31036
rect 19780 30980 19784 31036
rect 19720 30976 19784 30980
rect 5584 30492 5648 30496
rect 5584 30436 5588 30492
rect 5588 30436 5644 30492
rect 5644 30436 5648 30492
rect 5584 30432 5648 30436
rect 5664 30492 5728 30496
rect 5664 30436 5668 30492
rect 5668 30436 5724 30492
rect 5724 30436 5728 30492
rect 5664 30432 5728 30436
rect 5744 30492 5808 30496
rect 5744 30436 5748 30492
rect 5748 30436 5804 30492
rect 5804 30436 5808 30492
rect 5744 30432 5808 30436
rect 5824 30492 5888 30496
rect 5824 30436 5828 30492
rect 5828 30436 5884 30492
rect 5884 30436 5888 30492
rect 5824 30432 5888 30436
rect 14848 30492 14912 30496
rect 14848 30436 14852 30492
rect 14852 30436 14908 30492
rect 14908 30436 14912 30492
rect 14848 30432 14912 30436
rect 14928 30492 14992 30496
rect 14928 30436 14932 30492
rect 14932 30436 14988 30492
rect 14988 30436 14992 30492
rect 14928 30432 14992 30436
rect 15008 30492 15072 30496
rect 15008 30436 15012 30492
rect 15012 30436 15068 30492
rect 15068 30436 15072 30492
rect 15008 30432 15072 30436
rect 15088 30492 15152 30496
rect 15088 30436 15092 30492
rect 15092 30436 15148 30492
rect 15148 30436 15152 30492
rect 15088 30432 15152 30436
rect 24112 30492 24176 30496
rect 24112 30436 24116 30492
rect 24116 30436 24172 30492
rect 24172 30436 24176 30492
rect 24112 30432 24176 30436
rect 24192 30492 24256 30496
rect 24192 30436 24196 30492
rect 24196 30436 24252 30492
rect 24252 30436 24256 30492
rect 24192 30432 24256 30436
rect 24272 30492 24336 30496
rect 24272 30436 24276 30492
rect 24276 30436 24332 30492
rect 24332 30436 24336 30492
rect 24272 30432 24336 30436
rect 24352 30492 24416 30496
rect 24352 30436 24356 30492
rect 24356 30436 24412 30492
rect 24412 30436 24416 30492
rect 24352 30432 24416 30436
rect 10216 29948 10280 29952
rect 10216 29892 10220 29948
rect 10220 29892 10276 29948
rect 10276 29892 10280 29948
rect 10216 29888 10280 29892
rect 10296 29948 10360 29952
rect 10296 29892 10300 29948
rect 10300 29892 10356 29948
rect 10356 29892 10360 29948
rect 10296 29888 10360 29892
rect 10376 29948 10440 29952
rect 10376 29892 10380 29948
rect 10380 29892 10436 29948
rect 10436 29892 10440 29948
rect 10376 29888 10440 29892
rect 10456 29948 10520 29952
rect 10456 29892 10460 29948
rect 10460 29892 10516 29948
rect 10516 29892 10520 29948
rect 10456 29888 10520 29892
rect 19480 29948 19544 29952
rect 19480 29892 19484 29948
rect 19484 29892 19540 29948
rect 19540 29892 19544 29948
rect 19480 29888 19544 29892
rect 19560 29948 19624 29952
rect 19560 29892 19564 29948
rect 19564 29892 19620 29948
rect 19620 29892 19624 29948
rect 19560 29888 19624 29892
rect 19640 29948 19704 29952
rect 19640 29892 19644 29948
rect 19644 29892 19700 29948
rect 19700 29892 19704 29948
rect 19640 29888 19704 29892
rect 19720 29948 19784 29952
rect 19720 29892 19724 29948
rect 19724 29892 19780 29948
rect 19780 29892 19784 29948
rect 19720 29888 19784 29892
rect 5584 29404 5648 29408
rect 5584 29348 5588 29404
rect 5588 29348 5644 29404
rect 5644 29348 5648 29404
rect 5584 29344 5648 29348
rect 5664 29404 5728 29408
rect 5664 29348 5668 29404
rect 5668 29348 5724 29404
rect 5724 29348 5728 29404
rect 5664 29344 5728 29348
rect 5744 29404 5808 29408
rect 5744 29348 5748 29404
rect 5748 29348 5804 29404
rect 5804 29348 5808 29404
rect 5744 29344 5808 29348
rect 5824 29404 5888 29408
rect 5824 29348 5828 29404
rect 5828 29348 5884 29404
rect 5884 29348 5888 29404
rect 5824 29344 5888 29348
rect 14848 29404 14912 29408
rect 14848 29348 14852 29404
rect 14852 29348 14908 29404
rect 14908 29348 14912 29404
rect 14848 29344 14912 29348
rect 14928 29404 14992 29408
rect 14928 29348 14932 29404
rect 14932 29348 14988 29404
rect 14988 29348 14992 29404
rect 14928 29344 14992 29348
rect 15008 29404 15072 29408
rect 15008 29348 15012 29404
rect 15012 29348 15068 29404
rect 15068 29348 15072 29404
rect 15008 29344 15072 29348
rect 15088 29404 15152 29408
rect 15088 29348 15092 29404
rect 15092 29348 15148 29404
rect 15148 29348 15152 29404
rect 15088 29344 15152 29348
rect 24112 29404 24176 29408
rect 24112 29348 24116 29404
rect 24116 29348 24172 29404
rect 24172 29348 24176 29404
rect 24112 29344 24176 29348
rect 24192 29404 24256 29408
rect 24192 29348 24196 29404
rect 24196 29348 24252 29404
rect 24252 29348 24256 29404
rect 24192 29344 24256 29348
rect 24272 29404 24336 29408
rect 24272 29348 24276 29404
rect 24276 29348 24332 29404
rect 24332 29348 24336 29404
rect 24272 29344 24336 29348
rect 24352 29404 24416 29408
rect 24352 29348 24356 29404
rect 24356 29348 24412 29404
rect 24412 29348 24416 29404
rect 24352 29344 24416 29348
rect 10216 28860 10280 28864
rect 10216 28804 10220 28860
rect 10220 28804 10276 28860
rect 10276 28804 10280 28860
rect 10216 28800 10280 28804
rect 10296 28860 10360 28864
rect 10296 28804 10300 28860
rect 10300 28804 10356 28860
rect 10356 28804 10360 28860
rect 10296 28800 10360 28804
rect 10376 28860 10440 28864
rect 10376 28804 10380 28860
rect 10380 28804 10436 28860
rect 10436 28804 10440 28860
rect 10376 28800 10440 28804
rect 10456 28860 10520 28864
rect 10456 28804 10460 28860
rect 10460 28804 10516 28860
rect 10516 28804 10520 28860
rect 10456 28800 10520 28804
rect 19480 28860 19544 28864
rect 19480 28804 19484 28860
rect 19484 28804 19540 28860
rect 19540 28804 19544 28860
rect 19480 28800 19544 28804
rect 19560 28860 19624 28864
rect 19560 28804 19564 28860
rect 19564 28804 19620 28860
rect 19620 28804 19624 28860
rect 19560 28800 19624 28804
rect 19640 28860 19704 28864
rect 19640 28804 19644 28860
rect 19644 28804 19700 28860
rect 19700 28804 19704 28860
rect 19640 28800 19704 28804
rect 19720 28860 19784 28864
rect 19720 28804 19724 28860
rect 19724 28804 19780 28860
rect 19780 28804 19784 28860
rect 19720 28800 19784 28804
rect 5584 28316 5648 28320
rect 5584 28260 5588 28316
rect 5588 28260 5644 28316
rect 5644 28260 5648 28316
rect 5584 28256 5648 28260
rect 5664 28316 5728 28320
rect 5664 28260 5668 28316
rect 5668 28260 5724 28316
rect 5724 28260 5728 28316
rect 5664 28256 5728 28260
rect 5744 28316 5808 28320
rect 5744 28260 5748 28316
rect 5748 28260 5804 28316
rect 5804 28260 5808 28316
rect 5744 28256 5808 28260
rect 5824 28316 5888 28320
rect 5824 28260 5828 28316
rect 5828 28260 5884 28316
rect 5884 28260 5888 28316
rect 5824 28256 5888 28260
rect 14848 28316 14912 28320
rect 14848 28260 14852 28316
rect 14852 28260 14908 28316
rect 14908 28260 14912 28316
rect 14848 28256 14912 28260
rect 14928 28316 14992 28320
rect 14928 28260 14932 28316
rect 14932 28260 14988 28316
rect 14988 28260 14992 28316
rect 14928 28256 14992 28260
rect 15008 28316 15072 28320
rect 15008 28260 15012 28316
rect 15012 28260 15068 28316
rect 15068 28260 15072 28316
rect 15008 28256 15072 28260
rect 15088 28316 15152 28320
rect 15088 28260 15092 28316
rect 15092 28260 15148 28316
rect 15148 28260 15152 28316
rect 15088 28256 15152 28260
rect 24112 28316 24176 28320
rect 24112 28260 24116 28316
rect 24116 28260 24172 28316
rect 24172 28260 24176 28316
rect 24112 28256 24176 28260
rect 24192 28316 24256 28320
rect 24192 28260 24196 28316
rect 24196 28260 24252 28316
rect 24252 28260 24256 28316
rect 24192 28256 24256 28260
rect 24272 28316 24336 28320
rect 24272 28260 24276 28316
rect 24276 28260 24332 28316
rect 24332 28260 24336 28316
rect 24272 28256 24336 28260
rect 24352 28316 24416 28320
rect 24352 28260 24356 28316
rect 24356 28260 24412 28316
rect 24412 28260 24416 28316
rect 24352 28256 24416 28260
rect 10216 27772 10280 27776
rect 10216 27716 10220 27772
rect 10220 27716 10276 27772
rect 10276 27716 10280 27772
rect 10216 27712 10280 27716
rect 10296 27772 10360 27776
rect 10296 27716 10300 27772
rect 10300 27716 10356 27772
rect 10356 27716 10360 27772
rect 10296 27712 10360 27716
rect 10376 27772 10440 27776
rect 10376 27716 10380 27772
rect 10380 27716 10436 27772
rect 10436 27716 10440 27772
rect 10376 27712 10440 27716
rect 10456 27772 10520 27776
rect 10456 27716 10460 27772
rect 10460 27716 10516 27772
rect 10516 27716 10520 27772
rect 10456 27712 10520 27716
rect 19480 27772 19544 27776
rect 19480 27716 19484 27772
rect 19484 27716 19540 27772
rect 19540 27716 19544 27772
rect 19480 27712 19544 27716
rect 19560 27772 19624 27776
rect 19560 27716 19564 27772
rect 19564 27716 19620 27772
rect 19620 27716 19624 27772
rect 19560 27712 19624 27716
rect 19640 27772 19704 27776
rect 19640 27716 19644 27772
rect 19644 27716 19700 27772
rect 19700 27716 19704 27772
rect 19640 27712 19704 27716
rect 19720 27772 19784 27776
rect 19720 27716 19724 27772
rect 19724 27716 19780 27772
rect 19780 27716 19784 27772
rect 19720 27712 19784 27716
rect 5584 27228 5648 27232
rect 5584 27172 5588 27228
rect 5588 27172 5644 27228
rect 5644 27172 5648 27228
rect 5584 27168 5648 27172
rect 5664 27228 5728 27232
rect 5664 27172 5668 27228
rect 5668 27172 5724 27228
rect 5724 27172 5728 27228
rect 5664 27168 5728 27172
rect 5744 27228 5808 27232
rect 5744 27172 5748 27228
rect 5748 27172 5804 27228
rect 5804 27172 5808 27228
rect 5744 27168 5808 27172
rect 5824 27228 5888 27232
rect 5824 27172 5828 27228
rect 5828 27172 5884 27228
rect 5884 27172 5888 27228
rect 5824 27168 5888 27172
rect 14848 27228 14912 27232
rect 14848 27172 14852 27228
rect 14852 27172 14908 27228
rect 14908 27172 14912 27228
rect 14848 27168 14912 27172
rect 14928 27228 14992 27232
rect 14928 27172 14932 27228
rect 14932 27172 14988 27228
rect 14988 27172 14992 27228
rect 14928 27168 14992 27172
rect 15008 27228 15072 27232
rect 15008 27172 15012 27228
rect 15012 27172 15068 27228
rect 15068 27172 15072 27228
rect 15008 27168 15072 27172
rect 15088 27228 15152 27232
rect 15088 27172 15092 27228
rect 15092 27172 15148 27228
rect 15148 27172 15152 27228
rect 15088 27168 15152 27172
rect 24112 27228 24176 27232
rect 24112 27172 24116 27228
rect 24116 27172 24172 27228
rect 24172 27172 24176 27228
rect 24112 27168 24176 27172
rect 24192 27228 24256 27232
rect 24192 27172 24196 27228
rect 24196 27172 24252 27228
rect 24252 27172 24256 27228
rect 24192 27168 24256 27172
rect 24272 27228 24336 27232
rect 24272 27172 24276 27228
rect 24276 27172 24332 27228
rect 24332 27172 24336 27228
rect 24272 27168 24336 27172
rect 24352 27228 24416 27232
rect 24352 27172 24356 27228
rect 24356 27172 24412 27228
rect 24412 27172 24416 27228
rect 24352 27168 24416 27172
rect 10216 26684 10280 26688
rect 10216 26628 10220 26684
rect 10220 26628 10276 26684
rect 10276 26628 10280 26684
rect 10216 26624 10280 26628
rect 10296 26684 10360 26688
rect 10296 26628 10300 26684
rect 10300 26628 10356 26684
rect 10356 26628 10360 26684
rect 10296 26624 10360 26628
rect 10376 26684 10440 26688
rect 10376 26628 10380 26684
rect 10380 26628 10436 26684
rect 10436 26628 10440 26684
rect 10376 26624 10440 26628
rect 10456 26684 10520 26688
rect 10456 26628 10460 26684
rect 10460 26628 10516 26684
rect 10516 26628 10520 26684
rect 10456 26624 10520 26628
rect 19480 26684 19544 26688
rect 19480 26628 19484 26684
rect 19484 26628 19540 26684
rect 19540 26628 19544 26684
rect 19480 26624 19544 26628
rect 19560 26684 19624 26688
rect 19560 26628 19564 26684
rect 19564 26628 19620 26684
rect 19620 26628 19624 26684
rect 19560 26624 19624 26628
rect 19640 26684 19704 26688
rect 19640 26628 19644 26684
rect 19644 26628 19700 26684
rect 19700 26628 19704 26684
rect 19640 26624 19704 26628
rect 19720 26684 19784 26688
rect 19720 26628 19724 26684
rect 19724 26628 19780 26684
rect 19780 26628 19784 26684
rect 19720 26624 19784 26628
rect 5584 26140 5648 26144
rect 5584 26084 5588 26140
rect 5588 26084 5644 26140
rect 5644 26084 5648 26140
rect 5584 26080 5648 26084
rect 5664 26140 5728 26144
rect 5664 26084 5668 26140
rect 5668 26084 5724 26140
rect 5724 26084 5728 26140
rect 5664 26080 5728 26084
rect 5744 26140 5808 26144
rect 5744 26084 5748 26140
rect 5748 26084 5804 26140
rect 5804 26084 5808 26140
rect 5744 26080 5808 26084
rect 5824 26140 5888 26144
rect 5824 26084 5828 26140
rect 5828 26084 5884 26140
rect 5884 26084 5888 26140
rect 5824 26080 5888 26084
rect 14848 26140 14912 26144
rect 14848 26084 14852 26140
rect 14852 26084 14908 26140
rect 14908 26084 14912 26140
rect 14848 26080 14912 26084
rect 14928 26140 14992 26144
rect 14928 26084 14932 26140
rect 14932 26084 14988 26140
rect 14988 26084 14992 26140
rect 14928 26080 14992 26084
rect 15008 26140 15072 26144
rect 15008 26084 15012 26140
rect 15012 26084 15068 26140
rect 15068 26084 15072 26140
rect 15008 26080 15072 26084
rect 15088 26140 15152 26144
rect 15088 26084 15092 26140
rect 15092 26084 15148 26140
rect 15148 26084 15152 26140
rect 15088 26080 15152 26084
rect 24112 26140 24176 26144
rect 24112 26084 24116 26140
rect 24116 26084 24172 26140
rect 24172 26084 24176 26140
rect 24112 26080 24176 26084
rect 24192 26140 24256 26144
rect 24192 26084 24196 26140
rect 24196 26084 24252 26140
rect 24252 26084 24256 26140
rect 24192 26080 24256 26084
rect 24272 26140 24336 26144
rect 24272 26084 24276 26140
rect 24276 26084 24332 26140
rect 24332 26084 24336 26140
rect 24272 26080 24336 26084
rect 24352 26140 24416 26144
rect 24352 26084 24356 26140
rect 24356 26084 24412 26140
rect 24412 26084 24416 26140
rect 24352 26080 24416 26084
rect 10216 25596 10280 25600
rect 10216 25540 10220 25596
rect 10220 25540 10276 25596
rect 10276 25540 10280 25596
rect 10216 25536 10280 25540
rect 10296 25596 10360 25600
rect 10296 25540 10300 25596
rect 10300 25540 10356 25596
rect 10356 25540 10360 25596
rect 10296 25536 10360 25540
rect 10376 25596 10440 25600
rect 10376 25540 10380 25596
rect 10380 25540 10436 25596
rect 10436 25540 10440 25596
rect 10376 25536 10440 25540
rect 10456 25596 10520 25600
rect 10456 25540 10460 25596
rect 10460 25540 10516 25596
rect 10516 25540 10520 25596
rect 10456 25536 10520 25540
rect 19480 25596 19544 25600
rect 19480 25540 19484 25596
rect 19484 25540 19540 25596
rect 19540 25540 19544 25596
rect 19480 25536 19544 25540
rect 19560 25596 19624 25600
rect 19560 25540 19564 25596
rect 19564 25540 19620 25596
rect 19620 25540 19624 25596
rect 19560 25536 19624 25540
rect 19640 25596 19704 25600
rect 19640 25540 19644 25596
rect 19644 25540 19700 25596
rect 19700 25540 19704 25596
rect 19640 25536 19704 25540
rect 19720 25596 19784 25600
rect 19720 25540 19724 25596
rect 19724 25540 19780 25596
rect 19780 25540 19784 25596
rect 19720 25536 19784 25540
rect 5584 25052 5648 25056
rect 5584 24996 5588 25052
rect 5588 24996 5644 25052
rect 5644 24996 5648 25052
rect 5584 24992 5648 24996
rect 5664 25052 5728 25056
rect 5664 24996 5668 25052
rect 5668 24996 5724 25052
rect 5724 24996 5728 25052
rect 5664 24992 5728 24996
rect 5744 25052 5808 25056
rect 5744 24996 5748 25052
rect 5748 24996 5804 25052
rect 5804 24996 5808 25052
rect 5744 24992 5808 24996
rect 5824 25052 5888 25056
rect 5824 24996 5828 25052
rect 5828 24996 5884 25052
rect 5884 24996 5888 25052
rect 5824 24992 5888 24996
rect 14848 25052 14912 25056
rect 14848 24996 14852 25052
rect 14852 24996 14908 25052
rect 14908 24996 14912 25052
rect 14848 24992 14912 24996
rect 14928 25052 14992 25056
rect 14928 24996 14932 25052
rect 14932 24996 14988 25052
rect 14988 24996 14992 25052
rect 14928 24992 14992 24996
rect 15008 25052 15072 25056
rect 15008 24996 15012 25052
rect 15012 24996 15068 25052
rect 15068 24996 15072 25052
rect 15008 24992 15072 24996
rect 15088 25052 15152 25056
rect 15088 24996 15092 25052
rect 15092 24996 15148 25052
rect 15148 24996 15152 25052
rect 15088 24992 15152 24996
rect 24112 25052 24176 25056
rect 24112 24996 24116 25052
rect 24116 24996 24172 25052
rect 24172 24996 24176 25052
rect 24112 24992 24176 24996
rect 24192 25052 24256 25056
rect 24192 24996 24196 25052
rect 24196 24996 24252 25052
rect 24252 24996 24256 25052
rect 24192 24992 24256 24996
rect 24272 25052 24336 25056
rect 24272 24996 24276 25052
rect 24276 24996 24332 25052
rect 24332 24996 24336 25052
rect 24272 24992 24336 24996
rect 24352 25052 24416 25056
rect 24352 24996 24356 25052
rect 24356 24996 24412 25052
rect 24412 24996 24416 25052
rect 24352 24992 24416 24996
rect 10216 24508 10280 24512
rect 10216 24452 10220 24508
rect 10220 24452 10276 24508
rect 10276 24452 10280 24508
rect 10216 24448 10280 24452
rect 10296 24508 10360 24512
rect 10296 24452 10300 24508
rect 10300 24452 10356 24508
rect 10356 24452 10360 24508
rect 10296 24448 10360 24452
rect 10376 24508 10440 24512
rect 10376 24452 10380 24508
rect 10380 24452 10436 24508
rect 10436 24452 10440 24508
rect 10376 24448 10440 24452
rect 10456 24508 10520 24512
rect 10456 24452 10460 24508
rect 10460 24452 10516 24508
rect 10516 24452 10520 24508
rect 10456 24448 10520 24452
rect 19480 24508 19544 24512
rect 19480 24452 19484 24508
rect 19484 24452 19540 24508
rect 19540 24452 19544 24508
rect 19480 24448 19544 24452
rect 19560 24508 19624 24512
rect 19560 24452 19564 24508
rect 19564 24452 19620 24508
rect 19620 24452 19624 24508
rect 19560 24448 19624 24452
rect 19640 24508 19704 24512
rect 19640 24452 19644 24508
rect 19644 24452 19700 24508
rect 19700 24452 19704 24508
rect 19640 24448 19704 24452
rect 19720 24508 19784 24512
rect 19720 24452 19724 24508
rect 19724 24452 19780 24508
rect 19780 24452 19784 24508
rect 19720 24448 19784 24452
rect 5584 23964 5648 23968
rect 5584 23908 5588 23964
rect 5588 23908 5644 23964
rect 5644 23908 5648 23964
rect 5584 23904 5648 23908
rect 5664 23964 5728 23968
rect 5664 23908 5668 23964
rect 5668 23908 5724 23964
rect 5724 23908 5728 23964
rect 5664 23904 5728 23908
rect 5744 23964 5808 23968
rect 5744 23908 5748 23964
rect 5748 23908 5804 23964
rect 5804 23908 5808 23964
rect 5744 23904 5808 23908
rect 5824 23964 5888 23968
rect 5824 23908 5828 23964
rect 5828 23908 5884 23964
rect 5884 23908 5888 23964
rect 5824 23904 5888 23908
rect 14848 23964 14912 23968
rect 14848 23908 14852 23964
rect 14852 23908 14908 23964
rect 14908 23908 14912 23964
rect 14848 23904 14912 23908
rect 14928 23964 14992 23968
rect 14928 23908 14932 23964
rect 14932 23908 14988 23964
rect 14988 23908 14992 23964
rect 14928 23904 14992 23908
rect 15008 23964 15072 23968
rect 15008 23908 15012 23964
rect 15012 23908 15068 23964
rect 15068 23908 15072 23964
rect 15008 23904 15072 23908
rect 15088 23964 15152 23968
rect 15088 23908 15092 23964
rect 15092 23908 15148 23964
rect 15148 23908 15152 23964
rect 15088 23904 15152 23908
rect 24112 23964 24176 23968
rect 24112 23908 24116 23964
rect 24116 23908 24172 23964
rect 24172 23908 24176 23964
rect 24112 23904 24176 23908
rect 24192 23964 24256 23968
rect 24192 23908 24196 23964
rect 24196 23908 24252 23964
rect 24252 23908 24256 23964
rect 24192 23904 24256 23908
rect 24272 23964 24336 23968
rect 24272 23908 24276 23964
rect 24276 23908 24332 23964
rect 24332 23908 24336 23964
rect 24272 23904 24336 23908
rect 24352 23964 24416 23968
rect 24352 23908 24356 23964
rect 24356 23908 24412 23964
rect 24412 23908 24416 23964
rect 24352 23904 24416 23908
rect 10216 23420 10280 23424
rect 10216 23364 10220 23420
rect 10220 23364 10276 23420
rect 10276 23364 10280 23420
rect 10216 23360 10280 23364
rect 10296 23420 10360 23424
rect 10296 23364 10300 23420
rect 10300 23364 10356 23420
rect 10356 23364 10360 23420
rect 10296 23360 10360 23364
rect 10376 23420 10440 23424
rect 10376 23364 10380 23420
rect 10380 23364 10436 23420
rect 10436 23364 10440 23420
rect 10376 23360 10440 23364
rect 10456 23420 10520 23424
rect 10456 23364 10460 23420
rect 10460 23364 10516 23420
rect 10516 23364 10520 23420
rect 10456 23360 10520 23364
rect 19480 23420 19544 23424
rect 19480 23364 19484 23420
rect 19484 23364 19540 23420
rect 19540 23364 19544 23420
rect 19480 23360 19544 23364
rect 19560 23420 19624 23424
rect 19560 23364 19564 23420
rect 19564 23364 19620 23420
rect 19620 23364 19624 23420
rect 19560 23360 19624 23364
rect 19640 23420 19704 23424
rect 19640 23364 19644 23420
rect 19644 23364 19700 23420
rect 19700 23364 19704 23420
rect 19640 23360 19704 23364
rect 19720 23420 19784 23424
rect 19720 23364 19724 23420
rect 19724 23364 19780 23420
rect 19780 23364 19784 23420
rect 19720 23360 19784 23364
rect 5584 22876 5648 22880
rect 5584 22820 5588 22876
rect 5588 22820 5644 22876
rect 5644 22820 5648 22876
rect 5584 22816 5648 22820
rect 5664 22876 5728 22880
rect 5664 22820 5668 22876
rect 5668 22820 5724 22876
rect 5724 22820 5728 22876
rect 5664 22816 5728 22820
rect 5744 22876 5808 22880
rect 5744 22820 5748 22876
rect 5748 22820 5804 22876
rect 5804 22820 5808 22876
rect 5744 22816 5808 22820
rect 5824 22876 5888 22880
rect 5824 22820 5828 22876
rect 5828 22820 5884 22876
rect 5884 22820 5888 22876
rect 5824 22816 5888 22820
rect 14848 22876 14912 22880
rect 14848 22820 14852 22876
rect 14852 22820 14908 22876
rect 14908 22820 14912 22876
rect 14848 22816 14912 22820
rect 14928 22876 14992 22880
rect 14928 22820 14932 22876
rect 14932 22820 14988 22876
rect 14988 22820 14992 22876
rect 14928 22816 14992 22820
rect 15008 22876 15072 22880
rect 15008 22820 15012 22876
rect 15012 22820 15068 22876
rect 15068 22820 15072 22876
rect 15008 22816 15072 22820
rect 15088 22876 15152 22880
rect 15088 22820 15092 22876
rect 15092 22820 15148 22876
rect 15148 22820 15152 22876
rect 15088 22816 15152 22820
rect 24112 22876 24176 22880
rect 24112 22820 24116 22876
rect 24116 22820 24172 22876
rect 24172 22820 24176 22876
rect 24112 22816 24176 22820
rect 24192 22876 24256 22880
rect 24192 22820 24196 22876
rect 24196 22820 24252 22876
rect 24252 22820 24256 22876
rect 24192 22816 24256 22820
rect 24272 22876 24336 22880
rect 24272 22820 24276 22876
rect 24276 22820 24332 22876
rect 24332 22820 24336 22876
rect 24272 22816 24336 22820
rect 24352 22876 24416 22880
rect 24352 22820 24356 22876
rect 24356 22820 24412 22876
rect 24412 22820 24416 22876
rect 24352 22816 24416 22820
rect 10216 22332 10280 22336
rect 10216 22276 10220 22332
rect 10220 22276 10276 22332
rect 10276 22276 10280 22332
rect 10216 22272 10280 22276
rect 10296 22332 10360 22336
rect 10296 22276 10300 22332
rect 10300 22276 10356 22332
rect 10356 22276 10360 22332
rect 10296 22272 10360 22276
rect 10376 22332 10440 22336
rect 10376 22276 10380 22332
rect 10380 22276 10436 22332
rect 10436 22276 10440 22332
rect 10376 22272 10440 22276
rect 10456 22332 10520 22336
rect 10456 22276 10460 22332
rect 10460 22276 10516 22332
rect 10516 22276 10520 22332
rect 10456 22272 10520 22276
rect 19480 22332 19544 22336
rect 19480 22276 19484 22332
rect 19484 22276 19540 22332
rect 19540 22276 19544 22332
rect 19480 22272 19544 22276
rect 19560 22332 19624 22336
rect 19560 22276 19564 22332
rect 19564 22276 19620 22332
rect 19620 22276 19624 22332
rect 19560 22272 19624 22276
rect 19640 22332 19704 22336
rect 19640 22276 19644 22332
rect 19644 22276 19700 22332
rect 19700 22276 19704 22332
rect 19640 22272 19704 22276
rect 19720 22332 19784 22336
rect 19720 22276 19724 22332
rect 19724 22276 19780 22332
rect 19780 22276 19784 22332
rect 19720 22272 19784 22276
rect 5584 21788 5648 21792
rect 5584 21732 5588 21788
rect 5588 21732 5644 21788
rect 5644 21732 5648 21788
rect 5584 21728 5648 21732
rect 5664 21788 5728 21792
rect 5664 21732 5668 21788
rect 5668 21732 5724 21788
rect 5724 21732 5728 21788
rect 5664 21728 5728 21732
rect 5744 21788 5808 21792
rect 5744 21732 5748 21788
rect 5748 21732 5804 21788
rect 5804 21732 5808 21788
rect 5744 21728 5808 21732
rect 5824 21788 5888 21792
rect 5824 21732 5828 21788
rect 5828 21732 5884 21788
rect 5884 21732 5888 21788
rect 5824 21728 5888 21732
rect 14848 21788 14912 21792
rect 14848 21732 14852 21788
rect 14852 21732 14908 21788
rect 14908 21732 14912 21788
rect 14848 21728 14912 21732
rect 14928 21788 14992 21792
rect 14928 21732 14932 21788
rect 14932 21732 14988 21788
rect 14988 21732 14992 21788
rect 14928 21728 14992 21732
rect 15008 21788 15072 21792
rect 15008 21732 15012 21788
rect 15012 21732 15068 21788
rect 15068 21732 15072 21788
rect 15008 21728 15072 21732
rect 15088 21788 15152 21792
rect 15088 21732 15092 21788
rect 15092 21732 15148 21788
rect 15148 21732 15152 21788
rect 15088 21728 15152 21732
rect 10216 21244 10280 21248
rect 10216 21188 10220 21244
rect 10220 21188 10276 21244
rect 10276 21188 10280 21244
rect 10216 21184 10280 21188
rect 10296 21244 10360 21248
rect 10296 21188 10300 21244
rect 10300 21188 10356 21244
rect 10356 21188 10360 21244
rect 10296 21184 10360 21188
rect 10376 21244 10440 21248
rect 10376 21188 10380 21244
rect 10380 21188 10436 21244
rect 10436 21188 10440 21244
rect 10376 21184 10440 21188
rect 10456 21244 10520 21248
rect 10456 21188 10460 21244
rect 10460 21188 10516 21244
rect 10516 21188 10520 21244
rect 10456 21184 10520 21188
rect 24112 21788 24176 21792
rect 24112 21732 24116 21788
rect 24116 21732 24172 21788
rect 24172 21732 24176 21788
rect 24112 21728 24176 21732
rect 24192 21788 24256 21792
rect 24192 21732 24196 21788
rect 24196 21732 24252 21788
rect 24252 21732 24256 21788
rect 24192 21728 24256 21732
rect 24272 21788 24336 21792
rect 24272 21732 24276 21788
rect 24276 21732 24332 21788
rect 24332 21732 24336 21788
rect 24272 21728 24336 21732
rect 24352 21788 24416 21792
rect 24352 21732 24356 21788
rect 24356 21732 24412 21788
rect 24412 21732 24416 21788
rect 24352 21728 24416 21732
rect 19480 21244 19544 21248
rect 19480 21188 19484 21244
rect 19484 21188 19540 21244
rect 19540 21188 19544 21244
rect 19480 21184 19544 21188
rect 19560 21244 19624 21248
rect 19560 21188 19564 21244
rect 19564 21188 19620 21244
rect 19620 21188 19624 21244
rect 19560 21184 19624 21188
rect 19640 21244 19704 21248
rect 19640 21188 19644 21244
rect 19644 21188 19700 21244
rect 19700 21188 19704 21244
rect 19640 21184 19704 21188
rect 19720 21244 19784 21248
rect 19720 21188 19724 21244
rect 19724 21188 19780 21244
rect 19780 21188 19784 21244
rect 19720 21184 19784 21188
rect 5584 20700 5648 20704
rect 5584 20644 5588 20700
rect 5588 20644 5644 20700
rect 5644 20644 5648 20700
rect 5584 20640 5648 20644
rect 5664 20700 5728 20704
rect 5664 20644 5668 20700
rect 5668 20644 5724 20700
rect 5724 20644 5728 20700
rect 5664 20640 5728 20644
rect 5744 20700 5808 20704
rect 5744 20644 5748 20700
rect 5748 20644 5804 20700
rect 5804 20644 5808 20700
rect 5744 20640 5808 20644
rect 5824 20700 5888 20704
rect 5824 20644 5828 20700
rect 5828 20644 5884 20700
rect 5884 20644 5888 20700
rect 5824 20640 5888 20644
rect 14848 20700 14912 20704
rect 14848 20644 14852 20700
rect 14852 20644 14908 20700
rect 14908 20644 14912 20700
rect 14848 20640 14912 20644
rect 14928 20700 14992 20704
rect 14928 20644 14932 20700
rect 14932 20644 14988 20700
rect 14988 20644 14992 20700
rect 14928 20640 14992 20644
rect 15008 20700 15072 20704
rect 15008 20644 15012 20700
rect 15012 20644 15068 20700
rect 15068 20644 15072 20700
rect 15008 20640 15072 20644
rect 15088 20700 15152 20704
rect 15088 20644 15092 20700
rect 15092 20644 15148 20700
rect 15148 20644 15152 20700
rect 15088 20640 15152 20644
rect 24112 20700 24176 20704
rect 24112 20644 24116 20700
rect 24116 20644 24172 20700
rect 24172 20644 24176 20700
rect 24112 20640 24176 20644
rect 24192 20700 24256 20704
rect 24192 20644 24196 20700
rect 24196 20644 24252 20700
rect 24252 20644 24256 20700
rect 24192 20640 24256 20644
rect 24272 20700 24336 20704
rect 24272 20644 24276 20700
rect 24276 20644 24332 20700
rect 24332 20644 24336 20700
rect 24272 20640 24336 20644
rect 24352 20700 24416 20704
rect 24352 20644 24356 20700
rect 24356 20644 24412 20700
rect 24412 20644 24416 20700
rect 24352 20640 24416 20644
rect 10216 20156 10280 20160
rect 10216 20100 10220 20156
rect 10220 20100 10276 20156
rect 10276 20100 10280 20156
rect 10216 20096 10280 20100
rect 10296 20156 10360 20160
rect 10296 20100 10300 20156
rect 10300 20100 10356 20156
rect 10356 20100 10360 20156
rect 10296 20096 10360 20100
rect 10376 20156 10440 20160
rect 10376 20100 10380 20156
rect 10380 20100 10436 20156
rect 10436 20100 10440 20156
rect 10376 20096 10440 20100
rect 10456 20156 10520 20160
rect 10456 20100 10460 20156
rect 10460 20100 10516 20156
rect 10516 20100 10520 20156
rect 10456 20096 10520 20100
rect 19480 20156 19544 20160
rect 19480 20100 19484 20156
rect 19484 20100 19540 20156
rect 19540 20100 19544 20156
rect 19480 20096 19544 20100
rect 19560 20156 19624 20160
rect 19560 20100 19564 20156
rect 19564 20100 19620 20156
rect 19620 20100 19624 20156
rect 19560 20096 19624 20100
rect 19640 20156 19704 20160
rect 19640 20100 19644 20156
rect 19644 20100 19700 20156
rect 19700 20100 19704 20156
rect 19640 20096 19704 20100
rect 19720 20156 19784 20160
rect 19720 20100 19724 20156
rect 19724 20100 19780 20156
rect 19780 20100 19784 20156
rect 19720 20096 19784 20100
rect 5584 19612 5648 19616
rect 5584 19556 5588 19612
rect 5588 19556 5644 19612
rect 5644 19556 5648 19612
rect 5584 19552 5648 19556
rect 5664 19612 5728 19616
rect 5664 19556 5668 19612
rect 5668 19556 5724 19612
rect 5724 19556 5728 19612
rect 5664 19552 5728 19556
rect 5744 19612 5808 19616
rect 5744 19556 5748 19612
rect 5748 19556 5804 19612
rect 5804 19556 5808 19612
rect 5744 19552 5808 19556
rect 5824 19612 5888 19616
rect 5824 19556 5828 19612
rect 5828 19556 5884 19612
rect 5884 19556 5888 19612
rect 5824 19552 5888 19556
rect 14848 19612 14912 19616
rect 14848 19556 14852 19612
rect 14852 19556 14908 19612
rect 14908 19556 14912 19612
rect 14848 19552 14912 19556
rect 14928 19612 14992 19616
rect 14928 19556 14932 19612
rect 14932 19556 14988 19612
rect 14988 19556 14992 19612
rect 14928 19552 14992 19556
rect 15008 19612 15072 19616
rect 15008 19556 15012 19612
rect 15012 19556 15068 19612
rect 15068 19556 15072 19612
rect 15008 19552 15072 19556
rect 15088 19612 15152 19616
rect 15088 19556 15092 19612
rect 15092 19556 15148 19612
rect 15148 19556 15152 19612
rect 15088 19552 15152 19556
rect 10216 19068 10280 19072
rect 10216 19012 10220 19068
rect 10220 19012 10276 19068
rect 10276 19012 10280 19068
rect 10216 19008 10280 19012
rect 10296 19068 10360 19072
rect 10296 19012 10300 19068
rect 10300 19012 10356 19068
rect 10356 19012 10360 19068
rect 10296 19008 10360 19012
rect 10376 19068 10440 19072
rect 10376 19012 10380 19068
rect 10380 19012 10436 19068
rect 10436 19012 10440 19068
rect 10376 19008 10440 19012
rect 10456 19068 10520 19072
rect 10456 19012 10460 19068
rect 10460 19012 10516 19068
rect 10516 19012 10520 19068
rect 10456 19008 10520 19012
rect 5584 18524 5648 18528
rect 5584 18468 5588 18524
rect 5588 18468 5644 18524
rect 5644 18468 5648 18524
rect 5584 18464 5648 18468
rect 5664 18524 5728 18528
rect 5664 18468 5668 18524
rect 5668 18468 5724 18524
rect 5724 18468 5728 18524
rect 5664 18464 5728 18468
rect 5744 18524 5808 18528
rect 5744 18468 5748 18524
rect 5748 18468 5804 18524
rect 5804 18468 5808 18524
rect 5744 18464 5808 18468
rect 5824 18524 5888 18528
rect 5824 18468 5828 18524
rect 5828 18468 5884 18524
rect 5884 18468 5888 18524
rect 5824 18464 5888 18468
rect 24112 19612 24176 19616
rect 24112 19556 24116 19612
rect 24116 19556 24172 19612
rect 24172 19556 24176 19612
rect 24112 19552 24176 19556
rect 24192 19612 24256 19616
rect 24192 19556 24196 19612
rect 24196 19556 24252 19612
rect 24252 19556 24256 19612
rect 24192 19552 24256 19556
rect 24272 19612 24336 19616
rect 24272 19556 24276 19612
rect 24276 19556 24332 19612
rect 24332 19556 24336 19612
rect 24272 19552 24336 19556
rect 24352 19612 24416 19616
rect 24352 19556 24356 19612
rect 24356 19556 24412 19612
rect 24412 19556 24416 19612
rect 24352 19552 24416 19556
rect 19480 19068 19544 19072
rect 19480 19012 19484 19068
rect 19484 19012 19540 19068
rect 19540 19012 19544 19068
rect 19480 19008 19544 19012
rect 19560 19068 19624 19072
rect 19560 19012 19564 19068
rect 19564 19012 19620 19068
rect 19620 19012 19624 19068
rect 19560 19008 19624 19012
rect 19640 19068 19704 19072
rect 19640 19012 19644 19068
rect 19644 19012 19700 19068
rect 19700 19012 19704 19068
rect 19640 19008 19704 19012
rect 19720 19068 19784 19072
rect 19720 19012 19724 19068
rect 19724 19012 19780 19068
rect 19780 19012 19784 19068
rect 19720 19008 19784 19012
rect 14848 18524 14912 18528
rect 14848 18468 14852 18524
rect 14852 18468 14908 18524
rect 14908 18468 14912 18524
rect 14848 18464 14912 18468
rect 14928 18524 14992 18528
rect 14928 18468 14932 18524
rect 14932 18468 14988 18524
rect 14988 18468 14992 18524
rect 14928 18464 14992 18468
rect 15008 18524 15072 18528
rect 15008 18468 15012 18524
rect 15012 18468 15068 18524
rect 15068 18468 15072 18524
rect 15008 18464 15072 18468
rect 15088 18524 15152 18528
rect 15088 18468 15092 18524
rect 15092 18468 15148 18524
rect 15148 18468 15152 18524
rect 15088 18464 15152 18468
rect 24112 18524 24176 18528
rect 24112 18468 24116 18524
rect 24116 18468 24172 18524
rect 24172 18468 24176 18524
rect 24112 18464 24176 18468
rect 24192 18524 24256 18528
rect 24192 18468 24196 18524
rect 24196 18468 24252 18524
rect 24252 18468 24256 18524
rect 24192 18464 24256 18468
rect 24272 18524 24336 18528
rect 24272 18468 24276 18524
rect 24276 18468 24332 18524
rect 24332 18468 24336 18524
rect 24272 18464 24336 18468
rect 24352 18524 24416 18528
rect 24352 18468 24356 18524
rect 24356 18468 24412 18524
rect 24412 18468 24416 18524
rect 24352 18464 24416 18468
rect 10216 17980 10280 17984
rect 10216 17924 10220 17980
rect 10220 17924 10276 17980
rect 10276 17924 10280 17980
rect 10216 17920 10280 17924
rect 10296 17980 10360 17984
rect 10296 17924 10300 17980
rect 10300 17924 10356 17980
rect 10356 17924 10360 17980
rect 10296 17920 10360 17924
rect 10376 17980 10440 17984
rect 10376 17924 10380 17980
rect 10380 17924 10436 17980
rect 10436 17924 10440 17980
rect 10376 17920 10440 17924
rect 10456 17980 10520 17984
rect 10456 17924 10460 17980
rect 10460 17924 10516 17980
rect 10516 17924 10520 17980
rect 10456 17920 10520 17924
rect 19480 17980 19544 17984
rect 19480 17924 19484 17980
rect 19484 17924 19540 17980
rect 19540 17924 19544 17980
rect 19480 17920 19544 17924
rect 19560 17980 19624 17984
rect 19560 17924 19564 17980
rect 19564 17924 19620 17980
rect 19620 17924 19624 17980
rect 19560 17920 19624 17924
rect 19640 17980 19704 17984
rect 19640 17924 19644 17980
rect 19644 17924 19700 17980
rect 19700 17924 19704 17980
rect 19640 17920 19704 17924
rect 19720 17980 19784 17984
rect 19720 17924 19724 17980
rect 19724 17924 19780 17980
rect 19780 17924 19784 17980
rect 19720 17920 19784 17924
rect 5584 17436 5648 17440
rect 5584 17380 5588 17436
rect 5588 17380 5644 17436
rect 5644 17380 5648 17436
rect 5584 17376 5648 17380
rect 5664 17436 5728 17440
rect 5664 17380 5668 17436
rect 5668 17380 5724 17436
rect 5724 17380 5728 17436
rect 5664 17376 5728 17380
rect 5744 17436 5808 17440
rect 5744 17380 5748 17436
rect 5748 17380 5804 17436
rect 5804 17380 5808 17436
rect 5744 17376 5808 17380
rect 5824 17436 5888 17440
rect 5824 17380 5828 17436
rect 5828 17380 5884 17436
rect 5884 17380 5888 17436
rect 5824 17376 5888 17380
rect 14848 17436 14912 17440
rect 14848 17380 14852 17436
rect 14852 17380 14908 17436
rect 14908 17380 14912 17436
rect 14848 17376 14912 17380
rect 14928 17436 14992 17440
rect 14928 17380 14932 17436
rect 14932 17380 14988 17436
rect 14988 17380 14992 17436
rect 14928 17376 14992 17380
rect 15008 17436 15072 17440
rect 15008 17380 15012 17436
rect 15012 17380 15068 17436
rect 15068 17380 15072 17436
rect 15008 17376 15072 17380
rect 15088 17436 15152 17440
rect 15088 17380 15092 17436
rect 15092 17380 15148 17436
rect 15148 17380 15152 17436
rect 15088 17376 15152 17380
rect 24112 17436 24176 17440
rect 24112 17380 24116 17436
rect 24116 17380 24172 17436
rect 24172 17380 24176 17436
rect 24112 17376 24176 17380
rect 24192 17436 24256 17440
rect 24192 17380 24196 17436
rect 24196 17380 24252 17436
rect 24252 17380 24256 17436
rect 24192 17376 24256 17380
rect 24272 17436 24336 17440
rect 24272 17380 24276 17436
rect 24276 17380 24332 17436
rect 24332 17380 24336 17436
rect 24272 17376 24336 17380
rect 24352 17436 24416 17440
rect 24352 17380 24356 17436
rect 24356 17380 24412 17436
rect 24412 17380 24416 17436
rect 24352 17376 24416 17380
rect 10216 16892 10280 16896
rect 10216 16836 10220 16892
rect 10220 16836 10276 16892
rect 10276 16836 10280 16892
rect 10216 16832 10280 16836
rect 10296 16892 10360 16896
rect 10296 16836 10300 16892
rect 10300 16836 10356 16892
rect 10356 16836 10360 16892
rect 10296 16832 10360 16836
rect 10376 16892 10440 16896
rect 10376 16836 10380 16892
rect 10380 16836 10436 16892
rect 10436 16836 10440 16892
rect 10376 16832 10440 16836
rect 10456 16892 10520 16896
rect 10456 16836 10460 16892
rect 10460 16836 10516 16892
rect 10516 16836 10520 16892
rect 10456 16832 10520 16836
rect 19480 16892 19544 16896
rect 19480 16836 19484 16892
rect 19484 16836 19540 16892
rect 19540 16836 19544 16892
rect 19480 16832 19544 16836
rect 19560 16892 19624 16896
rect 19560 16836 19564 16892
rect 19564 16836 19620 16892
rect 19620 16836 19624 16892
rect 19560 16832 19624 16836
rect 19640 16892 19704 16896
rect 19640 16836 19644 16892
rect 19644 16836 19700 16892
rect 19700 16836 19704 16892
rect 19640 16832 19704 16836
rect 19720 16892 19784 16896
rect 19720 16836 19724 16892
rect 19724 16836 19780 16892
rect 19780 16836 19784 16892
rect 19720 16832 19784 16836
rect 5584 16348 5648 16352
rect 5584 16292 5588 16348
rect 5588 16292 5644 16348
rect 5644 16292 5648 16348
rect 5584 16288 5648 16292
rect 5664 16348 5728 16352
rect 5664 16292 5668 16348
rect 5668 16292 5724 16348
rect 5724 16292 5728 16348
rect 5664 16288 5728 16292
rect 5744 16348 5808 16352
rect 5744 16292 5748 16348
rect 5748 16292 5804 16348
rect 5804 16292 5808 16348
rect 5744 16288 5808 16292
rect 5824 16348 5888 16352
rect 5824 16292 5828 16348
rect 5828 16292 5884 16348
rect 5884 16292 5888 16348
rect 5824 16288 5888 16292
rect 14848 16348 14912 16352
rect 14848 16292 14852 16348
rect 14852 16292 14908 16348
rect 14908 16292 14912 16348
rect 14848 16288 14912 16292
rect 14928 16348 14992 16352
rect 14928 16292 14932 16348
rect 14932 16292 14988 16348
rect 14988 16292 14992 16348
rect 14928 16288 14992 16292
rect 15008 16348 15072 16352
rect 15008 16292 15012 16348
rect 15012 16292 15068 16348
rect 15068 16292 15072 16348
rect 15008 16288 15072 16292
rect 15088 16348 15152 16352
rect 15088 16292 15092 16348
rect 15092 16292 15148 16348
rect 15148 16292 15152 16348
rect 15088 16288 15152 16292
rect 24112 16348 24176 16352
rect 24112 16292 24116 16348
rect 24116 16292 24172 16348
rect 24172 16292 24176 16348
rect 24112 16288 24176 16292
rect 24192 16348 24256 16352
rect 24192 16292 24196 16348
rect 24196 16292 24252 16348
rect 24252 16292 24256 16348
rect 24192 16288 24256 16292
rect 24272 16348 24336 16352
rect 24272 16292 24276 16348
rect 24276 16292 24332 16348
rect 24332 16292 24336 16348
rect 24272 16288 24336 16292
rect 24352 16348 24416 16352
rect 24352 16292 24356 16348
rect 24356 16292 24412 16348
rect 24412 16292 24416 16348
rect 24352 16288 24416 16292
rect 10216 15804 10280 15808
rect 10216 15748 10220 15804
rect 10220 15748 10276 15804
rect 10276 15748 10280 15804
rect 10216 15744 10280 15748
rect 10296 15804 10360 15808
rect 10296 15748 10300 15804
rect 10300 15748 10356 15804
rect 10356 15748 10360 15804
rect 10296 15744 10360 15748
rect 10376 15804 10440 15808
rect 10376 15748 10380 15804
rect 10380 15748 10436 15804
rect 10436 15748 10440 15804
rect 10376 15744 10440 15748
rect 10456 15804 10520 15808
rect 10456 15748 10460 15804
rect 10460 15748 10516 15804
rect 10516 15748 10520 15804
rect 10456 15744 10520 15748
rect 19480 15804 19544 15808
rect 19480 15748 19484 15804
rect 19484 15748 19540 15804
rect 19540 15748 19544 15804
rect 19480 15744 19544 15748
rect 19560 15804 19624 15808
rect 19560 15748 19564 15804
rect 19564 15748 19620 15804
rect 19620 15748 19624 15804
rect 19560 15744 19624 15748
rect 19640 15804 19704 15808
rect 19640 15748 19644 15804
rect 19644 15748 19700 15804
rect 19700 15748 19704 15804
rect 19640 15744 19704 15748
rect 19720 15804 19784 15808
rect 19720 15748 19724 15804
rect 19724 15748 19780 15804
rect 19780 15748 19784 15804
rect 19720 15744 19784 15748
rect 5584 15260 5648 15264
rect 5584 15204 5588 15260
rect 5588 15204 5644 15260
rect 5644 15204 5648 15260
rect 5584 15200 5648 15204
rect 5664 15260 5728 15264
rect 5664 15204 5668 15260
rect 5668 15204 5724 15260
rect 5724 15204 5728 15260
rect 5664 15200 5728 15204
rect 5744 15260 5808 15264
rect 5744 15204 5748 15260
rect 5748 15204 5804 15260
rect 5804 15204 5808 15260
rect 5744 15200 5808 15204
rect 5824 15260 5888 15264
rect 5824 15204 5828 15260
rect 5828 15204 5884 15260
rect 5884 15204 5888 15260
rect 5824 15200 5888 15204
rect 14848 15260 14912 15264
rect 14848 15204 14852 15260
rect 14852 15204 14908 15260
rect 14908 15204 14912 15260
rect 14848 15200 14912 15204
rect 14928 15260 14992 15264
rect 14928 15204 14932 15260
rect 14932 15204 14988 15260
rect 14988 15204 14992 15260
rect 14928 15200 14992 15204
rect 15008 15260 15072 15264
rect 15008 15204 15012 15260
rect 15012 15204 15068 15260
rect 15068 15204 15072 15260
rect 15008 15200 15072 15204
rect 15088 15260 15152 15264
rect 15088 15204 15092 15260
rect 15092 15204 15148 15260
rect 15148 15204 15152 15260
rect 15088 15200 15152 15204
rect 24112 15260 24176 15264
rect 24112 15204 24116 15260
rect 24116 15204 24172 15260
rect 24172 15204 24176 15260
rect 24112 15200 24176 15204
rect 24192 15260 24256 15264
rect 24192 15204 24196 15260
rect 24196 15204 24252 15260
rect 24252 15204 24256 15260
rect 24192 15200 24256 15204
rect 24272 15260 24336 15264
rect 24272 15204 24276 15260
rect 24276 15204 24332 15260
rect 24332 15204 24336 15260
rect 24272 15200 24336 15204
rect 24352 15260 24416 15264
rect 24352 15204 24356 15260
rect 24356 15204 24412 15260
rect 24412 15204 24416 15260
rect 24352 15200 24416 15204
rect 10216 14716 10280 14720
rect 10216 14660 10220 14716
rect 10220 14660 10276 14716
rect 10276 14660 10280 14716
rect 10216 14656 10280 14660
rect 10296 14716 10360 14720
rect 10296 14660 10300 14716
rect 10300 14660 10356 14716
rect 10356 14660 10360 14716
rect 10296 14656 10360 14660
rect 10376 14716 10440 14720
rect 10376 14660 10380 14716
rect 10380 14660 10436 14716
rect 10436 14660 10440 14716
rect 10376 14656 10440 14660
rect 10456 14716 10520 14720
rect 10456 14660 10460 14716
rect 10460 14660 10516 14716
rect 10516 14660 10520 14716
rect 10456 14656 10520 14660
rect 19480 14716 19544 14720
rect 19480 14660 19484 14716
rect 19484 14660 19540 14716
rect 19540 14660 19544 14716
rect 19480 14656 19544 14660
rect 19560 14716 19624 14720
rect 19560 14660 19564 14716
rect 19564 14660 19620 14716
rect 19620 14660 19624 14716
rect 19560 14656 19624 14660
rect 19640 14716 19704 14720
rect 19640 14660 19644 14716
rect 19644 14660 19700 14716
rect 19700 14660 19704 14716
rect 19640 14656 19704 14660
rect 19720 14716 19784 14720
rect 19720 14660 19724 14716
rect 19724 14660 19780 14716
rect 19780 14660 19784 14716
rect 19720 14656 19784 14660
rect 5584 14172 5648 14176
rect 5584 14116 5588 14172
rect 5588 14116 5644 14172
rect 5644 14116 5648 14172
rect 5584 14112 5648 14116
rect 5664 14172 5728 14176
rect 5664 14116 5668 14172
rect 5668 14116 5724 14172
rect 5724 14116 5728 14172
rect 5664 14112 5728 14116
rect 5744 14172 5808 14176
rect 5744 14116 5748 14172
rect 5748 14116 5804 14172
rect 5804 14116 5808 14172
rect 5744 14112 5808 14116
rect 5824 14172 5888 14176
rect 5824 14116 5828 14172
rect 5828 14116 5884 14172
rect 5884 14116 5888 14172
rect 5824 14112 5888 14116
rect 14848 14172 14912 14176
rect 14848 14116 14852 14172
rect 14852 14116 14908 14172
rect 14908 14116 14912 14172
rect 14848 14112 14912 14116
rect 14928 14172 14992 14176
rect 14928 14116 14932 14172
rect 14932 14116 14988 14172
rect 14988 14116 14992 14172
rect 14928 14112 14992 14116
rect 15008 14172 15072 14176
rect 15008 14116 15012 14172
rect 15012 14116 15068 14172
rect 15068 14116 15072 14172
rect 15008 14112 15072 14116
rect 15088 14172 15152 14176
rect 15088 14116 15092 14172
rect 15092 14116 15148 14172
rect 15148 14116 15152 14172
rect 15088 14112 15152 14116
rect 24112 14172 24176 14176
rect 24112 14116 24116 14172
rect 24116 14116 24172 14172
rect 24172 14116 24176 14172
rect 24112 14112 24176 14116
rect 24192 14172 24256 14176
rect 24192 14116 24196 14172
rect 24196 14116 24252 14172
rect 24252 14116 24256 14172
rect 24192 14112 24256 14116
rect 24272 14172 24336 14176
rect 24272 14116 24276 14172
rect 24276 14116 24332 14172
rect 24332 14116 24336 14172
rect 24272 14112 24336 14116
rect 24352 14172 24416 14176
rect 24352 14116 24356 14172
rect 24356 14116 24412 14172
rect 24412 14116 24416 14172
rect 24352 14112 24416 14116
rect 10216 13628 10280 13632
rect 10216 13572 10220 13628
rect 10220 13572 10276 13628
rect 10276 13572 10280 13628
rect 10216 13568 10280 13572
rect 10296 13628 10360 13632
rect 10296 13572 10300 13628
rect 10300 13572 10356 13628
rect 10356 13572 10360 13628
rect 10296 13568 10360 13572
rect 10376 13628 10440 13632
rect 10376 13572 10380 13628
rect 10380 13572 10436 13628
rect 10436 13572 10440 13628
rect 10376 13568 10440 13572
rect 10456 13628 10520 13632
rect 10456 13572 10460 13628
rect 10460 13572 10516 13628
rect 10516 13572 10520 13628
rect 10456 13568 10520 13572
rect 19480 13628 19544 13632
rect 19480 13572 19484 13628
rect 19484 13572 19540 13628
rect 19540 13572 19544 13628
rect 19480 13568 19544 13572
rect 19560 13628 19624 13632
rect 19560 13572 19564 13628
rect 19564 13572 19620 13628
rect 19620 13572 19624 13628
rect 19560 13568 19624 13572
rect 19640 13628 19704 13632
rect 19640 13572 19644 13628
rect 19644 13572 19700 13628
rect 19700 13572 19704 13628
rect 19640 13568 19704 13572
rect 19720 13628 19784 13632
rect 19720 13572 19724 13628
rect 19724 13572 19780 13628
rect 19780 13572 19784 13628
rect 19720 13568 19784 13572
rect 5584 13084 5648 13088
rect 5584 13028 5588 13084
rect 5588 13028 5644 13084
rect 5644 13028 5648 13084
rect 5584 13024 5648 13028
rect 5664 13084 5728 13088
rect 5664 13028 5668 13084
rect 5668 13028 5724 13084
rect 5724 13028 5728 13084
rect 5664 13024 5728 13028
rect 5744 13084 5808 13088
rect 5744 13028 5748 13084
rect 5748 13028 5804 13084
rect 5804 13028 5808 13084
rect 5744 13024 5808 13028
rect 5824 13084 5888 13088
rect 5824 13028 5828 13084
rect 5828 13028 5884 13084
rect 5884 13028 5888 13084
rect 5824 13024 5888 13028
rect 14848 13084 14912 13088
rect 14848 13028 14852 13084
rect 14852 13028 14908 13084
rect 14908 13028 14912 13084
rect 14848 13024 14912 13028
rect 14928 13084 14992 13088
rect 14928 13028 14932 13084
rect 14932 13028 14988 13084
rect 14988 13028 14992 13084
rect 14928 13024 14992 13028
rect 15008 13084 15072 13088
rect 15008 13028 15012 13084
rect 15012 13028 15068 13084
rect 15068 13028 15072 13084
rect 15008 13024 15072 13028
rect 15088 13084 15152 13088
rect 15088 13028 15092 13084
rect 15092 13028 15148 13084
rect 15148 13028 15152 13084
rect 15088 13024 15152 13028
rect 24112 13084 24176 13088
rect 24112 13028 24116 13084
rect 24116 13028 24172 13084
rect 24172 13028 24176 13084
rect 24112 13024 24176 13028
rect 24192 13084 24256 13088
rect 24192 13028 24196 13084
rect 24196 13028 24252 13084
rect 24252 13028 24256 13084
rect 24192 13024 24256 13028
rect 24272 13084 24336 13088
rect 24272 13028 24276 13084
rect 24276 13028 24332 13084
rect 24332 13028 24336 13084
rect 24272 13024 24336 13028
rect 24352 13084 24416 13088
rect 24352 13028 24356 13084
rect 24356 13028 24412 13084
rect 24412 13028 24416 13084
rect 24352 13024 24416 13028
rect 10216 12540 10280 12544
rect 10216 12484 10220 12540
rect 10220 12484 10276 12540
rect 10276 12484 10280 12540
rect 10216 12480 10280 12484
rect 10296 12540 10360 12544
rect 10296 12484 10300 12540
rect 10300 12484 10356 12540
rect 10356 12484 10360 12540
rect 10296 12480 10360 12484
rect 10376 12540 10440 12544
rect 10376 12484 10380 12540
rect 10380 12484 10436 12540
rect 10436 12484 10440 12540
rect 10376 12480 10440 12484
rect 10456 12540 10520 12544
rect 10456 12484 10460 12540
rect 10460 12484 10516 12540
rect 10516 12484 10520 12540
rect 10456 12480 10520 12484
rect 19480 12540 19544 12544
rect 19480 12484 19484 12540
rect 19484 12484 19540 12540
rect 19540 12484 19544 12540
rect 19480 12480 19544 12484
rect 19560 12540 19624 12544
rect 19560 12484 19564 12540
rect 19564 12484 19620 12540
rect 19620 12484 19624 12540
rect 19560 12480 19624 12484
rect 19640 12540 19704 12544
rect 19640 12484 19644 12540
rect 19644 12484 19700 12540
rect 19700 12484 19704 12540
rect 19640 12480 19704 12484
rect 19720 12540 19784 12544
rect 19720 12484 19724 12540
rect 19724 12484 19780 12540
rect 19780 12484 19784 12540
rect 19720 12480 19784 12484
rect 5584 11996 5648 12000
rect 5584 11940 5588 11996
rect 5588 11940 5644 11996
rect 5644 11940 5648 11996
rect 5584 11936 5648 11940
rect 5664 11996 5728 12000
rect 5664 11940 5668 11996
rect 5668 11940 5724 11996
rect 5724 11940 5728 11996
rect 5664 11936 5728 11940
rect 5744 11996 5808 12000
rect 5744 11940 5748 11996
rect 5748 11940 5804 11996
rect 5804 11940 5808 11996
rect 5744 11936 5808 11940
rect 5824 11996 5888 12000
rect 5824 11940 5828 11996
rect 5828 11940 5884 11996
rect 5884 11940 5888 11996
rect 5824 11936 5888 11940
rect 14848 11996 14912 12000
rect 14848 11940 14852 11996
rect 14852 11940 14908 11996
rect 14908 11940 14912 11996
rect 14848 11936 14912 11940
rect 14928 11996 14992 12000
rect 14928 11940 14932 11996
rect 14932 11940 14988 11996
rect 14988 11940 14992 11996
rect 14928 11936 14992 11940
rect 15008 11996 15072 12000
rect 15008 11940 15012 11996
rect 15012 11940 15068 11996
rect 15068 11940 15072 11996
rect 15008 11936 15072 11940
rect 15088 11996 15152 12000
rect 15088 11940 15092 11996
rect 15092 11940 15148 11996
rect 15148 11940 15152 11996
rect 15088 11936 15152 11940
rect 24112 11996 24176 12000
rect 24112 11940 24116 11996
rect 24116 11940 24172 11996
rect 24172 11940 24176 11996
rect 24112 11936 24176 11940
rect 24192 11996 24256 12000
rect 24192 11940 24196 11996
rect 24196 11940 24252 11996
rect 24252 11940 24256 11996
rect 24192 11936 24256 11940
rect 24272 11996 24336 12000
rect 24272 11940 24276 11996
rect 24276 11940 24332 11996
rect 24332 11940 24336 11996
rect 24272 11936 24336 11940
rect 24352 11996 24416 12000
rect 24352 11940 24356 11996
rect 24356 11940 24412 11996
rect 24412 11940 24416 11996
rect 24352 11936 24416 11940
rect 10216 11452 10280 11456
rect 10216 11396 10220 11452
rect 10220 11396 10276 11452
rect 10276 11396 10280 11452
rect 10216 11392 10280 11396
rect 10296 11452 10360 11456
rect 10296 11396 10300 11452
rect 10300 11396 10356 11452
rect 10356 11396 10360 11452
rect 10296 11392 10360 11396
rect 10376 11452 10440 11456
rect 10376 11396 10380 11452
rect 10380 11396 10436 11452
rect 10436 11396 10440 11452
rect 10376 11392 10440 11396
rect 10456 11452 10520 11456
rect 10456 11396 10460 11452
rect 10460 11396 10516 11452
rect 10516 11396 10520 11452
rect 10456 11392 10520 11396
rect 19480 11452 19544 11456
rect 19480 11396 19484 11452
rect 19484 11396 19540 11452
rect 19540 11396 19544 11452
rect 19480 11392 19544 11396
rect 19560 11452 19624 11456
rect 19560 11396 19564 11452
rect 19564 11396 19620 11452
rect 19620 11396 19624 11452
rect 19560 11392 19624 11396
rect 19640 11452 19704 11456
rect 19640 11396 19644 11452
rect 19644 11396 19700 11452
rect 19700 11396 19704 11452
rect 19640 11392 19704 11396
rect 19720 11452 19784 11456
rect 19720 11396 19724 11452
rect 19724 11396 19780 11452
rect 19780 11396 19784 11452
rect 19720 11392 19784 11396
rect 5584 10908 5648 10912
rect 5584 10852 5588 10908
rect 5588 10852 5644 10908
rect 5644 10852 5648 10908
rect 5584 10848 5648 10852
rect 5664 10908 5728 10912
rect 5664 10852 5668 10908
rect 5668 10852 5724 10908
rect 5724 10852 5728 10908
rect 5664 10848 5728 10852
rect 5744 10908 5808 10912
rect 5744 10852 5748 10908
rect 5748 10852 5804 10908
rect 5804 10852 5808 10908
rect 5744 10848 5808 10852
rect 5824 10908 5888 10912
rect 5824 10852 5828 10908
rect 5828 10852 5884 10908
rect 5884 10852 5888 10908
rect 5824 10848 5888 10852
rect 14848 10908 14912 10912
rect 14848 10852 14852 10908
rect 14852 10852 14908 10908
rect 14908 10852 14912 10908
rect 14848 10848 14912 10852
rect 14928 10908 14992 10912
rect 14928 10852 14932 10908
rect 14932 10852 14988 10908
rect 14988 10852 14992 10908
rect 14928 10848 14992 10852
rect 15008 10908 15072 10912
rect 15008 10852 15012 10908
rect 15012 10852 15068 10908
rect 15068 10852 15072 10908
rect 15008 10848 15072 10852
rect 15088 10908 15152 10912
rect 15088 10852 15092 10908
rect 15092 10852 15148 10908
rect 15148 10852 15152 10908
rect 15088 10848 15152 10852
rect 24112 10908 24176 10912
rect 24112 10852 24116 10908
rect 24116 10852 24172 10908
rect 24172 10852 24176 10908
rect 24112 10848 24176 10852
rect 24192 10908 24256 10912
rect 24192 10852 24196 10908
rect 24196 10852 24252 10908
rect 24252 10852 24256 10908
rect 24192 10848 24256 10852
rect 24272 10908 24336 10912
rect 24272 10852 24276 10908
rect 24276 10852 24332 10908
rect 24332 10852 24336 10908
rect 24272 10848 24336 10852
rect 24352 10908 24416 10912
rect 24352 10852 24356 10908
rect 24356 10852 24412 10908
rect 24412 10852 24416 10908
rect 24352 10848 24416 10852
rect 10216 10364 10280 10368
rect 10216 10308 10220 10364
rect 10220 10308 10276 10364
rect 10276 10308 10280 10364
rect 10216 10304 10280 10308
rect 10296 10364 10360 10368
rect 10296 10308 10300 10364
rect 10300 10308 10356 10364
rect 10356 10308 10360 10364
rect 10296 10304 10360 10308
rect 10376 10364 10440 10368
rect 10376 10308 10380 10364
rect 10380 10308 10436 10364
rect 10436 10308 10440 10364
rect 10376 10304 10440 10308
rect 10456 10364 10520 10368
rect 10456 10308 10460 10364
rect 10460 10308 10516 10364
rect 10516 10308 10520 10364
rect 10456 10304 10520 10308
rect 19480 10364 19544 10368
rect 19480 10308 19484 10364
rect 19484 10308 19540 10364
rect 19540 10308 19544 10364
rect 19480 10304 19544 10308
rect 19560 10364 19624 10368
rect 19560 10308 19564 10364
rect 19564 10308 19620 10364
rect 19620 10308 19624 10364
rect 19560 10304 19624 10308
rect 19640 10364 19704 10368
rect 19640 10308 19644 10364
rect 19644 10308 19700 10364
rect 19700 10308 19704 10364
rect 19640 10304 19704 10308
rect 19720 10364 19784 10368
rect 19720 10308 19724 10364
rect 19724 10308 19780 10364
rect 19780 10308 19784 10364
rect 19720 10304 19784 10308
rect 5584 9820 5648 9824
rect 5584 9764 5588 9820
rect 5588 9764 5644 9820
rect 5644 9764 5648 9820
rect 5584 9760 5648 9764
rect 5664 9820 5728 9824
rect 5664 9764 5668 9820
rect 5668 9764 5724 9820
rect 5724 9764 5728 9820
rect 5664 9760 5728 9764
rect 5744 9820 5808 9824
rect 5744 9764 5748 9820
rect 5748 9764 5804 9820
rect 5804 9764 5808 9820
rect 5744 9760 5808 9764
rect 5824 9820 5888 9824
rect 5824 9764 5828 9820
rect 5828 9764 5884 9820
rect 5884 9764 5888 9820
rect 5824 9760 5888 9764
rect 14848 9820 14912 9824
rect 14848 9764 14852 9820
rect 14852 9764 14908 9820
rect 14908 9764 14912 9820
rect 14848 9760 14912 9764
rect 14928 9820 14992 9824
rect 14928 9764 14932 9820
rect 14932 9764 14988 9820
rect 14988 9764 14992 9820
rect 14928 9760 14992 9764
rect 15008 9820 15072 9824
rect 15008 9764 15012 9820
rect 15012 9764 15068 9820
rect 15068 9764 15072 9820
rect 15008 9760 15072 9764
rect 15088 9820 15152 9824
rect 15088 9764 15092 9820
rect 15092 9764 15148 9820
rect 15148 9764 15152 9820
rect 15088 9760 15152 9764
rect 24112 9820 24176 9824
rect 24112 9764 24116 9820
rect 24116 9764 24172 9820
rect 24172 9764 24176 9820
rect 24112 9760 24176 9764
rect 24192 9820 24256 9824
rect 24192 9764 24196 9820
rect 24196 9764 24252 9820
rect 24252 9764 24256 9820
rect 24192 9760 24256 9764
rect 24272 9820 24336 9824
rect 24272 9764 24276 9820
rect 24276 9764 24332 9820
rect 24332 9764 24336 9820
rect 24272 9760 24336 9764
rect 24352 9820 24416 9824
rect 24352 9764 24356 9820
rect 24356 9764 24412 9820
rect 24412 9764 24416 9820
rect 24352 9760 24416 9764
rect 10216 9276 10280 9280
rect 10216 9220 10220 9276
rect 10220 9220 10276 9276
rect 10276 9220 10280 9276
rect 10216 9216 10280 9220
rect 10296 9276 10360 9280
rect 10296 9220 10300 9276
rect 10300 9220 10356 9276
rect 10356 9220 10360 9276
rect 10296 9216 10360 9220
rect 10376 9276 10440 9280
rect 10376 9220 10380 9276
rect 10380 9220 10436 9276
rect 10436 9220 10440 9276
rect 10376 9216 10440 9220
rect 10456 9276 10520 9280
rect 10456 9220 10460 9276
rect 10460 9220 10516 9276
rect 10516 9220 10520 9276
rect 10456 9216 10520 9220
rect 19480 9276 19544 9280
rect 19480 9220 19484 9276
rect 19484 9220 19540 9276
rect 19540 9220 19544 9276
rect 19480 9216 19544 9220
rect 19560 9276 19624 9280
rect 19560 9220 19564 9276
rect 19564 9220 19620 9276
rect 19620 9220 19624 9276
rect 19560 9216 19624 9220
rect 19640 9276 19704 9280
rect 19640 9220 19644 9276
rect 19644 9220 19700 9276
rect 19700 9220 19704 9276
rect 19640 9216 19704 9220
rect 19720 9276 19784 9280
rect 19720 9220 19724 9276
rect 19724 9220 19780 9276
rect 19780 9220 19784 9276
rect 19720 9216 19784 9220
rect 5584 8732 5648 8736
rect 5584 8676 5588 8732
rect 5588 8676 5644 8732
rect 5644 8676 5648 8732
rect 5584 8672 5648 8676
rect 5664 8732 5728 8736
rect 5664 8676 5668 8732
rect 5668 8676 5724 8732
rect 5724 8676 5728 8732
rect 5664 8672 5728 8676
rect 5744 8732 5808 8736
rect 5744 8676 5748 8732
rect 5748 8676 5804 8732
rect 5804 8676 5808 8732
rect 5744 8672 5808 8676
rect 5824 8732 5888 8736
rect 5824 8676 5828 8732
rect 5828 8676 5884 8732
rect 5884 8676 5888 8732
rect 5824 8672 5888 8676
rect 14848 8732 14912 8736
rect 14848 8676 14852 8732
rect 14852 8676 14908 8732
rect 14908 8676 14912 8732
rect 14848 8672 14912 8676
rect 14928 8732 14992 8736
rect 14928 8676 14932 8732
rect 14932 8676 14988 8732
rect 14988 8676 14992 8732
rect 14928 8672 14992 8676
rect 15008 8732 15072 8736
rect 15008 8676 15012 8732
rect 15012 8676 15068 8732
rect 15068 8676 15072 8732
rect 15008 8672 15072 8676
rect 15088 8732 15152 8736
rect 15088 8676 15092 8732
rect 15092 8676 15148 8732
rect 15148 8676 15152 8732
rect 15088 8672 15152 8676
rect 24112 8732 24176 8736
rect 24112 8676 24116 8732
rect 24116 8676 24172 8732
rect 24172 8676 24176 8732
rect 24112 8672 24176 8676
rect 24192 8732 24256 8736
rect 24192 8676 24196 8732
rect 24196 8676 24252 8732
rect 24252 8676 24256 8732
rect 24192 8672 24256 8676
rect 24272 8732 24336 8736
rect 24272 8676 24276 8732
rect 24276 8676 24332 8732
rect 24332 8676 24336 8732
rect 24272 8672 24336 8676
rect 24352 8732 24416 8736
rect 24352 8676 24356 8732
rect 24356 8676 24412 8732
rect 24412 8676 24416 8732
rect 24352 8672 24416 8676
rect 10216 8188 10280 8192
rect 10216 8132 10220 8188
rect 10220 8132 10276 8188
rect 10276 8132 10280 8188
rect 10216 8128 10280 8132
rect 10296 8188 10360 8192
rect 10296 8132 10300 8188
rect 10300 8132 10356 8188
rect 10356 8132 10360 8188
rect 10296 8128 10360 8132
rect 10376 8188 10440 8192
rect 10376 8132 10380 8188
rect 10380 8132 10436 8188
rect 10436 8132 10440 8188
rect 10376 8128 10440 8132
rect 10456 8188 10520 8192
rect 10456 8132 10460 8188
rect 10460 8132 10516 8188
rect 10516 8132 10520 8188
rect 10456 8128 10520 8132
rect 19480 8188 19544 8192
rect 19480 8132 19484 8188
rect 19484 8132 19540 8188
rect 19540 8132 19544 8188
rect 19480 8128 19544 8132
rect 19560 8188 19624 8192
rect 19560 8132 19564 8188
rect 19564 8132 19620 8188
rect 19620 8132 19624 8188
rect 19560 8128 19624 8132
rect 19640 8188 19704 8192
rect 19640 8132 19644 8188
rect 19644 8132 19700 8188
rect 19700 8132 19704 8188
rect 19640 8128 19704 8132
rect 19720 8188 19784 8192
rect 19720 8132 19724 8188
rect 19724 8132 19780 8188
rect 19780 8132 19784 8188
rect 19720 8128 19784 8132
rect 5584 7644 5648 7648
rect 5584 7588 5588 7644
rect 5588 7588 5644 7644
rect 5644 7588 5648 7644
rect 5584 7584 5648 7588
rect 5664 7644 5728 7648
rect 5664 7588 5668 7644
rect 5668 7588 5724 7644
rect 5724 7588 5728 7644
rect 5664 7584 5728 7588
rect 5744 7644 5808 7648
rect 5744 7588 5748 7644
rect 5748 7588 5804 7644
rect 5804 7588 5808 7644
rect 5744 7584 5808 7588
rect 5824 7644 5888 7648
rect 5824 7588 5828 7644
rect 5828 7588 5884 7644
rect 5884 7588 5888 7644
rect 5824 7584 5888 7588
rect 14848 7644 14912 7648
rect 14848 7588 14852 7644
rect 14852 7588 14908 7644
rect 14908 7588 14912 7644
rect 14848 7584 14912 7588
rect 14928 7644 14992 7648
rect 14928 7588 14932 7644
rect 14932 7588 14988 7644
rect 14988 7588 14992 7644
rect 14928 7584 14992 7588
rect 15008 7644 15072 7648
rect 15008 7588 15012 7644
rect 15012 7588 15068 7644
rect 15068 7588 15072 7644
rect 15008 7584 15072 7588
rect 15088 7644 15152 7648
rect 15088 7588 15092 7644
rect 15092 7588 15148 7644
rect 15148 7588 15152 7644
rect 15088 7584 15152 7588
rect 24112 7644 24176 7648
rect 24112 7588 24116 7644
rect 24116 7588 24172 7644
rect 24172 7588 24176 7644
rect 24112 7584 24176 7588
rect 24192 7644 24256 7648
rect 24192 7588 24196 7644
rect 24196 7588 24252 7644
rect 24252 7588 24256 7644
rect 24192 7584 24256 7588
rect 24272 7644 24336 7648
rect 24272 7588 24276 7644
rect 24276 7588 24332 7644
rect 24332 7588 24336 7644
rect 24272 7584 24336 7588
rect 24352 7644 24416 7648
rect 24352 7588 24356 7644
rect 24356 7588 24412 7644
rect 24412 7588 24416 7644
rect 24352 7584 24416 7588
rect 10216 7100 10280 7104
rect 10216 7044 10220 7100
rect 10220 7044 10276 7100
rect 10276 7044 10280 7100
rect 10216 7040 10280 7044
rect 10296 7100 10360 7104
rect 10296 7044 10300 7100
rect 10300 7044 10356 7100
rect 10356 7044 10360 7100
rect 10296 7040 10360 7044
rect 10376 7100 10440 7104
rect 10376 7044 10380 7100
rect 10380 7044 10436 7100
rect 10436 7044 10440 7100
rect 10376 7040 10440 7044
rect 10456 7100 10520 7104
rect 10456 7044 10460 7100
rect 10460 7044 10516 7100
rect 10516 7044 10520 7100
rect 10456 7040 10520 7044
rect 19480 7100 19544 7104
rect 19480 7044 19484 7100
rect 19484 7044 19540 7100
rect 19540 7044 19544 7100
rect 19480 7040 19544 7044
rect 19560 7100 19624 7104
rect 19560 7044 19564 7100
rect 19564 7044 19620 7100
rect 19620 7044 19624 7100
rect 19560 7040 19624 7044
rect 19640 7100 19704 7104
rect 19640 7044 19644 7100
rect 19644 7044 19700 7100
rect 19700 7044 19704 7100
rect 19640 7040 19704 7044
rect 19720 7100 19784 7104
rect 19720 7044 19724 7100
rect 19724 7044 19780 7100
rect 19780 7044 19784 7100
rect 19720 7040 19784 7044
rect 5584 6556 5648 6560
rect 5584 6500 5588 6556
rect 5588 6500 5644 6556
rect 5644 6500 5648 6556
rect 5584 6496 5648 6500
rect 5664 6556 5728 6560
rect 5664 6500 5668 6556
rect 5668 6500 5724 6556
rect 5724 6500 5728 6556
rect 5664 6496 5728 6500
rect 5744 6556 5808 6560
rect 5744 6500 5748 6556
rect 5748 6500 5804 6556
rect 5804 6500 5808 6556
rect 5744 6496 5808 6500
rect 5824 6556 5888 6560
rect 5824 6500 5828 6556
rect 5828 6500 5884 6556
rect 5884 6500 5888 6556
rect 5824 6496 5888 6500
rect 14848 6556 14912 6560
rect 14848 6500 14852 6556
rect 14852 6500 14908 6556
rect 14908 6500 14912 6556
rect 14848 6496 14912 6500
rect 14928 6556 14992 6560
rect 14928 6500 14932 6556
rect 14932 6500 14988 6556
rect 14988 6500 14992 6556
rect 14928 6496 14992 6500
rect 15008 6556 15072 6560
rect 15008 6500 15012 6556
rect 15012 6500 15068 6556
rect 15068 6500 15072 6556
rect 15008 6496 15072 6500
rect 15088 6556 15152 6560
rect 15088 6500 15092 6556
rect 15092 6500 15148 6556
rect 15148 6500 15152 6556
rect 15088 6496 15152 6500
rect 24112 6556 24176 6560
rect 24112 6500 24116 6556
rect 24116 6500 24172 6556
rect 24172 6500 24176 6556
rect 24112 6496 24176 6500
rect 24192 6556 24256 6560
rect 24192 6500 24196 6556
rect 24196 6500 24252 6556
rect 24252 6500 24256 6556
rect 24192 6496 24256 6500
rect 24272 6556 24336 6560
rect 24272 6500 24276 6556
rect 24276 6500 24332 6556
rect 24332 6500 24336 6556
rect 24272 6496 24336 6500
rect 24352 6556 24416 6560
rect 24352 6500 24356 6556
rect 24356 6500 24412 6556
rect 24412 6500 24416 6556
rect 24352 6496 24416 6500
rect 10216 6012 10280 6016
rect 10216 5956 10220 6012
rect 10220 5956 10276 6012
rect 10276 5956 10280 6012
rect 10216 5952 10280 5956
rect 10296 6012 10360 6016
rect 10296 5956 10300 6012
rect 10300 5956 10356 6012
rect 10356 5956 10360 6012
rect 10296 5952 10360 5956
rect 10376 6012 10440 6016
rect 10376 5956 10380 6012
rect 10380 5956 10436 6012
rect 10436 5956 10440 6012
rect 10376 5952 10440 5956
rect 10456 6012 10520 6016
rect 10456 5956 10460 6012
rect 10460 5956 10516 6012
rect 10516 5956 10520 6012
rect 10456 5952 10520 5956
rect 19480 6012 19544 6016
rect 19480 5956 19484 6012
rect 19484 5956 19540 6012
rect 19540 5956 19544 6012
rect 19480 5952 19544 5956
rect 19560 6012 19624 6016
rect 19560 5956 19564 6012
rect 19564 5956 19620 6012
rect 19620 5956 19624 6012
rect 19560 5952 19624 5956
rect 19640 6012 19704 6016
rect 19640 5956 19644 6012
rect 19644 5956 19700 6012
rect 19700 5956 19704 6012
rect 19640 5952 19704 5956
rect 19720 6012 19784 6016
rect 19720 5956 19724 6012
rect 19724 5956 19780 6012
rect 19780 5956 19784 6012
rect 19720 5952 19784 5956
rect 5584 5468 5648 5472
rect 5584 5412 5588 5468
rect 5588 5412 5644 5468
rect 5644 5412 5648 5468
rect 5584 5408 5648 5412
rect 5664 5468 5728 5472
rect 5664 5412 5668 5468
rect 5668 5412 5724 5468
rect 5724 5412 5728 5468
rect 5664 5408 5728 5412
rect 5744 5468 5808 5472
rect 5744 5412 5748 5468
rect 5748 5412 5804 5468
rect 5804 5412 5808 5468
rect 5744 5408 5808 5412
rect 5824 5468 5888 5472
rect 5824 5412 5828 5468
rect 5828 5412 5884 5468
rect 5884 5412 5888 5468
rect 5824 5408 5888 5412
rect 14848 5468 14912 5472
rect 14848 5412 14852 5468
rect 14852 5412 14908 5468
rect 14908 5412 14912 5468
rect 14848 5408 14912 5412
rect 14928 5468 14992 5472
rect 14928 5412 14932 5468
rect 14932 5412 14988 5468
rect 14988 5412 14992 5468
rect 14928 5408 14992 5412
rect 15008 5468 15072 5472
rect 15008 5412 15012 5468
rect 15012 5412 15068 5468
rect 15068 5412 15072 5468
rect 15008 5408 15072 5412
rect 15088 5468 15152 5472
rect 15088 5412 15092 5468
rect 15092 5412 15148 5468
rect 15148 5412 15152 5468
rect 15088 5408 15152 5412
rect 24112 5468 24176 5472
rect 24112 5412 24116 5468
rect 24116 5412 24172 5468
rect 24172 5412 24176 5468
rect 24112 5408 24176 5412
rect 24192 5468 24256 5472
rect 24192 5412 24196 5468
rect 24196 5412 24252 5468
rect 24252 5412 24256 5468
rect 24192 5408 24256 5412
rect 24272 5468 24336 5472
rect 24272 5412 24276 5468
rect 24276 5412 24332 5468
rect 24332 5412 24336 5468
rect 24272 5408 24336 5412
rect 24352 5468 24416 5472
rect 24352 5412 24356 5468
rect 24356 5412 24412 5468
rect 24412 5412 24416 5468
rect 24352 5408 24416 5412
rect 10216 4924 10280 4928
rect 10216 4868 10220 4924
rect 10220 4868 10276 4924
rect 10276 4868 10280 4924
rect 10216 4864 10280 4868
rect 10296 4924 10360 4928
rect 10296 4868 10300 4924
rect 10300 4868 10356 4924
rect 10356 4868 10360 4924
rect 10296 4864 10360 4868
rect 10376 4924 10440 4928
rect 10376 4868 10380 4924
rect 10380 4868 10436 4924
rect 10436 4868 10440 4924
rect 10376 4864 10440 4868
rect 10456 4924 10520 4928
rect 10456 4868 10460 4924
rect 10460 4868 10516 4924
rect 10516 4868 10520 4924
rect 10456 4864 10520 4868
rect 19480 4924 19544 4928
rect 19480 4868 19484 4924
rect 19484 4868 19540 4924
rect 19540 4868 19544 4924
rect 19480 4864 19544 4868
rect 19560 4924 19624 4928
rect 19560 4868 19564 4924
rect 19564 4868 19620 4924
rect 19620 4868 19624 4924
rect 19560 4864 19624 4868
rect 19640 4924 19704 4928
rect 19640 4868 19644 4924
rect 19644 4868 19700 4924
rect 19700 4868 19704 4924
rect 19640 4864 19704 4868
rect 19720 4924 19784 4928
rect 19720 4868 19724 4924
rect 19724 4868 19780 4924
rect 19780 4868 19784 4924
rect 19720 4864 19784 4868
rect 5584 4380 5648 4384
rect 5584 4324 5588 4380
rect 5588 4324 5644 4380
rect 5644 4324 5648 4380
rect 5584 4320 5648 4324
rect 5664 4380 5728 4384
rect 5664 4324 5668 4380
rect 5668 4324 5724 4380
rect 5724 4324 5728 4380
rect 5664 4320 5728 4324
rect 5744 4380 5808 4384
rect 5744 4324 5748 4380
rect 5748 4324 5804 4380
rect 5804 4324 5808 4380
rect 5744 4320 5808 4324
rect 5824 4380 5888 4384
rect 5824 4324 5828 4380
rect 5828 4324 5884 4380
rect 5884 4324 5888 4380
rect 5824 4320 5888 4324
rect 14848 4380 14912 4384
rect 14848 4324 14852 4380
rect 14852 4324 14908 4380
rect 14908 4324 14912 4380
rect 14848 4320 14912 4324
rect 14928 4380 14992 4384
rect 14928 4324 14932 4380
rect 14932 4324 14988 4380
rect 14988 4324 14992 4380
rect 14928 4320 14992 4324
rect 15008 4380 15072 4384
rect 15008 4324 15012 4380
rect 15012 4324 15068 4380
rect 15068 4324 15072 4380
rect 15008 4320 15072 4324
rect 15088 4380 15152 4384
rect 15088 4324 15092 4380
rect 15092 4324 15148 4380
rect 15148 4324 15152 4380
rect 15088 4320 15152 4324
rect 24112 4380 24176 4384
rect 24112 4324 24116 4380
rect 24116 4324 24172 4380
rect 24172 4324 24176 4380
rect 24112 4320 24176 4324
rect 24192 4380 24256 4384
rect 24192 4324 24196 4380
rect 24196 4324 24252 4380
rect 24252 4324 24256 4380
rect 24192 4320 24256 4324
rect 24272 4380 24336 4384
rect 24272 4324 24276 4380
rect 24276 4324 24332 4380
rect 24332 4324 24336 4380
rect 24272 4320 24336 4324
rect 24352 4380 24416 4384
rect 24352 4324 24356 4380
rect 24356 4324 24412 4380
rect 24412 4324 24416 4380
rect 24352 4320 24416 4324
rect 10216 3836 10280 3840
rect 10216 3780 10220 3836
rect 10220 3780 10276 3836
rect 10276 3780 10280 3836
rect 10216 3776 10280 3780
rect 10296 3836 10360 3840
rect 10296 3780 10300 3836
rect 10300 3780 10356 3836
rect 10356 3780 10360 3836
rect 10296 3776 10360 3780
rect 10376 3836 10440 3840
rect 10376 3780 10380 3836
rect 10380 3780 10436 3836
rect 10436 3780 10440 3836
rect 10376 3776 10440 3780
rect 10456 3836 10520 3840
rect 10456 3780 10460 3836
rect 10460 3780 10516 3836
rect 10516 3780 10520 3836
rect 10456 3776 10520 3780
rect 19480 3836 19544 3840
rect 19480 3780 19484 3836
rect 19484 3780 19540 3836
rect 19540 3780 19544 3836
rect 19480 3776 19544 3780
rect 19560 3836 19624 3840
rect 19560 3780 19564 3836
rect 19564 3780 19620 3836
rect 19620 3780 19624 3836
rect 19560 3776 19624 3780
rect 19640 3836 19704 3840
rect 19640 3780 19644 3836
rect 19644 3780 19700 3836
rect 19700 3780 19704 3836
rect 19640 3776 19704 3780
rect 19720 3836 19784 3840
rect 19720 3780 19724 3836
rect 19724 3780 19780 3836
rect 19780 3780 19784 3836
rect 19720 3776 19784 3780
rect 5584 3292 5648 3296
rect 5584 3236 5588 3292
rect 5588 3236 5644 3292
rect 5644 3236 5648 3292
rect 5584 3232 5648 3236
rect 5664 3292 5728 3296
rect 5664 3236 5668 3292
rect 5668 3236 5724 3292
rect 5724 3236 5728 3292
rect 5664 3232 5728 3236
rect 5744 3292 5808 3296
rect 5744 3236 5748 3292
rect 5748 3236 5804 3292
rect 5804 3236 5808 3292
rect 5744 3232 5808 3236
rect 5824 3292 5888 3296
rect 5824 3236 5828 3292
rect 5828 3236 5884 3292
rect 5884 3236 5888 3292
rect 5824 3232 5888 3236
rect 14848 3292 14912 3296
rect 14848 3236 14852 3292
rect 14852 3236 14908 3292
rect 14908 3236 14912 3292
rect 14848 3232 14912 3236
rect 14928 3292 14992 3296
rect 14928 3236 14932 3292
rect 14932 3236 14988 3292
rect 14988 3236 14992 3292
rect 14928 3232 14992 3236
rect 15008 3292 15072 3296
rect 15008 3236 15012 3292
rect 15012 3236 15068 3292
rect 15068 3236 15072 3292
rect 15008 3232 15072 3236
rect 15088 3292 15152 3296
rect 15088 3236 15092 3292
rect 15092 3236 15148 3292
rect 15148 3236 15152 3292
rect 15088 3232 15152 3236
rect 24112 3292 24176 3296
rect 24112 3236 24116 3292
rect 24116 3236 24172 3292
rect 24172 3236 24176 3292
rect 24112 3232 24176 3236
rect 24192 3292 24256 3296
rect 24192 3236 24196 3292
rect 24196 3236 24252 3292
rect 24252 3236 24256 3292
rect 24192 3232 24256 3236
rect 24272 3292 24336 3296
rect 24272 3236 24276 3292
rect 24276 3236 24332 3292
rect 24332 3236 24336 3292
rect 24272 3232 24336 3236
rect 24352 3292 24416 3296
rect 24352 3236 24356 3292
rect 24356 3236 24412 3292
rect 24412 3236 24416 3292
rect 24352 3232 24416 3236
rect 10216 2748 10280 2752
rect 10216 2692 10220 2748
rect 10220 2692 10276 2748
rect 10276 2692 10280 2748
rect 10216 2688 10280 2692
rect 10296 2748 10360 2752
rect 10296 2692 10300 2748
rect 10300 2692 10356 2748
rect 10356 2692 10360 2748
rect 10296 2688 10360 2692
rect 10376 2748 10440 2752
rect 10376 2692 10380 2748
rect 10380 2692 10436 2748
rect 10436 2692 10440 2748
rect 10376 2688 10440 2692
rect 10456 2748 10520 2752
rect 10456 2692 10460 2748
rect 10460 2692 10516 2748
rect 10516 2692 10520 2748
rect 10456 2688 10520 2692
rect 19480 2748 19544 2752
rect 19480 2692 19484 2748
rect 19484 2692 19540 2748
rect 19540 2692 19544 2748
rect 19480 2688 19544 2692
rect 19560 2748 19624 2752
rect 19560 2692 19564 2748
rect 19564 2692 19620 2748
rect 19620 2692 19624 2748
rect 19560 2688 19624 2692
rect 19640 2748 19704 2752
rect 19640 2692 19644 2748
rect 19644 2692 19700 2748
rect 19700 2692 19704 2748
rect 19640 2688 19704 2692
rect 19720 2748 19784 2752
rect 19720 2692 19724 2748
rect 19724 2692 19780 2748
rect 19780 2692 19784 2748
rect 19720 2688 19784 2692
rect 5584 2204 5648 2208
rect 5584 2148 5588 2204
rect 5588 2148 5644 2204
rect 5644 2148 5648 2204
rect 5584 2144 5648 2148
rect 5664 2204 5728 2208
rect 5664 2148 5668 2204
rect 5668 2148 5724 2204
rect 5724 2148 5728 2204
rect 5664 2144 5728 2148
rect 5744 2204 5808 2208
rect 5744 2148 5748 2204
rect 5748 2148 5804 2204
rect 5804 2148 5808 2204
rect 5744 2144 5808 2148
rect 5824 2204 5888 2208
rect 5824 2148 5828 2204
rect 5828 2148 5884 2204
rect 5884 2148 5888 2204
rect 5824 2144 5888 2148
rect 14848 2204 14912 2208
rect 14848 2148 14852 2204
rect 14852 2148 14908 2204
rect 14908 2148 14912 2204
rect 14848 2144 14912 2148
rect 14928 2204 14992 2208
rect 14928 2148 14932 2204
rect 14932 2148 14988 2204
rect 14988 2148 14992 2204
rect 14928 2144 14992 2148
rect 15008 2204 15072 2208
rect 15008 2148 15012 2204
rect 15012 2148 15068 2204
rect 15068 2148 15072 2204
rect 15008 2144 15072 2148
rect 15088 2204 15152 2208
rect 15088 2148 15092 2204
rect 15092 2148 15148 2204
rect 15148 2148 15152 2204
rect 15088 2144 15152 2148
rect 24112 2204 24176 2208
rect 24112 2148 24116 2204
rect 24116 2148 24172 2204
rect 24172 2148 24176 2204
rect 24112 2144 24176 2148
rect 24192 2204 24256 2208
rect 24192 2148 24196 2204
rect 24196 2148 24252 2204
rect 24252 2148 24256 2204
rect 24192 2144 24256 2148
rect 24272 2204 24336 2208
rect 24272 2148 24276 2204
rect 24276 2148 24332 2204
rect 24332 2148 24336 2204
rect 24272 2144 24336 2148
rect 24352 2204 24416 2208
rect 24352 2148 24356 2204
rect 24356 2148 24412 2204
rect 24412 2148 24416 2204
rect 24352 2144 24416 2148
<< metal4 >>
rect 5576 53344 5896 53360
rect 5576 53280 5584 53344
rect 5648 53280 5664 53344
rect 5728 53280 5744 53344
rect 5808 53280 5824 53344
rect 5888 53280 5896 53344
rect 5576 52256 5896 53280
rect 5576 52192 5584 52256
rect 5648 52192 5664 52256
rect 5728 52192 5744 52256
rect 5808 52192 5824 52256
rect 5888 52192 5896 52256
rect 5576 51168 5896 52192
rect 5576 51104 5584 51168
rect 5648 51104 5664 51168
rect 5728 51104 5744 51168
rect 5808 51104 5824 51168
rect 5888 51104 5896 51168
rect 5576 50080 5896 51104
rect 5576 50016 5584 50080
rect 5648 50016 5664 50080
rect 5728 50016 5744 50080
rect 5808 50016 5824 50080
rect 5888 50016 5896 50080
rect 5576 48992 5896 50016
rect 5576 48928 5584 48992
rect 5648 48928 5664 48992
rect 5728 48928 5744 48992
rect 5808 48928 5824 48992
rect 5888 48928 5896 48992
rect 5576 47904 5896 48928
rect 5576 47840 5584 47904
rect 5648 47840 5664 47904
rect 5728 47840 5744 47904
rect 5808 47840 5824 47904
rect 5888 47840 5896 47904
rect 5576 46816 5896 47840
rect 5576 46752 5584 46816
rect 5648 46752 5664 46816
rect 5728 46752 5744 46816
rect 5808 46752 5824 46816
rect 5888 46752 5896 46816
rect 5576 45728 5896 46752
rect 5576 45664 5584 45728
rect 5648 45664 5664 45728
rect 5728 45664 5744 45728
rect 5808 45664 5824 45728
rect 5888 45664 5896 45728
rect 5576 44640 5896 45664
rect 5576 44576 5584 44640
rect 5648 44576 5664 44640
rect 5728 44576 5744 44640
rect 5808 44576 5824 44640
rect 5888 44576 5896 44640
rect 5576 43552 5896 44576
rect 5576 43488 5584 43552
rect 5648 43488 5664 43552
rect 5728 43488 5744 43552
rect 5808 43488 5824 43552
rect 5888 43488 5896 43552
rect 5576 42464 5896 43488
rect 5576 42400 5584 42464
rect 5648 42400 5664 42464
rect 5728 42400 5744 42464
rect 5808 42400 5824 42464
rect 5888 42400 5896 42464
rect 5576 41376 5896 42400
rect 5576 41312 5584 41376
rect 5648 41312 5664 41376
rect 5728 41312 5744 41376
rect 5808 41312 5824 41376
rect 5888 41312 5896 41376
rect 5576 40288 5896 41312
rect 5576 40224 5584 40288
rect 5648 40224 5664 40288
rect 5728 40224 5744 40288
rect 5808 40224 5824 40288
rect 5888 40224 5896 40288
rect 5576 39200 5896 40224
rect 5576 39136 5584 39200
rect 5648 39136 5664 39200
rect 5728 39136 5744 39200
rect 5808 39136 5824 39200
rect 5888 39136 5896 39200
rect 5576 38112 5896 39136
rect 5576 38048 5584 38112
rect 5648 38048 5664 38112
rect 5728 38048 5744 38112
rect 5808 38048 5824 38112
rect 5888 38048 5896 38112
rect 5576 37024 5896 38048
rect 5576 36960 5584 37024
rect 5648 36960 5664 37024
rect 5728 36960 5744 37024
rect 5808 36960 5824 37024
rect 5888 36960 5896 37024
rect 5576 35936 5896 36960
rect 5576 35872 5584 35936
rect 5648 35872 5664 35936
rect 5728 35872 5744 35936
rect 5808 35872 5824 35936
rect 5888 35872 5896 35936
rect 5576 34848 5896 35872
rect 5576 34784 5584 34848
rect 5648 34784 5664 34848
rect 5728 34784 5744 34848
rect 5808 34784 5824 34848
rect 5888 34784 5896 34848
rect 5576 33760 5896 34784
rect 5576 33696 5584 33760
rect 5648 33696 5664 33760
rect 5728 33696 5744 33760
rect 5808 33696 5824 33760
rect 5888 33696 5896 33760
rect 5576 32672 5896 33696
rect 5576 32608 5584 32672
rect 5648 32608 5664 32672
rect 5728 32608 5744 32672
rect 5808 32608 5824 32672
rect 5888 32608 5896 32672
rect 5576 31584 5896 32608
rect 5576 31520 5584 31584
rect 5648 31520 5664 31584
rect 5728 31520 5744 31584
rect 5808 31520 5824 31584
rect 5888 31520 5896 31584
rect 5576 30496 5896 31520
rect 5576 30432 5584 30496
rect 5648 30432 5664 30496
rect 5728 30432 5744 30496
rect 5808 30432 5824 30496
rect 5888 30432 5896 30496
rect 5576 29408 5896 30432
rect 5576 29344 5584 29408
rect 5648 29344 5664 29408
rect 5728 29344 5744 29408
rect 5808 29344 5824 29408
rect 5888 29344 5896 29408
rect 5576 28320 5896 29344
rect 5576 28256 5584 28320
rect 5648 28256 5664 28320
rect 5728 28256 5744 28320
rect 5808 28256 5824 28320
rect 5888 28256 5896 28320
rect 5576 27232 5896 28256
rect 5576 27168 5584 27232
rect 5648 27168 5664 27232
rect 5728 27168 5744 27232
rect 5808 27168 5824 27232
rect 5888 27168 5896 27232
rect 5576 26144 5896 27168
rect 5576 26080 5584 26144
rect 5648 26080 5664 26144
rect 5728 26080 5744 26144
rect 5808 26080 5824 26144
rect 5888 26080 5896 26144
rect 5576 25056 5896 26080
rect 5576 24992 5584 25056
rect 5648 24992 5664 25056
rect 5728 24992 5744 25056
rect 5808 24992 5824 25056
rect 5888 24992 5896 25056
rect 5576 23968 5896 24992
rect 5576 23904 5584 23968
rect 5648 23904 5664 23968
rect 5728 23904 5744 23968
rect 5808 23904 5824 23968
rect 5888 23904 5896 23968
rect 5576 22880 5896 23904
rect 5576 22816 5584 22880
rect 5648 22816 5664 22880
rect 5728 22816 5744 22880
rect 5808 22816 5824 22880
rect 5888 22816 5896 22880
rect 5576 21792 5896 22816
rect 5576 21728 5584 21792
rect 5648 21728 5664 21792
rect 5728 21728 5744 21792
rect 5808 21728 5824 21792
rect 5888 21728 5896 21792
rect 5576 20704 5896 21728
rect 5576 20640 5584 20704
rect 5648 20640 5664 20704
rect 5728 20640 5744 20704
rect 5808 20640 5824 20704
rect 5888 20640 5896 20704
rect 5576 19616 5896 20640
rect 5576 19552 5584 19616
rect 5648 19552 5664 19616
rect 5728 19552 5744 19616
rect 5808 19552 5824 19616
rect 5888 19552 5896 19616
rect 5576 18528 5896 19552
rect 5576 18464 5584 18528
rect 5648 18464 5664 18528
rect 5728 18464 5744 18528
rect 5808 18464 5824 18528
rect 5888 18464 5896 18528
rect 5576 17440 5896 18464
rect 5576 17376 5584 17440
rect 5648 17376 5664 17440
rect 5728 17376 5744 17440
rect 5808 17376 5824 17440
rect 5888 17376 5896 17440
rect 5576 16352 5896 17376
rect 5576 16288 5584 16352
rect 5648 16288 5664 16352
rect 5728 16288 5744 16352
rect 5808 16288 5824 16352
rect 5888 16288 5896 16352
rect 5576 15264 5896 16288
rect 5576 15200 5584 15264
rect 5648 15200 5664 15264
rect 5728 15200 5744 15264
rect 5808 15200 5824 15264
rect 5888 15200 5896 15264
rect 5576 14176 5896 15200
rect 5576 14112 5584 14176
rect 5648 14112 5664 14176
rect 5728 14112 5744 14176
rect 5808 14112 5824 14176
rect 5888 14112 5896 14176
rect 5576 13088 5896 14112
rect 5576 13024 5584 13088
rect 5648 13024 5664 13088
rect 5728 13024 5744 13088
rect 5808 13024 5824 13088
rect 5888 13024 5896 13088
rect 5576 12000 5896 13024
rect 5576 11936 5584 12000
rect 5648 11936 5664 12000
rect 5728 11936 5744 12000
rect 5808 11936 5824 12000
rect 5888 11936 5896 12000
rect 5576 10912 5896 11936
rect 5576 10848 5584 10912
rect 5648 10848 5664 10912
rect 5728 10848 5744 10912
rect 5808 10848 5824 10912
rect 5888 10848 5896 10912
rect 5576 9824 5896 10848
rect 5576 9760 5584 9824
rect 5648 9760 5664 9824
rect 5728 9760 5744 9824
rect 5808 9760 5824 9824
rect 5888 9760 5896 9824
rect 5576 8736 5896 9760
rect 5576 8672 5584 8736
rect 5648 8672 5664 8736
rect 5728 8672 5744 8736
rect 5808 8672 5824 8736
rect 5888 8672 5896 8736
rect 5576 7648 5896 8672
rect 5576 7584 5584 7648
rect 5648 7584 5664 7648
rect 5728 7584 5744 7648
rect 5808 7584 5824 7648
rect 5888 7584 5896 7648
rect 5576 6560 5896 7584
rect 5576 6496 5584 6560
rect 5648 6496 5664 6560
rect 5728 6496 5744 6560
rect 5808 6496 5824 6560
rect 5888 6496 5896 6560
rect 5576 5472 5896 6496
rect 5576 5408 5584 5472
rect 5648 5408 5664 5472
rect 5728 5408 5744 5472
rect 5808 5408 5824 5472
rect 5888 5408 5896 5472
rect 5576 4384 5896 5408
rect 5576 4320 5584 4384
rect 5648 4320 5664 4384
rect 5728 4320 5744 4384
rect 5808 4320 5824 4384
rect 5888 4320 5896 4384
rect 5576 3296 5896 4320
rect 5576 3232 5584 3296
rect 5648 3232 5664 3296
rect 5728 3232 5744 3296
rect 5808 3232 5824 3296
rect 5888 3232 5896 3296
rect 5576 2208 5896 3232
rect 5576 2144 5584 2208
rect 5648 2144 5664 2208
rect 5728 2144 5744 2208
rect 5808 2144 5824 2208
rect 5888 2144 5896 2208
rect 5576 2128 5896 2144
rect 10208 52800 10528 53360
rect 10208 52736 10216 52800
rect 10280 52736 10296 52800
rect 10360 52736 10376 52800
rect 10440 52736 10456 52800
rect 10520 52736 10528 52800
rect 10208 51712 10528 52736
rect 10208 51648 10216 51712
rect 10280 51648 10296 51712
rect 10360 51648 10376 51712
rect 10440 51648 10456 51712
rect 10520 51648 10528 51712
rect 10208 50624 10528 51648
rect 10208 50560 10216 50624
rect 10280 50560 10296 50624
rect 10360 50560 10376 50624
rect 10440 50560 10456 50624
rect 10520 50560 10528 50624
rect 10208 49536 10528 50560
rect 10208 49472 10216 49536
rect 10280 49472 10296 49536
rect 10360 49472 10376 49536
rect 10440 49472 10456 49536
rect 10520 49472 10528 49536
rect 10208 48448 10528 49472
rect 10208 48384 10216 48448
rect 10280 48384 10296 48448
rect 10360 48384 10376 48448
rect 10440 48384 10456 48448
rect 10520 48384 10528 48448
rect 10208 47360 10528 48384
rect 10208 47296 10216 47360
rect 10280 47296 10296 47360
rect 10360 47296 10376 47360
rect 10440 47296 10456 47360
rect 10520 47296 10528 47360
rect 10208 46272 10528 47296
rect 10208 46208 10216 46272
rect 10280 46208 10296 46272
rect 10360 46208 10376 46272
rect 10440 46208 10456 46272
rect 10520 46208 10528 46272
rect 10208 45184 10528 46208
rect 10208 45120 10216 45184
rect 10280 45120 10296 45184
rect 10360 45120 10376 45184
rect 10440 45120 10456 45184
rect 10520 45120 10528 45184
rect 10208 44096 10528 45120
rect 10208 44032 10216 44096
rect 10280 44032 10296 44096
rect 10360 44032 10376 44096
rect 10440 44032 10456 44096
rect 10520 44032 10528 44096
rect 10208 43008 10528 44032
rect 10208 42944 10216 43008
rect 10280 42944 10296 43008
rect 10360 42944 10376 43008
rect 10440 42944 10456 43008
rect 10520 42944 10528 43008
rect 10208 41920 10528 42944
rect 10208 41856 10216 41920
rect 10280 41856 10296 41920
rect 10360 41856 10376 41920
rect 10440 41856 10456 41920
rect 10520 41856 10528 41920
rect 10208 40832 10528 41856
rect 10208 40768 10216 40832
rect 10280 40768 10296 40832
rect 10360 40768 10376 40832
rect 10440 40768 10456 40832
rect 10520 40768 10528 40832
rect 10208 39744 10528 40768
rect 10208 39680 10216 39744
rect 10280 39680 10296 39744
rect 10360 39680 10376 39744
rect 10440 39680 10456 39744
rect 10520 39680 10528 39744
rect 10208 38656 10528 39680
rect 10208 38592 10216 38656
rect 10280 38592 10296 38656
rect 10360 38592 10376 38656
rect 10440 38592 10456 38656
rect 10520 38592 10528 38656
rect 10208 37568 10528 38592
rect 10208 37504 10216 37568
rect 10280 37504 10296 37568
rect 10360 37504 10376 37568
rect 10440 37504 10456 37568
rect 10520 37504 10528 37568
rect 10208 36480 10528 37504
rect 10208 36416 10216 36480
rect 10280 36416 10296 36480
rect 10360 36416 10376 36480
rect 10440 36416 10456 36480
rect 10520 36416 10528 36480
rect 10208 35392 10528 36416
rect 10208 35328 10216 35392
rect 10280 35328 10296 35392
rect 10360 35328 10376 35392
rect 10440 35328 10456 35392
rect 10520 35328 10528 35392
rect 10208 34304 10528 35328
rect 10208 34240 10216 34304
rect 10280 34240 10296 34304
rect 10360 34240 10376 34304
rect 10440 34240 10456 34304
rect 10520 34240 10528 34304
rect 10208 33216 10528 34240
rect 10208 33152 10216 33216
rect 10280 33152 10296 33216
rect 10360 33152 10376 33216
rect 10440 33152 10456 33216
rect 10520 33152 10528 33216
rect 10208 32128 10528 33152
rect 10208 32064 10216 32128
rect 10280 32064 10296 32128
rect 10360 32064 10376 32128
rect 10440 32064 10456 32128
rect 10520 32064 10528 32128
rect 10208 31040 10528 32064
rect 10208 30976 10216 31040
rect 10280 30976 10296 31040
rect 10360 30976 10376 31040
rect 10440 30976 10456 31040
rect 10520 30976 10528 31040
rect 10208 29952 10528 30976
rect 10208 29888 10216 29952
rect 10280 29888 10296 29952
rect 10360 29888 10376 29952
rect 10440 29888 10456 29952
rect 10520 29888 10528 29952
rect 10208 28864 10528 29888
rect 10208 28800 10216 28864
rect 10280 28800 10296 28864
rect 10360 28800 10376 28864
rect 10440 28800 10456 28864
rect 10520 28800 10528 28864
rect 10208 27776 10528 28800
rect 10208 27712 10216 27776
rect 10280 27712 10296 27776
rect 10360 27712 10376 27776
rect 10440 27712 10456 27776
rect 10520 27712 10528 27776
rect 10208 26688 10528 27712
rect 10208 26624 10216 26688
rect 10280 26624 10296 26688
rect 10360 26624 10376 26688
rect 10440 26624 10456 26688
rect 10520 26624 10528 26688
rect 10208 25600 10528 26624
rect 10208 25536 10216 25600
rect 10280 25536 10296 25600
rect 10360 25536 10376 25600
rect 10440 25536 10456 25600
rect 10520 25536 10528 25600
rect 10208 24512 10528 25536
rect 10208 24448 10216 24512
rect 10280 24448 10296 24512
rect 10360 24448 10376 24512
rect 10440 24448 10456 24512
rect 10520 24448 10528 24512
rect 10208 23424 10528 24448
rect 10208 23360 10216 23424
rect 10280 23360 10296 23424
rect 10360 23360 10376 23424
rect 10440 23360 10456 23424
rect 10520 23360 10528 23424
rect 10208 22336 10528 23360
rect 10208 22272 10216 22336
rect 10280 22272 10296 22336
rect 10360 22272 10376 22336
rect 10440 22272 10456 22336
rect 10520 22272 10528 22336
rect 10208 21248 10528 22272
rect 10208 21184 10216 21248
rect 10280 21184 10296 21248
rect 10360 21184 10376 21248
rect 10440 21184 10456 21248
rect 10520 21184 10528 21248
rect 10208 20160 10528 21184
rect 10208 20096 10216 20160
rect 10280 20096 10296 20160
rect 10360 20096 10376 20160
rect 10440 20096 10456 20160
rect 10520 20096 10528 20160
rect 10208 19072 10528 20096
rect 10208 19008 10216 19072
rect 10280 19008 10296 19072
rect 10360 19008 10376 19072
rect 10440 19008 10456 19072
rect 10520 19008 10528 19072
rect 10208 17984 10528 19008
rect 10208 17920 10216 17984
rect 10280 17920 10296 17984
rect 10360 17920 10376 17984
rect 10440 17920 10456 17984
rect 10520 17920 10528 17984
rect 10208 16896 10528 17920
rect 10208 16832 10216 16896
rect 10280 16832 10296 16896
rect 10360 16832 10376 16896
rect 10440 16832 10456 16896
rect 10520 16832 10528 16896
rect 10208 15808 10528 16832
rect 10208 15744 10216 15808
rect 10280 15744 10296 15808
rect 10360 15744 10376 15808
rect 10440 15744 10456 15808
rect 10520 15744 10528 15808
rect 10208 14720 10528 15744
rect 10208 14656 10216 14720
rect 10280 14656 10296 14720
rect 10360 14656 10376 14720
rect 10440 14656 10456 14720
rect 10520 14656 10528 14720
rect 10208 13632 10528 14656
rect 10208 13568 10216 13632
rect 10280 13568 10296 13632
rect 10360 13568 10376 13632
rect 10440 13568 10456 13632
rect 10520 13568 10528 13632
rect 10208 12544 10528 13568
rect 10208 12480 10216 12544
rect 10280 12480 10296 12544
rect 10360 12480 10376 12544
rect 10440 12480 10456 12544
rect 10520 12480 10528 12544
rect 10208 11456 10528 12480
rect 10208 11392 10216 11456
rect 10280 11392 10296 11456
rect 10360 11392 10376 11456
rect 10440 11392 10456 11456
rect 10520 11392 10528 11456
rect 10208 10368 10528 11392
rect 10208 10304 10216 10368
rect 10280 10304 10296 10368
rect 10360 10304 10376 10368
rect 10440 10304 10456 10368
rect 10520 10304 10528 10368
rect 10208 9280 10528 10304
rect 10208 9216 10216 9280
rect 10280 9216 10296 9280
rect 10360 9216 10376 9280
rect 10440 9216 10456 9280
rect 10520 9216 10528 9280
rect 10208 8192 10528 9216
rect 10208 8128 10216 8192
rect 10280 8128 10296 8192
rect 10360 8128 10376 8192
rect 10440 8128 10456 8192
rect 10520 8128 10528 8192
rect 10208 7104 10528 8128
rect 10208 7040 10216 7104
rect 10280 7040 10296 7104
rect 10360 7040 10376 7104
rect 10440 7040 10456 7104
rect 10520 7040 10528 7104
rect 10208 6016 10528 7040
rect 10208 5952 10216 6016
rect 10280 5952 10296 6016
rect 10360 5952 10376 6016
rect 10440 5952 10456 6016
rect 10520 5952 10528 6016
rect 10208 4928 10528 5952
rect 10208 4864 10216 4928
rect 10280 4864 10296 4928
rect 10360 4864 10376 4928
rect 10440 4864 10456 4928
rect 10520 4864 10528 4928
rect 10208 3840 10528 4864
rect 10208 3776 10216 3840
rect 10280 3776 10296 3840
rect 10360 3776 10376 3840
rect 10440 3776 10456 3840
rect 10520 3776 10528 3840
rect 10208 2752 10528 3776
rect 10208 2688 10216 2752
rect 10280 2688 10296 2752
rect 10360 2688 10376 2752
rect 10440 2688 10456 2752
rect 10520 2688 10528 2752
rect 10208 2128 10528 2688
rect 14840 53344 15160 53360
rect 14840 53280 14848 53344
rect 14912 53280 14928 53344
rect 14992 53280 15008 53344
rect 15072 53280 15088 53344
rect 15152 53280 15160 53344
rect 14840 52256 15160 53280
rect 14840 52192 14848 52256
rect 14912 52192 14928 52256
rect 14992 52192 15008 52256
rect 15072 52192 15088 52256
rect 15152 52192 15160 52256
rect 14840 51168 15160 52192
rect 14840 51104 14848 51168
rect 14912 51104 14928 51168
rect 14992 51104 15008 51168
rect 15072 51104 15088 51168
rect 15152 51104 15160 51168
rect 14840 50080 15160 51104
rect 14840 50016 14848 50080
rect 14912 50016 14928 50080
rect 14992 50016 15008 50080
rect 15072 50016 15088 50080
rect 15152 50016 15160 50080
rect 14840 48992 15160 50016
rect 14840 48928 14848 48992
rect 14912 48928 14928 48992
rect 14992 48928 15008 48992
rect 15072 48928 15088 48992
rect 15152 48928 15160 48992
rect 14840 47904 15160 48928
rect 14840 47840 14848 47904
rect 14912 47840 14928 47904
rect 14992 47840 15008 47904
rect 15072 47840 15088 47904
rect 15152 47840 15160 47904
rect 14840 46816 15160 47840
rect 14840 46752 14848 46816
rect 14912 46752 14928 46816
rect 14992 46752 15008 46816
rect 15072 46752 15088 46816
rect 15152 46752 15160 46816
rect 14840 45728 15160 46752
rect 14840 45664 14848 45728
rect 14912 45664 14928 45728
rect 14992 45664 15008 45728
rect 15072 45664 15088 45728
rect 15152 45664 15160 45728
rect 14840 44640 15160 45664
rect 14840 44576 14848 44640
rect 14912 44576 14928 44640
rect 14992 44576 15008 44640
rect 15072 44576 15088 44640
rect 15152 44576 15160 44640
rect 14840 43552 15160 44576
rect 14840 43488 14848 43552
rect 14912 43488 14928 43552
rect 14992 43488 15008 43552
rect 15072 43488 15088 43552
rect 15152 43488 15160 43552
rect 14840 42464 15160 43488
rect 14840 42400 14848 42464
rect 14912 42400 14928 42464
rect 14992 42400 15008 42464
rect 15072 42400 15088 42464
rect 15152 42400 15160 42464
rect 14840 41376 15160 42400
rect 14840 41312 14848 41376
rect 14912 41312 14928 41376
rect 14992 41312 15008 41376
rect 15072 41312 15088 41376
rect 15152 41312 15160 41376
rect 14840 40288 15160 41312
rect 14840 40224 14848 40288
rect 14912 40224 14928 40288
rect 14992 40224 15008 40288
rect 15072 40224 15088 40288
rect 15152 40224 15160 40288
rect 14840 39200 15160 40224
rect 14840 39136 14848 39200
rect 14912 39136 14928 39200
rect 14992 39136 15008 39200
rect 15072 39136 15088 39200
rect 15152 39136 15160 39200
rect 14840 38112 15160 39136
rect 14840 38048 14848 38112
rect 14912 38048 14928 38112
rect 14992 38048 15008 38112
rect 15072 38048 15088 38112
rect 15152 38048 15160 38112
rect 14840 37024 15160 38048
rect 14840 36960 14848 37024
rect 14912 36960 14928 37024
rect 14992 36960 15008 37024
rect 15072 36960 15088 37024
rect 15152 36960 15160 37024
rect 14840 35936 15160 36960
rect 14840 35872 14848 35936
rect 14912 35872 14928 35936
rect 14992 35872 15008 35936
rect 15072 35872 15088 35936
rect 15152 35872 15160 35936
rect 14840 34848 15160 35872
rect 14840 34784 14848 34848
rect 14912 34784 14928 34848
rect 14992 34784 15008 34848
rect 15072 34784 15088 34848
rect 15152 34784 15160 34848
rect 14840 33760 15160 34784
rect 14840 33696 14848 33760
rect 14912 33696 14928 33760
rect 14992 33696 15008 33760
rect 15072 33696 15088 33760
rect 15152 33696 15160 33760
rect 14840 32672 15160 33696
rect 14840 32608 14848 32672
rect 14912 32608 14928 32672
rect 14992 32608 15008 32672
rect 15072 32608 15088 32672
rect 15152 32608 15160 32672
rect 14840 31584 15160 32608
rect 14840 31520 14848 31584
rect 14912 31520 14928 31584
rect 14992 31520 15008 31584
rect 15072 31520 15088 31584
rect 15152 31520 15160 31584
rect 14840 30496 15160 31520
rect 14840 30432 14848 30496
rect 14912 30432 14928 30496
rect 14992 30432 15008 30496
rect 15072 30432 15088 30496
rect 15152 30432 15160 30496
rect 14840 29408 15160 30432
rect 14840 29344 14848 29408
rect 14912 29344 14928 29408
rect 14992 29344 15008 29408
rect 15072 29344 15088 29408
rect 15152 29344 15160 29408
rect 14840 28320 15160 29344
rect 14840 28256 14848 28320
rect 14912 28256 14928 28320
rect 14992 28256 15008 28320
rect 15072 28256 15088 28320
rect 15152 28256 15160 28320
rect 14840 27232 15160 28256
rect 14840 27168 14848 27232
rect 14912 27168 14928 27232
rect 14992 27168 15008 27232
rect 15072 27168 15088 27232
rect 15152 27168 15160 27232
rect 14840 26144 15160 27168
rect 14840 26080 14848 26144
rect 14912 26080 14928 26144
rect 14992 26080 15008 26144
rect 15072 26080 15088 26144
rect 15152 26080 15160 26144
rect 14840 25056 15160 26080
rect 14840 24992 14848 25056
rect 14912 24992 14928 25056
rect 14992 24992 15008 25056
rect 15072 24992 15088 25056
rect 15152 24992 15160 25056
rect 14840 23968 15160 24992
rect 14840 23904 14848 23968
rect 14912 23904 14928 23968
rect 14992 23904 15008 23968
rect 15072 23904 15088 23968
rect 15152 23904 15160 23968
rect 14840 22880 15160 23904
rect 14840 22816 14848 22880
rect 14912 22816 14928 22880
rect 14992 22816 15008 22880
rect 15072 22816 15088 22880
rect 15152 22816 15160 22880
rect 14840 21792 15160 22816
rect 14840 21728 14848 21792
rect 14912 21728 14928 21792
rect 14992 21728 15008 21792
rect 15072 21728 15088 21792
rect 15152 21728 15160 21792
rect 14840 20704 15160 21728
rect 14840 20640 14848 20704
rect 14912 20640 14928 20704
rect 14992 20640 15008 20704
rect 15072 20640 15088 20704
rect 15152 20640 15160 20704
rect 14840 19616 15160 20640
rect 14840 19552 14848 19616
rect 14912 19552 14928 19616
rect 14992 19552 15008 19616
rect 15072 19552 15088 19616
rect 15152 19552 15160 19616
rect 14840 18528 15160 19552
rect 14840 18464 14848 18528
rect 14912 18464 14928 18528
rect 14992 18464 15008 18528
rect 15072 18464 15088 18528
rect 15152 18464 15160 18528
rect 14840 17440 15160 18464
rect 14840 17376 14848 17440
rect 14912 17376 14928 17440
rect 14992 17376 15008 17440
rect 15072 17376 15088 17440
rect 15152 17376 15160 17440
rect 14840 16352 15160 17376
rect 14840 16288 14848 16352
rect 14912 16288 14928 16352
rect 14992 16288 15008 16352
rect 15072 16288 15088 16352
rect 15152 16288 15160 16352
rect 14840 15264 15160 16288
rect 14840 15200 14848 15264
rect 14912 15200 14928 15264
rect 14992 15200 15008 15264
rect 15072 15200 15088 15264
rect 15152 15200 15160 15264
rect 14840 14176 15160 15200
rect 14840 14112 14848 14176
rect 14912 14112 14928 14176
rect 14992 14112 15008 14176
rect 15072 14112 15088 14176
rect 15152 14112 15160 14176
rect 14840 13088 15160 14112
rect 14840 13024 14848 13088
rect 14912 13024 14928 13088
rect 14992 13024 15008 13088
rect 15072 13024 15088 13088
rect 15152 13024 15160 13088
rect 14840 12000 15160 13024
rect 14840 11936 14848 12000
rect 14912 11936 14928 12000
rect 14992 11936 15008 12000
rect 15072 11936 15088 12000
rect 15152 11936 15160 12000
rect 14840 10912 15160 11936
rect 14840 10848 14848 10912
rect 14912 10848 14928 10912
rect 14992 10848 15008 10912
rect 15072 10848 15088 10912
rect 15152 10848 15160 10912
rect 14840 9824 15160 10848
rect 14840 9760 14848 9824
rect 14912 9760 14928 9824
rect 14992 9760 15008 9824
rect 15072 9760 15088 9824
rect 15152 9760 15160 9824
rect 14840 8736 15160 9760
rect 14840 8672 14848 8736
rect 14912 8672 14928 8736
rect 14992 8672 15008 8736
rect 15072 8672 15088 8736
rect 15152 8672 15160 8736
rect 14840 7648 15160 8672
rect 14840 7584 14848 7648
rect 14912 7584 14928 7648
rect 14992 7584 15008 7648
rect 15072 7584 15088 7648
rect 15152 7584 15160 7648
rect 14840 6560 15160 7584
rect 14840 6496 14848 6560
rect 14912 6496 14928 6560
rect 14992 6496 15008 6560
rect 15072 6496 15088 6560
rect 15152 6496 15160 6560
rect 14840 5472 15160 6496
rect 14840 5408 14848 5472
rect 14912 5408 14928 5472
rect 14992 5408 15008 5472
rect 15072 5408 15088 5472
rect 15152 5408 15160 5472
rect 14840 4384 15160 5408
rect 14840 4320 14848 4384
rect 14912 4320 14928 4384
rect 14992 4320 15008 4384
rect 15072 4320 15088 4384
rect 15152 4320 15160 4384
rect 14840 3296 15160 4320
rect 14840 3232 14848 3296
rect 14912 3232 14928 3296
rect 14992 3232 15008 3296
rect 15072 3232 15088 3296
rect 15152 3232 15160 3296
rect 14840 2208 15160 3232
rect 14840 2144 14848 2208
rect 14912 2144 14928 2208
rect 14992 2144 15008 2208
rect 15072 2144 15088 2208
rect 15152 2144 15160 2208
rect 14840 2128 15160 2144
rect 19472 52800 19792 53360
rect 19472 52736 19480 52800
rect 19544 52736 19560 52800
rect 19624 52736 19640 52800
rect 19704 52736 19720 52800
rect 19784 52736 19792 52800
rect 19472 51712 19792 52736
rect 19472 51648 19480 51712
rect 19544 51648 19560 51712
rect 19624 51648 19640 51712
rect 19704 51648 19720 51712
rect 19784 51648 19792 51712
rect 19472 50624 19792 51648
rect 19472 50560 19480 50624
rect 19544 50560 19560 50624
rect 19624 50560 19640 50624
rect 19704 50560 19720 50624
rect 19784 50560 19792 50624
rect 19472 49536 19792 50560
rect 19472 49472 19480 49536
rect 19544 49472 19560 49536
rect 19624 49472 19640 49536
rect 19704 49472 19720 49536
rect 19784 49472 19792 49536
rect 19472 48448 19792 49472
rect 19472 48384 19480 48448
rect 19544 48384 19560 48448
rect 19624 48384 19640 48448
rect 19704 48384 19720 48448
rect 19784 48384 19792 48448
rect 19472 47360 19792 48384
rect 19472 47296 19480 47360
rect 19544 47296 19560 47360
rect 19624 47296 19640 47360
rect 19704 47296 19720 47360
rect 19784 47296 19792 47360
rect 19472 46272 19792 47296
rect 19472 46208 19480 46272
rect 19544 46208 19560 46272
rect 19624 46208 19640 46272
rect 19704 46208 19720 46272
rect 19784 46208 19792 46272
rect 19472 45184 19792 46208
rect 19472 45120 19480 45184
rect 19544 45120 19560 45184
rect 19624 45120 19640 45184
rect 19704 45120 19720 45184
rect 19784 45120 19792 45184
rect 19472 44096 19792 45120
rect 19472 44032 19480 44096
rect 19544 44032 19560 44096
rect 19624 44032 19640 44096
rect 19704 44032 19720 44096
rect 19784 44032 19792 44096
rect 19472 43008 19792 44032
rect 19472 42944 19480 43008
rect 19544 42944 19560 43008
rect 19624 42944 19640 43008
rect 19704 42944 19720 43008
rect 19784 42944 19792 43008
rect 19472 41920 19792 42944
rect 19472 41856 19480 41920
rect 19544 41856 19560 41920
rect 19624 41856 19640 41920
rect 19704 41856 19720 41920
rect 19784 41856 19792 41920
rect 19472 40832 19792 41856
rect 19472 40768 19480 40832
rect 19544 40768 19560 40832
rect 19624 40768 19640 40832
rect 19704 40768 19720 40832
rect 19784 40768 19792 40832
rect 19472 39744 19792 40768
rect 19472 39680 19480 39744
rect 19544 39680 19560 39744
rect 19624 39680 19640 39744
rect 19704 39680 19720 39744
rect 19784 39680 19792 39744
rect 19472 38656 19792 39680
rect 19472 38592 19480 38656
rect 19544 38592 19560 38656
rect 19624 38592 19640 38656
rect 19704 38592 19720 38656
rect 19784 38592 19792 38656
rect 19472 37568 19792 38592
rect 19472 37504 19480 37568
rect 19544 37504 19560 37568
rect 19624 37504 19640 37568
rect 19704 37504 19720 37568
rect 19784 37504 19792 37568
rect 19472 36480 19792 37504
rect 19472 36416 19480 36480
rect 19544 36416 19560 36480
rect 19624 36416 19640 36480
rect 19704 36416 19720 36480
rect 19784 36416 19792 36480
rect 19472 35392 19792 36416
rect 19472 35328 19480 35392
rect 19544 35328 19560 35392
rect 19624 35328 19640 35392
rect 19704 35328 19720 35392
rect 19784 35328 19792 35392
rect 19472 34304 19792 35328
rect 19472 34240 19480 34304
rect 19544 34240 19560 34304
rect 19624 34240 19640 34304
rect 19704 34240 19720 34304
rect 19784 34240 19792 34304
rect 19472 33216 19792 34240
rect 19472 33152 19480 33216
rect 19544 33152 19560 33216
rect 19624 33152 19640 33216
rect 19704 33152 19720 33216
rect 19784 33152 19792 33216
rect 19472 32128 19792 33152
rect 19472 32064 19480 32128
rect 19544 32064 19560 32128
rect 19624 32064 19640 32128
rect 19704 32064 19720 32128
rect 19784 32064 19792 32128
rect 19472 31040 19792 32064
rect 19472 30976 19480 31040
rect 19544 30976 19560 31040
rect 19624 30976 19640 31040
rect 19704 30976 19720 31040
rect 19784 30976 19792 31040
rect 19472 29952 19792 30976
rect 19472 29888 19480 29952
rect 19544 29888 19560 29952
rect 19624 29888 19640 29952
rect 19704 29888 19720 29952
rect 19784 29888 19792 29952
rect 19472 28864 19792 29888
rect 19472 28800 19480 28864
rect 19544 28800 19560 28864
rect 19624 28800 19640 28864
rect 19704 28800 19720 28864
rect 19784 28800 19792 28864
rect 19472 27776 19792 28800
rect 19472 27712 19480 27776
rect 19544 27712 19560 27776
rect 19624 27712 19640 27776
rect 19704 27712 19720 27776
rect 19784 27712 19792 27776
rect 19472 26688 19792 27712
rect 19472 26624 19480 26688
rect 19544 26624 19560 26688
rect 19624 26624 19640 26688
rect 19704 26624 19720 26688
rect 19784 26624 19792 26688
rect 19472 25600 19792 26624
rect 19472 25536 19480 25600
rect 19544 25536 19560 25600
rect 19624 25536 19640 25600
rect 19704 25536 19720 25600
rect 19784 25536 19792 25600
rect 19472 24512 19792 25536
rect 19472 24448 19480 24512
rect 19544 24448 19560 24512
rect 19624 24448 19640 24512
rect 19704 24448 19720 24512
rect 19784 24448 19792 24512
rect 19472 23424 19792 24448
rect 19472 23360 19480 23424
rect 19544 23360 19560 23424
rect 19624 23360 19640 23424
rect 19704 23360 19720 23424
rect 19784 23360 19792 23424
rect 19472 22336 19792 23360
rect 19472 22272 19480 22336
rect 19544 22272 19560 22336
rect 19624 22272 19640 22336
rect 19704 22272 19720 22336
rect 19784 22272 19792 22336
rect 19472 21248 19792 22272
rect 19472 21184 19480 21248
rect 19544 21184 19560 21248
rect 19624 21184 19640 21248
rect 19704 21184 19720 21248
rect 19784 21184 19792 21248
rect 19472 20160 19792 21184
rect 19472 20096 19480 20160
rect 19544 20096 19560 20160
rect 19624 20096 19640 20160
rect 19704 20096 19720 20160
rect 19784 20096 19792 20160
rect 19472 19072 19792 20096
rect 19472 19008 19480 19072
rect 19544 19008 19560 19072
rect 19624 19008 19640 19072
rect 19704 19008 19720 19072
rect 19784 19008 19792 19072
rect 19472 17984 19792 19008
rect 19472 17920 19480 17984
rect 19544 17920 19560 17984
rect 19624 17920 19640 17984
rect 19704 17920 19720 17984
rect 19784 17920 19792 17984
rect 19472 16896 19792 17920
rect 19472 16832 19480 16896
rect 19544 16832 19560 16896
rect 19624 16832 19640 16896
rect 19704 16832 19720 16896
rect 19784 16832 19792 16896
rect 19472 15808 19792 16832
rect 19472 15744 19480 15808
rect 19544 15744 19560 15808
rect 19624 15744 19640 15808
rect 19704 15744 19720 15808
rect 19784 15744 19792 15808
rect 19472 14720 19792 15744
rect 19472 14656 19480 14720
rect 19544 14656 19560 14720
rect 19624 14656 19640 14720
rect 19704 14656 19720 14720
rect 19784 14656 19792 14720
rect 19472 13632 19792 14656
rect 19472 13568 19480 13632
rect 19544 13568 19560 13632
rect 19624 13568 19640 13632
rect 19704 13568 19720 13632
rect 19784 13568 19792 13632
rect 19472 12544 19792 13568
rect 19472 12480 19480 12544
rect 19544 12480 19560 12544
rect 19624 12480 19640 12544
rect 19704 12480 19720 12544
rect 19784 12480 19792 12544
rect 19472 11456 19792 12480
rect 19472 11392 19480 11456
rect 19544 11392 19560 11456
rect 19624 11392 19640 11456
rect 19704 11392 19720 11456
rect 19784 11392 19792 11456
rect 19472 10368 19792 11392
rect 19472 10304 19480 10368
rect 19544 10304 19560 10368
rect 19624 10304 19640 10368
rect 19704 10304 19720 10368
rect 19784 10304 19792 10368
rect 19472 9280 19792 10304
rect 19472 9216 19480 9280
rect 19544 9216 19560 9280
rect 19624 9216 19640 9280
rect 19704 9216 19720 9280
rect 19784 9216 19792 9280
rect 19472 8192 19792 9216
rect 19472 8128 19480 8192
rect 19544 8128 19560 8192
rect 19624 8128 19640 8192
rect 19704 8128 19720 8192
rect 19784 8128 19792 8192
rect 19472 7104 19792 8128
rect 19472 7040 19480 7104
rect 19544 7040 19560 7104
rect 19624 7040 19640 7104
rect 19704 7040 19720 7104
rect 19784 7040 19792 7104
rect 19472 6016 19792 7040
rect 19472 5952 19480 6016
rect 19544 5952 19560 6016
rect 19624 5952 19640 6016
rect 19704 5952 19720 6016
rect 19784 5952 19792 6016
rect 19472 4928 19792 5952
rect 19472 4864 19480 4928
rect 19544 4864 19560 4928
rect 19624 4864 19640 4928
rect 19704 4864 19720 4928
rect 19784 4864 19792 4928
rect 19472 3840 19792 4864
rect 19472 3776 19480 3840
rect 19544 3776 19560 3840
rect 19624 3776 19640 3840
rect 19704 3776 19720 3840
rect 19784 3776 19792 3840
rect 19472 2752 19792 3776
rect 19472 2688 19480 2752
rect 19544 2688 19560 2752
rect 19624 2688 19640 2752
rect 19704 2688 19720 2752
rect 19784 2688 19792 2752
rect 19472 2128 19792 2688
rect 24104 53344 24424 53360
rect 24104 53280 24112 53344
rect 24176 53280 24192 53344
rect 24256 53280 24272 53344
rect 24336 53280 24352 53344
rect 24416 53280 24424 53344
rect 24104 52256 24424 53280
rect 24104 52192 24112 52256
rect 24176 52192 24192 52256
rect 24256 52192 24272 52256
rect 24336 52192 24352 52256
rect 24416 52192 24424 52256
rect 24104 51168 24424 52192
rect 24104 51104 24112 51168
rect 24176 51104 24192 51168
rect 24256 51104 24272 51168
rect 24336 51104 24352 51168
rect 24416 51104 24424 51168
rect 24104 50080 24424 51104
rect 24104 50016 24112 50080
rect 24176 50016 24192 50080
rect 24256 50016 24272 50080
rect 24336 50016 24352 50080
rect 24416 50016 24424 50080
rect 24104 48992 24424 50016
rect 24104 48928 24112 48992
rect 24176 48928 24192 48992
rect 24256 48928 24272 48992
rect 24336 48928 24352 48992
rect 24416 48928 24424 48992
rect 24104 47904 24424 48928
rect 24104 47840 24112 47904
rect 24176 47840 24192 47904
rect 24256 47840 24272 47904
rect 24336 47840 24352 47904
rect 24416 47840 24424 47904
rect 24104 46816 24424 47840
rect 24104 46752 24112 46816
rect 24176 46752 24192 46816
rect 24256 46752 24272 46816
rect 24336 46752 24352 46816
rect 24416 46752 24424 46816
rect 24104 45728 24424 46752
rect 24104 45664 24112 45728
rect 24176 45664 24192 45728
rect 24256 45664 24272 45728
rect 24336 45664 24352 45728
rect 24416 45664 24424 45728
rect 24104 44640 24424 45664
rect 24104 44576 24112 44640
rect 24176 44576 24192 44640
rect 24256 44576 24272 44640
rect 24336 44576 24352 44640
rect 24416 44576 24424 44640
rect 24104 43552 24424 44576
rect 24104 43488 24112 43552
rect 24176 43488 24192 43552
rect 24256 43488 24272 43552
rect 24336 43488 24352 43552
rect 24416 43488 24424 43552
rect 24104 42464 24424 43488
rect 24104 42400 24112 42464
rect 24176 42400 24192 42464
rect 24256 42400 24272 42464
rect 24336 42400 24352 42464
rect 24416 42400 24424 42464
rect 24104 41376 24424 42400
rect 24104 41312 24112 41376
rect 24176 41312 24192 41376
rect 24256 41312 24272 41376
rect 24336 41312 24352 41376
rect 24416 41312 24424 41376
rect 24104 40288 24424 41312
rect 24104 40224 24112 40288
rect 24176 40224 24192 40288
rect 24256 40224 24272 40288
rect 24336 40224 24352 40288
rect 24416 40224 24424 40288
rect 24104 39200 24424 40224
rect 24104 39136 24112 39200
rect 24176 39136 24192 39200
rect 24256 39136 24272 39200
rect 24336 39136 24352 39200
rect 24416 39136 24424 39200
rect 24104 38112 24424 39136
rect 24104 38048 24112 38112
rect 24176 38048 24192 38112
rect 24256 38048 24272 38112
rect 24336 38048 24352 38112
rect 24416 38048 24424 38112
rect 24104 37024 24424 38048
rect 24104 36960 24112 37024
rect 24176 36960 24192 37024
rect 24256 36960 24272 37024
rect 24336 36960 24352 37024
rect 24416 36960 24424 37024
rect 24104 35936 24424 36960
rect 24104 35872 24112 35936
rect 24176 35872 24192 35936
rect 24256 35872 24272 35936
rect 24336 35872 24352 35936
rect 24416 35872 24424 35936
rect 24104 34848 24424 35872
rect 24104 34784 24112 34848
rect 24176 34784 24192 34848
rect 24256 34784 24272 34848
rect 24336 34784 24352 34848
rect 24416 34784 24424 34848
rect 24104 33760 24424 34784
rect 24104 33696 24112 33760
rect 24176 33696 24192 33760
rect 24256 33696 24272 33760
rect 24336 33696 24352 33760
rect 24416 33696 24424 33760
rect 24104 32672 24424 33696
rect 24104 32608 24112 32672
rect 24176 32608 24192 32672
rect 24256 32608 24272 32672
rect 24336 32608 24352 32672
rect 24416 32608 24424 32672
rect 24104 31584 24424 32608
rect 24104 31520 24112 31584
rect 24176 31520 24192 31584
rect 24256 31520 24272 31584
rect 24336 31520 24352 31584
rect 24416 31520 24424 31584
rect 24104 30496 24424 31520
rect 24104 30432 24112 30496
rect 24176 30432 24192 30496
rect 24256 30432 24272 30496
rect 24336 30432 24352 30496
rect 24416 30432 24424 30496
rect 24104 29408 24424 30432
rect 24104 29344 24112 29408
rect 24176 29344 24192 29408
rect 24256 29344 24272 29408
rect 24336 29344 24352 29408
rect 24416 29344 24424 29408
rect 24104 28320 24424 29344
rect 24104 28256 24112 28320
rect 24176 28256 24192 28320
rect 24256 28256 24272 28320
rect 24336 28256 24352 28320
rect 24416 28256 24424 28320
rect 24104 27232 24424 28256
rect 24104 27168 24112 27232
rect 24176 27168 24192 27232
rect 24256 27168 24272 27232
rect 24336 27168 24352 27232
rect 24416 27168 24424 27232
rect 24104 26144 24424 27168
rect 24104 26080 24112 26144
rect 24176 26080 24192 26144
rect 24256 26080 24272 26144
rect 24336 26080 24352 26144
rect 24416 26080 24424 26144
rect 24104 25056 24424 26080
rect 24104 24992 24112 25056
rect 24176 24992 24192 25056
rect 24256 24992 24272 25056
rect 24336 24992 24352 25056
rect 24416 24992 24424 25056
rect 24104 23968 24424 24992
rect 24104 23904 24112 23968
rect 24176 23904 24192 23968
rect 24256 23904 24272 23968
rect 24336 23904 24352 23968
rect 24416 23904 24424 23968
rect 24104 22880 24424 23904
rect 24104 22816 24112 22880
rect 24176 22816 24192 22880
rect 24256 22816 24272 22880
rect 24336 22816 24352 22880
rect 24416 22816 24424 22880
rect 24104 21792 24424 22816
rect 24104 21728 24112 21792
rect 24176 21728 24192 21792
rect 24256 21728 24272 21792
rect 24336 21728 24352 21792
rect 24416 21728 24424 21792
rect 24104 20704 24424 21728
rect 24104 20640 24112 20704
rect 24176 20640 24192 20704
rect 24256 20640 24272 20704
rect 24336 20640 24352 20704
rect 24416 20640 24424 20704
rect 24104 19616 24424 20640
rect 24104 19552 24112 19616
rect 24176 19552 24192 19616
rect 24256 19552 24272 19616
rect 24336 19552 24352 19616
rect 24416 19552 24424 19616
rect 24104 18528 24424 19552
rect 24104 18464 24112 18528
rect 24176 18464 24192 18528
rect 24256 18464 24272 18528
rect 24336 18464 24352 18528
rect 24416 18464 24424 18528
rect 24104 17440 24424 18464
rect 24104 17376 24112 17440
rect 24176 17376 24192 17440
rect 24256 17376 24272 17440
rect 24336 17376 24352 17440
rect 24416 17376 24424 17440
rect 24104 16352 24424 17376
rect 24104 16288 24112 16352
rect 24176 16288 24192 16352
rect 24256 16288 24272 16352
rect 24336 16288 24352 16352
rect 24416 16288 24424 16352
rect 24104 15264 24424 16288
rect 24104 15200 24112 15264
rect 24176 15200 24192 15264
rect 24256 15200 24272 15264
rect 24336 15200 24352 15264
rect 24416 15200 24424 15264
rect 24104 14176 24424 15200
rect 24104 14112 24112 14176
rect 24176 14112 24192 14176
rect 24256 14112 24272 14176
rect 24336 14112 24352 14176
rect 24416 14112 24424 14176
rect 24104 13088 24424 14112
rect 24104 13024 24112 13088
rect 24176 13024 24192 13088
rect 24256 13024 24272 13088
rect 24336 13024 24352 13088
rect 24416 13024 24424 13088
rect 24104 12000 24424 13024
rect 24104 11936 24112 12000
rect 24176 11936 24192 12000
rect 24256 11936 24272 12000
rect 24336 11936 24352 12000
rect 24416 11936 24424 12000
rect 24104 10912 24424 11936
rect 24104 10848 24112 10912
rect 24176 10848 24192 10912
rect 24256 10848 24272 10912
rect 24336 10848 24352 10912
rect 24416 10848 24424 10912
rect 24104 9824 24424 10848
rect 24104 9760 24112 9824
rect 24176 9760 24192 9824
rect 24256 9760 24272 9824
rect 24336 9760 24352 9824
rect 24416 9760 24424 9824
rect 24104 8736 24424 9760
rect 24104 8672 24112 8736
rect 24176 8672 24192 8736
rect 24256 8672 24272 8736
rect 24336 8672 24352 8736
rect 24416 8672 24424 8736
rect 24104 7648 24424 8672
rect 24104 7584 24112 7648
rect 24176 7584 24192 7648
rect 24256 7584 24272 7648
rect 24336 7584 24352 7648
rect 24416 7584 24424 7648
rect 24104 6560 24424 7584
rect 24104 6496 24112 6560
rect 24176 6496 24192 6560
rect 24256 6496 24272 6560
rect 24336 6496 24352 6560
rect 24416 6496 24424 6560
rect 24104 5472 24424 6496
rect 24104 5408 24112 5472
rect 24176 5408 24192 5472
rect 24256 5408 24272 5472
rect 24336 5408 24352 5472
rect 24416 5408 24424 5472
rect 24104 4384 24424 5408
rect 24104 4320 24112 4384
rect 24176 4320 24192 4384
rect 24256 4320 24272 4384
rect 24336 4320 24352 4384
rect 24416 4320 24424 4384
rect 24104 3296 24424 4320
rect 24104 3232 24112 3296
rect 24176 3232 24192 3296
rect 24256 3232 24272 3296
rect 24336 3232 24352 3296
rect 24416 3232 24424 3296
rect 24104 2208 24424 3232
rect 24104 2144 24112 2208
rect 24176 2144 24192 2208
rect 24256 2144 24272 2208
rect 24336 2144 24352 2208
rect 24416 2144 24424 2208
rect 24104 2128 24424 2144
use sky130_fd_sc_hd__fill_2  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input156 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input147
timestamp 1623621585
transform 1 0 1564 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1623621585
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1623621585
transform 1 0 1932 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11
timestamp 1623621585
transform 1 0 2116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output248
timestamp 1623621585
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 2300 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_1_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 2944 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19
timestamp 1623621585
transform 1 0 2852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1623621585
transform 1 0 3864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 3680 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1623621585
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1623621585
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 3772 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1623621585
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1790_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 4232 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1770_
timestamp 1623621585
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 4508 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44
timestamp 1623621585
transform 1 0 5152 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37
timestamp 1623621585
transform 1 0 4508 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 4876 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _2221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 5060 0 1 2720
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2222_
timestamp 1623621585
transform 1 0 6992 0 1 2720
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1623621585
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 5704 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1623621585
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59
timestamp 1623621585
transform 1 0 6532 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67
timestamp 1623621585
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_60
timestamp 1623621585
transform 1 0 6624 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1623621585
transform 1 0 8004 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 8372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 7452 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_87
timestamp 1623621585
transform 1 0 9108 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_85
timestamp 1623621585
transform 1 0 8924 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1623621585
transform 1 0 8556 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1623621585
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1623621585
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82
timestamp 1623621585
transform 1 0 8648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1623621585
transform 1 0 9016 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1623621585
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 9476 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1789_
timestamp 1623621585
transform 1 0 11132 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2011_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 11500 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1623621585
transform 1 0 9568 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1623621585
transform 1 0 10212 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95
timestamp 1623621585
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102
timestamp 1623621585
transform 1 0 10488 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108
timestamp 1623621585
transform 1 0 11040 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1623621585
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_107
timestamp 1623621585
transform 1 0 10948 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1623621585
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1623621585
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1623621585
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_122
timestamp 1623621585
transform 1 0 12328 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124
timestamp 1623621585
transform 1 0 12512 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1623621585
transform 1 0 12696 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_129
timestamp 1623621585
transform 1 0 12972 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_131
timestamp 1623621585
transform 1 0 13156 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1813_
timestamp 1623621585
transform 1 0 12880 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_135
timestamp 1623621585
transform 1 0 13524 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137
timestamp 1623621585
transform 1 0 13708 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1623621585
transform 1 0 13616 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_144
timestamp 1623621585
transform 1 0 14352 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1623621585
transform 1 0 13892 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1623621585
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1623621585
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1623621585
transform 1 0 14260 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1623621585
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1812_
timestamp 1623621585
transform 1 0 13800 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_148
timestamp 1623621585
transform 1 0 14720 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1623621585
transform 1 0 15180 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2005_
timestamp 1623621585
transform 1 0 14812 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1623621585
transform 1 0 14904 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_158
timestamp 1623621585
transform 1 0 15640 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1623621585
transform 1 0 15548 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_168
timestamp 1623621585
transform 1 0 16560 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_164
timestamp 1623621585
transform 1 0 16192 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_167
timestamp 1623621585
transform 1 0 16468 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_160
timestamp 1623621585
transform 1 0 15824 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1623621585
transform 1 0 16192 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1623621585
transform 1 0 16284 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_172
timestamp 1623621585
transform 1 0 16928 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1623621585
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1623621585
transform 1 0 17020 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1623621585
transform 1 0 17572 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1623621585
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _2003_
timestamp 1623621585
transform 1 0 17020 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_182
timestamp 1623621585
transform 1 0 17848 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1623621585
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_189
timestamp 1623621585
transform 1 0 18492 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1623621585
transform 1 0 18492 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1623621585
transform 1 0 18216 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1623621585
transform 1 0 18216 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_196
timestamp 1623621585
transform 1 0 19136 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1623621585
transform 1 0 19044 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1623621585
transform 1 0 19136 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1623621585
transform 1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1623621585
transform 1 0 19596 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1623621585
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1623621585
transform 1 0 19504 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1623621585
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1623621585
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1623621585
transform 1 0 19964 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1079_
timestamp 1623621585
transform 1 0 21528 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _2272_
timestamp 1623621585
transform 1 0 20976 0 1 2720
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1623621585
transform 1 0 20884 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1623621585
transform 1 0 20240 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_211
timestamp 1623621585
transform 1 0 20516 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1623621585
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225
timestamp 1623621585
transform 1 0 21804 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_208
timestamp 1623621585
transform 1 0 20240 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_233
timestamp 1623621585
transform 1 0 22540 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_237
timestamp 1623621585
transform 1 0 22908 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1623621585
transform 1 0 22540 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_231
timestamp 1623621585
transform 1 0 22356 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1623621585
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 22908 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_245
timestamp 1623621585
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1623621585
transform 1 0 23276 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output221
timestamp 1623621585
transform 1 0 23644 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1811_
timestamp 1623621585
transform 1 0 23000 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_249
timestamp 1623621585
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output230
timestamp 1623621585
transform 1 0 24012 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_258
timestamp 1623621585
transform 1 0 24840 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_253
timestamp 1623621585
transform 1 0 24380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1623621585
transform 1 0 24748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output212
timestamp 1623621585
transform 1 0 24380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1623621585
transform 1 0 24748 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_262
timestamp 1623621585
transform 1 0 25208 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1623621585
transform 1 0 25208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output194
timestamp 1623621585
transform 1 0 25576 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1623621585
transform 1 0 25116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1121_
timestamp 1623621585
transform 1 0 25300 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_271
timestamp 1623621585
transform 1 0 26036 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_270
timestamp 1623621585
transform 1 0 25944 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output185
timestamp 1623621585
transform 1 0 26312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_282
timestamp 1623621585
transform 1 0 27048 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_277
timestamp 1623621585
transform 1 0 26588 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_278
timestamp 1623621585
transform 1 0 26680 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output203
timestamp 1623621585
transform 1 0 26680 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output176
timestamp 1623621585
transform 1 0 27048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_291
timestamp 1623621585
transform 1 0 27876 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1623621585
transform 1 0 27416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1623621585
transform 1 0 27784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1997_
timestamp 1623621585
transform 1 0 27416 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_295
timestamp 1623621585
transform 1 0 28244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1623621585
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1623621585
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1703_
timestamp 1623621585
transform 1 0 1564 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _2230_
timestamp 1623621585
transform 1 0 2760 0 -1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1623621585
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1623621585
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_8
timestamp 1623621585
transform 1 0 1840 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_16
timestamp 1623621585
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1017_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 4692 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_35
timestamp 1623621585
transform 1 0 4324 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1351_
timestamp 1623621585
transform 1 0 6808 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1623621585
transform 1 0 6348 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_48
timestamp 1623621585
transform 1 0 5520 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_56
timestamp 1623621585
transform 1 0 6256 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_58
timestamp 1623621585
transform 1 0 6440 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1623621585
transform 1 0 9384 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1352_
timestamp 1623621585
transform 1 0 8188 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_2_71
timestamp 1623621585
transform 1 0 7636 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_84
timestamp 1623621585
transform 1 0 8832 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1623621585
transform 1 0 10580 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1623621585
transform 1 0 11592 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_93
timestamp 1623621585
transform 1 0 9660 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1623621585
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_106
timestamp 1623621585
transform 1 0 10856 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2260_
timestamp 1623621585
transform 1 0 12420 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_2_115
timestamp 1623621585
transform 1 0 11684 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2266_
timestamp 1623621585
transform 1 0 14352 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_139
timestamp 1623621585
transform 1 0 13892 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_143
timestamp 1623621585
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1089_
timestamp 1623621585
transform 1 0 17296 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1136_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 16192 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1623621585
transform 1 0 16836 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_160
timestamp 1623621585
transform 1 0 15824 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1623621585
transform 1 0 16468 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1623621585
transform 1 0 16928 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1623621585
transform 1 0 17572 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2001_
timestamp 1623621585
transform 1 0 19872 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _2270_
timestamp 1623621585
transform 1 0 17940 0 -1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 19688 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_200
timestamp 1623621585
transform 1 0 19504 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _1125_
timestamp 1623621585
transform 1 0 21068 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1623621585
transform 1 0 22080 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_213
timestamp 1623621585
transform 1 0 20700 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_220
timestamp 1623621585
transform 1 0 21344 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1118_
timestamp 1623621585
transform 1 0 22540 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _2273_
timestamp 1623621585
transform 1 0 23184 0 -1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_2_229
timestamp 1623621585
transform 1 0 22172 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_236
timestamp 1623621585
transform 1 0 22816 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1119_
timestamp 1623621585
transform 1 0 25300 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_257
timestamp 1623621585
transform 1 0 24748 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_271
timestamp 1623621585
transform 1 0 26036 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1623621585
transform 1 0 27324 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output177
timestamp 1623621585
transform 1 0 27876 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output195
timestamp 1623621585
transform 1 0 26588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_281
timestamp 1623621585
transform 1 0 26956 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_286
timestamp 1623621585
transform 1 0 27416 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_290
timestamp 1623621585
transform 1 0 27784 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1623621585
transform 1 0 28244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1623621585
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1281_
timestamp 1623621585
transform 1 0 2576 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1746_
timestamp 1623621585
transform 1 0 1564 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1623621585
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1623621585
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_8
timestamp 1623621585
transform 1 0 1840 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _2231_
timestamp 1623621585
transform 1 0 4232 0 1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1623621585
transform 1 0 3772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_25
timestamp 1623621585
transform 1 0 3404 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1623621585
transform 1 0 3864 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1353_
timestamp 1623621585
transform 1 0 6164 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1623621585
transform 1 0 5796 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_64
timestamp 1623621585
transform 1 0 6992 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_68
timestamp 1623621585
transform 1 0 7360 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_2  _1298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 7452 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1623621585
transform 1 0 9016 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_82
timestamp 1623621585
transform 1 0 8648 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_87
timestamp 1623621585
transform 1 0 9108 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_91
timestamp 1623621585
transform 1 0 9476 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1295_
timestamp 1623621585
transform 1 0 10764 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1450_
timestamp 1623621585
transform 1 0 9568 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1623621585
transform 1 0 11500 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_101
timestamp 1623621585
transform 1 0 10396 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1623621585
transform 1 0 11040 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_112
timestamp 1623621585
transform 1 0 11408 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1155_
timestamp 1623621585
transform 1 0 12236 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1156_
timestamp 1623621585
transform 1 0 12880 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_116
timestamp 1623621585
transform 1 0 11776 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_120
timestamp 1623621585
transform 1 0 12144 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_124
timestamp 1623621585
transform 1 0 12512 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_136
timestamp 1623621585
transform 1 0 13616 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1142_
timestamp 1623621585
transform 1 0 14720 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1623621585
transform 1 0 14260 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_142
timestamp 1623621585
transform 1 0 14168 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_144
timestamp 1623621585
transform 1 0 14352 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_156
timestamp 1623621585
transform 1 0 15456 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2268_
timestamp 1623621585
transform 1 0 15916 0 1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_3_160
timestamp 1623621585
transform 1 0 15824 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_178
timestamp 1623621585
transform 1 0 17480 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1129_
timestamp 1623621585
transform 1 0 18400 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _2271_
timestamp 1623621585
transform 1 0 19964 0 1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1623621585
transform 1 0 19504 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_186
timestamp 1623621585
transform 1 0 18216 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_196
timestamp 1623621585
transform 1 0 19136 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_201
timestamp 1623621585
transform 1 0 19596 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1123_
timestamp 1623621585
transform 1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_222
timestamp 1623621585
transform 1 0 21528 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1623621585
transform 1 0 24104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1999_
timestamp 1623621585
transform 1 0 22540 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_1
timestamp 1623621585
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_229
timestamp 1623621585
transform 1 0 22172 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_242
timestamp 1623621585
transform 1 0 23368 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _2274_
timestamp 1623621585
transform 1 0 26036 0 1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1623621585
transform 1 0 24748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output239
timestamp 1623621585
transform 1 0 25300 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_253
timestamp 1623621585
transform 1 0 24380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_258
timestamp 1623621585
transform 1 0 24840 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_262
timestamp 1623621585
transform 1 0 25208 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_267
timestamp 1623621585
transform 1 0 25668 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1623621585
transform 1 0 27968 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_288
timestamp 1623621585
transform 1 0 27600 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_295
timestamp 1623621585
transform 1 0 28244 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1623621585
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1623621585
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1623621585
transform 1 0 1748 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1623621585
transform 1 0 2392 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1623621585
transform 1 0 3036 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1623621585
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1623621585
transform 1 0 2024 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1623621585
transform 1 0 2668 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1279_
timestamp 1623621585
transform 1 0 4140 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_24
timestamp 1623621585
transform 1 0 3312 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_32
timestamp 1623621585
transform 1 0 4048 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_42
timestamp 1623621585
transform 1 0 4968 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1350_
timestamp 1623621585
transform 1 0 6808 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1623621585
transform 1 0 6348 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1623621585
transform 1 0 5336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_49
timestamp 1623621585
transform 1 0 5612 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_58
timestamp 1623621585
transform 1 0 6440 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_4  _1300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 8096 0 -1 4896
box -38 -48 1418 592
use sky130_fd_sc_hd__decap_6  FILLER_4_69
timestamp 1623621585
transform 1 0 7452 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_75
timestamp 1623621585
transform 1 0 8004 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_91
timestamp 1623621585
transform 1 0 9476 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1297_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 9936 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1623621585
transform 1 0 11592 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_95
timestamp 1623621585
transform 1 0 9844 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_109
timestamp 1623621585
transform 1 0 11132 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_113
timestamp 1623621585
transform 1 0 11500 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1117_
timestamp 1623621585
transform 1 0 13708 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1788_
timestamp 1623621585
transform 1 0 12328 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_115
timestamp 1623621585
transform 1 0 11684 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_121
timestamp 1623621585
transform 1 0 12236 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_125 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 12604 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__o211a_1  _1137_
timestamp 1623621585
transform 1 0 15732 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1141_
timestamp 1623621585
transform 1 0 14444 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1702_
timestamp 1623621585
transform 1 0 15088 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1623621585
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1623621585
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_155
timestamp 1623621585
transform 1 0 15364 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1132_
timestamp 1623621585
transform 1 0 17848 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1623621585
transform 1 0 16836 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_167
timestamp 1623621585
transform 1 0 16468 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_172
timestamp 1623621585
transform 1 0 16928 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_180
timestamp 1623621585
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _1128_
timestamp 1623621585
transform 1 0 18952 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2002_
timestamp 1623621585
transform 1 0 19596 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_190
timestamp 1623621585
transform 1 0 18584 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_197
timestamp 1623621585
transform 1 0 19228 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1126_
timestamp 1623621585
transform 1 0 20976 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1623621585
transform 1 0 22080 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_210
timestamp 1623621585
transform 1 0 20424 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_224
timestamp 1623621585
transform 1 0 21712 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _2000_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 23000 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_229
timestamp 1623621585
transform 1 0 22172 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_237
timestamp 1623621585
transform 1 0 22908 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_247
timestamp 1623621585
transform 1 0 23828 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1623621585
transform 1 0 24472 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _2275_
timestamp 1623621585
transform 1 0 25392 0 -1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_4_253
timestamp 1623621585
transform 1 0 24380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_257
timestamp 1623621585
transform 1 0 24748 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_263
timestamp 1623621585
transform 1 0 25300 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1623621585
transform 1 0 27324 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output186
timestamp 1623621585
transform 1 0 27876 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_281
timestamp 1623621585
transform 1 0 26956 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_286
timestamp 1623621585
transform 1 0 27416 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_290
timestamp 1623621585
transform 1 0 27784 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_295
timestamp 1623621585
transform 1 0 28244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1623621585
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 2668 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1623621585
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1623621585
transform 1 0 1748 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1623621585
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_10
timestamp 1623621585
transform 1 0 2024 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_16
timestamp 1623621585
transform 1 0 2576 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _2228_
timestamp 1623621585
transform 1 0 4416 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1623621585
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_23
timestamp 1623621585
transform 1 0 3220 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_30
timestamp 1623621585
transform 1 0 3864 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input139
timestamp 1623621585
transform 1 0 6348 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input158
timestamp 1623621585
transform 1 0 6992 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_53
timestamp 1623621585
transform 1 0 5980 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_60
timestamp 1623621585
transform 1 0 6624 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_67
timestamp 1623621585
transform 1 0 7268 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 8188 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1623621585
transform 1 0 9016 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_75
timestamp 1623621585
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_80
timestamp 1623621585
transform 1 0 8464 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_87
timestamp 1623621585
transform 1 0 9108 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1296_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 9936 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1356_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 11132 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_95
timestamp 1623621585
transform 1 0 9844 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_105
timestamp 1623621585
transform 1 0 10764 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1140_
timestamp 1623621585
transform 1 0 13524 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1355_
timestamp 1623621585
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_115
timestamp 1623621585
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_122
timestamp 1623621585
transform 1 0 12328 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_134
timestamp 1623621585
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1623621585
transform 1 0 14260 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp 1623621585
transform 1 0 13892 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_144
timestamp 1623621585
transform 1 0 14352 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_156
timestamp 1623621585
transform 1 0 15456 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1130_
timestamp 1623621585
transform 1 0 16284 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1131_
timestamp 1623621585
transform 1 0 17572 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_164
timestamp 1623621585
transform 1 0 16192 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1623621585
transform 1 0 16652 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1623621585
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_182
timestamp 1623621585
transform 1 0 17848 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1116_
timestamp 1623621585
transform 1 0 18216 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1623621585
transform 1 0 19504 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1623621585
transform 1 0 19964 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_190
timestamp 1623621585
transform 1 0 18584 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_198
timestamp 1623621585
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_201
timestamp 1623621585
transform 1 0 19596 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1623621585
transform 1 0 21068 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_208
timestamp 1623621585
transform 1 0 20240 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_216
timestamp 1623621585
transform 1 0 20976 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1623621585
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1120_
timestamp 1623621585
transform 1 0 24104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1623621585
transform 1 0 23460 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_232
timestamp 1623621585
transform 1 0 22448 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_240
timestamp 1623621585
transform 1 0 23184 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_246
timestamp 1623621585
transform 1 0 23736 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1066_
timestamp 1623621585
transform 1 0 25668 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1623621585
transform 1 0 24748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output213
timestamp 1623621585
transform 1 0 26312 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_253
timestamp 1623621585
transform 1 0 24380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_258
timestamp 1623621585
transform 1 0 24840 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_266
timestamp 1623621585
transform 1 0 25576 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_270
timestamp 1623621585
transform 1 0 25944 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1998_
timestamp 1623621585
transform 1 0 27048 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_278
timestamp 1623621585
transform 1 0 26680 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_291
timestamp 1623621585
transform 1 0 27876 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1623621585
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_8
timestamp 1623621585
transform 1 0 1840 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1623621585
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1623621585
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1623621585
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1766_
timestamp 1623621585
transform 1 0 1564 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_21
timestamp 1623621585
transform 1 0 3036 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_22
timestamp 1623621585
transform 1 0 3128 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_18
timestamp 1623621585
transform 1 0 2760 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 2208 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _2105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1380 0 1 5984
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_7_30
timestamp 1623621585
transform 1 0 3864 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_30
timestamp 1623621585
transform 1 0 3864 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1623621585
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _1278_
timestamp 1623621585
transform 1 0 3220 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 1623621585
transform 1 0 4508 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_37
timestamp 1623621585
transform 1 0 4508 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input121
timestamp 1623621585
transform 1 0 4232 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input103
timestamp 1623621585
transform 1 0 4232 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_44
timestamp 1623621585
transform 1 0 5152 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_45
timestamp 1623621585
transform 1 0 5244 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input129
timestamp 1623621585
transform 1 0 4876 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_54
timestamp 1623621585
transform 1 0 6072 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_50
timestamp 1623621585
transform 1 0 5704 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_49
timestamp 1623621585
transform 1 0 5612 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input112
timestamp 1623621585
transform 1 0 5336 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1623621585
transform 1 0 6348 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1765_
timestamp 1623621585
transform 1 0 5796 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1623621585
transform 1 0 6440 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input138
timestamp 1623621585
transform 1 0 6808 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1989_
timestamp 1623621585
transform 1 0 6440 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_7_67
timestamp 1623621585
transform 1 0 7268 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1623621585
transform 1 0 7084 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1623621585
transform 1 0 9016 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input120
timestamp 1623621585
transform 1 0 8372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_77
timestamp 1623621585
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_82
timestamp 1623621585
transform 1 0 8648 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_90
timestamp 1623621585
transform 1 0 9384 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_79
timestamp 1623621585
transform 1 0 8372 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_85
timestamp 1623621585
transform 1 0 8924 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_87
timestamp 1623621585
transform 1 0 9108 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _1294_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 9660 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _1358_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 10488 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _1359_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 11040 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1623621585
transform 1 0 11592 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_98
timestamp 1623621585
transform 1 0 10120 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_108
timestamp 1623621585
transform 1 0 11040 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_99
timestamp 1623621585
transform 1 0 10212 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_107
timestamp 1623621585
transform 1 0 10948 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_113
timestamp 1623621585
transform 1 0 11500 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _1114_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 12696 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1623621585
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2220_
timestamp 1623621585
transform 1 0 12052 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_115
timestamp 1623621585
transform 1 0 11684 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1623621585
transform 1 0 13524 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_122
timestamp 1623621585
transform 1 0 12328 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_148
timestamp 1623621585
transform 1 0 14720 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_144
timestamp 1623621585
transform 1 0 14352 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_139
timestamp 1623621585
transform 1 0 13892 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_143
timestamp 1623621585
transform 1 0 14260 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1623621585
transform 1 0 14260 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1127_
timestamp 1623621585
transform 1 0 14628 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1115_
timestamp 1623621585
transform 1 0 13892 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_152
timestamp 1623621585
transform 1 0 15088 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1138_
timestamp 1623621585
transform 1 0 14812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_151
timestamp 1623621585
transform 1 0 14996 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1623621585
transform 1 0 16192 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_163
timestamp 1623621585
transform 1 0 16100 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1135_
timestamp 1623621585
transform 1 0 15824 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1104_
timestamp 1623621585
transform 1 0 16560 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1623621585
transform 1 0 17112 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_172
timestamp 1623621585
transform 1 0 16928 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1623621585
transform 1 0 16836 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1133_
timestamp 1623621585
transform 1 0 17296 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_182
timestamp 1623621585
transform 1 0 17848 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_179
timestamp 1623621585
transform 1 0 17572 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1122_
timestamp 1623621585
transform 1 0 17480 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1354_
timestamp 1623621585
transform 1 0 18676 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2188_
timestamp 1623621585
transform 1 0 19964 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1623621585
transform 1 0 19504 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1623621585
transform 1 0 18308 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1623621585
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1623621585
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_190
timestamp 1623621585
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_194
timestamp 1623621585
transform 1 0 18952 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_201
timestamp 1623621585
transform 1 0 19596 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2156_
timestamp 1623621585
transform 1 0 21988 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1623621585
transform 1 0 22080 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_214
timestamp 1623621585
transform 1 0 20792 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_226
timestamp 1623621585
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_221
timestamp 1623621585
transform 1 0 21436 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1869_
timestamp 1623621585
transform 1 0 24104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1623621585
transform 1 0 23828 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_229
timestamp 1623621585
transform 1 0 22172 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_241
timestamp 1623621585
transform 1 0 23276 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_250
timestamp 1623621585
transform 1 0 24104 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_243
timestamp 1623621585
transform 1 0 23460 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_249
timestamp 1623621585
transform 1 0 24012 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_258
timestamp 1623621585
transform 1 0 24840 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_253
timestamp 1623621585
transform 1 0 24380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_257
timestamp 1623621585
transform 1 0 24748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1623621585
transform 1 0 24472 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1623621585
transform 1 0 24748 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_266
timestamp 1623621585
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_265
timestamp 1623621585
transform 1 0 25484 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output240
timestamp 1623621585
transform 1 0 25116 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1656_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 25760 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_273
timestamp 1623621585
transform 1 0 26220 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output231
timestamp 1623621585
transform 1 0 25852 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_275
timestamp 1623621585
transform 1 0 26404 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_281
timestamp 1623621585
transform 1 0 26956 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output222
timestamp 1623621585
transform 1 0 26588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1623621585
transform 1 0 27324 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_295
timestamp 1623621585
transform 1 0 28244 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_295
timestamp 1623621585
transform 1 0 28244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_290
timestamp 1623621585
transform 1 0 27784 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_286
timestamp 1623621585
transform 1 0 27416 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output204
timestamp 1623621585
transform 1 0 27876 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2140_
timestamp 1623621585
transform 1 0 26772 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1623621585
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1623621585
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1220_
timestamp 1623621585
transform 1 0 2116 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1221_
timestamp 1623621585
transform 1 0 3128 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1699_
timestamp 1623621585
transform 1 0 1472 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1623621585
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1623621585
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1623621585
transform 1 0 1748 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_18
timestamp 1623621585
transform 1 0 2760 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2031_
timestamp 1623621585
transform 1 0 5152 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input130
timestamp 1623621585
transform 1 0 3772 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input148
timestamp 1623621585
transform 1 0 4416 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_25
timestamp 1623621585
transform 1 0 3404 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1623621585
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_39
timestamp 1623621585
transform 1 0 4692 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_43
timestamp 1623621585
transform 1 0 5060 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2197_
timestamp 1623621585
transform 1 0 7360 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1623621585
transform 1 0 6348 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_53
timestamp 1623621585
transform 1 0 5980 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_58
timestamp 1623621585
transform 1 0 6440 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_66
timestamp 1623621585
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1449_
timestamp 1623621585
transform 1 0 9200 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_84
timestamp 1623621585
transform 1 0 8832 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1767_
timestamp 1623621585
transform 1 0 10396 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1623621585
transform 1 0 11592 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_97
timestamp 1623621585
transform 1 0 10028 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_104
timestamp 1623621585
transform 1 0 10672 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_112
timestamp 1623621585
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 1623621585
transform 1 0 12236 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2049_
timestamp 1623621585
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_115
timestamp 1623621585
transform 1 0 11684 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_124
timestamp 1623621585
transform 1 0 12512 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_137
timestamp 1623621585
transform 1 0 13708 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _2267_
timestamp 1623621585
transform 1 0 14260 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__o211a_1  _1134_
timestamp 1623621585
transform 1 0 17296 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1623621585
transform 1 0 16836 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_160
timestamp 1623621585
transform 1 0 15824 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_168
timestamp 1623621585
transform 1 0 16560 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_172
timestamp 1623621585
transform 1 0 16928 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _2103_
timestamp 1623621585
transform 1 0 18492 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_8_184
timestamp 1623621585
transform 1 0 18032 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_188
timestamp 1623621585
transform 1 0 18400 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _1597_
timestamp 1623621585
transform 1 0 20608 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1623621585
transform 1 0 22080 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_207
timestamp 1623621585
transform 1 0 20148 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_211
timestamp 1623621585
transform 1 0 20516 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_219
timestamp 1623621585
transform 1 0 21252 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_227
timestamp 1623621585
transform 1 0 21988 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1808_
timestamp 1623621585
transform 1 0 23000 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _2101_
timestamp 1623621585
transform 1 0 23644 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_8_229
timestamp 1623621585
transform 1 0 22172 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_237
timestamp 1623621585
transform 1 0 22908 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_241
timestamp 1623621585
transform 1 0 23276 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1628_
timestamp 1623621585
transform 1 0 25668 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_263
timestamp 1623621585
transform 1 0 25300 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1623621585
transform 1 0 27324 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output178
timestamp 1623621585
transform 1 0 27876 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_276
timestamp 1623621585
transform 1 0 26496 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_284
timestamp 1623621585
transform 1 0 27232 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_286
timestamp 1623621585
transform 1 0 27416 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_290
timestamp 1623621585
transform 1 0 27784 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_295
timestamp 1623621585
transform 1 0 28244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1623621585
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1742_
timestamp 1623621585
transform 1 0 2208 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1803_
timestamp 1623621585
transform 1 0 1564 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1623621585
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1623621585
transform 1 0 2852 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1623621585
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1623621585
transform 1 0 1840 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1623621585
transform 1 0 2484 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_22
timestamp 1623621585
transform 1 0 3128 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2034_
timestamp 1623621585
transform 1 0 4968 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1623621585
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_28
timestamp 1623621585
transform 1 0 3680 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_30
timestamp 1623621585
transform 1 0 3864 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1988_
timestamp 1623621585
transform 1 0 6716 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1623621585
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1623621585
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1764_
timestamp 1623621585
transform 1 0 9476 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1623621585
transform 1 0 9016 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1623621585
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_82
timestamp 1623621585
transform 1 0 8648 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_87
timestamp 1623621585
transform 1 0 9108 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1768_
timestamp 1623621585
transform 1 0 11592 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2029_
timestamp 1623621585
transform 1 0 10396 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_94
timestamp 1623621585
transform 1 0 9752 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_100
timestamp 1623621585
transform 1 0 10304 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_110
timestamp 1623621585
transform 1 0 11224 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1816_
timestamp 1623621585
transform 1 0 13432 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_117
timestamp 1623621585
transform 1 0 11868 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_129
timestamp 1623621585
transform 1 0 12972 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_133
timestamp 1623621585
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1139_
timestamp 1623621585
transform 1 0 14720 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1623621585
transform 1 0 14260 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_138
timestamp 1623621585
transform 1 0 13800 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_142
timestamp 1623621585
transform 1 0 14168 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_144
timestamp 1623621585
transform 1 0 14352 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_156
timestamp 1623621585
transform 1 0 15456 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1952_
timestamp 1623621585
transform 1 0 15916 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _2269_
timestamp 1623621585
transform 1 0 17112 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_9_160
timestamp 1623621585
transform 1 0 15824 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_170
timestamp 1623621585
transform 1 0 16744 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1623621585
transform 1 0 19504 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_191
timestamp 1623621585
transform 1 0 18676 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_199
timestamp 1623621585
transform 1 0 19412 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_201
timestamp 1623621585
transform 1 0 19596 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1567_
timestamp 1623621585
transform 1 0 20516 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _2102_
timestamp 1623621585
transform 1 0 21160 0 1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_9_209
timestamp 1623621585
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_214
timestamp 1623621585
transform 1 0 20792 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _1512_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 23736 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_9_236
timestamp 1623621585
transform 1 0 22816 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_244
timestamp 1623621585
transform 1 0 23552 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2148_
timestamp 1623621585
transform 1 0 25300 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1623621585
transform 1 0 24748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_253
timestamp 1623621585
transform 1 0 24380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_258
timestamp 1623621585
transform 1 0 24840 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_262
timestamp 1623621585
transform 1 0 25208 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1657_
timestamp 1623621585
transform 1 0 27416 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_279
timestamp 1623621585
transform 1 0 26772 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_285
timestamp 1623621585
transform 1 0 27324 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_295
timestamp 1623621585
transform 1 0 28244 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1623621585
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1623621585
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1623621585
transform 1 0 1748 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 1623621585
transform 1 0 2392 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input140
timestamp 1623621585
transform 1 0 3036 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1623621585
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_10
timestamp 1623621585
transform 1 0 2024 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_17
timestamp 1623621585
transform 1 0 2668 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1738_
timestamp 1623621585
transform 1 0 4140 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2052_
timestamp 1623621585
transform 1 0 4784 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_24
timestamp 1623621585
transform 1 0 3312 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp 1623621585
transform 1 0 4048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_36
timestamp 1623621585
transform 1 0 4416 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1762_
timestamp 1623621585
transform 1 0 6808 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1623621585
transform 1 0 6348 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_49
timestamp 1623621585
transform 1 0 5612 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_58
timestamp 1623621585
transform 1 0 6440 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_65
timestamp 1623621585
transform 1 0 7084 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1763_
timestamp 1623621585
transform 1 0 7912 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2033_
timestamp 1623621585
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_73
timestamp 1623621585
transform 1 0 7820 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_77
timestamp 1623621585
transform 1 0 8188 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_90
timestamp 1623621585
transform 1 0 9384 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _2030_
timestamp 1623621585
transform 1 0 9844 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1623621585
transform 1 0 11592 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_94
timestamp 1623621585
transform 1 0 9752 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_104
timestamp 1623621585
transform 1 0 10672 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_112
timestamp 1623621585
transform 1 0 11408 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _2009_
timestamp 1623621585
transform 1 0 12052 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_115
timestamp 1623621585
transform 1 0 11684 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_128
timestamp 1623621585
transform 1 0 12880 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _2073_
timestamp 1623621585
transform 1 0 15640 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2076_
timestamp 1623621585
transform 1 0 14444 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_140
timestamp 1623621585
transform 1 0 13984 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_144
timestamp 1623621585
transform 1 0 14352 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1623621585
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _2004_
timestamp 1623621585
transform 1 0 17296 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1623621585
transform 1 0 16836 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_167
timestamp 1623621585
transform 1 0 16468 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_172
timestamp 1623621585
transform 1 0 16928 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1757_
timestamp 1623621585
transform 1 0 18676 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1804_
timestamp 1623621585
transform 1 0 19320 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_185
timestamp 1623621585
transform 1 0 18124 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_194
timestamp 1623621585
transform 1 0 18952 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_201
timestamp 1623621585
transform 1 0 19596 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1578_
timestamp 1623621585
transform 1 0 20608 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1623621585
transform 1 0 22080 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_209
timestamp 1623621585
transform 1 0 20332 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_216
timestamp 1623621585
transform 1 0 20976 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1598_
timestamp 1623621585
transform 1 0 22540 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1627_
timestamp 1623621585
transform 1 0 23736 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_10_229
timestamp 1623621585
transform 1 0 22172 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_242
timestamp 1623621585
transform 1 0 23368 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1629_
timestamp 1623621585
transform 1 0 25208 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output232
timestamp 1623621585
transform 1 0 25852 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_253
timestamp 1623621585
transform 1 0 24380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_261
timestamp 1623621585
transform 1 0 25116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_265
timestamp 1623621585
transform 1 0 25484 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_273
timestamp 1623621585
transform 1 0 26220 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1623621585
transform 1 0 27324 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output187
timestamp 1623621585
transform 1 0 27876 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output196
timestamp 1623621585
transform 1 0 26588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_281
timestamp 1623621585
transform 1 0 26956 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_286
timestamp 1623621585
transform 1 0 27416 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_290
timestamp 1623621585
transform 1 0 27784 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_295
timestamp 1623621585
transform 1 0 28244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1623621585
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1623621585
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1623621585
transform 1 0 1748 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input122
timestamp 1623621585
transform 1 0 2392 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1623621585
transform 1 0 3036 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1623621585
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_10
timestamp 1623621585
transform 1 0 2024 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_17
timestamp 1623621585
transform 1 0 2668 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2229_
timestamp 1623621585
transform 1 0 4232 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1623621585
transform 1 0 3772 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1623621585
transform 1 0 3312 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_28
timestamp 1623621585
transform 1 0 3680 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1623621585
transform 1 0 3864 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_51
timestamp 1623621585
transform 1 0 5796 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_63
timestamp 1623621585
transform 1 0 6900 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _2032_
timestamp 1623621585
transform 1 0 9476 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1623621585
transform 1 0 9016 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_75
timestamp 1623621585
transform 1 0 8004 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_83
timestamp 1623621585
transform 1 0 8740 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_87
timestamp 1623621585
transform 1 0 9108 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_100
timestamp 1623621585
transform 1 0 10304 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_112
timestamp 1623621585
transform 1 0 11408 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1741_
timestamp 1623621585
transform 1 0 13248 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2010_
timestamp 1623621585
transform 1 0 11684 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_124
timestamp 1623621585
transform 1 0 12512 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_135
timestamp 1623621585
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1694_
timestamp 1623621585
transform 1 0 14720 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1623621585
transform 1 0 14260 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_144
timestamp 1623621585
transform 1 0 14352 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_151
timestamp 1623621585
transform 1 0 14996 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_159
timestamp 1623621585
transform 1 0 15732 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _1953_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 15824 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_172
timestamp 1623621585
transform 1 0 16928 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1623621585
transform 1 0 19504 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1623621585
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_196
timestamp 1623621585
transform 1 0 19136 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_201
timestamp 1623621585
transform 1 0 19596 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_213
timestamp 1623621585
transform 1 0 20700 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1623621585
transform 1 0 21804 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1632_
timestamp 1623621585
transform 1 0 24104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1623621585
transform 1 0 22908 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_249
timestamp 1623621585
transform 1 0 24012 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _1653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 26312 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1623621585
transform 1 0 24748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output214
timestamp 1623621585
transform 1 0 25576 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_253
timestamp 1623621585
transform 1 0 24380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_258
timestamp 1623621585
transform 1 0 24840 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_270
timestamp 1623621585
transform 1 0 25944 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1655_
timestamp 1623621585
transform 1 0 27508 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_282
timestamp 1623621585
transform 1 0 27048 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_286
timestamp 1623621585
transform 1 0 27416 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_295
timestamp 1623621585
transform 1 0 28244 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1623621585
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _1284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 3128 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1754_
timestamp 1623621585
transform 1 0 2484 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1623621585
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input149
timestamp 1623621585
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1623621585
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1623621585
transform 1 0 2116 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_18
timestamp 1623621585
transform 1 0 2760 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1658_
timestamp 1623621585
transform 1 0 4232 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_27
timestamp 1623621585
transform 1 0 3588 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_33
timestamp 1623621585
transform 1 0 4140 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_37
timestamp 1623621585
transform 1 0 4508 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1349_
timestamp 1623621585
transform 1 0 6808 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1623621585
transform 1 0 6348 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_49
timestamp 1623621585
transform 1 0 5612 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1623621585
transform 1 0 6440 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1991_
timestamp 1623621585
transform 1 0 8372 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_71
timestamp 1623621585
transform 1 0 7636 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1623621585
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1747_
timestamp 1623621585
transform 1 0 9568 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1990_
timestamp 1623621585
transform 1 0 10396 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1623621585
transform 1 0 11592 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_96
timestamp 1623621585
transform 1 0 9936 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_100
timestamp 1623621585
transform 1 0 10304 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1623621585
transform 1 0 11224 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1695_
timestamp 1623621585
transform 1 0 12052 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1769_
timestamp 1623621585
transform 1 0 12696 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _1971_
timestamp 1623621585
transform 1 0 13340 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_115
timestamp 1623621585
transform 1 0 11684 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_122
timestamp 1623621585
transform 1 0 12328 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_129
timestamp 1623621585
transform 1 0 12972 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1970_
timestamp 1623621585
transform 1 0 14812 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_145
timestamp 1623621585
transform 1 0 14444 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_158
timestamp 1623621585
transform 1 0 15640 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1698_
timestamp 1623621585
transform 1 0 16008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1623621585
transform 1 0 16836 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_165
timestamp 1623621585
transform 1 0 16284 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_172
timestamp 1623621585
transform 1 0 16928 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_184
timestamp 1623621585
transform 1 0 18032 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_196
timestamp 1623621585
transform 1 0 19136 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1568_
timestamp 1623621585
transform 1 0 20424 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1623621585
transform 1 0 22080 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_208
timestamp 1623621585
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_213
timestamp 1623621585
transform 1 0 20700 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_225
timestamp 1623621585
transform 1 0 21804 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1602_
timestamp 1623621585
transform 1 0 23276 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1659_
timestamp 1623621585
transform 1 0 22540 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output241
timestamp 1623621585
transform 1 0 23920 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_229
timestamp 1623621585
transform 1 0 22172 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_236
timestamp 1623621585
transform 1 0 22816 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_240
timestamp 1623621585
transform 1 0 23184 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_244
timestamp 1623621585
transform 1 0 23552 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1996_
timestamp 1623621585
transform 1 0 25392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output223
timestamp 1623621585
transform 1 0 24656 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_252
timestamp 1623621585
transform 1 0 24288 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_260
timestamp 1623621585
transform 1 0 25024 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_273
timestamp 1623621585
transform 1 0 26220 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 26588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1623621585
transform 1 0 27324 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output205
timestamp 1623621585
transform 1 0 27876 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_281
timestamp 1623621585
transform 1 0 26956 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_286
timestamp 1623621585
transform 1 0 27416 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_290
timestamp 1623621585
transform 1 0 27784 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_295
timestamp 1623621585
transform 1 0 28244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1623621585
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1226_
timestamp 1623621585
transform 1 0 2024 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _1228_
timestamp 1623621585
transform 1 0 2852 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__mux4_2  _2106_
timestamp 1623621585
transform 1 0 1380 0 1 9248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1623621585
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1623621585
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1623621585
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_21
timestamp 1623621585
transform 1 0 3036 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_6
timestamp 1623621585
transform 1 0 1656 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 1623621585
transform 1 0 2484 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2ai_1  _1286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 4232 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _1973_
timestamp 1623621585
transform 1 0 4784 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1623621585
transform 1 0 3772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_30
timestamp 1623621585
transform 1 0 3864 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_41
timestamp 1623621585
transform 1 0 4876 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_32
timestamp 1623621585
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1347_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 6900 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2223_
timestamp 1623621585
transform 1 0 5612 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1623621585
transform 1 0 6348 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_66
timestamp 1623621585
transform 1 0 7176 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_52
timestamp 1623621585
transform 1 0 5888 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_56
timestamp 1623621585
transform 1 0 6256 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1623621585
transform 1 0 6440 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_62
timestamp 1623621585
transform 1 0 6808 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_67
timestamp 1623621585
transform 1 0 7268 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_77
timestamp 1623621585
transform 1 0 8188 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_77
timestamp 1623621585
transform 1 0 8188 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1348_
timestamp 1623621585
transform 1 0 7544 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1346_
timestamp 1623621585
transform 1 0 7636 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1623621585
transform 1 0 8924 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_85
timestamp 1623621585
transform 1 0 8924 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1623621585
transform 1 0 9016 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1760_
timestamp 1623621585
transform 1 0 9016 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_89
timestamp 1623621585
transform 1 0 9292 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_87
timestamp 1623621585
transform 1 0 9108 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1954_
timestamp 1623621585
transform 1 0 11132 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1623621585
transform 1 0 11592 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_99
timestamp 1623621585
transform 1 0 10212 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_107
timestamp 1623621585
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_101
timestamp 1623621585
transform 1 0 10396 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_113
timestamp 1623621585
transform 1 0 11500 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1151_
timestamp 1623621585
transform 1 0 12328 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2262_
timestamp 1623621585
transform 1 0 12420 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1623621585
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1623621585
transform 1 0 12604 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_137
timestamp 1623621585
transform 1 0 13708 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_115
timestamp 1623621585
transform 1 0 11684 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_4  _1955_
timestamp 1623621585
transform 1 0 14720 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1623621585
transform 1 0 14260 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_144
timestamp 1623621585
transform 1 0 14352 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_139
timestamp 1623621585
transform 1 0 13892 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_151
timestamp 1623621585
transform 1 0 14996 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_1  _1554_
timestamp 1623621585
transform 1 0 17296 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2172_
timestamp 1623621585
transform 1 0 17296 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1623621585
transform 1 0 16836 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_160
timestamp 1623621585
transform 1 0 15824 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_172
timestamp 1623621585
transform 1 0 16928 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_163
timestamp 1623621585
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_172
timestamp 1623621585
transform 1 0 16928 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _2126_
timestamp 1623621585
transform 1 0 18400 0 -1 10336
box -38 -48 1694 592
use sky130_fd_sc_hd__dfxtp_1  _2173_
timestamp 1623621585
transform 1 0 19964 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1623621585
transform 1 0 19504 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_192
timestamp 1623621585
transform 1 0 18768 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_201
timestamp 1623621585
transform 1 0 19596 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_183
timestamp 1623621585
transform 1 0 17940 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_187
timestamp 1623621585
transform 1 0 18308 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1550_
timestamp 1623621585
transform 1 0 21804 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  _1569_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 20424 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1623621585
transform 1 0 22080 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_221
timestamp 1623621585
transform 1 0 21436 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_228
timestamp 1623621585
transform 1 0 22080 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_206
timestamp 1623621585
transform 1 0 20056 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_218
timestamp 1623621585
transform 1 0 21160 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_226
timestamp 1623621585
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1507_
timestamp 1623621585
transform 1 0 22724 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_4  _1603_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 23552 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _1994_
timestamp 1623621585
transform 1 0 22908 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_236
timestamp 1623621585
transform 1 0 22816 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_246
timestamp 1623621585
transform 1 0 23736 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_229
timestamp 1623621585
transform 1 0 22172 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_238
timestamp 1623621585
transform 1 0 23000 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1995_
timestamp 1623621585
transform 1 0 25300 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2149_
timestamp 1623621585
transform 1 0 25392 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1623621585
transform 1 0 24748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_254
timestamp 1623621585
transform 1 0 24472 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_258
timestamp 1623621585
transform 1 0 24840 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_262
timestamp 1623621585
transform 1 0 25208 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_272
timestamp 1623621585
transform 1 0 26128 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_260
timestamp 1623621585
transform 1 0 25024 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1630_
timestamp 1623621585
transform 1 0 27876 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_4  _1633_
timestamp 1623621585
transform 1 0 26496 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1623621585
transform 1 0 27324 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_292
timestamp 1623621585
transform 1 0 27968 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_280
timestamp 1623621585
transform 1 0 26864 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_284
timestamp 1623621585
transform 1 0 27232 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_286
timestamp 1623621585
transform 1 0 27416 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_290
timestamp 1623621585
transform 1 0 27784 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_295
timestamp 1623621585
transform 1 0 28244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1623621585
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1623621585
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_298
timestamp 1623621585
transform 1 0 28520 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 1623621585
transform 1 0 1932 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1227_
timestamp 1623621585
transform 1 0 2576 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1623621585
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1623621585
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_12
timestamp 1623621585
transform 1 0 2208 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_22
timestamp 1623621585
transform 1 0 3128 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1972_
timestamp 1623621585
transform 1 0 4784 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1623621585
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_28
timestamp 1623621585
transform 1 0 3680 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_30
timestamp 1623621585
transform 1 0 3864 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_38
timestamp 1623621585
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_49
timestamp 1623621585
transform 1 0 5612 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_61
timestamp 1623621585
transform 1 0 6716 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2198_
timestamp 1623621585
transform 1 0 9476 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1623621585
transform 1 0 9016 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_73
timestamp 1623621585
transform 1 0 7820 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_85
timestamp 1623621585
transform 1 0 8924 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_87
timestamp 1623621585
transform 1 0 9108 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_wb_clk_i
timestamp 1623621585
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1623621585
transform 1 0 10948 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_114
timestamp 1623621585
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1152_
timestamp 1623621585
transform 1 0 12512 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_122
timestamp 1623621585
transform 1 0 12328 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_132
timestamp 1623621585
transform 1 0 13248 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_2  _2104_
timestamp 1623621585
transform 1 0 14904 0 1 10336
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1623621585
transform 1 0 14260 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_140
timestamp 1623621585
transform 1 0 13984 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_144
timestamp 1623621585
transform 1 0 14352 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _2119_
timestamp 1623621585
transform 1 0 16928 0 1 10336
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_15_168
timestamp 1623621585
transform 1 0 16560 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1623621585
transform 1 0 19504 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_190
timestamp 1623621585
transform 1 0 18584 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_198
timestamp 1623621585
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_201
timestamp 1623621585
transform 1 0 19596 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux4_2  _2133_
timestamp 1623621585
transform 1 0 21252 0 1 10336
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_15_213
timestamp 1623621585
transform 1 0 20700 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1611_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 23552 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_237
timestamp 1623621585
transform 1 0 22908 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_243
timestamp 1623621585
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_1  _1625_
timestamp 1623621585
transform 1 0 25208 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1872_
timestamp 1623621585
transform 1 0 26128 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1623621585
transform 1 0 24748 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_252
timestamp 1623621585
transform 1 0 24288 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_256
timestamp 1623621585
transform 1 0 24656 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_258
timestamp 1623621585
transform 1 0 24840 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_268
timestamp 1623621585
transform 1 0 25760 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2141_
timestamp 1623621585
transform 1 0 26772 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1623621585
transform 1 0 26404 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_295
timestamp 1623621585
transform 1 0 28244 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1623621585
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 3036 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1623621585
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1623621585
transform 1 0 1748 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1623621585
transform 1 0 2392 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1623621585
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_10
timestamp 1623621585
transform 1 0 2024 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_17
timestamp 1623621585
transform 1 0 2668 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1282_
timestamp 1623621585
transform 1 0 3956 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1285_
timestamp 1623621585
transform 1 0 4968 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1623621585
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_34
timestamp 1623621585
transform 1 0 4232 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_45
timestamp 1623621585
transform 1 0 5244 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_4  _1301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 7084 0 -1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1623621585
transform 1 0 6348 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_58
timestamp 1623621585
transform 1 0 6440 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_64
timestamp 1623621585
transform 1 0 6992 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1448_
timestamp 1623621585
transform 1 0 9476 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1623621585
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1690_
timestamp 1623621585
transform 1 0 10672 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1623621585
transform 1 0 11592 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_100
timestamp 1623621585
transform 1 0 10304 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_107
timestamp 1623621585
transform 1 0 10948 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_113
timestamp 1623621585
transform 1 0 11500 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1143_
timestamp 1623621585
transform 1 0 13524 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2079_
timestamp 1623621585
transform 1 0 12052 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_115
timestamp 1623621585
transform 1 0 11684 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_128
timestamp 1623621585
transform 1 0 12880 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_134
timestamp 1623621585
transform 1 0 13432 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_139
timestamp 1623621585
transform 1 0 13892 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_151
timestamp 1623621585
transform 1 0 14996 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1555_
timestamp 1623621585
transform 1 0 17664 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1623621585
transform 1 0 16836 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_163
timestamp 1623621585
transform 1 0 16100 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_172
timestamp 1623621585
transform 1 0 16928 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1526_
timestamp 1623621585
transform 1 0 19596 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1553_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 18860 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_189
timestamp 1623621585
transform 1 0 18492 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1623621585
transform 1 0 19228 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_204
timestamp 1623621585
transform 1 0 19872 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1623621585
transform 1 0 22080 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_wb_clk_i
timestamp 1623621585
transform 1 0 20240 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_211
timestamp 1623621585
transform 1 0 20516 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_223
timestamp 1623621585
transform 1 0 21620 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_227
timestamp 1623621585
transform 1 0 21988 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _1624_
timestamp 1623621585
transform 1 0 23552 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_229
timestamp 1623621585
transform 1 0 22172 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_241
timestamp 1623621585
transform 1 0 23276 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1626_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 24656 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output206
timestamp 1623621585
transform 1 0 25852 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_252
timestamp 1623621585
transform 1 0 24288 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_263
timestamp 1623621585
transform 1 0 25300 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_273
timestamp 1623621585
transform 1 0 26220 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1623621585
transform 1 0 27324 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output179
timestamp 1623621585
transform 1 0 27876 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output188
timestamp 1623621585
transform 1 0 26588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_281
timestamp 1623621585
transform 1 0 26956 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_286
timestamp 1623621585
transform 1 0 27416 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_290
timestamp 1623621585
transform 1 0 27784 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_295
timestamp 1623621585
transform 1 0 28244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1623621585
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1623621585
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1623621585
transform 1 0 1748 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input123
timestamp 1623621585
transform 1 0 2392 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1623621585
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_10
timestamp 1623621585
transform 1 0 2024 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_17
timestamp 1623621585
transform 1 0 2668 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux4_2  _2113_
timestamp 1623621585
transform 1 0 4324 0 1 11424
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1623621585
transform 1 0 3772 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_30
timestamp 1623621585
transform 1 0 3864 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_34
timestamp 1623621585
transform 1 0 4232 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _2055_
timestamp 1623621585
transform 1 0 6348 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_53
timestamp 1623621585
transform 1 0 5980 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_66
timestamp 1623621585
transform 1 0 7176 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1304_
timestamp 1623621585
transform 1 0 7544 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1447_
timestamp 1623621585
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1623621585
transform 1 0 9016 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_74
timestamp 1623621585
transform 1 0 7912 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_78
timestamp 1623621585
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1623621585
transform 1 0 8648 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_87
timestamp 1623621585
transform 1 0 9108 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_91
timestamp 1623621585
transform 1 0 9476 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1956_
timestamp 1623621585
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2035_
timestamp 1623621585
transform 1 0 9568 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_101
timestamp 1623621585
transform 1 0 10396 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_114
timestamp 1623621585
transform 1 0 11592 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1153_
timestamp 1623621585
transform 1 0 12236 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1688_
timestamp 1623621585
transform 1 0 12880 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_wb_clk_i
timestamp 1623621585
transform 1 0 13524 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_120
timestamp 1623621585
transform 1 0 12144 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_124
timestamp 1623621585
transform 1 0 12512 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_131
timestamp 1623621585
transform 1 0 13156 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1623621585
transform 1 0 14260 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_wb_clk_i
timestamp 1623621585
transform 1 0 14720 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_138
timestamp 1623621585
transform 1 0 13800 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_142
timestamp 1623621585
transform 1 0 14168 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1623621585
transform 1 0 14352 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_151
timestamp 1623621585
transform 1 0 14996 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_163
timestamp 1623621585
transform 1 0 16100 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_175
timestamp 1623621585
transform 1 0 17204 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1623621585
transform 1 0 19504 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_187
timestamp 1623621585
transform 1 0 18308 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_199
timestamp 1623621585
transform 1 0 19412 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_201
timestamp 1623621585
transform 1 0 19596 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1594_
timestamp 1623621585
transform 1 0 20516 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2157_
timestamp 1623621585
transform 1 0 21436 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_209
timestamp 1623621585
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_217
timestamp 1623621585
transform 1 0 21068 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1595_
timestamp 1623621585
transform 1 0 23276 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_237
timestamp 1623621585
transform 1 0 22908 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_247
timestamp 1623621585
transform 1 0 23828 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1623621585
transform 1 0 24748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output215
timestamp 1623621585
transform 1 0 26036 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output233
timestamp 1623621585
transform 1 0 25300 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_255
timestamp 1623621585
transform 1 0 24564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_258
timestamp 1623621585
transform 1 0 24840 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_262
timestamp 1623621585
transform 1 0 25208 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_267
timestamp 1623621585
transform 1 0 25668 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2142_
timestamp 1623621585
transform 1 0 26772 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 1623621585
transform 1 0 26404 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_295
timestamp 1623621585
transform 1 0 28244 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1623621585
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _2107_
timestamp 1623621585
transform 1 0 1380 0 -1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1623621585
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_21
timestamp 1623621585
transform 1 0 3036 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_4  _1232_
timestamp 1623621585
transform 1 0 3404 0 -1 12512
box -38 -48 1418 592
use sky130_fd_sc_hd__decap_8  FILLER_18_40
timestamp 1623621585
transform 1 0 4784 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1306_
timestamp 1623621585
transform 1 0 7176 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1732_
timestamp 1623621585
transform 1 0 5704 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1623621585
transform 1 0 6348 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1623621585
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_53
timestamp 1623621585
transform 1 0 5980 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_58
timestamp 1623621585
transform 1 0 6440 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _2036_
timestamp 1623621585
transform 1 0 8832 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_73
timestamp 1623621585
transform 1 0 7820 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 1623621585
transform 1 0 8556 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1689_
timestamp 1623621585
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1761_
timestamp 1623621585
transform 1 0 10212 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1623621585
transform 1 0 11592 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_93
timestamp 1623621585
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_102
timestamp 1623621585
transform 1 0 10488 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_106
timestamp 1623621585
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_110
timestamp 1623621585
transform 1 0 11224 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1150_
timestamp 1623621585
transform 1 0 12328 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_115
timestamp 1623621585
transform 1 0 11684 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 1623621585
transform 1 0 12236 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_130
timestamp 1623621585
transform 1 0 13064 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1145_
timestamp 1623621585
transform 1 0 13800 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_4  _2006_
timestamp 1623621585
transform 1 0 14996 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_146
timestamp 1623621585
transform 1 0 14536 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_150
timestamp 1623621585
transform 1 0 14904 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1623621585
transform 1 0 16836 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_163
timestamp 1623621585
transform 1 0 16100 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_172
timestamp 1623621585
transform 1 0 16928 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux4_2  _2127_
timestamp 1623621585
transform 1 0 18952 0 -1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_18_184
timestamp 1623621585
transform 1 0 18032 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_192
timestamp 1623621585
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__a31o_1  _1596_
timestamp 1623621585
transform 1 0 20976 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1623621585
transform 1 0 22080 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_212
timestamp 1623621585
transform 1 0 20608 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_223
timestamp 1623621585
transform 1 0 21620 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_227
timestamp 1623621585
transform 1 0 21988 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _1622_
timestamp 1623621585
transform 1 0 23920 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_wb_clk_i
timestamp 1623621585
transform 1 0 22540 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_229
timestamp 1623621585
transform 1 0 22172 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_236
timestamp 1623621585
transform 1 0 22816 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1623_
timestamp 1623621585
transform 1 0 24932 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1651_
timestamp 1623621585
transform 1 0 26312 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_18_255
timestamp 1623621585
transform 1 0 24564 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_268
timestamp 1623621585
transform 1 0 25760 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1623621585
transform 1 0 27324 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output197
timestamp 1623621585
transform 1 0 27876 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_281
timestamp 1623621585
transform 1 0 26956 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_286
timestamp 1623621585
transform 1 0 27416 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_290
timestamp 1623621585
transform 1 0 27784 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_295
timestamp 1623621585
transform 1 0 28244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1623621585
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1623621585
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1623621585
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input150
timestamp 1623621585
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input141
timestamp 1623621585
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1623621585
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1623621585
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_15
timestamp 1623621585
transform 1 0 2484 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_11
timestamp 1623621585
transform 1 0 2116 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_11
timestamp 1623621585
transform 1 0 2116 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input132
timestamp 1623621585
transform 1 0 2484 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1230_
timestamp 1623621585
transform 1 0 2576 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_19
timestamp 1623621585
transform 1 0 2852 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_18
timestamp 1623621585
transform 1 0 2760 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1623621585
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_26
timestamp 1623621585
transform 1 0 3496 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_30
timestamp 1623621585
transform 1 0 3864 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_26
timestamp 1623621585
transform 1 0 3496 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1623621585
transform 1 0 3220 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1623621585
transform 1 0 3772 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 1623621585
transform 1 0 3956 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_38
timestamp 1623621585
transform 1 0 4600 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_34
timestamp 1623621585
transform 1 0 4232 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_41
timestamp 1623621585
transform 1 0 4876 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_37
timestamp 1623621585
transform 1 0 4508 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1974_
timestamp 1623621585
transform 1 0 4692 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1734_
timestamp 1623621585
transform 1 0 4232 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1733_
timestamp 1623621585
transform 1 0 4968 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_45
timestamp 1623621585
transform 1 0 5244 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_4  _1321_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 7084 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_4  _1975_
timestamp 1623621585
transform 1 0 5612 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1623621585
transform 1 0 6348 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_61
timestamp 1623621585
transform 1 0 6716 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_48
timestamp 1623621585
transform 1 0 5520 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_56
timestamp 1623621585
transform 1 0 6256 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_58
timestamp 1623621585
transform 1 0 6440 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_66
timestamp 1623621585
transform 1 0 7176 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_2  _1305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 7452 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1758_
timestamp 1623621585
transform 1 0 8924 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1623621585
transform 1 0 9016 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1623621585
transform 1 0 8648 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_87
timestamp 1623621585
transform 1 0 9108 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_81
timestamp 1623621585
transform 1 0 8556 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_88
timestamp 1623621585
transform 1 0 9200 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1684_
timestamp 1623621585
transform 1 0 10396 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_8  _1957_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 10948 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1623621585
transform 1 0 11592 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_99
timestamp 1623621585
transform 1 0 10212 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_100
timestamp 1623621585
transform 1 0 10304 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_104
timestamp 1623621585
transform 1 0 10672 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_112
timestamp 1623621585
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _1144_
timestamp 1623621585
transform 1 0 13616 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2263_
timestamp 1623621585
transform 1 0 12144 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_19_128
timestamp 1623621585
transform 1 0 12880 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_115
timestamp 1623621585
transform 1 0 11684 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_119
timestamp 1623621585
transform 1 0 12052 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1623621585
transform 1 0 13616 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _2120_
timestamp 1623621585
transform 1 0 15272 0 1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__dfxtp_1  _2265_
timestamp 1623621585
transform 1 0 14076 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1623621585
transform 1 0 14260 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_139
timestamp 1623621585
transform 1 0 13892 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_144
timestamp 1623621585
transform 1 0 14352 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1623621585
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_140
timestamp 1623621585
transform 1 0 13984 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_157
timestamp 1623621585
transform 1 0 15548 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_2  _1547_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 17296 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1548_
timestamp 1623621585
transform 1 0 17572 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1551_
timestamp 1623621585
transform 1 0 15916 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1623621585
transform 1 0 16836 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_172
timestamp 1623621585
transform 1 0 16928 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_167
timestamp 1623621585
transform 1 0 16468 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_172
timestamp 1623621585
transform 1 0 16928 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_178
timestamp 1623621585
transform 1 0 17480 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _1552_
timestamp 1623621585
transform 1 0 18492 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2174_
timestamp 1623621585
transform 1 0 18584 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1623621585
transform 1 0 19504 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_185
timestamp 1623621585
transform 1 0 18124 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_193
timestamp 1623621585
transform 1 0 18860 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_199
timestamp 1623621585
transform 1 0 19412 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_201
timestamp 1623621585
transform 1 0 19596 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_186
timestamp 1623621585
transform 1 0 18216 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_212
timestamp 1623621585
transform 1 0 20608 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_206
timestamp 1623621585
transform 1 0 20056 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_213
timestamp 1623621585
transform 1 0 20700 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _1591_
timestamp 1623621585
transform 1 0 20700 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_20_218
timestamp 1623621585
transform 1 0 21160 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_221
timestamp 1623621585
transform 1 0 21436 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_wb_clk_i
timestamp 1623621585
transform 1 0 21528 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_226
timestamp 1623621585
transform 1 0 21896 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_225
timestamp 1623621585
transform 1 0 21804 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1623621585
transform 1 0 22080 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_2  _1604_
timestamp 1623621585
transform 1 0 23736 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _2134_
timestamp 1623621585
transform 1 0 22356 0 1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_19_249
timestamp 1623621585
transform 1 0 24012 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_229
timestamp 1623621585
transform 1 0 22172 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_241
timestamp 1623621585
transform 1 0 23276 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_245
timestamp 1623621585
transform 1 0 23644 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_2  _2100_
timestamp 1623621585
transform 1 0 25208 0 1 12512
box -38 -48 1694 592
use sky130_fd_sc_hd__dfxtp_1  _2150_
timestamp 1623621585
transform 1 0 24932 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1623621585
transform 1 0 24748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_258
timestamp 1623621585
transform 1 0 24840 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_255
timestamp 1623621585
transform 1 0 24564 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_283
timestamp 1623621585
transform 1 0 27140 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_275
timestamp 1623621585
transform 1 0 26404 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_280
timestamp 1623621585
transform 1 0 26864 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_290
timestamp 1623621585
transform 1 0 27784 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_286
timestamp 1623621585
transform 1 0 27416 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output180
timestamp 1623621585
transform 1 0 27876 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1623621585
transform 1 0 27324 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1652_
timestamp 1623621585
transform 1 0 27416 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_295
timestamp 1623621585
transform 1 0 28244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1623621585
transform 1 0 28244 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1623621585
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1623621585
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _1231_
timestamp 1623621585
transform 1 0 1840 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1623621585
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1623621585
transform 1 0 2852 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1623621585
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1623621585
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_15
timestamp 1623621585
transform 1 0 2484 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_22
timestamp 1623621585
transform 1 0 3128 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2ai_1  _1292_
timestamp 1623621585
transform 1 0 4232 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1623621585
transform 1 0 3772 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_28
timestamp 1623621585
transform 1 0 3680 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_30
timestamp 1623621585
transform 1 0 3864 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_41
timestamp 1623621585
transform 1 0 4876 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_4  _1302_
timestamp 1623621585
transform 1 0 6624 0 1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_6  FILLER_21_53
timestamp 1623621585
transform 1 0 5980 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_59
timestamp 1623621585
transform 1 0 6532 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _2038_
timestamp 1623621585
transform 1 0 9476 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1623621585
transform 1 0 9016 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_82
timestamp 1623621585
transform 1 0 8648 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_87
timestamp 1623621585
transform 1 0 9108 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2082_
timestamp 1623621585
transform 1 0 10948 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_103
timestamp 1623621585
transform 1 0 10580 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1149_
timestamp 1623621585
transform 1 0 12144 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_116
timestamp 1623621585
transform 1 0 11776 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1623621585
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_135
timestamp 1623621585
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1623621585
transform 1 0 14260 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_144
timestamp 1623621585
transform 1 0 14352 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_156
timestamp 1623621585
transform 1 0 15456 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _1529_
timestamp 1623621585
transform 1 0 16652 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1538_
timestamp 1623621585
transform 1 0 17572 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_168
timestamp 1623621585
transform 1 0 16560 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_175
timestamp 1623621585
transform 1 0 17204 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_182
timestamp 1623621585
transform 1 0 17848 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1549_
timestamp 1623621585
transform 1 0 18308 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1623621585
transform 1 0 19504 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_186
timestamp 1623621585
transform 1 0 18216 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_196
timestamp 1623621585
transform 1 0 19136 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_201
timestamp 1623621585
transform 1 0 19596 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1588_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 20516 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_209
timestamp 1623621585
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_219
timestamp 1623621585
transform 1 0 21252 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2158_
timestamp 1623621585
transform 1 0 22356 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_21_247
timestamp 1623621585
transform 1 0 23828 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1623621585
transform 1 0 24748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output242
timestamp 1623621585
transform 1 0 25668 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_255
timestamp 1623621585
transform 1 0 24564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_258
timestamp 1623621585
transform 1 0 24840 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_266
timestamp 1623621585
transform 1 0 25576 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_271
timestamp 1623621585
transform 1 0 26036 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output189
timestamp 1623621585
transform 1 0 27876 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output216
timestamp 1623621585
transform 1 0 27140 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output224
timestamp 1623621585
transform 1 0 26404 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_279
timestamp 1623621585
transform 1 0 26772 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_287
timestamp 1623621585
transform 1 0 27508 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_295
timestamp 1623621585
transform 1 0 28244 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1623621585
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1623621585
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1623621585
transform 1 0 1748 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1623621585
transform 1 0 2392 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1623621585
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_10
timestamp 1623621585
transform 1 0 2024 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_17
timestamp 1623621585
transform 1 0 2668 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 3312 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _1289_
timestamp 1623621585
transform 1 0 4876 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_23
timestamp 1623621585
transform 1 0 3220 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_37
timestamp 1623621585
transform 1 0 4508 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1623621585
transform 1 0 6348 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_47
timestamp 1623621585
transform 1 0 5428 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_55
timestamp 1623621585
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_58
timestamp 1623621585
transform 1 0 6440 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_66
timestamp 1623621585
transform 1 0 7176 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1303_
timestamp 1623621585
transform 1 0 7452 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1759_
timestamp 1623621585
transform 1 0 9016 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_72
timestamp 1623621585
transform 1 0 7728 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1623621585
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_89
timestamp 1623621585
transform 1 0 9292 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1682_
timestamp 1623621585
transform 1 0 10856 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2037_
timestamp 1623621585
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1623621585
transform 1 0 11592 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1623621585
transform 1 0 10488 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_109
timestamp 1623621585
transform 1 0 11132 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_113
timestamp 1623621585
transform 1 0 11500 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1146_
timestamp 1623621585
transform 1 0 13340 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2012_
timestamp 1623621585
transform 1 0 12052 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_115
timestamp 1623621585
transform 1 0 11684 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_128
timestamp 1623621585
transform 1 0 12880 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_132
timestamp 1623621585
transform 1 0 13248 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_136
timestamp 1623621585
transform 1 0 13616 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_148
timestamp 1623621585
transform 1 0 14720 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _1539_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 17296 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1623621585
transform 1 0 16836 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_160
timestamp 1623621585
transform 1 0 15824 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_168
timestamp 1623621585
transform 1 0 16560 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_172
timestamp 1623621585
transform 1 0 16928 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_183
timestamp 1623621585
transform 1 0 17940 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_195
timestamp 1623621585
transform 1 0 19044 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _1579_
timestamp 1623621585
transform 1 0 20792 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1623621585
transform 1 0 22080 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_207
timestamp 1623621585
transform 1 0 20148 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_213
timestamp 1623621585
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_221
timestamp 1623621585
transform 1 0 21436 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_227
timestamp 1623621585
transform 1 0 21988 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1592_
timestamp 1623621585
transform 1 0 22540 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_229
timestamp 1623621585
transform 1 0 22172 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_236
timestamp 1623621585
transform 1 0 22816 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_248
timestamp 1623621585
transform 1 0 23920 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output234
timestamp 1623621585
transform 1 0 25668 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_260
timestamp 1623621585
transform 1 0 25024 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_266
timestamp 1623621585
transform 1 0 25576 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1623621585
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1648_
timestamp 1623621585
transform 1 0 26404 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1623621585
transform 1 0 27324 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output198
timestamp 1623621585
transform 1 0 27876 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_281
timestamp 1623621585
transform 1 0 26956 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_286
timestamp 1623621585
transform 1 0 27416 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_290
timestamp 1623621585
transform 1 0 27784 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_295
timestamp 1623621585
transform 1 0 28244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1623621585
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _2108_
timestamp 1623621585
transform 1 0 1380 0 1 14688
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1623621585
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_21
timestamp 1623621585
transform 1 0 3036 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1623621585
transform 1 0 4232 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _2114_
timestamp 1623621585
transform 1 0 4968 0 1 14688
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1623621585
transform 1 0 3772 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_30
timestamp 1623621585
transform 1 0 3864 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_37
timestamp 1623621585
transform 1 0 4508 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_41
timestamp 1623621585
transform 1 0 4876 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _2058_
timestamp 1623621585
transform 1 0 6992 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_60
timestamp 1623621585
transform 1 0 6624 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1446_
timestamp 1623621585
transform 1 0 9476 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1623621585
transform 1 0 9016 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_73
timestamp 1623621585
transform 1 0 7820 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_85
timestamp 1623621585
transform 1 0 8924 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_87
timestamp 1623621585
transform 1 0 9108 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1958_
timestamp 1623621585
transform 1 0 10672 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_100
timestamp 1623621585
transform 1 0 10304 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1623621585
transform 1 0 11500 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1147_
timestamp 1623621585
transform 1 0 13156 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1154_
timestamp 1623621585
transform 1 0 12052 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_127
timestamp 1623621585
transform 1 0 12788 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1623621585
transform 1 0 14260 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_139
timestamp 1623621585
transform 1 0 13892 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_144
timestamp 1623621585
transform 1 0 14352 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_156
timestamp 1623621585
transform 1 0 15456 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_2  _1530_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 17112 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_168
timestamp 1623621585
transform 1 0 16560 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_182
timestamp 1623621585
transform 1 0 17848 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1623621585
transform 1 0 19504 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_194
timestamp 1623621585
transform 1 0 18952 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_201
timestamp 1623621585
transform 1 0 19596 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__o31ai_1  _1593_
timestamp 1623621585
transform 1 0 21620 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_213
timestamp 1623621585
transform 1 0 20700 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1623621585
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_229
timestamp 1623621585
transform 1 0 22172 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_241
timestamp 1623621585
transform 1 0 23276 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__xor2_1  _1649_
timestamp 1623621585
transform 1 0 25760 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1623621585
transform 1 0 24748 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_253
timestamp 1623621585
transform 1 0 24380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_258
timestamp 1623621585
transform 1 0 24840 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_266
timestamp 1623621585
transform 1 0 25576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2143_
timestamp 1623621585
transform 1 0 26772 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_275
timestamp 1623621585
transform 1 0 26404 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_295
timestamp 1623621585
transform 1 0 28244 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1623621585
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _1223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 2944 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1623621585
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input142
timestamp 1623621585
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1623621585
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_11
timestamp 1623621585
transform 1 0 2116 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_19
timestamp 1623621585
transform 1 0 2852 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a31oi_1  _1290_
timestamp 1623621585
transform 1 0 3956 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  input124
timestamp 1623621585
transform 1 0 4784 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1623621585
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_36
timestamp 1623621585
transform 1 0 4416 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_43
timestamp 1623621585
transform 1 0 5060 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1623621585
transform 1 0 6348 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_55
timestamp 1623621585
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_58
timestamp 1623621585
transform 1 0 6440 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2199_
timestamp 1623621585
transform 1 0 8280 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_70
timestamp 1623621585
transform 1 0 7544 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _1959_
timestamp 1623621585
transform 1 0 10396 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1623621585
transform 1 0 11592 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_94
timestamp 1623621585
transform 1 0 9752 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_100
timestamp 1623621585
transform 1 0 10304 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_110
timestamp 1623621585
transform 1 0 11224 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2261_
timestamp 1623621585
transform 1 0 12052 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1623621585
transform 1 0 11684 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1623621585
transform 1 0 13524 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2264_
timestamp 1623621585
transform 1 0 13892 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_24_155
timestamp 1623621585
transform 1 0 15364 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1148_
timestamp 1623621585
transform 1 0 16008 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1623621585
transform 1 0 16836 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_161
timestamp 1623621585
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_166
timestamp 1623621585
transform 1 0 16376 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_170
timestamp 1623621585
transform 1 0 16744 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_172
timestamp 1623621585
transform 1 0 16928 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux4_2  _2128_
timestamp 1623621585
transform 1 0 18768 0 -1 15776
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_24_184
timestamp 1623621585
transform 1 0 18032 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1623621585
transform 1 0 22080 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_210
timestamp 1623621585
transform 1 0 20424 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_222
timestamp 1623621585
transform 1 0 21528 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_229
timestamp 1623621585
transform 1 0 22172 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_241
timestamp 1623621585
transform 1 0 23276 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux4_2  _2099_
timestamp 1623621585
transform 1 0 24932 0 -1 15776
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_24_253
timestamp 1623621585
transform 1 0 24380 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1623621585
transform 1 0 27324 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output207
timestamp 1623621585
transform 1 0 27876 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_277
timestamp 1623621585
transform 1 0 26588 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_286
timestamp 1623621585
transform 1 0 27416 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_290
timestamp 1623621585
transform 1 0 27784 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_295
timestamp 1623621585
transform 1 0 28244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1623621585
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1222_
timestamp 1623621585
transform 1 0 2760 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1623621585
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input151
timestamp 1623621585
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1623621585
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_11
timestamp 1623621585
transform 1 0 2116 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_17
timestamp 1623621585
transform 1 0 2668 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1728_
timestamp 1623621585
transform 1 0 4876 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1623621585
transform 1 0 3772 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_24
timestamp 1623621585
transform 1 0 3312 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_28
timestamp 1623621585
transform 1 0 3680 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_30
timestamp 1623621585
transform 1 0 3864 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_38
timestamp 1623621585
transform 1 0 4600 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_44
timestamp 1623621585
transform 1 0 5152 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_56
timestamp 1623621585
transform 1 0 6256 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_68
timestamp 1623621585
transform 1 0 7360 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1623621585
transform 1 0 9016 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_80
timestamp 1623621585
transform 1 0 8464 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_87
timestamp 1623621585
transform 1 0 9108 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1683_
timestamp 1623621585
transform 1 0 10764 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_99
timestamp 1623621585
transform 1 0 10212 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_108
timestamp 1623621585
transform 1 0 11040 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_wb_clk_i
timestamp 1623621585
transform 1 0 13248 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_120
timestamp 1623621585
transform 1 0 12144 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1623621585
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_2  _2121_
timestamp 1623621585
transform 1 0 15456 0 1 15776
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1623621585
transform 1 0 14260 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_144
timestamp 1623621585
transform 1 0 14352 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1439_
timestamp 1623621585
transform 1 0 17480 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_174
timestamp 1623621585
transform 1 0 17112 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1623621585
transform 1 0 17756 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1623621585
transform 1 0 19504 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_193
timestamp 1623621585
transform 1 0 18860 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_199
timestamp 1623621585
transform 1 0 19412 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_201
timestamp 1623621585
transform 1 0 19596 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _2135_
timestamp 1623621585
transform 1 0 22080 0 1 15776
box -38 -48 1694 592
use sky130_fd_sc_hd__dfxtp_1  _2159_
timestamp 1623621585
transform 1 0 20240 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_207
timestamp 1623621585
transform 1 0 20148 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_224
timestamp 1623621585
transform 1 0 21712 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_246
timestamp 1623621585
transform 1 0 23736 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1621_
timestamp 1623621585
transform 1 0 25208 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1623621585
transform 1 0 24748 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_254
timestamp 1623621585
transform 1 0 24472 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_258
timestamp 1623621585
transform 1 0 24840 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_271
timestamp 1623621585
transform 1 0 26036 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_4  _1634_
timestamp 1623621585
transform 1 0 26588 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp 1623621585
transform 1 0 28060 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1623621585
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1623621585
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1623621585
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1623621585
transform 1 0 1748 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1623621585
transform 1 0 1748 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1623621585
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1623621585
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_10
timestamp 1623621585
transform 1 0 2024 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_17
timestamp 1623621585
transform 1 0 2668 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_10
timestamp 1623621585
transform 1 0 2024 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1623621585
transform 1 0 2392 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_18
timestamp 1623621585
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input116
timestamp 1623621585
transform 1 0 3036 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1783_
timestamp 1623621585
transform 1 0 2944 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_23
timestamp 1623621585
transform 1 0 3220 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_31
timestamp 1623621585
transform 1 0 3956 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1623621585
transform 1 0 3312 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input133
timestamp 1623621585
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1623621585
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_42
timestamp 1623621585
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_45
timestamp 1623621585
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_39
timestamp 1623621585
transform 1 0 4692 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1976_
timestamp 1623621585
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1727_
timestamp 1623621585
transform 1 0 4968 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_30
timestamp 1623621585
transform 1 0 3864 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_53
timestamp 1623621585
transform 1 0 5980 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_56
timestamp 1623621585
transform 1 0 6256 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_52
timestamp 1623621585
transform 1 0 5888 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1623621585
transform 1 0 6348 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1726_
timestamp 1623621585
transform 1 0 5612 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_61
timestamp 1623621585
transform 1 0 6716 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_62
timestamp 1623621585
transform 1 0 6808 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_58
timestamp 1623621585
transform 1 0 6440 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1345_
timestamp 1623621585
transform 1 0 6900 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _2224_
timestamp 1623621585
transform 1 0 6900 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1623621585
transform 1 0 9016 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1623621585
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_72
timestamp 1623621585
transform 1 0 7728 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1623621585
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_87
timestamp 1623621585
transform 1 0 9108 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_91
timestamp 1623621585
transform 1 0 9476 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1213_
timestamp 1623621585
transform 1 0 10948 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1357_
timestamp 1623621585
transform 1 0 10304 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1756_
timestamp 1623621585
transform 1 0 9568 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1623621585
transform 1 0 11592 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_92
timestamp 1623621585
transform 1 0 9568 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_104
timestamp 1623621585
transform 1 0 10672 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_112
timestamp 1623621585
transform 1 0 11408 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_95
timestamp 1623621585
transform 1 0 9844 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_111
timestamp 1623621585
transform 1 0 11316 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_115
timestamp 1623621585
transform 1 0 11684 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_127
timestamp 1623621585
transform 1 0 12788 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1623621585
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_135
timestamp 1623621585
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _2204_
timestamp 1623621585
transform 1 0 14812 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1623621585
transform 1 0 14260 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_139
timestamp 1623621585
transform 1 0 13892 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_147
timestamp 1623621585
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_144
timestamp 1623621585
transform 1 0 14352 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_156
timestamp 1623621585
transform 1 0 15456 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__xor2_1  _1545_
timestamp 1623621585
transform 1 0 17388 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1623621585
transform 1 0 16836 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_166
timestamp 1623621585
transform 1 0 16376 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_170
timestamp 1623621585
transform 1 0 16744 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_172
timestamp 1623621585
transform 1 0 16928 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_176
timestamp 1623621585
transform 1 0 17296 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_168
timestamp 1623621585
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_180
timestamp 1623621585
transform 1 0 17664 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_186
timestamp 1623621585
transform 1 0 18216 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_188
timestamp 1623621585
transform 1 0 18400 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_184
timestamp 1623621585
transform 1 0 18032 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1546_
timestamp 1623621585
transform 1 0 18308 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_201
timestamp 1623621585
transform 1 0 19596 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_196
timestamp 1623621585
transform 1 0 19136 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_205
timestamp 1623621585
transform 1 0 19964 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_wb_clk_i
timestamp 1623621585
transform 1 0 19964 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1623621585
transform 1 0 19504 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2175_
timestamp 1623621585
transform 1 0 18492 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__and2b_1  _1589_
timestamp 1623621585
transform 1 0 21252 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1590_
timestamp 1623621585
transform 1 0 20700 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1623621585
transform 1 0 22080 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_220
timestamp 1623621585
transform 1 0 21344 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_208
timestamp 1623621585
transform 1 0 20240 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_216
timestamp 1623621585
transform 1 0 20976 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1623621585
transform 1 0 21804 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__xor2_1  _1620_
timestamp 1623621585
transform 1 0 23644 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_26_229
timestamp 1623621585
transform 1 0 22172 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_241
timestamp 1623621585
transform 1 0 23276 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1623621585
transform 1 0 22908 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_249
timestamp 1623621585
transform 1 0 24012 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2151_
timestamp 1623621585
transform 1 0 24656 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1623621585
transform 1 0 24748 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output243
timestamp 1623621585
transform 1 0 25944 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_252
timestamp 1623621585
transform 1 0 24288 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_272
timestamp 1623621585
transform 1 0 26128 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_258
timestamp 1623621585
transform 1 0 24840 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_274
timestamp 1623621585
transform 1 0 26312 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_282
timestamp 1623621585
transform 1 0 27048 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_281
timestamp 1623621585
transform 1 0 26956 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1623621585
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output225
timestamp 1623621585
transform 1 0 26588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output199
timestamp 1623621585
transform 1 0 26680 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_290
timestamp 1623621585
transform 1 0 27784 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_286
timestamp 1623621585
transform 1 0 27416 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output181
timestamp 1623621585
transform 1 0 27876 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1623621585
transform 1 0 27324 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1650_
timestamp 1623621585
transform 1 0 27416 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_295
timestamp 1623621585
transform 1 0 28244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_295
timestamp 1623621585
transform 1 0 28244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1623621585
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1623621585
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2214_
timestamp 1623621585
transform 1 0 1380 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1623621585
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_19
timestamp 1623621585
transform 1 0 2852 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1373_
timestamp 1623621585
transform 1 0 4416 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1977_
timestamp 1623621585
transform 1 0 5152 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2017_
timestamp 1623621585
transform 1 0 3220 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_32
timestamp 1623621585
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_39
timestamp 1623621585
transform 1 0 4692 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_43
timestamp 1623621585
transform 1 0 5060 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _1344_
timestamp 1623621585
transform 1 0 6808 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1623621585
transform 1 0 6348 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_53
timestamp 1623621585
transform 1 0 5980 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1623621585
transform 1 0 6440 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2200_
timestamp 1623621585
transform 1 0 8280 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_28_69
timestamp 1623621585
transform 1 0 7452 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_77
timestamp 1623621585
transform 1 0 8188 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _2085_
timestamp 1623621585
transform 1 0 10212 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1623621585
transform 1 0 11592 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_94
timestamp 1623621585
transform 1 0 9752 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_98
timestamp 1623621585
transform 1 0 10120 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_108
timestamp 1623621585
transform 1 0 11040 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 12052 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_28_115
timestamp 1623621585
transform 1 0 11684 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2007_
timestamp 1623621585
transform 1 0 14168 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_138
timestamp 1623621585
transform 1 0 13800 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_151
timestamp 1623621585
transform 1 0 14996 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _1540_
timestamp 1623621585
transform 1 0 17480 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1623621585
transform 1 0 16836 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_163
timestamp 1623621585
transform 1 0 16100 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_172
timestamp 1623621585
transform 1 0 16928 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_185
timestamp 1623621585
transform 1 0 18124 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1623621585
transform 1 0 19228 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1623621585
transform 1 0 22080 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1623621585
transform 1 0 20332 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_221
timestamp 1623621585
transform 1 0 21436 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_227
timestamp 1623621585
transform 1 0 21988 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1586_
timestamp 1623621585
transform 1 0 22540 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_229
timestamp 1623621585
transform 1 0 22172 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_236
timestamp 1623621585
transform 1 0 22816 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_248
timestamp 1623621585
transform 1 0 23920 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1631_
timestamp 1623621585
transform 1 0 25944 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_260
timestamp 1623621585
transform 1 0 25024 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_268
timestamp 1623621585
transform 1 0 25760 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_273
timestamp 1623621585
transform 1 0 26220 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1623621585
transform 1 0 27324 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output190
timestamp 1623621585
transform 1 0 27876 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output208
timestamp 1623621585
transform 1 0 26588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_281
timestamp 1623621585
transform 1 0 26956 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_286
timestamp 1623621585
transform 1 0 27416 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_290
timestamp 1623621585
transform 1 0 27784 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_295
timestamp 1623621585
transform 1 0 28244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1623621585
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1371_
timestamp 1623621585
transform 1 0 1840 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1782_
timestamp 1623621585
transform 1 0 3036 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1623621585
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1623621585
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1623621585
transform 1 0 1748 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_17
timestamp 1623621585
transform 1 0 2668 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _2018_
timestamp 1623621585
transform 1 0 4232 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1623621585
transform 1 0 3772 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_24
timestamp 1623621585
transform 1 0 3312 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_28
timestamp 1623621585
transform 1 0 3680 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_30
timestamp 1623621585
transform 1 0 3864 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_43
timestamp 1623621585
transform 1 0 5060 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2061_
timestamp 1623621585
transform 1 0 5428 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_56
timestamp 1623621585
transform 1 0 6256 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_68
timestamp 1623621585
transform 1 0 7360 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1336_
timestamp 1623621585
transform 1 0 9476 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1623621585
transform 1 0 9016 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_80
timestamp 1623621585
transform 1 0 8464 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_87
timestamp 1623621585
transform 1 0 9108 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1676_
timestamp 1623621585
transform 1 0 10212 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_8  _1961_
timestamp 1623621585
transform 1 0 10856 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_29_95
timestamp 1623621585
transform 1 0 9844 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_102
timestamp 1623621585
transform 1 0 10488 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_127
timestamp 1623621585
transform 1 0 12788 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1745_
timestamp 1623621585
transform 1 0 14720 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _2122_
timestamp 1623621585
transform 1 0 15640 0 1 17952
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1623621585
transform 1 0 14260 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_139
timestamp 1623621585
transform 1 0 13892 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_144
timestamp 1623621585
transform 1 0 14352 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_151
timestamp 1623621585
transform 1 0 14996 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_157
timestamp 1623621585
transform 1 0 15548 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_176
timestamp 1623621585
transform 1 0 17296 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1544_
timestamp 1623621585
transform 1 0 18308 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1623621585
transform 1 0 19504 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_184
timestamp 1623621585
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1623621585
transform 1 0 19136 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_201
timestamp 1623621585
transform 1 0 19596 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_2  _1573_
timestamp 1623621585
transform 1 0 20608 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_209
timestamp 1623621585
transform 1 0 20332 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_221
timestamp 1623621585
transform 1 0 21436 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1605_
timestamp 1623621585
transform 1 0 24104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2160_
timestamp 1623621585
transform 1 0 22264 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_29_229
timestamp 1623621585
transform 1 0 22172 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_246
timestamp 1623621585
transform 1 0 23736 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2152_
timestamp 1623621585
transform 1 0 25208 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1623621585
transform 1 0 24748 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_253
timestamp 1623621585
transform 1 0 24380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_258
timestamp 1623621585
transform 1 0 24840 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1647_
timestamp 1623621585
transform 1 0 27416 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_278
timestamp 1623621585
transform 1 0 26680 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_295
timestamp 1623621585
transform 1 0 28244 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1623621585
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _2109_
timestamp 1623621585
transform 1 0 1380 0 -1 19040
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1623621585
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_21
timestamp 1623621585
transform 1 0 3036 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _2115_
timestamp 1623621585
transform 1 0 4140 0 -1 19040
box -38 -48 1694 592
use sky130_fd_sc_hd__buf_1  input134
timestamp 1623621585
transform 1 0 3404 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_28
timestamp 1623621585
transform 1 0 3680 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_32
timestamp 1623621585
transform 1 0 4048 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1323_
timestamp 1623621585
transform 1 0 6808 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1623621585
transform 1 0 6348 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_51
timestamp 1623621585
transform 1 0 5796 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1623621585
transform 1 0 6440 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_65
timestamp 1623621585
transform 1 0 7084 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1445_
timestamp 1623621585
transform 1 0 8556 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1755_
timestamp 1623621585
transform 1 0 7912 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_73
timestamp 1623621585
transform 1 0 7820 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_77
timestamp 1623621585
transform 1 0 8188 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_90
timestamp 1623621585
transform 1 0 9384 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1678_
timestamp 1623621585
transform 1 0 9752 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1960_
timestamp 1623621585
transform 1 0 10396 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1623621585
transform 1 0 11592 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1623621585
transform 1 0 10028 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_110
timestamp 1623621585
transform 1 0 11224 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2246_
timestamp 1623621585
transform 1 0 12236 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_30_115
timestamp 1623621585
transform 1 0 11684 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _2008_
timestamp 1623621585
transform 1 0 14352 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_140
timestamp 1623621585
transform 1 0 13984 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_153
timestamp 1623621585
transform 1 0 15180 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _1531_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 17388 0 -1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1623621585
transform 1 0 16836 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_wb_clk_i
timestamp 1623621585
transform 1 0 16100 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_161
timestamp 1623621585
transform 1 0 15916 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_166
timestamp 1623621585
transform 1 0 16376 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_170
timestamp 1623621585
transform 1 0 16744 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1623621585
transform 1 0 16928 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_176
timestamp 1623621585
transform 1 0 17296 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_2  _2129_
timestamp 1623621585
transform 1 0 19044 0 -1 19040
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 1623621585
transform 1 0 18676 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1587_
timestamp 1623621585
transform 1 0 21160 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1623621585
transform 1 0 22080 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1623621585
transform 1 0 20700 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_217
timestamp 1623621585
transform 1 0 21068 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_224
timestamp 1623621585
transform 1 0 21712 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _2136_
timestamp 1623621585
transform 1 0 22540 0 -1 19040
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_30_229
timestamp 1623621585
transform 1 0 22172 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_251
timestamp 1623621585
transform 1 0 24196 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1601_
timestamp 1623621585
transform 1 0 24564 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _2098_
timestamp 1623621585
transform 1 0 25208 0 -1 19040
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1623621585
transform 1 0 24840 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1623621585
transform 1 0 27324 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output217
timestamp 1623621585
transform 1 0 27876 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_280
timestamp 1623621585
transform 1 0 26864 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_284
timestamp 1623621585
transform 1 0 27232 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_286
timestamp 1623621585
transform 1 0 27416 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_290
timestamp 1623621585
transform 1 0 27784 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_295
timestamp 1623621585
transform 1 0 28244 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1623621585
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1786_
timestamp 1623621585
transform 1 0 3128 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1623621585
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input125
timestamp 1623621585
transform 1 0 2484 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input143
timestamp 1623621585
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1623621585
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_11
timestamp 1623621585
transform 1 0 2116 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_18
timestamp 1623621585
transform 1 0 2760 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2014_
timestamp 1623621585
transform 1 0 4232 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1623621585
transform 1 0 3772 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_25
timestamp 1623621585
transform 1 0 3404 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_30
timestamp 1623621585
transform 1 0 3864 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_43
timestamp 1623621585
transform 1 0 5060 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1313_
timestamp 1623621585
transform 1 0 5980 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _1340_
timestamp 1623621585
transform 1 0 6900 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_51
timestamp 1623621585
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_59
timestamp 1623621585
transform 1 0 6532 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1320_
timestamp 1623621585
transform 1 0 7820 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2039_
timestamp 1623621585
transform 1 0 9476 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1623621585
transform 1 0 9016 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_69
timestamp 1623621585
transform 1 0 7452 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_76
timestamp 1623621585
transform 1 0 8096 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_84
timestamp 1623621585
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_87
timestamp 1623621585
transform 1 0 9108 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1677_
timestamp 1623621585
transform 1 0 11224 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_100
timestamp 1623621585
transform 1 0 10304 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_108
timestamp 1623621585
transform 1 0 11040 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1623621585
transform 1 0 11500 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_wb_clk_i
timestamp 1623621585
transform 1 0 11868 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_120
timestamp 1623621585
transform 1 0 12144 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_132
timestamp 1623621585
transform 1 0 13248 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2249_
timestamp 1623621585
transform 1 0 14720 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1623621585
transform 1 0 14260 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_140
timestamp 1623621585
transform 1 0 13984 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_144
timestamp 1623621585
transform 1 0 14352 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2250_
timestamp 1623621585
transform 1 0 16836 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_31_167
timestamp 1623621585
transform 1 0 16468 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1623621585
transform 1 0 19504 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_190
timestamp 1623621585
transform 1 0 18584 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_198
timestamp 1623621585
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_201
timestamp 1623621585
transform 1 0 19596 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_1  _1570_
timestamp 1623621585
transform 1 0 20792 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1585_
timestamp 1623621585
transform 1 0 21896 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_213
timestamp 1623621585
transform 1 0 20700 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_222
timestamp 1623621585
transform 1 0 21528 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1618_
timestamp 1623621585
transform 1 0 23736 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_31_230
timestamp 1623621585
transform 1 0 22264 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_242
timestamp 1623621585
transform 1 0 23368 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1619_
timestamp 1623621585
transform 1 0 25208 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1623621585
transform 1 0 24748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_253
timestamp 1623621585
transform 1 0 24380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_258
timestamp 1623621585
transform 1 0 24840 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_271
timestamp 1623621585
transform 1 0 26036 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2144_
timestamp 1623621585
transform 1 0 26772 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_295
timestamp 1623621585
transform 1 0 28244 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1623621585
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1623621585
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1623621585
transform 1 0 2484 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input126
timestamp 1623621585
transform 1 0 3128 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input152
timestamp 1623621585
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1623621585
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_11
timestamp 1623621585
transform 1 0 2116 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_18
timestamp 1623621585
transform 1 0 2760 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2013_
timestamp 1623621585
transform 1 0 4140 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_25
timestamp 1623621585
transform 1 0 3404 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_42
timestamp 1623621585
transform 1 0 4968 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_4  _1309_
timestamp 1623621585
transform 1 0 7084 0 -1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1623621585
transform 1 0 6348 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_54
timestamp 1623621585
transform 1 0 6072 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_58
timestamp 1623621585
transform 1 0 6440 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_64
timestamp 1623621585
transform 1 0 6992 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _2040_
timestamp 1623621585
transform 1 0 8740 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1623621585
transform 1 0 8372 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1342_
timestamp 1623621585
transform 1 0 9936 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1623621585
transform 1 0 11592 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_92
timestamp 1623621585
transform 1 0 9568 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_99
timestamp 1623621585
transform 1 0 10212 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_111
timestamp 1623621585
transform 1 0 11316 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_115
timestamp 1623621585
transform 1 0 11684 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_127
timestamp 1623621585
transform 1 0 12788 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_139
timestamp 1623621585
transform 1 0 13892 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_151
timestamp 1623621585
transform 1 0 14996 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__xor2_1  _1543_
timestamp 1623621585
transform 1 0 17388 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1623621585
transform 1 0 16836 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_163
timestamp 1623621585
transform 1 0 16100 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_172
timestamp 1623621585
transform 1 0 16928 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_176
timestamp 1623621585
transform 1 0 17296 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2176_
timestamp 1623621585
transform 1 0 18584 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_32_184
timestamp 1623621585
transform 1 0 18032 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1623621585
transform 1 0 22080 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_206
timestamp 1623621585
transform 1 0 20056 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_218
timestamp 1623621585
transform 1 0 21160 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_226
timestamp 1623621585
transform 1 0 21896 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_229
timestamp 1623621585
transform 1 0 22172 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_241
timestamp 1623621585
transform 1 0 23276 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1599_
timestamp 1623621585
transform 1 0 24932 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1646_
timestamp 1623621585
transform 1 0 26312 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output235
timestamp 1623621585
transform 1 0 25576 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_253
timestamp 1623621585
transform 1 0 24380 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_262
timestamp 1623621585
transform 1 0 25208 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_270
timestamp 1623621585
transform 1 0 25944 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1623621585
transform 1 0 27324 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output182
timestamp 1623621585
transform 1 0 27876 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_281
timestamp 1623621585
transform 1 0 26956 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_286
timestamp 1623621585
transform 1 0 27416 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_290
timestamp 1623621585
transform 1 0 27784 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_295
timestamp 1623621585
transform 1 0 28244 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1623621585
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_7
timestamp 1623621585
transform 1 0 1748 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_3
timestamp 1623621585
transform 1 0 1380 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1623621585
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1623621585
transform 1 0 1472 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1623621585
transform 1 0 1748 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1623621585
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1623621585
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_18
timestamp 1623621585
transform 1 0 2760 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_10
timestamp 1623621585
transform 1 0 2024 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _2016_
timestamp 1623621585
transform 1 0 2116 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1784_
timestamp 1623621585
transform 1 0 2852 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_20
timestamp 1623621585
transform 1 0 2944 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_22
timestamp 1623621585
transform 1 0 3128 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1721_
timestamp 1623621585
transform 1 0 4416 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2015_
timestamp 1623621585
transform 1 0 3312 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1623621585
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_28
timestamp 1623621585
transform 1 0 3680 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_30
timestamp 1623621585
transform 1 0 3864 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_39
timestamp 1623621585
transform 1 0 4692 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_33
timestamp 1623621585
transform 1 0 4140 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_45
timestamp 1623621585
transform 1 0 5244 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_2  _1307_
timestamp 1623621585
transform 1 0 5612 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__o21bai_1  _1325_
timestamp 1623621585
transform 1 0 6808 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1623621585
transform 1 0 6348 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_47
timestamp 1623621585
transform 1 0 5428 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_62
timestamp 1623621585
transform 1 0 6808 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_58
timestamp 1623621585
transform 1 0 6440 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1623621585
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__xor2_1  _1341_
timestamp 1623621585
transform 1 0 7544 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1623621585
transform 1 0 9016 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_wb_clk_i
timestamp 1623621585
transform 1 0 9016 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_77
timestamp 1623621585
transform 1 0 8188 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_85
timestamp 1623621585
transform 1 0 8924 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_87
timestamp 1623621585
transform 1 0 9108 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_80
timestamp 1623621585
transform 1 0 8464 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_89
timestamp 1623621585
transform 1 0 9292 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 10672 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1343_
timestamp 1623621585
transform 1 0 9660 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2225_
timestamp 1623621585
transform 1 0 9936 0 1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1623621585
transform 1 0 11592 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_95
timestamp 1623621585
transform 1 0 9844 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1623621585
transform 1 0 11500 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_97
timestamp 1623621585
transform 1 0 10028 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_103
timestamp 1623621585
transform 1 0 10580 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_110
timestamp 1623621585
transform 1 0 11224 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_115
timestamp 1623621585
transform 1 0 11684 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1623621585
transform 1 0 12052 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1199_
timestamp 1623621585
transform 1 0 12144 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1197_
timestamp 1623621585
transform 1 0 12052 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_127
timestamp 1623621585
transform 1 0 12788 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_128
timestamp 1623621585
transform 1 0 12880 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_133
timestamp 1623621585
transform 1 0 13340 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_135
timestamp 1623621585
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_wb_clk_i
timestamp 1623621585
transform 1 0 13248 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1191_
timestamp 1623621585
transform 1 0 13432 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _1187_
timestamp 1623621585
transform 1 0 14904 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1192_
timestamp 1623621585
transform 1 0 14720 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1623621585
transform 1 0 14260 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_144
timestamp 1623621585
transform 1 0 14352 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_156
timestamp 1623621585
transform 1 0 15456 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_140
timestamp 1623621585
transform 1 0 13984 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_148
timestamp 1623621585
transform 1 0 14720 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_156
timestamp 1623621585
transform 1 0 15456 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1186_
timestamp 1623621585
transform 1 0 15824 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _2123_
timestamp 1623621585
transform 1 0 16100 0 1 20128
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1623621585
transform 1 0 16836 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_162
timestamp 1623621585
transform 1 0 16008 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1623621585
transform 1 0 17756 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_163
timestamp 1623621585
transform 1 0 16100 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_172
timestamp 1623621585
transform 1 0 16928 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_180
timestamp 1623621585
transform 1 0 17664 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1541_
timestamp 1623621585
transform 1 0 17940 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1623621585
transform 1 0 19504 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_193
timestamp 1623621585
transform 1 0 18860 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_199
timestamp 1623621585
transform 1 0 19412 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_201
timestamp 1623621585
transform 1 0 19596 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_187
timestamp 1623621585
transform 1 0 18308 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_199
timestamp 1623621585
transform 1 0 19412 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_1  _1574_
timestamp 1623621585
transform 1 0 20792 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1583_
timestamp 1623621585
transform 1 0 21436 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1623621585
transform 1 0 22080 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_wb_clk_i
timestamp 1623621585
transform 1 0 20792 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_213
timestamp 1623621585
transform 1 0 20700 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_217
timestamp 1623621585
transform 1 0 21068 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_228
timestamp 1623621585
transform 1 0 22080 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_211
timestamp 1623621585
transform 1 0 20516 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_222
timestamp 1623621585
transform 1 0 21528 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1584_
timestamp 1623621585
transform 1 0 22540 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1612_
timestamp 1623621585
transform 1 0 23920 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_wb_clk_i
timestamp 1623621585
transform 1 0 22448 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_235
timestamp 1623621585
transform 1 0 22724 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_247
timestamp 1623621585
transform 1 0 23828 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_229
timestamp 1623621585
transform 1 0 22172 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_242
timestamp 1623621585
transform 1 0 23368 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1600_
timestamp 1623621585
transform 1 0 25300 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1623621585
transform 1 0 24748 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output244
timestamp 1623621585
transform 1 0 25668 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_255
timestamp 1623621585
transform 1 0 24564 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_258
timestamp 1623621585
transform 1 0 24840 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_266
timestamp 1623621585
transform 1 0 25576 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_271
timestamp 1623621585
transform 1 0 26036 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_255
timestamp 1623621585
transform 1 0 24564 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_267
timestamp 1623621585
transform 1 0 25668 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_275
timestamp 1623621585
transform 1 0 26404 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output226
timestamp 1623621585
transform 1 0 26404 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output209
timestamp 1623621585
transform 1 0 26588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_281
timestamp 1623621585
transform 1 0 26956 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_279
timestamp 1623621585
transform 1 0 26772 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output218
timestamp 1623621585
transform 1 0 27140 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_286
timestamp 1623621585
transform 1 0 27416 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_287
timestamp 1623621585
transform 1 0 27508 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1623621585
transform 1 0 27324 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_290
timestamp 1623621585
transform 1 0 27784 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output200
timestamp 1623621585
transform 1 0 27876 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output191
timestamp 1623621585
transform 1 0 27876 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_295
timestamp 1623621585
transform 1 0 28244 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_295
timestamp 1623621585
transform 1 0 28244 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1623621585
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1623621585
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _2110_
timestamp 1623621585
transform 1 0 1380 0 1 21216
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1623621585
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_21
timestamp 1623621585
transform 1 0 3036 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2064_
timestamp 1623621585
transform 1 0 4692 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1623621585
transform 1 0 3772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_30
timestamp 1623621585
transform 1 0 3864 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_38
timestamp 1623621585
transform 1 0 4600 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__o22ai_1  _1324_
timestamp 1623621585
transform 1 0 6716 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_35_48
timestamp 1623621585
transform 1 0 5520 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_60
timestamp 1623621585
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_66
timestamp 1623621585
transform 1 0 7176 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1623621585
transform 1 0 9016 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_78
timestamp 1623621585
transform 1 0 8280 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_87
timestamp 1623621585
transform 1 0 9108 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _2088_
timestamp 1623621585
transform 1 0 10212 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_35_108
timestamp 1623621585
transform 1 0 11040 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1194_
timestamp 1623621585
transform 1 0 12052 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1195_
timestamp 1623621585
transform 1 0 12972 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_116
timestamp 1623621585
transform 1 0 11776 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp 1623621585
transform 1 0 12604 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_137
timestamp 1623621585
transform 1 0 13708 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1188_
timestamp 1623621585
transform 1 0 15272 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1623621585
transform 1 0 14260 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_144
timestamp 1623621585
transform 1 0 14352 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_152
timestamp 1623621585
transform 1 0 15088 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_162
timestamp 1623621585
transform 1 0 16008 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_174
timestamp 1623621585
transform 1 0 17112 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_1  _1542_
timestamp 1623621585
transform 1 0 18400 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_2  _2130_
timestamp 1623621585
transform 1 0 19964 0 1 21216
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1623621585
transform 1 0 19504 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_186
timestamp 1623621585
transform 1 0 18216 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_196
timestamp 1623621585
transform 1 0 19136 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_201
timestamp 1623621585
transform 1 0 19596 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_223
timestamp 1623621585
transform 1 0 21620 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2161_
timestamp 1623621585
transform 1 0 22356 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_35_247
timestamp 1623621585
transform 1 0 23828 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2153_
timestamp 1623621585
transform 1 0 25208 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1623621585
transform 1 0 24748 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_255
timestamp 1623621585
transform 1 0 24564 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_258
timestamp 1623621585
transform 1 0 24840 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1645_
timestamp 1623621585
transform 1 0 27416 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_35_278
timestamp 1623621585
transform 1 0 26680 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_295
timestamp 1623621585
transform 1 0 28244 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1623621585
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1372_
timestamp 1623621585
transform 1 0 2024 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1623621585
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1623621585
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_6
timestamp 1623621585
transform 1 0 1656 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_19
timestamp 1623621585
transform 1 0 2852 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1785_
timestamp 1623621585
transform 1 0 3220 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _2116_
timestamp 1623621585
transform 1 0 4232 0 -1 22304
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_36_26
timestamp 1623621585
transform 1 0 3496 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1322_
timestamp 1623621585
transform 1 0 6992 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1623621585
transform 1 0 6348 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_52
timestamp 1623621585
transform 1 0 5888 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_56
timestamp 1623621585
transform 1 0 6256 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_58
timestamp 1623621585
transform 1 0 6440 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_67
timestamp 1623621585
transform 1 0 7268 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1444_
timestamp 1623621585
transform 1 0 8096 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_36_75
timestamp 1623621585
transform 1 0 8004 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1623621585
transform 1 0 8924 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1339_
timestamp 1623621585
transform 1 0 10120 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1671_
timestamp 1623621585
transform 1 0 10764 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1623621585
transform 1 0 11592 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_97
timestamp 1623621585
transform 1 0 10028 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_101
timestamp 1623621585
transform 1 0 10396 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_108
timestamp 1623621585
transform 1 0 11040 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _1196_
timestamp 1623621585
transform 1 0 12052 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2248_
timestamp 1623621585
transform 1 0 13248 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_36_115
timestamp 1623621585
transform 1 0 11684 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_125
timestamp 1623621585
transform 1 0 12604 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_131
timestamp 1623621585
transform 1 0 13156 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1181_
timestamp 1623621585
transform 1 0 15732 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_151
timestamp 1623621585
transform 1 0 14996 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1623621585
transform 1 0 16836 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_167
timestamp 1623621585
transform 1 0 16468 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_172
timestamp 1623621585
transform 1 0 16928 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2177_
timestamp 1623621585
transform 1 0 18308 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_36_184
timestamp 1623621585
transform 1 0 18032 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_203
timestamp 1623621585
transform 1 0 19780 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a41oi_2  _1580_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 20516 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1623621585
transform 1 0 22080 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_224
timestamp 1623621585
transform 1 0 21712 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _2137_
timestamp 1623621585
transform 1 0 22540 0 -1 22304
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_36_229
timestamp 1623621585
transform 1 0 22172 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_251
timestamp 1623621585
transform 1 0 24196 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_2  _2097_
timestamp 1623621585
transform 1 0 25116 0 -1 22304
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_36_259
timestamp 1623621585
transform 1 0 24932 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_2  _1635_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 27784 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1623621585
transform 1 0 27324 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_279
timestamp 1623621585
transform 1 0 26772 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_286
timestamp 1623621585
transform 1 0 27416 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_295
timestamp 1623621585
transform 1 0 28244 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1623621585
transform -1 0 28888 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2213_
timestamp 1623621585
transform 1 0 1380 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1623621585
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_19
timestamp 1623621585
transform 1 0 2852 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1787_
timestamp 1623621585
transform 1 0 4232 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1623621585
transform 1 0 3772 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_27
timestamp 1623621585
transform 1 0 3588 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_30
timestamp 1623621585
transform 1 0 3864 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_37
timestamp 1623621585
transform 1 0 4508 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_2  _1308_
timestamp 1623621585
transform 1 0 6348 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_37_49
timestamp 1623621585
transform 1 0 5612 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1752_
timestamp 1623621585
transform 1 0 8372 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1753_
timestamp 1623621585
transform 1 0 9476 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1623621585
transform 1 0 9016 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_70
timestamp 1623621585
transform 1 0 7544 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_78
timestamp 1623621585
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_82
timestamp 1623621585
transform 1 0 8648 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_87
timestamp 1623621585
transform 1 0 9108 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_4  _1963_
timestamp 1623621585
transform 1 0 10580 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_94
timestamp 1623621585
transform 1 0 9752 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_102
timestamp 1623621585
transform 1 0 10488 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1962_
timestamp 1623621585
transform 1 0 12052 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_37_115
timestamp 1623621585
transform 1 0 11684 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_128
timestamp 1623621585
transform 1 0 12880 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3b_1  _1180_
timestamp 1623621585
transform 1 0 15456 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1623621585
transform 1 0 14260 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_140
timestamp 1623621585
transform 1 0 13984 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_144
timestamp 1623621585
transform 1 0 14352 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _2253_
timestamp 1623621585
transform 1 0 16376 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_37_162
timestamp 1623621585
transform 1 0 16008 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1623621585
transform 1 0 19504 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_185
timestamp 1623621585
transform 1 0 18124 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_197
timestamp 1623621585
transform 1 0 19228 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_201
timestamp 1623621585
transform 1 0 19596 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1571_
timestamp 1623621585
transform 1 0 21344 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_wb_clk_i
timestamp 1623621585
transform 1 0 20148 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_210
timestamp 1623621585
transform 1 0 20424 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_218
timestamp 1623621585
transform 1 0 21160 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_227
timestamp 1623621585
transform 1 0 21988 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1572_
timestamp 1623621585
transform 1 0 22448 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _1615_
timestamp 1623621585
transform 1 0 23828 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_37_231
timestamp 1623621585
transform 1 0 22356 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_236
timestamp 1623621585
transform 1 0 22816 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_244
timestamp 1623621585
transform 1 0 23552 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1616_
timestamp 1623621585
transform 1 0 26128 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1617_
timestamp 1623621585
transform 1 0 25208 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1623621585
transform 1 0 24748 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_252
timestamp 1623621585
transform 1 0 24288 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_256
timestamp 1623621585
transform 1 0 24656 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_258
timestamp 1623621585
transform 1 0 24840 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_268
timestamp 1623621585
transform 1 0 25760 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2145_
timestamp 1623621585
transform 1 0 26772 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1623621585
transform 1 0 26404 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_295
timestamp 1623621585
transform 1 0 28244 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1623621585
transform -1 0 28888 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1623621585
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1623621585
transform 1 0 2484 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input144
timestamp 1623621585
transform 1 0 1748 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1623621585
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_11
timestamp 1623621585
transform 1 0 2116 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_18
timestamp 1623621585
transform 1 0 2760 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_22
timestamp 1623621585
transform 1 0 3128 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1374_
timestamp 1623621585
transform 1 0 3220 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1716_
timestamp 1623621585
transform 1 0 4692 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_32
timestamp 1623621585
transform 1 0 4048 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_38
timestamp 1623621585
transform 1 0 4600 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_42
timestamp 1623621585
transform 1 0 4968 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _1314_
timestamp 1623621585
transform 1 0 6808 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1623621585
transform 1 0 6348 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_54
timestamp 1623621585
transform 1 0 6072 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_58
timestamp 1623621585
transform 1 0 6440 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_68
timestamp 1623621585
transform 1 0 7360 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2201_
timestamp 1623621585
transform 1 0 7820 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_38_72
timestamp 1623621585
transform 1 0 7728 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_89
timestamp 1623621585
transform 1 0 9292 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1672_
timestamp 1623621585
transform 1 0 10856 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2041_
timestamp 1623621585
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1623621585
transform 1 0 11592 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_102
timestamp 1623621585
transform 1 0 10488 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_109
timestamp 1623621585
transform 1 0 11132 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_113
timestamp 1623621585
transform 1 0 11500 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1190_
timestamp 1623621585
transform 1 0 13432 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_115
timestamp 1623621585
transform 1 0 11684 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_127
timestamp 1623621585
transform 1 0 12788 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_133
timestamp 1623621585
transform 1 0 13340 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1172_
timestamp 1623621585
transform 1 0 15640 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1179_
timestamp 1623621585
transform 1 0 14904 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1193_
timestamp 1623621585
transform 1 0 14168 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_138
timestamp 1623621585
transform 1 0 13800 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_146
timestamp 1623621585
transform 1 0 14536 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_154
timestamp 1623621585
transform 1 0 15272 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1165_
timestamp 1623621585
transform 1 0 17572 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1623621585
transform 1 0 16836 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_161
timestamp 1623621585
transform 1 0 15916 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_169
timestamp 1623621585
transform 1 0 16652 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_172
timestamp 1623621585
transform 1 0 16928 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_178
timestamp 1623621585
transform 1 0 17480 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_183
timestamp 1623621585
transform 1 0 17940 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_195
timestamp 1623621585
transform 1 0 19044 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1623621585
transform 1 0 22080 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_207
timestamp 1623621585
transform 1 0 20148 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_219
timestamp 1623621585
transform 1 0 21252 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_227
timestamp 1623621585
transform 1 0 21988 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_229
timestamp 1623621585
transform 1 0 22172 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_241
timestamp 1623621585
transform 1 0 23276 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__xor2_1  _1644_
timestamp 1623621585
transform 1 0 26312 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output227
timestamp 1623621585
transform 1 0 25576 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output245
timestamp 1623621585
transform 1 0 24840 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_253
timestamp 1623621585
transform 1 0 24380 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_257
timestamp 1623621585
transform 1 0 24748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_262
timestamp 1623621585
transform 1 0 25208 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_270
timestamp 1623621585
transform 1 0 25944 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1623621585
transform 1 0 27324 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output183
timestamp 1623621585
transform 1 0 27876 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_281
timestamp 1623621585
transform 1 0 26956 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_286
timestamp 1623621585
transform 1 0 27416 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_290
timestamp 1623621585
transform 1 0 27784 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_295
timestamp 1623621585
transform 1 0 28244 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1623621585
transform -1 0 28888 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_10
timestamp 1623621585
transform 1 0 2024 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1623621585
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_11
timestamp 1623621585
transform 1 0 2116 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1623621585
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input153
timestamp 1623621585
transform 1 0 1748 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1623621585
transform 1 0 1748 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1623621585
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1623621585
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_18
timestamp 1623621585
transform 1 0 2760 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_18
timestamp 1623621585
transform 1 0 2760 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1623621585
transform 1 0 3128 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1623621585
transform 1 0 2484 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2212_
timestamp 1623621585
transform 1 0 2852 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _2067_
timestamp 1623621585
transform 1 0 4784 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1623621585
transform 1 0 3772 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input135
timestamp 1623621585
transform 1 0 4232 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_25
timestamp 1623621585
transform 1 0 3404 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_30
timestamp 1623621585
transform 1 0 3864 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_37
timestamp 1623621585
transform 1 0 4508 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_35
timestamp 1623621585
transform 1 0 4324 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_39
timestamp 1623621585
transform 1 0 4692 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_49
timestamp 1623621585
transform 1 0 5612 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_53
timestamp 1623621585
transform 1 0 5980 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_49
timestamp 1623621585
transform 1 0 5612 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1623621585
transform 1 0 6348 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_1  _1311_
timestamp 1623621585
transform 1 0 6072 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_58
timestamp 1623621585
transform 1 0 6440 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_67
timestamp 1623621585
transform 1 0 7268 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_60
timestamp 1623621585
transform 1 0 6624 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1312_
timestamp 1623621585
transform 1 0 6992 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1315_
timestamp 1623621585
transform 1 0 6808 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _2042_
timestamp 1623621585
transform 1 0 7820 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1623621585
transform 1 0 9016 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_82
timestamp 1623621585
transform 1 0 8648 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_87
timestamp 1623621585
transform 1 0 9108 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_75
timestamp 1623621585
transform 1 0 8004 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_87
timestamp 1623621585
transform 1 0 9108 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _2245_
timestamp 1623621585
transform 1 0 11408 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1623621585
transform 1 0 11592 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_99
timestamp 1623621585
transform 1 0 10212 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1623621585
transform 1 0 11316 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_99
timestamp 1623621585
transform 1 0 10212 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_111
timestamp 1623621585
transform 1 0 11316 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1160_
timestamp 1623621585
transform 1 0 13156 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1189_
timestamp 1623621585
transform 1 0 13524 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1201_
timestamp 1623621585
transform 1 0 12052 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_131
timestamp 1623621585
transform 1 0 13156 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_115
timestamp 1623621585
transform 1 0 11684 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_127
timestamp 1623621585
transform 1 0 12788 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_134
timestamp 1623621585
transform 1 0 13432 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1103_
timestamp 1623621585
transform 1 0 15364 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2244_
timestamp 1623621585
transform 1 0 13800 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1623621585
transform 1 0 14260 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_139
timestamp 1623621585
transform 1 0 13892 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_144
timestamp 1623621585
transform 1 0 14352 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_152
timestamp 1623621585
transform 1 0 15088 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1623621585
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_157
timestamp 1623621585
transform 1 0 15548 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1177_
timestamp 1623621585
transform 1 0 16836 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1178_
timestamp 1623621585
transform 1 0 17756 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1182_
timestamp 1623621585
transform 1 0 15916 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1623621585
transform 1 0 16836 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_177
timestamp 1623621585
transform 1 0 17388 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_167
timestamp 1623621585
transform 1 0 16468 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_172
timestamp 1623621585
transform 1 0 16928 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _2254_
timestamp 1623621585
transform 1 0 18032 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1623621585
transform 1 0 19504 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_189
timestamp 1623621585
transform 1 0 18492 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_197
timestamp 1623621585
transform 1 0 19228 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_201
timestamp 1623621585
transform 1 0 19596 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_203
timestamp 1623621585
transform 1 0 19780 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__o21bai_1  _1576_
timestamp 1623621585
transform 1 0 21160 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1582_
timestamp 1623621585
transform 1 0 20884 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1623621585
transform 1 0 22080 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_213
timestamp 1623621585
transform 1 0 20700 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_221
timestamp 1623621585
transform 1 0 21436 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_215
timestamp 1623621585
transform 1 0 20884 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_224
timestamp 1623621585
transform 1 0 21712 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1581_
timestamp 1623621585
transform 1 0 22540 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1613_
timestamp 1623621585
transform 1 0 23920 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_39_233
timestamp 1623621585
transform 1 0 22540 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1623621585
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_229
timestamp 1623621585
transform 1 0 22172 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_236
timestamp 1623621585
transform 1 0 22816 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1623621585
transform 1 0 24748 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output219
timestamp 1623621585
transform 1 0 25852 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output236
timestamp 1623621585
transform 1 0 25944 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_258
timestamp 1623621585
transform 1 0 24840 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_274
timestamp 1623621585
transform 1 0 26312 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_255
timestamp 1623621585
transform 1 0 24564 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_267
timestamp 1623621585
transform 1 0 25668 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_273
timestamp 1623621585
transform 1 0 26220 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_4  _1641_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 26680 0 1 23392
box -38 -48 1418 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1623621585
transform 1 0 27324 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output192
timestamp 1623621585
transform 1 0 27876 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output201
timestamp 1623621585
transform 1 0 26588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1623621585
transform 1 0 28060 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_281
timestamp 1623621585
transform 1 0 26956 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_286
timestamp 1623621585
transform 1 0 27416 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_290
timestamp 1623621585
transform 1 0 27784 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_295
timestamp 1623621585
transform 1 0 28244 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1623621585
transform -1 0 28888 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1623621585
transform -1 0 28888 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _2111_
timestamp 1623621585
transform 1 0 1380 0 1 24480
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1623621585
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_21
timestamp 1623621585
transform 1 0 3036 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_2  _2117_
timestamp 1623621585
transform 1 0 4508 0 1 24480
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1623621585
transform 1 0 3772 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_30
timestamp 1623621585
transform 1 0 3864 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_36
timestamp 1623621585
transform 1 0 4416 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_55
timestamp 1623621585
transform 1 0 6164 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_67
timestamp 1623621585
transform 1 0 7268 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1623621585
transform 1 0 9016 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_79
timestamp 1623621585
transform 1 0 8372 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_85
timestamp 1623621585
transform 1 0 8924 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_87
timestamp 1623621585
transform 1 0 9108 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _2091_
timestamp 1623621585
transform 1 0 10212 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_41_108
timestamp 1623621585
transform 1 0 11040 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1200_
timestamp 1623621585
transform 1 0 11868 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _1203_
timestamp 1623621585
transform 1 0 13248 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_116
timestamp 1623621585
transform 1 0 11776 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_123
timestamp 1623621585
transform 1 0 12420 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_131
timestamp 1623621585
transform 1 0 13156 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _1184_
timestamp 1623621585
transform 1 0 15088 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1623621585
transform 1 0 14260 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_138
timestamp 1623621585
transform 1 0 13800 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_142
timestamp 1623621585
transform 1 0 14168 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_144
timestamp 1623621585
transform 1 0 14352 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_158
timestamp 1623621585
transform 1 0 15640 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1175_
timestamp 1623621585
transform 1 0 17480 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1183_
timestamp 1623621585
transform 1 0 16100 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_162
timestamp 1623621585
transform 1 0 16008 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_171
timestamp 1623621585
transform 1 0 16836 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_177
timestamp 1623621585
transform 1 0 17388 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_182
timestamp 1623621585
transform 1 0 17848 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__mux4_2  _2131_
timestamp 1623621585
transform 1 0 19964 0 1 24480
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1623621585
transform 1 0 19504 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_194
timestamp 1623621585
transform 1 0 18952 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_201
timestamp 1623621585
transform 1 0 19596 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1566_
timestamp 1623621585
transform 1 0 21988 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_223
timestamp 1623621585
transform 1 0 21620 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2163_
timestamp 1623621585
transform 1 0 22724 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_231
timestamp 1623621585
transform 1 0 22356 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_251
timestamp 1623621585
transform 1 0 24196 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2154_
timestamp 1623621585
transform 1 0 25208 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1623621585
transform 1 0 24748 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_258
timestamp 1623621585
transform 1 0 24840 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1643_
timestamp 1623621585
transform 1 0 27416 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_41_278
timestamp 1623621585
transform 1 0 26680 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_295
timestamp 1623621585
transform 1 0 28244 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1623621585
transform -1 0 28888 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1275_
timestamp 1623621585
transform 1 0 2392 0 -1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1623621585
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input145
timestamp 1623621585
transform 1 0 1656 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_3
timestamp 1623621585
transform 1 0 1380 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_10
timestamp 1623621585
transform 1 0 2024 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1216_
timestamp 1623621585
transform 1 0 3956 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1720_
timestamp 1623621585
transform 1 0 4692 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1623621585
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_35
timestamp 1623621585
transform 1 0 4324 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_42
timestamp 1623621585
transform 1 0 4968 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1623621585
transform 1 0 6348 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_54
timestamp 1623621585
transform 1 0 6072 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_58
timestamp 1623621585
transform 1 0 6440 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1333_
timestamp 1623621585
transform 1 0 7728 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1334_
timestamp 1623621585
transform 1 0 8372 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1337_
timestamp 1623621585
transform 1 0 9200 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_70
timestamp 1623621585
transform 1 0 7544 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_75
timestamp 1623621585
transform 1 0 8004 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_82
timestamp 1623621585
transform 1 0 8648 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_91
timestamp 1623621585
transform 1 0 9476 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1666_
timestamp 1623621585
transform 1 0 10580 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1623621585
transform 1 0 11592 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_106
timestamp 1623621585
transform 1 0 10856 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1161_
timestamp 1623621585
transform 1 0 12972 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1204_
timestamp 1623621585
transform 1 0 13708 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_115
timestamp 1623621585
transform 1 0 11684 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_127
timestamp 1623621585
transform 1 0 12788 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_133
timestamp 1623621585
transform 1 0 13340 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1185_
timestamp 1623621585
transform 1 0 15364 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_145
timestamp 1623621585
transform 1 0 14444 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_153
timestamp 1623621585
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1623621585
transform 1 0 16836 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_163
timestamp 1623621585
transform 1 0 16100 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_172
timestamp 1623621585
transform 1 0 16928 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1537_
timestamp 1623621585
transform 1 0 18308 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2178_
timestamp 1623621585
transform 1 0 19504 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_42_184
timestamp 1623621585
transform 1 0 18032 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_196
timestamp 1623621585
transform 1 0 19136 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1575_
timestamp 1623621585
transform 1 0 21344 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1623621585
transform 1 0 22080 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_216
timestamp 1623621585
transform 1 0 20976 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_224
timestamp 1623621585
transform 1 0 21712 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2ai_1  _1577_
timestamp 1623621585
transform 1 0 22540 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1614_
timestamp 1623621585
transform 1 0 24104 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_229
timestamp 1623621585
transform 1 0 22172 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_240
timestamp 1623621585
transform 1 0 23184 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_248
timestamp 1623621585
transform 1 0 23920 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux4_2  _2096_
timestamp 1623621585
transform 1 0 25300 0 -1 25568
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_42_259
timestamp 1623621585
transform 1 0 24932 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1623621585
transform 1 0 27324 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output210
timestamp 1623621585
transform 1 0 27876 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_281
timestamp 1623621585
transform 1 0 26956 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_286
timestamp 1623621585
transform 1 0 27416 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_290
timestamp 1623621585
transform 1 0 27784 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_295
timestamp 1623621585
transform 1 0 28244 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1623621585
transform -1 0 28888 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1365_
timestamp 1623621585
transform 1 0 2944 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1623621585
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input154
timestamp 1623621585
transform 1 0 1748 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1623621585
transform 1 0 1380 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_11
timestamp 1623621585
transform 1 0 2116 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_19
timestamp 1623621585
transform 1 0 2852 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_8  _1979_
timestamp 1623621585
transform 1 0 4324 0 1 25568
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1623621585
transform 1 0 3772 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_24
timestamp 1623621585
transform 1 0 3312 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_28
timestamp 1623621585
transform 1 0 3680 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_30
timestamp 1623621585
transform 1 0 3864 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_34
timestamp 1623621585
transform 1 0 4232 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1316_
timestamp 1623621585
transform 1 0 7360 0 1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__nand3_1  _1326_
timestamp 1623621585
transform 1 0 6624 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_56
timestamp 1623621585
transform 1 0 6256 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_64
timestamp 1623621585
transform 1 0 6992 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2226_
timestamp 1623621585
transform 1 0 9476 0 1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1623621585
transform 1 0 9016 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_82
timestamp 1623621585
transform 1 0 8648 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_87
timestamp 1623621585
transform 1 0 9108 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1964_
timestamp 1623621585
transform 1 0 11408 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1623621585
transform 1 0 11040 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1202_
timestamp 1623621585
transform 1 0 13064 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_121
timestamp 1623621585
transform 1 0 12236 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_129
timestamp 1623621585
transform 1 0 12972 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_134
timestamp 1623621585
transform 1 0 13432 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1053_
timestamp 1623621585
transform 1 0 14720 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1176_
timestamp 1623621585
transform 1 0 15548 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1623621585
transform 1 0 14260 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_142
timestamp 1623621585
transform 1 0 14168 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_144
timestamp 1623621585
transform 1 0 14352 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_152
timestamp 1623621585
transform 1 0 15088 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_156
timestamp 1623621585
transform 1 0 15456 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2252_
timestamp 1623621585
transform 1 0 16284 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_43_161
timestamp 1623621585
transform 1 0 15916 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1536_
timestamp 1623621585
transform 1 0 18400 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1623621585
transform 1 0 19504 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_184
timestamp 1623621585
transform 1 0 18032 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_195
timestamp 1623621585
transform 1 0 19044 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_199
timestamp 1623621585
transform 1 0 19412 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_201
timestamp 1623621585
transform 1 0 19596 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2162_
timestamp 1623621585
transform 1 0 21160 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_43_213
timestamp 1623621585
transform 1 0 20700 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_217
timestamp 1623621585
transform 1 0 21068 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output246
timestamp 1623621585
transform 1 0 24012 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_234
timestamp 1623621585
transform 1 0 22632 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_246
timestamp 1623621585
transform 1 0 23736 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1642_
timestamp 1623621585
transform 1 0 25760 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1623621585
transform 1 0 24748 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_253
timestamp 1623621585
transform 1 0 24380 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_258
timestamp 1623621585
transform 1 0 24840 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_266
timestamp 1623621585
transform 1 0 25576 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2146_
timestamp 1623621585
transform 1 0 26772 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 1623621585
transform 1 0 26404 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_295
timestamp 1623621585
transform 1 0 28244 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1623621585
transform -1 0 28888 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1229_
timestamp 1623621585
transform 1 0 2392 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1623621585
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1623621585
transform 1 0 1748 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input127
timestamp 1623621585
transform 1 0 3036 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1623621585
transform 1 0 1380 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_10
timestamp 1623621585
transform 1 0 2024 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_17
timestamp 1623621585
transform 1 0 2668 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1978_
timestamp 1623621585
transform 1 0 4140 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_44_24
timestamp 1623621585
transform 1 0 3312 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_32
timestamp 1623621585
transform 1 0 4048 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_42
timestamp 1623621585
transform 1 0 4968 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1623621585
transform 1 0 6348 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input136
timestamp 1623621585
transform 1 0 5336 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_49
timestamp 1623621585
transform 1 0 5612 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_58
timestamp 1623621585
transform 1 0 6440 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__xor2_1  _1335_
timestamp 1623621585
transform 1 0 7820 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1338_
timestamp 1623621585
transform 1 0 9016 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_70
timestamp 1623621585
transform 1 0 7544 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_80
timestamp 1623621585
transform 1 0 8464 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_90
timestamp 1623621585
transform 1 0 9384 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1668_
timestamp 1623621585
transform 1 0 9752 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1965_
timestamp 1623621585
transform 1 0 10396 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1623621585
transform 1 0 11592 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_97
timestamp 1623621585
transform 1 0 10028 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_110
timestamp 1623621585
transform 1 0 11224 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1015_
timestamp 1623621585
transform 1 0 12788 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_115
timestamp 1623621585
transform 1 0 11684 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_130
timestamp 1623621585
transform 1 0 13064 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1018_
timestamp 1623621585
transform 1 0 14352 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1836_
timestamp 1623621585
transform 1 0 15088 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_142
timestamp 1623621585
transform 1 0 14168 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_148
timestamp 1623621585
transform 1 0 14720 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_156
timestamp 1623621585
transform 1 0 15456 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1842_
timestamp 1623621585
transform 1 0 15824 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1623621585
transform 1 0 16836 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_164
timestamp 1623621585
transform 1 0 16192 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_170
timestamp 1623621585
transform 1 0 16744 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_172
timestamp 1623621585
transform 1 0 16928 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1533_
timestamp 1623621585
transform 1 0 18400 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_184
timestamp 1623621585
transform 1 0 18032 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_191
timestamp 1623621585
transform 1 0 18676 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_203
timestamp 1623621585
transform 1 0 19780 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1623621585
transform 1 0 22080 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_215
timestamp 1623621585
transform 1 0 20884 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_227
timestamp 1623621585
transform 1 0 21988 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_229
timestamp 1623621585
transform 1 0 22172 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_241
timestamp 1623621585
transform 1 0 23276 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output228
timestamp 1623621585
transform 1 0 25852 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output237
timestamp 1623621585
transform 1 0 25116 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1623621585
transform 1 0 24380 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_265
timestamp 1623621585
transform 1 0 25484 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_273
timestamp 1623621585
transform 1 0 26220 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1623621585
transform 1 0 27324 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output184
timestamp 1623621585
transform 1 0 27876 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output211
timestamp 1623621585
transform 1 0 26588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_281
timestamp 1623621585
transform 1 0 26956 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_286
timestamp 1623621585
transform 1 0 27416 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_290
timestamp 1623621585
transform 1 0 27784 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_295
timestamp 1623621585
transform 1 0 28244 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1623621585
transform -1 0 28888 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1623621585
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1623621585
transform 1 0 1748 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1623621585
transform 1 0 2392 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input128
timestamp 1623621585
transform 1 0 3036 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1623621585
transform 1 0 1380 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_10
timestamp 1623621585
transform 1 0 2024 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_17
timestamp 1623621585
transform 1 0 2668 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _2118_
timestamp 1623621585
transform 1 0 4508 0 1 26656
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1623621585
transform 1 0 3772 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_24
timestamp 1623621585
transform 1 0 3312 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_28
timestamp 1623621585
transform 1 0 3680 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_30
timestamp 1623621585
transform 1 0 3864 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_36
timestamp 1623621585
transform 1 0 4416 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_55
timestamp 1623621585
transform 1 0 6164 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_67
timestamp 1623621585
transform 1 0 7268 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1623621585
transform 1 0 9016 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_79
timestamp 1623621585
transform 1 0 8372 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_85
timestamp 1623621585
transform 1 0 8924 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_87
timestamp 1623621585
transform 1 0 9108 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1667_
timestamp 1623621585
transform 1 0 10856 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_99
timestamp 1623621585
transform 1 0 10212 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_105
timestamp 1623621585
transform 1 0 10764 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_109
timestamp 1623621585
transform 1 0 11132 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1826_
timestamp 1623621585
transform 1 0 11868 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1831_
timestamp 1623621585
transform 1 0 12788 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1837_
timestamp 1623621585
transform 1 0 13524 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_123
timestamp 1623621585
transform 1 0 12420 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_131
timestamp 1623621585
transform 1 0 13156 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1830_
timestamp 1623621585
transform 1 0 14720 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1623621585
transform 1 0 14260 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_139
timestamp 1623621585
transform 1 0 13892 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_144
timestamp 1623621585
transform 1 0 14352 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_152
timestamp 1623621585
transform 1 0 15088 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_2  _2124_
timestamp 1623621585
transform 1 0 16008 0 1 26656
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_45_160
timestamp 1623621585
transform 1 0 15824 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_180
timestamp 1623621585
transform 1 0 17664 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _1534_
timestamp 1623621585
transform 1 0 18492 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1623621585
transform 1 0 19504 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_188
timestamp 1623621585
transform 1 0 18400 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_195
timestamp 1623621585
transform 1 0 19044 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_199
timestamp 1623621585
transform 1 0 19412 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_201
timestamp 1623621585
transform 1 0 19596 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__mux4_2  _2138_
timestamp 1623621585
transform 1 0 22080 0 1 26656
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_45_213
timestamp 1623621585
transform 1 0 20700 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_225
timestamp 1623621585
transform 1 0 21804 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_246
timestamp 1623621585
transform 1 0 23736 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1608_
timestamp 1623621585
transform 1 0 25208 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1623621585
transform 1 0 24748 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_254
timestamp 1623621585
transform 1 0 24472 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_258
timestamp 1623621585
transform 1 0 24840 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_266
timestamp 1623621585
transform 1 0 25576 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_274
timestamp 1623621585
transform 1 0 26312 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__o21bai_1  _1639_
timestamp 1623621585
transform 1 0 27232 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output193
timestamp 1623621585
transform 1 0 26496 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_280
timestamp 1623621585
transform 1 0 26864 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_290
timestamp 1623621585
transform 1 0 27784 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1623621585
transform -1 0 28888 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_298
timestamp 1623621585
transform 1 0 28520 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _2020_
timestamp 1623621585
transform 1 0 2576 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _2112_
timestamp 1623621585
transform 1 0 1380 0 -1 27744
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1623621585
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1623621585
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1623621585
transform 1 0 1748 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_21
timestamp 1623621585
transform 1 0 3036 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1623621585
transform 1 0 1380 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_10
timestamp 1623621585
transform 1 0 2024 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1781_
timestamp 1623621585
transform 1 0 4232 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2019_
timestamp 1623621585
transform 1 0 3404 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1623621585
transform 1 0 3772 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input137
timestamp 1623621585
transform 1 0 4876 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_34
timestamp 1623621585
transform 1 0 4232 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_25
timestamp 1623621585
transform 1 0 3404 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_30
timestamp 1623621585
transform 1 0 3864 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_37
timestamp 1623621585
transform 1 0 4508 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_44
timestamp 1623621585
transform 1 0 5152 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_52
timestamp 1623621585
transform 1 0 5888 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_54
timestamp 1623621585
transform 1 0 6072 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_46
timestamp 1623621585
transform 1 0 5336 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1331_
timestamp 1623621585
transform 1 0 6072 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1623621585
transform 1 0 6348 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_62
timestamp 1623621585
transform 1 0 6808 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_58
timestamp 1623621585
transform 1 0 6440 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1623621585
transform 1 0 6348 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_1  _1329_
timestamp 1623621585
transform 1 0 6716 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1327_
timestamp 1623621585
transform 1 0 6900 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_67
timestamp 1623621585
transform 1 0 7268 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_67
timestamp 1623621585
transform 1 0 7268 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_78
timestamp 1623621585
transform 1 0 8280 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_75
timestamp 1623621585
transform 1 0 8004 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1330_
timestamp 1623621585
transform 1 0 7636 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1317_
timestamp 1623621585
transform 1 0 8372 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _1310_
timestamp 1623621585
transform 1 0 7636 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_47_87
timestamp 1623621585
transform 1 0 9108 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_82
timestamp 1623621585
transform 1 0 8648 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1623621585
transform 1 0 9016 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1750_
timestamp 1623621585
transform 1 0 9016 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1328_
timestamp 1623621585
transform 1 0 9476 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_89
timestamp 1623621585
transform 1 0 9292 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_1  _1827_
timestamp 1623621585
transform 1 0 11592 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2094_
timestamp 1623621585
transform 1 0 10120 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1623621585
transform 1 0 11592 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_101
timestamp 1623621585
transform 1 0 10396 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_113
timestamp 1623621585
transform 1 0 11500 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_94
timestamp 1623621585
transform 1 0 9752 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_107
timestamp 1623621585
transform 1 0 10948 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_113
timestamp 1623621585
transform 1 0 11500 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _1051_
timestamp 1623621585
transform 1 0 12972 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _1833_
timestamp 1623621585
transform 1 0 13156 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1834_
timestamp 1623621585
transform 1 0 12052 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_115
timestamp 1623621585
transform 1 0 11684 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_127
timestamp 1623621585
transform 1 0 12788 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_137
timestamp 1623621585
transform 1 0 13708 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_122
timestamp 1623621585
transform 1 0 12328 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_128
timestamp 1623621585
transform 1 0 12880 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_135
timestamp 1623621585
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2251_
timestamp 1623621585
transform 1 0 15272 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1623621585
transform 1 0 14260 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 14628 0 -1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_46_145
timestamp 1623621585
transform 1 0 14444 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_144
timestamp 1623621585
transform 1 0 14352 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_152
timestamp 1623621585
transform 1 0 15088 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1528_
timestamp 1623621585
transform 1 0 17664 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _2125_
timestamp 1623621585
transform 1 0 17388 0 1 27744
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1623621585
transform 1 0 16836 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_2
timestamp 1623621585
transform 1 0 17204 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_167
timestamp 1623621585
transform 1 0 16468 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_172
timestamp 1623621585
transform 1 0 16928 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_173
timestamp 1623621585
transform 1 0 17020 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__nor3b_4  _1532_
timestamp 1623621585
transform 1 0 18308 0 -1 27744
box -38 -48 1418 592
use sky130_fd_sc_hd__mux4_2  _2132_
timestamp 1623621585
transform 1 0 19964 0 1 27744
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1623621585
transform 1 0 19504 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_183
timestamp 1623621585
transform 1 0 17940 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_202
timestamp 1623621585
transform 1 0 19688 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_195
timestamp 1623621585
transform 1 0 19044 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_199
timestamp 1623621585
transform 1 0 19412 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_201
timestamp 1623621585
transform 1 0 19596 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2ai_1  _1535_
timestamp 1623621585
transform 1 0 20056 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1623621585
transform 1 0 22080 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_213
timestamp 1623621585
transform 1 0 20700 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_225
timestamp 1623621585
transform 1 0 21804 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_223
timestamp 1623621585
transform 1 0 21620 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__o31ai_1  _1610_
timestamp 1623621585
transform 1 0 23828 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _2139_
timestamp 1623621585
transform 1 0 22540 0 -1 27744
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_46_229
timestamp 1623621585
transform 1 0 22172 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_251
timestamp 1623621585
transform 1 0 24196 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_235
timestamp 1623621585
transform 1 0 22724 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__a31oi_1  _1606_
timestamp 1623621585
transform 1 0 25576 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1607_
timestamp 1623621585
transform 1 0 24564 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_2  _2095_
timestamp 1623621585
transform 1 0 25392 0 1 27744
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1623621585
transform 1 0 24748 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_262
timestamp 1623621585
transform 1 0 25208 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_271
timestamp 1623621585
transform 1 0 26036 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_253
timestamp 1623621585
transform 1 0 24380 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_258
timestamp 1623621585
transform 1 0 24840 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1636_
timestamp 1623621585
transform 1 0 27416 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1638_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 27784 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1623621585
transform 1 0 27324 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output202
timestamp 1623621585
transform 1 0 26588 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_281
timestamp 1623621585
transform 1 0 26956 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_286
timestamp 1623621585
transform 1 0 27416 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_295
timestamp 1623621585
transform 1 0 28244 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_282
timestamp 1623621585
transform 1 0 27048 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_293
timestamp 1623621585
transform 1 0 28060 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1623621585
transform -1 0 28888 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1623621585
transform -1 0 28888 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1369_
timestamp 1623621585
transform 1 0 2484 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1780_
timestamp 1623621585
transform 1 0 3128 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1623621585
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input146
timestamp 1623621585
transform 1 0 1748 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1623621585
transform 1 0 1380 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_11
timestamp 1623621585
transform 1 0 2116 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_18
timestamp 1623621585
transform 1 0 2760 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1266_
timestamp 1623621585
transform 1 0 4324 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1715_
timestamp 1623621585
transform 1 0 4968 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_25
timestamp 1623621585
transform 1 0 3404 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_33
timestamp 1623621585
transform 1 0 4140 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_38
timestamp 1623621585
transform 1 0 4600 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_45
timestamp 1623621585
transform 1 0 5244 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1319_
timestamp 1623621585
transform 1 0 6992 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1332_
timestamp 1623621585
transform 1 0 5704 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1623621585
transform 1 0 6348 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_49
timestamp 1623621585
transform 1 0 5612 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_53
timestamp 1623621585
transform 1 0 5980 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_58
timestamp 1623621585
transform 1 0 6440 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2043_
timestamp 1623621585
transform 1 0 9108 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2044_
timestamp 1623621585
transform 1 0 7912 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_70
timestamp 1623621585
transform 1 0 7544 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_83
timestamp 1623621585
transform 1 0 8740 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1966_
timestamp 1623621585
transform 1 0 10304 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1623621585
transform 1 0 11592 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_96
timestamp 1623621585
transform 1 0 9936 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_109
timestamp 1623621585
transform 1 0 11132 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_113
timestamp 1623621585
transform 1 0 11500 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1660_
timestamp 1623621585
transform 1 0 12052 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  _1817_
timestamp 1623621585
transform 1 0 13708 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_115
timestamp 1623621585
transform 1 0 11684 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_122
timestamp 1623621585
transform 1 0 12328 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_134
timestamp 1623621585
transform 1 0 13432 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1843_
timestamp 1623621585
transform 1 0 15180 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_145
timestamp 1623621585
transform 1 0 14444 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_157
timestamp 1623621585
transform 1 0 15548 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1623621585
transform 1 0 16836 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_169
timestamp 1623621585
transform 1 0 16652 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_172
timestamp 1623621585
transform 1 0 16928 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1527_
timestamp 1623621585
transform 1 0 18860 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2179_
timestamp 1623621585
transform 1 0 19964 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_48_184
timestamp 1623621585
transform 1 0 18032 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_192
timestamp 1623621585
transform 1 0 18768 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp 1623621585
transform 1 0 19228 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1623621585
transform 1 0 22080 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_221
timestamp 1623621585
transform 1 0 21436 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_227
timestamp 1623621585
transform 1 0 21988 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_229
timestamp 1623621585
transform 1 0 22172 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_241
timestamp 1623621585
transform 1 0 23276 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1609_
timestamp 1623621585
transform 1 0 24748 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2155_
timestamp 1623621585
transform 1 0 25392 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1623621585
transform 1 0 24380 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_260
timestamp 1623621585
transform 1 0 25024 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1637_
timestamp 1623621585
transform 1 0 27876 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1623621585
transform 1 0 27324 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_280
timestamp 1623621585
transform 1 0 26864 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_284
timestamp 1623621585
transform 1 0 27232 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_286
timestamp 1623621585
transform 1 0 27416 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_290
timestamp 1623621585
transform 1 0 27784 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_295
timestamp 1623621585
transform 1 0 28244 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1623621585
transform -1 0 28888 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2215_
timestamp 1623621585
transform 1 0 1380 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1623621585
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_19
timestamp 1623621585
transform 1 0 2852 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1980_
timestamp 1623621585
transform 1 0 4232 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1623621585
transform 1 0 3772 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_27
timestamp 1623621585
transform 1 0 3588 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_30
timestamp 1623621585
transform 1 0 3864 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_43
timestamp 1623621585
transform 1 0 5060 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2227_
timestamp 1623621585
transform 1 0 5428 0 1 28832
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_49_64
timestamp 1623621585
transform 1 0 6992 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1318_
timestamp 1623621585
transform 1 0 7912 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1623621585
transform 1 0 9016 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_72
timestamp 1623621585
transform 1 0 7728 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_79
timestamp 1623621585
transform 1 0 8372 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_85
timestamp 1623621585
transform 1 0 8924 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_87
timestamp 1623621585
transform 1 0 9108 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1661_
timestamp 1623621585
transform 1 0 9752 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _1967_
timestamp 1623621585
transform 1 0 10396 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_93
timestamp 1623621585
transform 1 0 9660 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_97
timestamp 1623621585
transform 1 0 10028 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_113
timestamp 1623621585
transform 1 0 11500 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1662_
timestamp 1623621585
transform 1 0 11868 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_120
timestamp 1623621585
transform 1 0 12144 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_132
timestamp 1623621585
transform 1 0 13248 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _1845_
timestamp 1623621585
transform 1 0 14996 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1623621585
transform 1 0 14260 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_140
timestamp 1623621585
transform 1 0 13984 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_144
timestamp 1623621585
transform 1 0 14352 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_150
timestamp 1623621585
transform 1 0 14904 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_155
timestamp 1623621585
transform 1 0 15364 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_167
timestamp 1623621585
transform 1 0 16468 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_179
timestamp 1623621585
transform 1 0 17572 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1623621585
transform 1 0 19504 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_191
timestamp 1623621585
transform 1 0 18676 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_199
timestamp 1623621585
transform 1 0 19412 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_201
timestamp 1623621585
transform 1 0 19596 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_213
timestamp 1623621585
transform 1 0 20700 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1623621585
transform 1 0 21804 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1623621585
transform 1 0 22908 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_249
timestamp 1623621585
transform 1 0 24012 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1623621585
transform 1 0 24748 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output229
timestamp 1623621585
transform 1 0 26128 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output247
timestamp 1623621585
transform 1 0 25392 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_258
timestamp 1623621585
transform 1 0 24840 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_268
timestamp 1623621585
transform 1 0 25760 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2ai_1  _1640_
timestamp 1623621585
transform 1 0 27600 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output220
timestamp 1623621585
transform 1 0 26864 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1623621585
transform 1 0 26496 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_284
timestamp 1623621585
transform 1 0 27232 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_295
timestamp 1623621585
transform 1 0 28244 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1623621585
transform -1 0 28888 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1370_
timestamp 1623621585
transform 1 0 1748 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _2233_
timestamp 1623621585
transform 1 0 3128 0 -1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1623621585
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1623621585
transform 1 0 1380 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_16
timestamp 1623621585
transform 1 0 2576 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2070_
timestamp 1623621585
transform 1 0 5152 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_39
timestamp 1623621585
transform 1 0 4692 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_43
timestamp 1623621585
transform 1 0 5060 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1623621585
transform 1 0 6348 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_53
timestamp 1623621585
transform 1 0 5980 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_58
timestamp 1623621585
transform 1 0 6440 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2202_
timestamp 1623621585
transform 1 0 8188 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_50_70
timestamp 1623621585
transform 1 0 7544 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_76
timestamp 1623621585
transform 1 0 8096 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1443_
timestamp 1623621585
transform 1 0 10028 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1623621585
transform 1 0 11592 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_93
timestamp 1623621585
transform 1 0 9660 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_106
timestamp 1623621585
transform 1 0 10856 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _1158_
timestamp 1623621585
transform 1 0 13432 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_50_115
timestamp 1623621585
transform 1 0 11684 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_127
timestamp 1623621585
transform 1 0 12788 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_133
timestamp 1623621585
transform 1 0 13340 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _1846_
timestamp 1623621585
transform 1 0 14996 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_147
timestamp 1623621585
transform 1 0 14628 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_157
timestamp 1623621585
transform 1 0 15548 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1847_
timestamp 1623621585
transform 1 0 15916 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1623621585
transform 1 0 16836 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_164
timestamp 1623621585
transform 1 0 16192 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_170
timestamp 1623621585
transform 1 0 16744 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_172
timestamp 1623621585
transform 1 0 16928 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_184
timestamp 1623621585
transform 1 0 18032 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_196
timestamp 1623621585
transform 1 0 19136 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1623621585
transform 1 0 22080 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_208
timestamp 1623621585
transform 1 0 20240 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_220
timestamp 1623621585
transform 1 0 21344 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_229
timestamp 1623621585
transform 1 0 22172 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_241
timestamp 1623621585
transform 1 0 23276 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1623621585
transform 1 0 25944 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1623621585
transform 1 0 24380 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_265
timestamp 1623621585
transform 1 0 25484 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_269
timestamp 1623621585
transform 1 0 25852 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_273
timestamp 1623621585
transform 1 0 26220 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1878_
timestamp 1623621585
transform 1 0 27876 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1623621585
transform 1 0 27324 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output238
timestamp 1623621585
transform 1 0 26588 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_281
timestamp 1623621585
transform 1 0 26956 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_286
timestamp 1623621585
transform 1 0 27416 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_290
timestamp 1623621585
transform 1 0 27784 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_295
timestamp 1623621585
transform 1 0 28244 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1623621585
transform -1 0 28888 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1271_
timestamp 1623621585
transform 1 0 3036 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1623621585
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input155
timestamp 1623621585
transform 1 0 1748 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1623621585
transform 1 0 1380 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_11
timestamp 1623621585
transform 1 0 2116 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_19
timestamp 1623621585
transform 1 0 2852 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_4  _1981_
timestamp 1623621585
transform 1 0 4508 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1623621585
transform 1 0 3772 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_25
timestamp 1623621585
transform 1 0 3404 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_30
timestamp 1623621585
transform 1 0 3864 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_36
timestamp 1623621585
transform 1 0 4416 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1710_
timestamp 1623621585
transform 1 0 5980 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1711_
timestamp 1623621585
transform 1 0 6624 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_49
timestamp 1623621585
transform 1 0 5612 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_56
timestamp 1623621585
transform 1 0 6256 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_63
timestamp 1623621585
transform 1 0 6900 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1623621585
transform 1 0 9016 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_75
timestamp 1623621585
transform 1 0 8004 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_83
timestamp 1623621585
transform 1 0 8740 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_87
timestamp 1623621585
transform 1 0 9108 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_91
timestamp 1623621585
transform 1 0 9476 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1751_
timestamp 1623621585
transform 1 0 9568 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_95
timestamp 1623621585
transform 1 0 9844 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_107
timestamp 1623621585
transform 1 0 10948 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__o2111ai_4  _1822_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 11868 0 1 29920
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_51_115
timestamp 1623621585
transform 1 0 11684 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_2  _1814_
timestamp 1623621585
transform 1 0 14720 0 1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1829_
timestamp 1623621585
transform 1 0 15548 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1623621585
transform 1 0 14260 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_138
timestamp 1623621585
transform 1 0 13800 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_142
timestamp 1623621585
transform 1 0 14168 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_144
timestamp 1623621585
transform 1 0 14352 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_153
timestamp 1623621585
transform 1 0 15180 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1110_
timestamp 1623621585
transform 1 0 17480 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1849_
timestamp 1623621585
transform 1 0 16284 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_161
timestamp 1623621585
transform 1 0 15916 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1623621585
transform 1 0 16652 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_177
timestamp 1623621585
transform 1 0 17388 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_181
timestamp 1623621585
transform 1 0 17756 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1173_
timestamp 1623621585
transform 1 0 18492 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1623621585
transform 1 0 19504 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_195
timestamp 1623621585
transform 1 0 19044 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_199
timestamp 1623621585
transform 1 0 19412 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_201
timestamp 1623621585
transform 1 0 19596 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1171_
timestamp 1623621585
transform 1 0 20332 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2256_
timestamp 1623621585
transform 1 0 21436 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_51_217
timestamp 1623621585
transform 1 0 21068 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1163_
timestamp 1623621585
transform 1 0 23552 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_240
timestamp 1623621585
transform 1 0 23184 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_250
timestamp 1623621585
transform 1 0 24104 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1623621585
transform 1 0 24748 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1623621585
transform 1 0 26128 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1623621585
transform 1 0 25484 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_256
timestamp 1623621585
transform 1 0 24656 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_258
timestamp 1623621585
transform 1 0 24840 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_264
timestamp 1623621585
transform 1 0 25392 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_268
timestamp 1623621585
transform 1 0 25760 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1879_
timestamp 1623621585
transform 1 0 27876 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1880_
timestamp 1623621585
transform 1 0 26772 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_275
timestamp 1623621585
transform 1 0 26404 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_283
timestamp 1623621585
transform 1 0 27140 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_295
timestamp 1623621585
transform 1 0 28244 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1623621585
transform -1 0 28888 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_7
timestamp 1623621585
transform 1 0 1748 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1623621585
transform 1 0 1380 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output271
timestamp 1623621585
transform 1 0 1380 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output249
timestamp 1623621585
transform 1 0 1748 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1623621585
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1623621585
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_17
timestamp 1623621585
transform 1 0 2668 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_11
timestamp 1623621585
transform 1 0 2116 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output260
timestamp 1623621585
transform 1 0 2484 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1234_
timestamp 1623621585
transform 1 0 2116 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_19
timestamp 1623621585
transform 1 0 2852 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output282
timestamp 1623621585
transform 1 0 3036 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_30
timestamp 1623621585
transform 1 0 3864 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_25
timestamp 1623621585
transform 1 0 3404 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_27
timestamp 1623621585
transform 1 0 3588 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1623621585
transform 1 0 3772 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1047_
timestamp 1623621585
transform 1 0 3772 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_40
timestamp 1623621585
transform 1 0 4784 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_33
timestamp 1623621585
transform 1 0 4140 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output293
timestamp 1623621585
transform 1 0 4508 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1273_
timestamp 1623621585
transform 1 0 4232 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_41
timestamp 1623621585
transform 1 0 4876 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output304
timestamp 1623621585
transform 1 0 5244 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1623621585
transform 1 0 5888 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_48
timestamp 1623621585
transform 1 0 5520 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_49
timestamp 1623621585
transform 1 0 5612 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1623621585
transform 1 0 6348 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1705_
timestamp 1623621585
transform 1 0 6256 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1704_
timestamp 1623621585
transform 1 0 5612 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_59
timestamp 1623621585
transform 1 0 6532 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_66
timestamp 1623621585
transform 1 0 7176 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_58
timestamp 1623621585
transform 1 0 6440 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1795_
timestamp 1623621585
transform 1 0 6900 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_4  _1798_
timestamp 1623621585
transform 1 0 7268 0 -1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1796_
timestamp 1623621585
transform 1 0 7820 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1623621585
transform 1 0 9016 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_84
timestamp 1623621585
transform 1 0 8832 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_69
timestamp 1623621585
transform 1 0 7452 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_76
timestamp 1623621585
transform 1 0 8096 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_84
timestamp 1623621585
transform 1 0 8832 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_87
timestamp 1623621585
transform 1 0 9108 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2293_
timestamp 1623621585
transform 1 0 9752 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1623621585
transform 1 0 11592 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_96
timestamp 1623621585
transform 1 0 9936 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_108
timestamp 1623621585
transform 1 0 11040 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_93
timestamp 1623621585
transform 1 0 9660 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_113
timestamp 1623621585
transform 1 0 11500 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1054_
timestamp 1623621585
transform 1 0 13432 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1157_
timestamp 1623621585
transform 1 0 12972 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_2  _1819_
timestamp 1623621585
transform 1 0 12052 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_2  _1821_
timestamp 1623621585
transform 1 0 11868 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_115
timestamp 1623621585
transform 1 0 11684 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_128
timestamp 1623621585
transform 1 0 12880 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_125
timestamp 1623621585
transform 1 0 12604 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_133
timestamp 1623621585
transform 1 0 13340 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1111_
timestamp 1623621585
transform 1 0 15088 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _2276_
timestamp 1623621585
transform 1 0 15364 0 1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1623621585
transform 1 0 14260 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_147
timestamp 1623621585
transform 1 0 14628 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_151
timestamp 1623621585
transform 1 0 14996 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_158
timestamp 1623621585
transform 1 0 15640 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_141
timestamp 1623621585
transform 1 0 14076 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_144
timestamp 1623621585
transform 1 0 14352 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_152
timestamp 1623621585
transform 1 0 15088 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1815_
timestamp 1623621585
transform 1 0 16008 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1850_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 17296 0 1 31008
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1852_
timestamp 1623621585
transform 1 0 17296 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1623621585
transform 1 0 16836 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_166
timestamp 1623621585
transform 1 0 16376 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_170
timestamp 1623621585
transform 1 0 16744 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_172
timestamp 1623621585
transform 1 0 16928 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_172
timestamp 1623621585
transform 1 0 16928 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_186
timestamp 1623621585
transform 1 0 18216 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1623621585
transform 1 0 18768 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_187
timestamp 1623621585
transform 1 0 18308 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_183
timestamp 1623621585
transform 1 0 17940 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1162_
timestamp 1623621585
transform 1 0 18768 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1159_
timestamp 1623621585
transform 1 0 18400 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_201
timestamp 1623621585
transform 1 0 19596 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_196
timestamp 1623621585
transform 1 0 19136 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_204
timestamp 1623621585
transform 1 0 19872 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1623621585
transform 1 0 19504 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1174_
timestamp 1623621585
transform 1 0 19136 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2255_
timestamp 1623621585
transform 1 0 19964 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__nand3b_1  _1170_
timestamp 1623621585
transform 1 0 20700 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1623621585
transform 1 0 22080 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_212
timestamp 1623621585
transform 1 0 20608 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_219
timestamp 1623621585
transform 1 0 21252 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_227
timestamp 1623621585
transform 1 0 21988 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_224
timestamp 1623621585
transform 1 0 21712 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_228
timestamp 1623621585
transform 1 0 22080 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1164_
timestamp 1623621585
transform 1 0 23644 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1167_
timestamp 1623621585
transform 1 0 22816 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1169_
timestamp 1623621585
transform 1 0 22172 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2258_
timestamp 1623621585
transform 1 0 23920 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_52_229
timestamp 1623621585
transform 1 0 22172 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_235
timestamp 1623621585
transform 1 0 22724 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_244
timestamp 1623621585
transform 1 0 23552 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_237
timestamp 1623621585
transform 1 0 22908 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2259_
timestamp 1623621585
transform 1 0 25208 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1623621585
transform 1 0 24748 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_267
timestamp 1623621585
transform 1 0 25668 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_253
timestamp 1623621585
transform 1 0 24380 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_258
timestamp 1623621585
transform 1 0 24840 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_281
timestamp 1623621585
transform 1 0 26956 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_281
timestamp 1623621585
transform 1 0 26956 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_275
timestamp 1623621585
transform 1 0 26404 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  _1881_
timestamp 1623621585
transform 1 0 26588 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_289
timestamp 1623621585
transform 1 0 27692 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_286
timestamp 1623621585
transform 1 0 27416 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1623621585
transform 1 0 27324 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1882_
timestamp 1623621585
transform 1 0 27324 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_295
timestamp 1623621585
transform 1 0 28244 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1623621585
transform 1 0 27968 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1623621585
transform -1 0 28888 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1623621585
transform -1 0 28888 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_297
timestamp 1623621585
transform 1 0 28428 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1235_
timestamp 1623621585
transform 1 0 1380 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1272_
timestamp 1623621585
transform 1 0 2024 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _2232_
timestamp 1623621585
transform 1 0 2944 0 -1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1623621585
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_6
timestamp 1623621585
transform 1 0 1656 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_16
timestamp 1623621585
transform 1 0 2576 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1982_
timestamp 1623621585
transform 1 0 4876 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_54_37
timestamp 1623621585
transform 1 0 4508 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1293_
timestamp 1623621585
transform 1 0 6808 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1623621585
transform 1 0 6348 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_50
timestamp 1623621585
transform 1 0 5704 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_56
timestamp 1623621585
transform 1 0 6256 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_58
timestamp 1623621585
transform 1 0 6440 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1748_
timestamp 1623621585
transform 1 0 8740 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1797_
timestamp 1623621585
transform 1 0 7820 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_69
timestamp 1623621585
transform 1 0 7452 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_79
timestamp 1623621585
transform 1 0 8372 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_86
timestamp 1623621585
transform 1 0 9016 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1049_
timestamp 1623621585
transform 1 0 10488 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1623621585
transform 1 0 11592 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_98
timestamp 1623621585
transform 1 0 10120 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_105
timestamp 1623621585
transform 1 0 10764 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_113
timestamp 1623621585
transform 1 0 11500 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1014_
timestamp 1623621585
transform 1 0 12144 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1623621585
transform 1 0 13524 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1818_
timestamp 1623621585
transform 1 0 12788 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_115
timestamp 1623621585
transform 1 0 11684 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_119
timestamp 1623621585
transform 1 0 12052 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_123
timestamp 1623621585
transform 1 0 12420 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_131
timestamp 1623621585
transform 1 0 13156 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1112_
timestamp 1623621585
transform 1 0 15548 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_2  _1839_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 14260 0 -1 32096
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_54_138
timestamp 1623621585
transform 1 0 13800 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_142
timestamp 1623621585
transform 1 0 14168 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_153
timestamp 1623621585
transform 1 0 15180 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 17296 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1623621585
transform 1 0 16836 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_165
timestamp 1623621585
transform 1 0 16284 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_172
timestamp 1623621585
transform 1 0 16928 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1854_
timestamp 1623621585
transform 1 0 18308 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_54_183
timestamp 1623621585
transform 1 0 17940 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_194
timestamp 1623621585
transform 1 0 18952 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3b_1  _1168_
timestamp 1623621585
transform 1 0 21160 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1623621585
transform 1 0 22080 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_206
timestamp 1623621585
transform 1 0 20056 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_224
timestamp 1623621585
transform 1 0 21712 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1166_
timestamp 1623621585
transform 1 0 22816 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1623621585
transform 1 0 24104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_229
timestamp 1623621585
transform 1 0 22172 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_235
timestamp 1623621585
transform 1 0 22724 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_242
timestamp 1623621585
transform 1 0 23368 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1855_
timestamp 1623621585
transform 1 0 24748 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1623621585
transform 1 0 25944 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1623621585
transform 1 0 24380 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_261
timestamp 1623621585
transform 1 0 25116 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_269
timestamp 1623621585
transform 1 0 25852 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_273
timestamp 1623621585
transform 1 0 26220 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1883_
timestamp 1623621585
transform 1 0 27784 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1884_
timestamp 1623621585
transform 1 0 26588 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1623621585
transform 1 0 27324 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_281
timestamp 1623621585
transform 1 0 26956 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_286
timestamp 1623621585
transform 1 0 27416 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_294
timestamp 1623621585
transform 1 0 28152 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1623621585
transform -1 0 28888 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_298
timestamp 1623621585
transform 1 0 28520 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o2111ai_4  _1250_
timestamp 1623621585
transform 1 0 1472 0 1 32096
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1623621585
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_3
timestamp 1623621585
transform 1 0 1380 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _1983_
timestamp 1623621585
transform 1 0 4692 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1623621585
transform 1 0 3772 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_25
timestamp 1623621585
transform 1 0 3404 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_30
timestamp 1623621585
transform 1 0 3864 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_38
timestamp 1623621585
transform 1 0 4600 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1984_
timestamp 1623621585
transform 1 0 5888 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1985_
timestamp 1623621585
transform 1 0 7084 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_55_48
timestamp 1623621585
transform 1 0 5520 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_61
timestamp 1623621585
transform 1 0 6716 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1441_
timestamp 1623621585
transform 1 0 8280 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2045_
timestamp 1623621585
transform 1 0 9476 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1623621585
transform 1 0 9016 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_74
timestamp 1623621585
transform 1 0 7912 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_81
timestamp 1623621585
transform 1 0 8556 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_85
timestamp 1623621585
transform 1 0 8924 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_87
timestamp 1623621585
transform 1 0 9108 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1046_
timestamp 1623621585
transform 1 0 10672 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_100
timestamp 1623621585
transform 1 0 10304 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_112
timestamp 1623621585
transform 1 0 11408 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1050_
timestamp 1623621585
transform 1 0 11776 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1057_
timestamp 1623621585
transform 1 0 13340 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_124
timestamp 1623621585
transform 1 0 12512 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_132
timestamp 1623621585
transform 1 0 13248 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1623621585
transform 1 0 14260 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_139
timestamp 1623621585
transform 1 0 13892 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_144
timestamp 1623621585
transform 1 0 14352 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_156
timestamp 1623621585
transform 1 0 15456 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1820_
timestamp 1623621585
transform 1 0 15824 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1853_
timestamp 1623621585
transform 1 0 17388 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_55_164
timestamp 1623621585
transform 1 0 16192 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_176
timestamp 1623621585
transform 1 0 17296 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _1857_
timestamp 1623621585
transform 1 0 18492 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1623621585
transform 1 0 19504 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_184
timestamp 1623621585
transform 1 0 18032 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_188
timestamp 1623621585
transform 1 0 18400 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_196
timestamp 1623621585
transform 1 0 19136 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_201
timestamp 1623621585
transform 1 0 19596 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1859_
timestamp 1623621585
transform 1 0 20240 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1862_
timestamp 1623621585
transform 1 0 21252 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_55_207
timestamp 1623621585
transform 1 0 20148 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_215
timestamp 1623621585
transform 1 0 20884 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_226
timestamp 1623621585
transform 1 0 21896 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _1864_
timestamp 1623621585
transform 1 0 23644 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1623621585
transform 1 0 23000 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_241
timestamp 1623621585
transform 1 0 23276 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1867_
timestamp 1623621585
transform 1 0 25208 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1623621585
transform 1 0 24748 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_252
timestamp 1623621585
transform 1 0 24288 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_256
timestamp 1623621585
transform 1 0 24656 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_258
timestamp 1623621585
transform 1 0 24840 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_269
timestamp 1623621585
transform 1 0 25852 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2147_
timestamp 1623621585
transform 1 0 26772 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_55_277
timestamp 1623621585
transform 1 0 26588 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_295
timestamp 1623621585
transform 1 0 28244 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1623621585
transform -1 0 28888 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _1233_
timestamp 1623621585
transform 1 0 1380 0 -1 33184
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1623621585
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1274_
timestamp 1623621585
transform 1 0 3772 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1722_
timestamp 1623621585
transform 1 0 4784 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_25
timestamp 1623621585
transform 1 0 3404 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_36
timestamp 1623621585
transform 1 0 4416 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_43
timestamp 1623621585
transform 1 0 5060 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1623621585
transform 1 0 6348 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_55
timestamp 1623621585
transform 1 0 6164 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_58
timestamp 1623621585
transform 1 0 6440 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1749_
timestamp 1623621585
transform 1 0 9476 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2046_
timestamp 1623621585
transform 1 0 8280 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_56_70
timestamp 1623621585
transform 1 0 7544 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_87
timestamp 1623621585
transform 1 0 9108 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1045_
timestamp 1623621585
transform 1 0 10672 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1623621585
transform 1 0 11592 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_94
timestamp 1623621585
transform 1 0 9752 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_102
timestamp 1623621585
transform 1 0 10488 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_107
timestamp 1623621585
transform 1 0 10948 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_113
timestamp 1623621585
transform 1 0 11500 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1016_
timestamp 1623621585
transform 1 0 12972 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1108_
timestamp 1623621585
transform 1 0 12052 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_115
timestamp 1623621585
transform 1 0 11684 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_125
timestamp 1623621585
transform 1 0 12604 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_132
timestamp 1623621585
transform 1 0 13248 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_2  _1841_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 13984 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_56_149
timestamp 1623621585
transform 1 0 14812 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1623621585
transform 1 0 16836 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_161
timestamp 1623621585
transform 1 0 15916 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_169
timestamp 1623621585
transform 1 0 16652 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_172
timestamp 1623621585
transform 1 0 16928 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1107_
timestamp 1623621585
transform 1 0 18032 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1856_
timestamp 1623621585
transform 1 0 18768 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_56_188
timestamp 1623621585
transform 1 0 18400 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_199
timestamp 1623621585
transform 1 0 19412 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1860_
timestamp 1623621585
transform 1 0 20240 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1623621585
transform 1 0 22080 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_207
timestamp 1623621585
transform 1 0 20148 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_215
timestamp 1623621585
transform 1 0 20884 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_227
timestamp 1623621585
transform 1 0 21988 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2257_
timestamp 1623621585
transform 1 0 22540 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_56_229
timestamp 1623621585
transform 1 0 22172 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1865_
timestamp 1623621585
transform 1 0 25024 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1866_
timestamp 1623621585
transform 1 0 26036 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_56_252
timestamp 1623621585
transform 1 0 24288 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_267
timestamp 1623621585
transform 1 0 25668 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1885_
timestamp 1623621585
transform 1 0 27784 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1623621585
transform 1 0 27324 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_278
timestamp 1623621585
transform 1 0 26680 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_284
timestamp 1623621585
transform 1 0 27232 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_286
timestamp 1623621585
transform 1 0 27416 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_294
timestamp 1623621585
transform 1 0 28152 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1623621585
transform -1 0 28888 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_298
timestamp 1623621585
transform 1 0 28520 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1236_
timestamp 1623621585
transform 1 0 2116 0 1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1623621585
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output250
timestamp 1623621585
transform 1 0 1380 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_7
timestamp 1623621585
transform 1 0 1748 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1267_
timestamp 1623621585
transform 1 0 4968 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1623621585
transform 1 0 3772 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output312
timestamp 1623621585
transform 1 0 4232 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_25
timestamp 1623621585
transform 1 0 3404 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_30
timestamp 1623621585
transform 1 0 3864 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_38
timestamp 1623621585
transform 1 0 4600 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_45
timestamp 1623621585
transform 1 0 5244 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1712_
timestamp 1623621585
transform 1 0 5612 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_52
timestamp 1623621585
transform 1 0 5888 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_64
timestamp 1623621585
transform 1 0 6992 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1442_
timestamp 1623621585
transform 1 0 7820 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1623621585
transform 1 0 9016 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_72
timestamp 1623621585
transform 1 0 7728 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_82
timestamp 1623621585
transform 1 0 8648 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_87
timestamp 1623621585
transform 1 0 9108 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1039_
timestamp 1623621585
transform 1 0 9660 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_97
timestamp 1623621585
transform 1 0 10028 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_109
timestamp 1623621585
transform 1 0 11132 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1019_
timestamp 1623621585
transform 1 0 12696 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1823_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 13340 0 1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_57_121
timestamp 1623621585
transform 1 0 12236 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_125
timestamp 1623621585
transform 1 0 12604 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_129
timestamp 1623621585
transform 1 0 12972 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1058_
timestamp 1623621585
transform 1 0 14996 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1623621585
transform 1 0 14260 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_138
timestamp 1623621585
transform 1 0 13800 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_142
timestamp 1623621585
transform 1 0 14168 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_144
timestamp 1623621585
transform 1 0 14352 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_150
timestamp 1623621585
transform 1 0 14904 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_154
timestamp 1623621585
transform 1 0 15272 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1073_
timestamp 1623621585
transform 1 0 16008 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1078_
timestamp 1623621585
transform 1 0 16744 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_165
timestamp 1623621585
transform 1 0 16284 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_169
timestamp 1623621585
transform 1 0 16652 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_173
timestamp 1623621585
transform 1 0 17020 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1056_
timestamp 1623621585
transform 1 0 18124 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1858_
timestamp 1623621585
transform 1 0 19964 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1623621585
transform 1 0 19504 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_188
timestamp 1623621585
transform 1 0 18400 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_201
timestamp 1623621585
transform 1 0 19596 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1861_
timestamp 1623621585
transform 1 0 21436 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_57_209
timestamp 1623621585
transform 1 0 20332 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_228
timestamp 1623621585
transform 1 0 22080 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1863_
timestamp 1623621585
transform 1 0 23644 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_57_240
timestamp 1623621585
transform 1 0 23184 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_244
timestamp 1623621585
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _1868_
timestamp 1623621585
transform 1 0 25576 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1623621585
transform 1 0 24748 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_252
timestamp 1623621585
transform 1 0 24288 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_256
timestamp 1623621585
transform 1 0 24656 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_258
timestamp 1623621585
transform 1 0 24840 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_273
timestamp 1623621585
transform 1 0 26220 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1886_
timestamp 1623621585
transform 1 0 27048 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1887_
timestamp 1623621585
transform 1 0 27784 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_281
timestamp 1623621585
transform 1 0 26956 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_286
timestamp 1623621585
transform 1 0 27416 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_294
timestamp 1623621585
transform 1 0 28152 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1623621585
transform -1 0 28888 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_298
timestamp 1623621585
transform 1 0 28520 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1623621585
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output251
timestamp 1623621585
transform 1 0 1748 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output309
timestamp 1623621585
transform 1 0 2484 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_3
timestamp 1623621585
transform 1 0 1380 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_11
timestamp 1623621585
transform 1 0 2116 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_19
timestamp 1623621585
transform 1 0 2852 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1255_
timestamp 1623621585
transform 1 0 3680 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1264_
timestamp 1623621585
transform 1 0 5152 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output311
timestamp 1623621585
transform 1 0 4416 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1623621585
transform 1 0 3588 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_32
timestamp 1623621585
transform 1 0 4048 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_40
timestamp 1623621585
transform 1 0 4784 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2203_
timestamp 1623621585
transform 1 0 7360 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1623621585
transform 1 0 6348 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_47
timestamp 1623621585
transform 1 0 5428 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_55
timestamp 1623621585
transform 1 0 6164 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_58
timestamp 1623621585
transform 1 0 6440 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_66
timestamp 1623621585
transform 1 0 7176 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_84
timestamp 1623621585
transform 1 0 8832 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1041_
timestamp 1623621585
transform 1 0 10948 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1623621585
transform 1 0 11592 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_96
timestamp 1623621585
transform 1 0 9936 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_104
timestamp 1623621585
transform 1 0 10672 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_110
timestamp 1623621585
transform 1 0 11224 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1024_
timestamp 1623621585
transform 1 0 13248 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1032_
timestamp 1623621585
transform 1 0 12512 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_115
timestamp 1623621585
transform 1 0 11684 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_123
timestamp 1623621585
transform 1 0 12420 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_128
timestamp 1623621585
transform 1 0 12880 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1623621585
transform 1 0 13616 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1096_
timestamp 1623621585
transform 1 0 13984 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1876_
timestamp 1623621585
transform 1 0 14628 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_143
timestamp 1623621585
transform 1 0 14260 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_153
timestamp 1623621585
transform 1 0 15180 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1080_
timestamp 1623621585
transform 1 0 17572 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _1090_
timestamp 1623621585
transform 1 0 15916 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1623621585
transform 1 0 16836 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_167
timestamp 1623621585
transform 1 0 16468 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_172
timestamp 1623621585
transform 1 0 16928 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_178
timestamp 1623621585
transform 1 0 17480 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _1075_
timestamp 1623621585
transform 1 0 18768 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_185
timestamp 1623621585
transform 1 0 18124 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_191
timestamp 1623621585
transform 1 0 18676 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_198
timestamp 1623621585
transform 1 0 19320 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3b_1  _1071_
timestamp 1623621585
transform 1 0 20792 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1623621585
transform 1 0 22080 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_210
timestamp 1623621585
transform 1 0 20424 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_220
timestamp 1623621585
transform 1 0 21344 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_229
timestamp 1623621585
transform 1 0 22172 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_241
timestamp 1623621585
transform 1 0 23276 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1623621585
transform 1 0 25944 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1623621585
transform 1 0 25300 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1623621585
transform 1 0 24656 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_253
timestamp 1623621585
transform 1 0 24380 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_259
timestamp 1623621585
transform 1 0 24932 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_266
timestamp 1623621585
transform 1 0 25576 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_273
timestamp 1623621585
transform 1 0 26220 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1888_
timestamp 1623621585
transform 1 0 26588 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1889_
timestamp 1623621585
transform 1 0 27784 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1623621585
transform 1 0 27324 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_281
timestamp 1623621585
transform 1 0 26956 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_286
timestamp 1623621585
transform 1 0 27416 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_294
timestamp 1623621585
transform 1 0 28152 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1623621585
transform -1 0 28888 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_298
timestamp 1623621585
transform 1 0 28520 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_8
timestamp 1623621585
transform 1 0 1840 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_3
timestamp 1623621585
transform 1 0 1380 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1623621585
transform 1 0 1380 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_3
timestamp 1623621585
transform 1 0 1564 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output253
timestamp 1623621585
transform 1 0 1472 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output252
timestamp 1623621585
transform 1 0 1748 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1623621585
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1623621585
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_11
timestamp 1623621585
transform 1 0 2116 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output310
timestamp 1623621585
transform 1 0 2484 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1268_
timestamp 1623621585
transform 1 0 2208 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_18
timestamp 1623621585
transform 1 0 2760 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_19
timestamp 1623621585
transform 1 0 2852 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1269_
timestamp 1623621585
transform 1 0 3128 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1215_
timestamp 1623621585
transform 1 0 4232 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1265_
timestamp 1623621585
transform 1 0 4968 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2234_
timestamp 1623621585
transform 1 0 4416 0 -1 35360
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1623621585
transform 1 0 3772 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_27
timestamp 1623621585
transform 1 0 3588 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_30
timestamp 1623621585
transform 1 0 3864 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_38
timestamp 1623621585
transform 1 0 4600 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_28
timestamp 1623621585
transform 1 0 3680 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2292_
timestamp 1623621585
transform 1 0 5888 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1623621585
transform 1 0 6348 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_46
timestamp 1623621585
transform 1 0 5336 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_53
timestamp 1623621585
transform 1 0 5980 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_58
timestamp 1623621585
transform 1 0 6440 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _2294_
timestamp 1623621585
transform 1 0 9476 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1623621585
transform 1 0 9016 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_wb_clk_i
timestamp 1623621585
transform 1 0 7728 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_71
timestamp 1623621585
transform 1 0 7636 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_83
timestamp 1623621585
transform 1 0 8740 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_87
timestamp 1623621585
transform 1 0 9108 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_70
timestamp 1623621585
transform 1 0 7544 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_75
timestamp 1623621585
transform 1 0 8004 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_87
timestamp 1623621585
transform 1 0 9108 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1037_
timestamp 1623621585
transform 1 0 9752 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1042_
timestamp 1623621585
transform 1 0 10396 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1623621585
transform 1 0 11592 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_110
timestamp 1623621585
transform 1 0 11224 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_114
timestamp 1623621585
transform 1 0 11592 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_93
timestamp 1623621585
transform 1 0 9660 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_97
timestamp 1623621585
transform 1 0 10028 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_109
timestamp 1623621585
transform 1 0 11132 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_113
timestamp 1623621585
transform 1 0 11500 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_121
timestamp 1623621585
transform 1 0 12236 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_115
timestamp 1623621585
transform 1 0 11684 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_121
timestamp 1623621585
transform 1 0 12236 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1105_
timestamp 1623621585
transform 1 0 11684 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _1099_
timestamp 1623621585
transform 1 0 12328 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_128
timestamp 1623621585
transform 1 0 12880 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_129
timestamp 1623621585
transform 1 0 12972 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_135
timestamp 1623621585
transform 1 0 13524 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_136
timestamp 1623621585
transform 1 0 13616 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1034_
timestamp 1623621585
transform 1 0 13248 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1020_
timestamp 1623621585
transform 1 0 13248 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_143
timestamp 1623621585
transform 1 0 14260 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_142
timestamp 1623621585
transform 1 0 14168 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1623621585
transform 1 0 14260 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1026_
timestamp 1623621585
transform 1 0 14536 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_157
timestamp 1623621585
transform 1 0 15548 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_149
timestamp 1623621585
transform 1 0 14812 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_156
timestamp 1623621585
transform 1 0 15456 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1093_
timestamp 1623621585
transform 1 0 15732 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1092_
timestamp 1623621585
transform 1 0 15180 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_144
timestamp 1623621585
transform 1 0 14352 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_164
timestamp 1623621585
transform 1 0 16192 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_165
timestamp 1623621585
transform 1 0 16284 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1022_
timestamp 1623621585
transform 1 0 15916 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_172
timestamp 1623621585
transform 1 0 16928 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_170
timestamp 1623621585
transform 1 0 16744 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_177
timestamp 1623621585
transform 1 0 17388 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1623621585
transform 1 0 16836 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _1083_
timestamp 1623621585
transform 1 0 16836 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1087_
timestamp 1623621585
transform 1 0 17664 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1086_
timestamp 1623621585
transform 1 0 17756 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_192
timestamp 1623621585
transform 1 0 18768 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_188
timestamp 1623621585
transform 1 0 18400 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1055_
timestamp 1623621585
transform 1 0 18860 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_197
timestamp 1623621585
transform 1 0 19228 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_201
timestamp 1623621585
transform 1 0 19596 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_199
timestamp 1623621585
transform 1 0 19412 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1623621585
transform 1 0 19504 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1076_
timestamp 1623621585
transform 1 0 19596 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_187
timestamp 1623621585
transform 1 0 18308 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2287_
timestamp 1623621585
transform 1 0 19964 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__o211a_1  _1072_
timestamp 1623621585
transform 1 0 20884 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1623621585
transform 1 0 22080 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_221
timestamp 1623621585
transform 1 0 21436 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_60_209
timestamp 1623621585
transform 1 0 20332 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_223
timestamp 1623621585
transform 1 0 21620 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_227
timestamp 1623621585
transform 1 0 21988 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_237
timestamp 1623621585
transform 1 0 22908 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_229
timestamp 1623621585
transform 1 0 22172 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_237
timestamp 1623621585
transform 1 0 22908 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_229
timestamp 1623621585
transform 1 0 22172 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__nand3b_1  _1067_
timestamp 1623621585
transform 1 0 22356 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_244
timestamp 1623621585
transform 1 0 23552 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_241
timestamp 1623621585
transform 1 0 23276 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _1064_
timestamp 1623621585
transform 1 0 23368 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _1061_
timestamp 1623621585
transform 1 0 23000 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_248
timestamp 1623621585
transform 1 0 23920 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1065_
timestamp 1623621585
transform 1 0 23920 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2290_
timestamp 1623621585
transform 1 0 25024 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1623621585
transform 1 0 24748 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1623621585
transform 1 0 25852 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1623621585
transform 1 0 25208 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_256
timestamp 1623621585
transform 1 0 24656 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_258
timestamp 1623621585
transform 1 0 24840 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_265
timestamp 1623621585
transform 1 0 25484 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_272
timestamp 1623621585
transform 1 0 26128 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_256
timestamp 1623621585
transform 1 0 24656 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_276
timestamp 1623621585
transform 1 0 26496 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_279
timestamp 1623621585
transform 1 0 26772 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1623621585
transform 1 0 26496 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_290
timestamp 1623621585
transform 1 0 27784 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_286
timestamp 1623621585
transform 1 0 27416 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_284
timestamp 1623621585
transform 1 0 27232 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_287
timestamp 1623621585
transform 1 0 27508 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1623621585
transform 1 0 27324 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1892_
timestamp 1623621585
transform 1 0 27876 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1891_
timestamp 1623621585
transform 1 0 27876 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1890_
timestamp 1623621585
transform 1 0 27140 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_295
timestamp 1623621585
transform 1 0 28244 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_295
timestamp 1623621585
transform 1 0 28244 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1623621585
transform -1 0 28888 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1623621585
transform -1 0 28888 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _1237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1564 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1270_
timestamp 1623621585
transform 1 0 2852 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1623621585
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1623621585
transform 1 0 1380 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_12
timestamp 1623621585
transform 1 0 2208 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_18
timestamp 1623621585
transform 1 0 2760 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1258_
timestamp 1623621585
transform 1 0 4232 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1623621585
transform 1 0 3772 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_25
timestamp 1623621585
transform 1 0 3404 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_30
timestamp 1623621585
transform 1 0 3864 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_38
timestamp 1623621585
transform 1 0 4600 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2b_1  _1218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 6992 0 1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_61_50
timestamp 1623621585
transform 1 0 5704 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_62
timestamp 1623621585
transform 1 0 6808 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2295_
timestamp 1623621585
transform 1 0 9476 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1623621585
transform 1 0 9016 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1623621585
transform 1 0 7452 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_81
timestamp 1623621585
transform 1 0 8556 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_85
timestamp 1623621585
transform 1 0 8924 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_87
timestamp 1623621585
transform 1 0 9108 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1101_
timestamp 1623621585
transform 1 0 11592 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_110
timestamp 1623621585
transform 1 0 11224 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1097_
timestamp 1623621585
transform 1 0 13156 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_120
timestamp 1623621585
transform 1 0 12144 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_128
timestamp 1623621585
transform 1 0 12880 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_61_137
timestamp 1623621585
transform 1 0 13708 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1623621585
transform 1 0 14720 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1623621585
transform 1 0 14260 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_144
timestamp 1623621585
transform 1 0 14352 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_151
timestamp 1623621585
transform 1 0 14996 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_159
timestamp 1623621585
transform 1 0 15732 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1043_
timestamp 1623621585
transform 1 0 15824 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1069_
timestamp 1623621585
transform 1 0 16652 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1623621585
transform 1 0 16192 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_168
timestamp 1623621585
transform 1 0 16560 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_173
timestamp 1623621585
transform 1 0 17020 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__o211a_1  _1081_
timestamp 1623621585
transform 1 0 18216 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1623621585
transform 1 0 19504 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_185
timestamp 1623621585
transform 1 0 18124 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_194
timestamp 1623621585
transform 1 0 18952 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_201
timestamp 1623621585
transform 1 0 19596 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2288_
timestamp 1623621585
transform 1 0 21160 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_61_213
timestamp 1623621585
transform 1 0 20700 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_217
timestamp 1623621585
transform 1 0 21068 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1062_
timestamp 1623621585
transform 1 0 23644 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_wb_clk_i
timestamp 1623621585
transform 1 0 23000 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_234
timestamp 1623621585
transform 1 0 22632 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_241
timestamp 1623621585
transform 1 0 23276 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2291_
timestamp 1623621585
transform 1 0 25208 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1623621585
transform 1 0 24748 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_253
timestamp 1623621585
transform 1 0 24380 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_258
timestamp 1623621585
transform 1 0 24840 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1893_
timestamp 1623621585
transform 1 0 27876 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1894_
timestamp 1623621585
transform 1 0 27140 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_278
timestamp 1623621585
transform 1 0 26680 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_282
timestamp 1623621585
transform 1 0 27048 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_287
timestamp 1623621585
transform 1 0 27508 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_295
timestamp 1623621585
transform 1 0 28244 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1623621585
transform -1 0 28888 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1239_
timestamp 1623621585
transform 1 0 2944 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1249_
timestamp 1623621585
transform 1 0 1380 0 -1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1623621585
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_16
timestamp 1623621585
transform 1 0 2576 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1257_
timestamp 1623621585
transform 1 0 3772 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1259_
timestamp 1623621585
transform 1 0 4692 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_23
timestamp 1623621585
transform 1 0 3220 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_32
timestamp 1623621585
transform 1 0 4048 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_38
timestamp 1623621585
transform 1 0 4600 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_42
timestamp 1623621585
transform 1 0 4968 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1706_
timestamp 1623621585
transform 1 0 5428 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2237_
timestamp 1623621585
transform 1 0 6900 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1623621585
transform 1 0 6348 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_46
timestamp 1623621585
transform 1 0 5336 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_50
timestamp 1623621585
transform 1 0 5704 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_56
timestamp 1623621585
transform 1 0 6256 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_58
timestamp 1623621585
transform 1 0 6440 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_62
timestamp 1623621585
transform 1 0 6808 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1992_
timestamp 1623621585
transform 1 0 8740 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_62_79
timestamp 1623621585
transform 1 0 8372 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1038_
timestamp 1623621585
transform 1 0 10488 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1623621585
transform 1 0 11592 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_92
timestamp 1623621585
transform 1 0 9568 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_100
timestamp 1623621585
transform 1 0 10304 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_110
timestamp 1623621585
transform 1 0 11224 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_wb_clk_i
timestamp 1623621585
transform 1 0 12052 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_115
timestamp 1623621585
transform 1 0 11684 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_122
timestamp 1623621585
transform 1 0 12328 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_134
timestamp 1623621585
transform 1 0 13432 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1029_
timestamp 1623621585
transform 1 0 13892 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1877_
timestamp 1623621585
transform 1 0 15180 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_138
timestamp 1623621585
transform 1 0 13800 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_142
timestamp 1623621585
transform 1 0 14168 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_150
timestamp 1623621585
transform 1 0 14904 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1084_
timestamp 1623621585
transform 1 0 17388 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1623621585
transform 1 0 16836 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_161
timestamp 1623621585
transform 1 0 15916 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_169
timestamp 1623621585
transform 1 0 16652 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_172
timestamp 1623621585
transform 1 0 16928 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_176
timestamp 1623621585
transform 1 0 17296 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2286_
timestamp 1623621585
transform 1 0 18676 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_62_185
timestamp 1623621585
transform 1 0 18124 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1623621585
transform 1 0 22080 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_207
timestamp 1623621585
transform 1 0 20148 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_219
timestamp 1623621585
transform 1 0 21252 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_227
timestamp 1623621585
transform 1 0 21988 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1068_
timestamp 1623621585
transform 1 0 22724 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_62_229
timestamp 1623621585
transform 1 0 22172 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_243
timestamp 1623621585
transform 1 0 23460 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1623621585
transform 1 0 26036 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1623621585
transform 1 0 25392 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_255
timestamp 1623621585
transform 1 0 24564 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_263
timestamp 1623621585
transform 1 0 25300 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_267
timestamp 1623621585
transform 1 0 25668 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_274
timestamp 1623621585
transform 1 0 26312 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1895_
timestamp 1623621585
transform 1 0 27876 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1623621585
transform 1 0 27324 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1623621585
transform 1 0 26680 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_281
timestamp 1623621585
transform 1 0 26956 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_286
timestamp 1623621585
transform 1 0 27416 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_290
timestamp 1623621585
transform 1 0 27784 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_295
timestamp 1623621585
transform 1 0 28244 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1623621585
transform -1 0 28888 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1623621585
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output254
timestamp 1623621585
transform 1 0 1748 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output256
timestamp 1623621585
transform 1 0 2484 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1623621585
transform 1 0 1380 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_11
timestamp 1623621585
transform 1 0 2116 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_19
timestamp 1623621585
transform 1 0 2852 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__nor2b_1  _1217_
timestamp 1623621585
transform 1 0 4968 0 1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1262_
timestamp 1623621585
transform 1 0 4232 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1623621585
transform 1 0 3772 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_27
timestamp 1623621585
transform 1 0 3588 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_30
timestamp 1623621585
transform 1 0 3864 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_37
timestamp 1623621585
transform 1 0 4508 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_41
timestamp 1623621585
transform 1 0 4876 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2238_
timestamp 1623621585
transform 1 0 5796 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_63_47
timestamp 1623621585
transform 1 0 5428 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_67
timestamp 1623621585
transform 1 0 7268 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1623621585
transform 1 0 9016 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_wb_clk_i
timestamp 1623621585
transform 1 0 9476 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_79
timestamp 1623621585
transform 1 0 8372 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_85
timestamp 1623621585
transform 1 0 8924 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_87
timestamp 1623621585
transform 1 0 9108 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_94
timestamp 1623621585
transform 1 0 9752 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_106
timestamp 1623621585
transform 1 0 10856 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_114
timestamp 1623621585
transform 1 0 11592 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1095_
timestamp 1623621585
transform 1 0 13524 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1109_
timestamp 1623621585
transform 1 0 11684 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1623621585
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1023_
timestamp 1623621585
transform 1 0 14904 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2299_
timestamp 1623621585
transform 1 0 15640 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1623621585
transform 1 0 14260 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_139
timestamp 1623621585
transform 1 0 13892 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_144
timestamp 1623621585
transform 1 0 14352 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_154
timestamp 1623621585
transform 1 0 15272 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1077_
timestamp 1623621585
transform 1 0 17756 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_177
timestamp 1623621585
transform 1 0 17388 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1623621585
transform 1 0 19504 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_wb_clk_i
timestamp 1623621585
transform 1 0 18492 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_185
timestamp 1623621585
transform 1 0 18124 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_192
timestamp 1623621585
transform 1 0 18768 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_201
timestamp 1623621585
transform 1 0 19596 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1565_
timestamp 1623621585
transform 1 0 21436 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_wb_clk_i
timestamp 1623621585
transform 1 0 20516 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_209
timestamp 1623621585
transform 1 0 20332 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_214
timestamp 1623621585
transform 1 0 20792 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_220
timestamp 1623621585
transform 1 0 21344 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_224
timestamp 1623621585
transform 1 0 21712 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_236
timestamp 1623621585
transform 1 0 22816 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_248
timestamp 1623621585
transform 1 0 23920 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1875_
timestamp 1623621585
transform 1 0 25852 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1623621585
transform 1 0 24748 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1623621585
transform 1 0 25208 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_256
timestamp 1623621585
transform 1 0 24656 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_258
timestamp 1623621585
transform 1 0 24840 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_265
timestamp 1623621585
transform 1 0 25484 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_272
timestamp 1623621585
transform 1 0 26128 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1896_
timestamp 1623621585
transform 1 0 27876 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1623621585
transform 1 0 27232 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1623621585
transform 1 0 26588 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_276
timestamp 1623621585
transform 1 0 26496 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_280
timestamp 1623621585
transform 1 0 26864 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_287
timestamp 1623621585
transform 1 0 27508 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_295
timestamp 1623621585
transform 1 0 28244 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1623621585
transform -1 0 28888 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1623621585
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output255
timestamp 1623621585
transform 1 0 1748 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output258
timestamp 1623621585
transform 1 0 2484 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1623621585
transform 1 0 1380 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_11
timestamp 1623621585
transform 1 0 2116 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_19
timestamp 1623621585
transform 1 0 2852 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1256_
timestamp 1623621585
transform 1 0 4600 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1260_
timestamp 1623621585
transform 1 0 5244 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1263_
timestamp 1623621585
transform 1 0 3312 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_64_23
timestamp 1623621585
transform 1 0 3220 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_31
timestamp 1623621585
transform 1 0 3956 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_37
timestamp 1623621585
transform 1 0 4508 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_41
timestamp 1623621585
transform 1 0 4876 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1623621585
transform 1 0 6348 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_48
timestamp 1623621585
transform 1 0 5520 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_56
timestamp 1623621585
transform 1 0 6256 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_58
timestamp 1623621585
transform 1 0 6440 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _1993_
timestamp 1623621585
transform 1 0 8648 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_64_70
timestamp 1623621585
transform 1 0 7544 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_91
timestamp 1623621585
transform 1 0 9476 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1807_
timestamp 1623621585
transform 1 0 9844 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1623621585
transform 1 0 11592 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_98
timestamp 1623621585
transform 1 0 10120 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_110
timestamp 1623621585
transform 1 0 11224 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1098_
timestamp 1623621585
transform 1 0 13156 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1106_
timestamp 1623621585
transform 1 0 12052 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_115
timestamp 1623621585
transform 1 0 11684 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_127
timestamp 1623621585
transform 1 0 12788 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1059_
timestamp 1623621585
transform 1 0 15640 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1840_
timestamp 1623621585
transform 1 0 14352 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_64_139
timestamp 1623621585
transform 1 0 13892 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_143
timestamp 1623621585
transform 1 0 14260 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_151
timestamp 1623621585
transform 1 0 14996 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_157
timestamp 1623621585
transform 1 0 15548 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1623621585
transform 1 0 16836 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_162
timestamp 1623621585
transform 1 0 16008 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_170
timestamp 1623621585
transform 1 0 16744 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_172
timestamp 1623621585
transform 1 0 16928 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1947_
timestamp 1623621585
transform 1 0 19964 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2284_
timestamp 1623621585
transform 1 0 18032 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_64_200
timestamp 1623621585
transform 1 0 19504 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_204
timestamp 1623621585
transform 1 0 19872 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1207_
timestamp 1623621585
transform 1 0 21160 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1623621585
transform 1 0 22080 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_214
timestamp 1623621585
transform 1 0 20792 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_222
timestamp 1623621585
transform 1 0 21528 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2289_
timestamp 1623621585
transform 1 0 22816 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_64_229
timestamp 1623621585
transform 1 0 22172 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_235
timestamp 1623621585
transform 1 0 22724 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__nor2b_1  _1206_
timestamp 1623621585
transform 1 0 24656 0 -1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _1943_
timestamp 1623621585
transform 1 0 25484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_252
timestamp 1623621585
transform 1 0 24288 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_261
timestamp 1623621585
transform 1 0 25116 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1897_
timestamp 1623621585
transform 1 0 27876 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1623621585
transform 1 0 27324 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_277
timestamp 1623621585
transform 1 0 26588 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_286
timestamp 1623621585
transform 1 0 27416 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_290
timestamp 1623621585
transform 1 0 27784 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_295
timestamp 1623621585
transform 1 0 28244 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1623621585
transform -1 0 28888 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1251_
timestamp 1623621585
transform 1 0 2208 0 1 37536
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1623621585
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output257
timestamp 1623621585
transform 1 0 1472 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_3
timestamp 1623621585
transform 1 0 1380 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_8
timestamp 1623621585
transform 1 0 1840 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1240_
timestamp 1623621585
transform 1 0 4232 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _2235_
timestamp 1623621585
transform 1 0 5060 0 1 37536
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1623621585
transform 1 0 3772 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_25
timestamp 1623621585
transform 1 0 3404 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_30
timestamp 1623621585
transform 1 0 3864 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_37
timestamp 1623621585
transform 1 0 4508 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_60
timestamp 1623621585
transform 1 0 6624 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1623621585
transform 1 0 9016 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_72
timestamp 1623621585
transform 1 0 7728 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_84
timestamp 1623621585
transform 1 0 8832 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_87
timestamp 1623621585
transform 1 0 9108 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2277_
timestamp 1623621585
transform 1 0 10120 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_65_95
timestamp 1623621585
transform 1 0 9844 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_114
timestamp 1623621585
transform 1 0 11592 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2278_
timestamp 1623621585
transform 1 0 11960 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_65_134
timestamp 1623621585
transform 1 0 13432 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1824_
timestamp 1623621585
transform 1 0 14720 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1848_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 15456 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1623621585
transform 1 0 14260 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_142
timestamp 1623621585
transform 1 0 14168 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_144
timestamp 1623621585
transform 1 0 14352 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_152
timestamp 1623621585
transform 1 0 15088 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1088_
timestamp 1623621585
transform 1 0 16560 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_164
timestamp 1623621585
transform 1 0 16192 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_172
timestamp 1623621585
transform 1 0 16928 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1623621585
transform 1 0 19504 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_184
timestamp 1623621585
transform 1 0 18032 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_196
timestamp 1623621585
transform 1 0 19136 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_201
timestamp 1623621585
transform 1 0 19596 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_205
timestamp 1623621585
transform 1 0 19964 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1874_
timestamp 1623621585
transform 1 0 20056 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2242_
timestamp 1623621585
transform 1 0 20792 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_65_209
timestamp 1623621585
transform 1 0 20332 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_213
timestamp 1623621585
transform 1 0 20700 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _1945_
timestamp 1623621585
transform 1 0 22724 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_230
timestamp 1623621585
transform 1 0 22264 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_234
timestamp 1623621585
transform 1 0 22632 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_247
timestamp 1623621585
transform 1 0 23828 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1942_
timestamp 1623621585
transform 1 0 25392 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1623621585
transform 1 0 24748 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_255
timestamp 1623621585
transform 1 0 24564 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_258
timestamp 1623621585
transform 1 0 24840 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_65_273
timestamp 1623621585
transform 1 0 26220 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1898_
timestamp 1623621585
transform 1 0 27048 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1899_
timestamp 1623621585
transform 1 0 27784 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_281
timestamp 1623621585
transform 1 0 26956 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_286
timestamp 1623621585
transform 1 0 27416 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_294
timestamp 1623621585
transform 1 0 28152 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1623621585
transform -1 0 28888 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_65_298
timestamp 1623621585
transform 1 0 28520 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_3
timestamp 1623621585
transform 1 0 1380 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_3
timestamp 1623621585
transform 1 0 1380 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1623621585
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1623621585
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1243_
timestamp 1623621585
transform 1 0 1472 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1238_
timestamp 1623621585
transform 1 0 1656 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_10
timestamp 1623621585
transform 1 0 2024 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_12
timestamp 1623621585
transform 1 0 2208 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output261
timestamp 1623621585
transform 1 0 2576 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_18
timestamp 1623621585
transform 1 0 2760 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_20
timestamp 1623621585
transform 1 0 2944 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1245_
timestamp 1623621585
transform 1 0 2944 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_30
timestamp 1623621585
transform 1 0 3864 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_28
timestamp 1623621585
transform 1 0 3680 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_24
timestamp 1623621585
transform 1 0 3312 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1623621585
transform 1 0 3772 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _1253_
timestamp 1623621585
transform 1 0 4232 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_40
timestamp 1623621585
transform 1 0 4784 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_45
timestamp 1623621585
transform 1 0 5244 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_38
timestamp 1623621585
transform 1 0 4600 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1254_
timestamp 1623621585
transform 1 0 5152 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1244_
timestamp 1623621585
transform 1 0 4968 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _1252_
timestamp 1623621585
transform 1 0 3312 0 -1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_67_54
timestamp 1623621585
transform 1 0 6072 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_47
timestamp 1623621585
transform 1 0 5428 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_56
timestamp 1623621585
transform 1 0 6256 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_52
timestamp 1623621585
transform 1 0 5888 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1623621585
transform 1 0 6348 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1792_
timestamp 1623621585
transform 1 0 5612 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1367_
timestamp 1623621585
transform 1 0 5796 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_68
timestamp 1623621585
transform 1 0 7360 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_58
timestamp 1623621585
transform 1 0 6440 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1403_
timestamp 1623621585
transform 1 0 6532 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_58
timestamp 1623621585
transform 1 0 6440 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_75
timestamp 1623621585
transform 1 0 8004 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_78
timestamp 1623621585
transform 1 0 8280 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_70
timestamp 1623621585
transform 1 0 7544 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1799_
timestamp 1623621585
transform 1 0 8372 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1405_
timestamp 1623621585
transform 1 0 7728 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_87
timestamp 1623621585
transform 1 0 9108 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_82
timestamp 1623621585
transform 1 0 8648 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_90
timestamp 1623621585
transform 1 0 9384 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1623621585
transform 1 0 9016 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1986_
timestamp 1623621585
transform 1 0 8556 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1987_
timestamp 1623621585
transform 1 0 9476 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _1828_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 10396 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _1832_
timestamp 1623621585
transform 1 0 10948 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1623621585
transform 1 0 11592 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_98
timestamp 1623621585
transform 1 0 10120 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_110
timestamp 1623621585
transform 1 0 11224 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_103
timestamp 1623621585
transform 1 0 10580 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2281_
timestamp 1623621585
transform 1 0 13156 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_115
timestamp 1623621585
transform 1 0 11684 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_127
timestamp 1623621585
transform 1 0 12788 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_116
timestamp 1623621585
transform 1 0 11776 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_128
timestamp 1623621585
transform 1 0 12880 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1825_
timestamp 1623621585
transform 1 0 14996 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1623621585
transform 1 0 14260 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_wb_clk_i
timestamp 1623621585
transform 1 0 14720 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_147
timestamp 1623621585
transform 1 0 14628 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_155
timestamp 1623621585
transform 1 0 15364 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_140
timestamp 1623621585
transform 1 0 13984 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_144
timestamp 1623621585
transform 1 0 14352 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_151
timestamp 1623621585
transform 1 0 14996 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__o211a_1  _1091_
timestamp 1623621585
transform 1 0 16376 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2283_
timestamp 1623621585
transform 1 0 17296 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2285_
timestamp 1623621585
transform 1 0 17572 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1623621585
transform 1 0 16836 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_167
timestamp 1623621585
transform 1 0 16468 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_172
timestamp 1623621585
transform 1 0 16928 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_163
timestamp 1623621585
transform 1 0 16100 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_174
timestamp 1623621585
transform 1 0 17112 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_178
timestamp 1623621585
transform 1 0 17480 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1946_
timestamp 1623621585
transform 1 0 19596 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1623621585
transform 1 0 19504 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_192
timestamp 1623621585
transform 1 0 18768 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_200
timestamp 1623621585
transform 1 0 19504 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_195
timestamp 1623621585
transform 1 0 19044 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_199
timestamp 1623621585
transform 1 0 19412 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_201
timestamp 1623621585
transform 1 0 19596 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2b_1  _1208_
timestamp 1623621585
transform 1 0 20792 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1623621585
transform 1 0 22080 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_210
timestamp 1623621585
transform 1 0 20424 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_219
timestamp 1623621585
transform 1 0 21252 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_227
timestamp 1623621585
transform 1 0 21988 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_213
timestamp 1623621585
transform 1 0 20700 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_225
timestamp 1623621585
transform 1 0 21804 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1873_
timestamp 1623621585
transform 1 0 22540 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1944_
timestamp 1623621585
transform 1 0 22540 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2243_
timestamp 1623621585
transform 1 0 24196 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_66_229
timestamp 1623621585
transform 1 0 22172 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_242
timestamp 1623621585
transform 1 0 23368 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_250
timestamp 1623621585
transform 1 0 24104 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_236
timestamp 1623621585
transform 1 0 22816 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_248
timestamp 1623621585
transform 1 0 23920 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1623621585
transform 1 0 24748 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1623621585
transform 1 0 26036 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1623621585
transform 1 0 25852 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_267
timestamp 1623621585
transform 1 0 25668 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_274
timestamp 1623621585
transform 1 0 26312 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_256
timestamp 1623621585
transform 1 0 24656 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_258
timestamp 1623621585
transform 1 0 24840 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_266
timestamp 1623621585
transform 1 0 25576 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_272
timestamp 1623621585
transform 1 0 26128 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1623621585
transform 1 0 26496 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1623621585
transform 1 0 26680 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_279
timestamp 1623621585
transform 1 0 26772 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_281
timestamp 1623621585
transform 1 0 26956 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1902_
timestamp 1623621585
transform 1 0 27140 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_287
timestamp 1623621585
transform 1 0 27508 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_286
timestamp 1623621585
transform 1 0 27416 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1623621585
transform 1 0 27324 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1901_
timestamp 1623621585
transform 1 0 27876 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1900_
timestamp 1623621585
transform 1 0 27784 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_295
timestamp 1623621585
transform 1 0 28244 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_294
timestamp 1623621585
transform 1 0 28152 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1623621585
transform -1 0 28888 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1623621585
transform -1 0 28888 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_298
timestamp 1623621585
transform 1 0 28520 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1623621585
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output259
timestamp 1623621585
transform 1 0 1748 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output263
timestamp 1623621585
transform 1 0 2484 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_3
timestamp 1623621585
transform 1 0 1380 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_11
timestamp 1623621585
transform 1 0 2116 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_19
timestamp 1623621585
transform 1 0 2852 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _1248_
timestamp 1623621585
transform 1 0 3680 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output266
timestamp 1623621585
transform 1 0 4416 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output267
timestamp 1623621585
transform 1 0 5152 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1623621585
transform 1 0 3588 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_32
timestamp 1623621585
transform 1 0 4048 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_40
timestamp 1623621585
transform 1 0 4784 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1404_
timestamp 1623621585
transform 1 0 6808 0 -1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1623621585
transform 1 0 6348 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_48
timestamp 1623621585
transform 1 0 5520 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_56
timestamp 1623621585
transform 1 0 6256 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_58
timestamp 1623621585
transform 1 0 6440 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_67
timestamp 1623621585
transform 1 0 7268 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_4  _1800_
timestamp 1623621585
transform 1 0 7728 0 -1 39712
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_68_71
timestamp 1623621585
transform 1 0 7636 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_89
timestamp 1623621585
transform 1 0 9292 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1810_
timestamp 1623621585
transform 1 0 9660 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1835_
timestamp 1623621585
transform 1 0 10304 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1623621585
transform 1 0 11592 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_96
timestamp 1623621585
transform 1 0 9936 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_108
timestamp 1623621585
transform 1 0 11040 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1102_
timestamp 1623621585
transform 1 0 12052 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_115
timestamp 1623621585
transform 1 0 11684 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_127
timestamp 1623621585
transform 1 0 12788 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__o211a_1  _1030_
timestamp 1623621585
transform 1 0 13892 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1844_
timestamp 1623621585
transform 1 0 14996 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_147
timestamp 1623621585
transform 1 0 14628 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_159
timestamp 1623621585
transform 1 0 15732 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1623621585
transform 1 0 16836 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_172
timestamp 1623621585
transform 1 0 16928 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2236_
timestamp 1623621585
transform 1 0 18676 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_wb_clk_i
timestamp 1623621585
transform 1 0 18032 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_187
timestamp 1623621585
transform 1 0 18308 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1623621585
transform 1 0 22080 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_207
timestamp 1623621585
transform 1 0 20148 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_219
timestamp 1623621585
transform 1 0 21252 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_227
timestamp 1623621585
transform 1 0 21988 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1680_
timestamp 1623621585
transform 1 0 22540 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_229
timestamp 1623621585
transform 1 0 22172 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_236
timestamp 1623621585
transform 1 0 22816 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1623621585
transform 1 0 23920 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1499_
timestamp 1623621585
transform 1 0 24288 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_68_259
timestamp 1623621585
transform 1 0 24932 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_271
timestamp 1623621585
transform 1 0 26036 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1903_
timestamp 1623621585
transform 1 0 27876 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1623621585
transform 1 0 27324 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1623621585
transform 1 0 26680 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_68_277
timestamp 1623621585
transform 1 0 26588 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_281
timestamp 1623621585
transform 1 0 26956 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_286
timestamp 1623621585
transform 1 0 27416 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_290
timestamp 1623621585
transform 1 0 27784 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_295
timestamp 1623621585
transform 1 0 28244 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1623621585
transform -1 0 28888 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1623621585
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output262
timestamp 1623621585
transform 1 0 1748 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output265
timestamp 1623621585
transform 1 0 2484 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_3
timestamp 1623621585
transform 1 0 1380 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_11
timestamp 1623621585
transform 1 0 2116 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_19
timestamp 1623621585
transform 1 0 2852 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_4  _1794_
timestamp 1623621585
transform 1 0 4416 0 1 39712
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1623621585
transform 1 0 3772 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_27
timestamp 1623621585
transform 1 0 3588 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_30
timestamp 1623621585
transform 1 0 3864 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1708_
timestamp 1623621585
transform 1 0 6348 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_53
timestamp 1623621585
transform 1 0 5980 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_60
timestamp 1623621585
transform 1 0 6624 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__o211a_1  _1407_
timestamp 1623621585
transform 1 0 7912 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1623621585
transform 1 0 9016 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_72
timestamp 1623621585
transform 1 0 7728 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_82
timestamp 1623621585
transform 1 0 8648 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_87
timestamp 1623621585
transform 1 0 9108 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2279_
timestamp 1623621585
transform 1 0 10672 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_99
timestamp 1623621585
transform 1 0 10212 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_103
timestamp 1623621585
transform 1 0 10580 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1035_
timestamp 1623621585
transform 1 0 13156 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_69_120
timestamp 1623621585
transform 1 0 12144 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_128
timestamp 1623621585
transform 1 0 12880 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1027_
timestamp 1623621585
transform 1 0 14904 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1623621585
transform 1 0 14260 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_139
timestamp 1623621585
transform 1 0 13892 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_144
timestamp 1623621585
transform 1 0 14352 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_158
timestamp 1623621585
transform 1 0 15640 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1094_
timestamp 1623621585
transform 1 0 16192 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_172
timestamp 1623621585
transform 1 0 16928 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2b_1  _1219_
timestamp 1623621585
transform 1 0 18216 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1806_
timestamp 1623621585
transform 1 0 19964 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1623621585
transform 1 0 19504 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_184
timestamp 1623621585
transform 1 0 18032 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_191
timestamp 1623621585
transform 1 0 18676 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_199
timestamp 1623621585
transform 1 0 19412 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_201
timestamp 1623621585
transform 1 0 19596 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2083_
timestamp 1623621585
transform 1 0 20700 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _2084_
timestamp 1623621585
transform 1 0 21896 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_209
timestamp 1623621585
transform 1 0 20332 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_222
timestamp 1623621585
transform 1 0 21528 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1494_
timestamp 1623621585
transform 1 0 23368 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1495_
timestamp 1623621585
transform 1 0 24012 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_238
timestamp 1623621585
transform 1 0 23000 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_245
timestamp 1623621585
transform 1 0 23644 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2192_
timestamp 1623621585
transform 1 0 25852 0 1 39712
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1623621585
transform 1 0 24748 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1623621585
transform 1 0 25208 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_253
timestamp 1623621585
transform 1 0 24380 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_258
timestamp 1623621585
transform 1 0 24840 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_265
timestamp 1623621585
transform 1 0 25484 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1904_
timestamp 1623621585
transform 1 0 27784 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_286
timestamp 1623621585
transform 1 0 27416 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_294
timestamp 1623621585
transform 1 0 28152 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1623621585
transform -1 0 28888 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_69_298
timestamp 1623621585
transform 1 0 28520 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _2021_
timestamp 1623621585
transform 1 0 2484 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1623621585
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output264
timestamp 1623621585
transform 1 0 1748 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1623621585
transform 1 0 1380 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_11
timestamp 1623621585
transform 1 0 2116 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_2  _1247_
timestamp 1623621585
transform 1 0 3680 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1793_
timestamp 1623621585
transform 1 0 4692 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_24
timestamp 1623621585
transform 1 0 3312 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_35
timestamp 1623621585
transform 1 0 4324 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_45
timestamp 1623621585
transform 1 0 5244 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1778_
timestamp 1623621585
transform 1 0 5612 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2069_
timestamp 1623621585
transform 1 0 6808 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1623621585
transform 1 0 6348 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_52
timestamp 1623621585
transform 1 0 5888 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_56
timestamp 1623621585
transform 1 0 6256 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_58
timestamp 1623621585
transform 1 0 6440 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_71
timestamp 1623621585
transform 1 0 7636 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_83
timestamp 1623621585
transform 1 0 8740 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1623621585
transform 1 0 11592 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_wb_clk_i
timestamp 1623621585
transform 1 0 10948 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_95
timestamp 1623621585
transform 1 0 9844 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_110
timestamp 1623621585
transform 1 0 11224 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1100_
timestamp 1623621585
transform 1 0 12420 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_70_115
timestamp 1623621585
transform 1 0 11684 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_70_131
timestamp 1623621585
transform 1 0 13156 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2297_
timestamp 1623621585
transform 1 0 13984 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1623621585
transform 1 0 13892 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_159
timestamp 1623621585
transform 1 0 15732 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1870_
timestamp 1623621585
transform 1 0 17848 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1623621585
transform 1 0 16836 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_172
timestamp 1623621585
transform 1 0 16928 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_180
timestamp 1623621585
transform 1 0 17664 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_4  _1949_
timestamp 1623621585
transform 1 0 18492 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2168_
timestamp 1623621585
transform 1 0 19964 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_70_185
timestamp 1623621585
transform 1 0 18124 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_201
timestamp 1623621585
transform 1 0 19596 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1623621585
transform 1 0 22080 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_221
timestamp 1623621585
transform 1 0 21436 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_227
timestamp 1623621585
transform 1 0 21988 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_4  _1467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 22908 0 -1 40800
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_70_229
timestamp 1623621585
transform 1 0 22172 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1500_
timestamp 1623621585
transform 1 0 25576 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_70_259
timestamp 1623621585
transform 1 0 24932 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_265
timestamp 1623621585
transform 1 0 25484 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1905_
timestamp 1623621585
transform 1 0 27784 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1623621585
transform 1 0 27324 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_275
timestamp 1623621585
transform 1 0 26404 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_283
timestamp 1623621585
transform 1 0 27140 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_286
timestamp 1623621585
transform 1 0 27416 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_294
timestamp 1623621585
transform 1 0 28152 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1623621585
transform -1 0 28888 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_298
timestamp 1623621585
transform 1 0 28520 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _2022_
timestamp 1623621585
transform 1 0 1748 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1623621585
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output268
timestamp 1623621585
transform 1 0 2944 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_3
timestamp 1623621585
transform 1 0 1380 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_16
timestamp 1623621585
transform 1 0 2576 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1242_
timestamp 1623621585
transform 1 0 4232 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2187_
timestamp 1623621585
transform 1 0 4968 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1623621585
transform 1 0 3772 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_24
timestamp 1623621585
transform 1 0 3312 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_28
timestamp 1623621585
transform 1 0 3680 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_30
timestamp 1623621585
transform 1 0 3864 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_37
timestamp 1623621585
transform 1 0 4508 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_41
timestamp 1623621585
transform 1 0 4876 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1518_
timestamp 1623621585
transform 1 0 6808 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_71_58
timestamp 1623621585
transform 1 0 6440 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1709_
timestamp 1623621585
transform 1 0 8004 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _2211_
timestamp 1623621585
transform 1 0 9476 0 1 40800
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1623621585
transform 1 0 9016 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_71
timestamp 1623621585
transform 1 0 7636 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_78
timestamp 1623621585
transform 1 0 8280 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_87
timestamp 1623621585
transform 1 0 9108 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_108
timestamp 1623621585
transform 1 0 11040 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _1838_
timestamp 1623621585
transform 1 0 12880 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_71_120
timestamp 1623621585
transform 1 0 12144 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_71_136
timestamp 1623621585
transform 1 0 13616 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2298_
timestamp 1623621585
transform 1 0 15456 0 1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1623621585
transform 1 0 14260 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_142
timestamp 1623621585
transform 1 0 14168 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_144
timestamp 1623621585
transform 1 0 14352 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2282_
timestamp 1623621585
transform 1 0 17572 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_175
timestamp 1623621585
transform 1 0 17204 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1623621585
transform 1 0 19504 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_195
timestamp 1623621585
transform 1 0 19044 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_199
timestamp 1623621585
transform 1 0 19412 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_201
timestamp 1623621585
transform 1 0 19596 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1560_
timestamp 1623621585
transform 1 0 20516 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1679_
timestamp 1623621585
transform 1 0 21988 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_209
timestamp 1623621585
transform 1 0 20332 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_220
timestamp 1623621585
transform 1 0 21344 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_226
timestamp 1623621585
transform 1 0 21896 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__a211oi_4  _1474_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 22724 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_230
timestamp 1623621585
transform 1 0 22264 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_234
timestamp 1623621585
transform 1 0 22632 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_251
timestamp 1623621585
transform 1 0 24196 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1623621585
transform 1 0 24748 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1623621585
transform 1 0 25944 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1623621585
transform 1 0 25300 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_258
timestamp 1623621585
transform 1 0 24840 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_262
timestamp 1623621585
transform 1 0 25208 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_266
timestamp 1623621585
transform 1 0 25576 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_273
timestamp 1623621585
transform 1 0 26220 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1906_
timestamp 1623621585
transform 1 0 27232 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1623621585
transform 1 0 27968 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1623621585
transform 1 0 26588 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_280
timestamp 1623621585
transform 1 0 26864 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_288
timestamp 1623621585
transform 1 0 27600 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_295
timestamp 1623621585
transform 1 0 28244 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1623621585
transform -1 0 28888 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1261_
timestamp 1623621585
transform 1 0 2668 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1368_
timestamp 1623621585
transform 1 0 1472 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2216_
timestamp 1623621585
transform 1 0 1380 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1623621585
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1623621585
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_72_3
timestamp 1623621585
transform 1 0 1380 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_13
timestamp 1623621585
transform 1 0 2300 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_19
timestamp 1623621585
transform 1 0 2852 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_30
timestamp 1623621585
transform 1 0 3864 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_27
timestamp 1623621585
transform 1 0 3588 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_34
timestamp 1623621585
transform 1 0 4232 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1623621585
transform 1 0 3312 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1623621585
transform 1 0 3772 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1776_
timestamp 1623621585
transform 1 0 4232 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1241_
timestamp 1623621585
transform 1 0 3680 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_37
timestamp 1623621585
transform 1 0 4508 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1791_
timestamp 1623621585
transform 1 0 4600 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1779_
timestamp 1623621585
transform 1 0 4876 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_44
timestamp 1623621585
transform 1 0 5152 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_44
timestamp 1623621585
transform 1 0 5152 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _2068_
timestamp 1623621585
transform 1 0 7176 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1623621585
transform 1 0 6348 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_56
timestamp 1623621585
transform 1 0 6256 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_58
timestamp 1623621585
transform 1 0 6440 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_56
timestamp 1623621585
transform 1 0 6256 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_68
timestamp 1623621585
transform 1 0 7360 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__a21boi_1  _1406_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 8372 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _1409_
timestamp 1623621585
transform 1 0 9292 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1410_
timestamp 1623621585
transform 1 0 9476 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1623621585
transform 1 0 9016 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_75
timestamp 1623621585
transform 1 0 8004 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_85
timestamp 1623621585
transform 1 0 8924 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_80
timestamp 1623621585
transform 1 0 8464 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_87
timestamp 1623621585
transform 1 0 9108 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1375_
timestamp 1623621585
transform 1 0 10212 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1623621585
transform 1 0 11592 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_95
timestamp 1623621585
transform 1 0 9844 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_102
timestamp 1623621585
transform 1 0 10488 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_95
timestamp 1623621585
transform 1 0 9844 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_107
timestamp 1623621585
transform 1 0 10948 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _1969_
timestamp 1623621585
transform 1 0 12604 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2280_
timestamp 1623621585
transform 1 0 12236 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_72_115
timestamp 1623621585
transform 1 0 11684 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_123
timestamp 1623621585
transform 1 0 12420 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_134
timestamp 1623621585
transform 1 0 13432 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_119
timestamp 1623621585
transform 1 0 12052 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_137
timestamp 1623621585
transform 1 0 13708 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__nor2b_1  _1212_
timestamp 1623621585
transform 1 0 14904 0 1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1809_
timestamp 1623621585
transform 1 0 13800 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1623621585
transform 1 0 14260 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1623621585
transform 1 0 14076 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1623621585
transform 1 0 15180 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_144
timestamp 1623621585
transform 1 0 14352 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_73_155
timestamp 1623621585
transform 1 0 15364 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1871_
timestamp 1623621585
transform 1 0 17296 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1950_
timestamp 1623621585
transform 1 0 16008 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1951_
timestamp 1623621585
transform 1 0 17204 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1623621585
transform 1 0 16836 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_165
timestamp 1623621585
transform 1 0 16284 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_172
timestamp 1623621585
transform 1 0 16928 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_179
timestamp 1623621585
transform 1 0 17572 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_161
timestamp 1623621585
transform 1 0 15916 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_171
timestamp 1623621585
transform 1 0 16836 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1205_
timestamp 1623621585
transform 1 0 18400 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1948_
timestamp 1623621585
transform 1 0 19136 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1623621585
transform 1 0 19504 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_191
timestamp 1623621585
transform 1 0 18676 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1623621585
transform 1 0 19044 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_205
timestamp 1623621585
transform 1 0 19964 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_184
timestamp 1623621585
transform 1 0 18032 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_192
timestamp 1623621585
transform 1 0 18768 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_201
timestamp 1623621585
transform 1 0 19596 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1673_
timestamp 1623621585
transform 1 0 22080 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1681_
timestamp 1623621585
transform 1 0 21436 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1623621585
transform 1 0 22080 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_217
timestamp 1623621585
transform 1 0 21068 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_224
timestamp 1623621585
transform 1 0 21712 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_213
timestamp 1623621585
transform 1 0 20700 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_225
timestamp 1623621585
transform 1 0 21804 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1468_
timestamp 1623621585
transform 1 0 23092 0 1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1469_
timestamp 1623621585
transform 1 0 23920 0 1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _1471_
timestamp 1623621585
transform 1 0 24012 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_229
timestamp 1623621585
transform 1 0 22172 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_241
timestamp 1623621585
transform 1 0 23276 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_231
timestamp 1623621585
transform 1 0 22356 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_244
timestamp 1623621585
transform 1 0 23552 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_258
timestamp 1623621585
transform 1 0 24840 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_253
timestamp 1623621585
transform 1 0 24380 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_257
timestamp 1623621585
transform 1 0 24748 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1623621585
transform 1 0 24748 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _1496_
timestamp 1623621585
transform 1 0 25116 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1475_
timestamp 1623621585
transform 1 0 25208 0 1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_73_267
timestamp 1623621585
transform 1 0 25668 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_268
timestamp 1623621585
transform 1 0 25760 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1498_
timestamp 1623621585
transform 1 0 26128 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _2193_
timestamp 1623621585
transform 1 0 26036 0 1 41888
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_72_278
timestamp 1623621585
transform 1 0 26680 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_286
timestamp 1623621585
transform 1 0 27416 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_284
timestamp 1623621585
transform 1 0 27232 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1623621585
transform 1 0 27324 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_288
timestamp 1623621585
transform 1 0 27600 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_290
timestamp 1623621585
transform 1 0 27784 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1623621585
transform 1 0 27968 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1907_
timestamp 1623621585
transform 1 0 27876 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_295
timestamp 1623621585
transform 1 0 28244 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_295
timestamp 1623621585
transform 1 0 28244 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1623621585
transform -1 0 28888 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1623621585
transform -1 0 28888 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1623621585
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output269
timestamp 1623621585
transform 1 0 1748 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output272
timestamp 1623621585
transform 1 0 2484 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_3
timestamp 1623621585
transform 1 0 1380 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_11
timestamp 1623621585
transform 1 0 2116 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_19
timestamp 1623621585
transform 1 0 2852 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1246_
timestamp 1623621585
transform 1 0 3496 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1774_
timestamp 1623621585
transform 1 0 4508 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_74_25
timestamp 1623621585
transform 1 0 3404 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_33
timestamp 1623621585
transform 1 0 4140 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_40
timestamp 1623621585
transform 1 0 4784 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1623621585
transform 1 0 6348 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_52
timestamp 1623621585
transform 1 0 5888 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_56
timestamp 1623621585
transform 1 0 6256 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_58
timestamp 1623621585
transform 1 0 6440 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1402_
timestamp 1623621585
transform 1 0 7636 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1517_
timestamp 1623621585
transform 1 0 8832 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_70
timestamp 1623621585
transform 1 0 7544 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_74
timestamp 1623621585
transform 1 0 7912 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_82
timestamp 1623621585
transform 1 0 8648 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_88
timestamp 1623621585
transform 1 0 9200 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1211_
timestamp 1623621585
transform 1 0 9752 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_1  _1214_
timestamp 1623621585
transform 1 0 10764 0 -1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1623621585
transform 1 0 11592 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_98
timestamp 1623621585
transform 1 0 10120 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_104
timestamp 1623621585
transform 1 0 10672 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_110
timestamp 1623621585
transform 1 0 11224 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1968_
timestamp 1623621585
transform 1 0 12052 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _2296_
timestamp 1623621585
transform 1 0 13708 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_74_115
timestamp 1623621585
transform 1 0 11684 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_128
timestamp 1623621585
transform 1 0 12880 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_136
timestamp 1623621585
transform 1 0 13616 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_156
timestamp 1623621585
transform 1 0 15456 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1623621585
transform 1 0 16836 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_168
timestamp 1623621585
transform 1 0 16560 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_172
timestamp 1623621585
transform 1 0 16928 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2241_
timestamp 1623621585
transform 1 0 18400 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_74_184
timestamp 1623621585
transform 1 0 18032 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_204
timestamp 1623621585
transform 1 0 19872 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1674_
timestamp 1623621585
transform 1 0 21436 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1623621585
transform 1 0 22080 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_216
timestamp 1623621585
transform 1 0 20976 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_220
timestamp 1623621585
transform 1 0 21344 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_224
timestamp 1623621585
transform 1 0 21712 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1470_
timestamp 1623621585
transform 1 0 23736 0 -1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _2087_
timestamp 1623621585
transform 1 0 22540 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_74_229
timestamp 1623621585
transform 1 0 22172 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_242
timestamp 1623621585
transform 1 0 23368 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_251
timestamp 1623621585
transform 1 0 24196 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1497_
timestamp 1623621585
transform 1 0 25116 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_259
timestamp 1623621585
transform 1 0 24932 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_267
timestamp 1623621585
transform 1 0 25668 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1908_
timestamp 1623621585
transform 1 0 27876 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1911_
timestamp 1623621585
transform 1 0 26588 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1623621585
transform 1 0 27324 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_275
timestamp 1623621585
transform 1 0 26404 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_281
timestamp 1623621585
transform 1 0 26956 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_286
timestamp 1623621585
transform 1 0 27416 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_290
timestamp 1623621585
transform 1 0 27784 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_295
timestamp 1623621585
transform 1 0 28244 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1623621585
transform -1 0 28888 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1623621585
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output270
timestamp 1623621585
transform 1 0 1748 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output274
timestamp 1623621585
transform 1 0 2484 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_3
timestamp 1623621585
transform 1 0 1380 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_11
timestamp 1623621585
transform 1 0 2116 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_19
timestamp 1623621585
transform 1 0 2852 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1360_
timestamp 1623621585
transform 1 0 4232 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1364_
timestamp 1623621585
transform 1 0 4876 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1623621585
transform 1 0 3772 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_27
timestamp 1623621585
transform 1 0 3588 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_30
timestamp 1623621585
transform 1 0 3864 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_37
timestamp 1623621585
transform 1 0 4508 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_44
timestamp 1623621585
transform 1 0 5152 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1713_
timestamp 1623621585
transform 1 0 5704 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_53
timestamp 1623621585
transform 1 0 5980 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_65
timestamp 1623621585
transform 1 0 7084 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1408_
timestamp 1623621585
transform 1 0 9476 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1623621585
transform 1 0 9016 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_77
timestamp 1623621585
transform 1 0 8188 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_85
timestamp 1623621585
transform 1 0 8924 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_87
timestamp 1623621585
transform 1 0 9108 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2239_
timestamp 1623621585
transform 1 0 10856 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_wb_clk_i
timestamp 1623621585
transform 1 0 10120 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_94
timestamp 1623621585
transform 1 0 9752 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_101
timestamp 1623621585
transform 1 0 10396 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_105
timestamp 1623621585
transform 1 0 10764 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_122
timestamp 1623621585
transform 1 0 12328 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_134
timestamp 1623621585
transform 1 0 13432 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2240_
timestamp 1623621585
transform 1 0 14996 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1623621585
transform 1 0 14260 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_142
timestamp 1623621585
transform 1 0 14168 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_144
timestamp 1623621585
transform 1 0 14352 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_150
timestamp 1623621585
transform 1 0 14904 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_wb_clk_i
timestamp 1623621585
transform 1 0 17388 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_167
timestamp 1623621585
transform 1 0 16468 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_175
timestamp 1623621585
transform 1 0 17204 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_180
timestamp 1623621585
transform 1 0 17664 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__nor2b_1  _1210_
timestamp 1623621585
transform 1 0 18584 0 1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2169_
timestamp 1623621585
transform 1 0 19964 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1623621585
transform 1 0 19504 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_188
timestamp 1623621585
transform 1 0 18400 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_195
timestamp 1623621585
transform 1 0 19044 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_199
timestamp 1623621585
transform 1 0 19412 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_201
timestamp 1623621585
transform 1 0 19596 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2086_
timestamp 1623621585
transform 1 0 21804 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_75_221
timestamp 1623621585
transform 1 0 21436 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1675_
timestamp 1623621585
transform 1 0 23000 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1623621585
transform 1 0 24104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_234
timestamp 1623621585
transform 1 0 22632 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_241
timestamp 1623621585
transform 1 0 23276 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_249
timestamp 1623621585
transform 1 0 24012 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1484_
timestamp 1623621585
transform 1 0 25208 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1623621585
transform 1 0 24748 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1623621585
transform 1 0 25852 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_253
timestamp 1623621585
transform 1 0 24380 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_258
timestamp 1623621585
transform 1 0 24840 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_265
timestamp 1623621585
transform 1 0 25484 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_272
timestamp 1623621585
transform 1 0 26128 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1909_
timestamp 1623621585
transform 1 0 27876 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1910_
timestamp 1623621585
transform 1 0 27140 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1623621585
transform 1 0 26496 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_279
timestamp 1623621585
transform 1 0 26772 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_287
timestamp 1623621585
transform 1 0 27508 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_295
timestamp 1623621585
transform 1 0 28244 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1623621585
transform -1 0 28888 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1623621585
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output273
timestamp 1623621585
transform 1 0 1748 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output275
timestamp 1623621585
transform 1 0 2484 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  INSDIODE3_0
timestamp 1623621585
transform 1 0 3036 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_3
timestamp 1623621585
transform 1 0 1380 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_11
timestamp 1623621585
transform 1 0 2116 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_19
timestamp 1623621585
transform 1 0 2852 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2186_
timestamp 1623621585
transform 1 0 4232 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output277
timestamp 1623621585
transform 1 0 3220 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_27
timestamp 1623621585
transform 1 0 3588 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_33
timestamp 1623621585
transform 1 0 4140 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _1401_
timestamp 1623621585
transform 1 0 6808 0 -1 44064
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1623621585
transform 1 0 6348 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_50
timestamp 1623621585
transform 1 0 5704 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_56
timestamp 1623621585
transform 1 0 6256 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_58
timestamp 1623621585
transform 1 0 6440 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_67
timestamp 1623621585
transform 1 0 7268 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1397_
timestamp 1623621585
transform 1 0 7636 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1412_
timestamp 1623621585
transform 1 0 8280 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_wb_clk_i
timestamp 1623621585
transform 1 0 8924 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_74
timestamp 1623621585
transform 1 0 7912 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_81
timestamp 1623621585
transform 1 0 8556 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_88
timestamp 1623621585
transform 1 0 9200 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2210_
timestamp 1623621585
transform 1 0 9568 0 -1 44064
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1623621585
transform 1 0 11592 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_109
timestamp 1623621585
transform 1 0 11132 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_113
timestamp 1623621585
transform 1 0 11500 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1378_
timestamp 1623621585
transform 1 0 13248 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_115
timestamp 1623621585
transform 1 0 11684 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_127
timestamp 1623621585
transform 1 0 12788 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_131
timestamp 1623621585
transform 1 0 13156 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_135
timestamp 1623621585
transform 1 0 13524 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1421_
timestamp 1623621585
transform 1 0 14720 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_147
timestamp 1623621585
transform 1 0 14628 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_152
timestamp 1623621585
transform 1 0 15088 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1454_
timestamp 1623621585
transform 1 0 17572 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1623621585
transform 1 0 16836 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_164
timestamp 1623621585
transform 1 0 16192 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_170
timestamp 1623621585
transform 1 0 16744 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_172
timestamp 1623621585
transform 1 0 16928 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_178
timestamp 1623621585
transform 1 0 17480 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_182
timestamp 1623621585
transform 1 0 17848 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_4  _1516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 18400 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_76_204
timestamp 1623621585
transform 1 0 19872 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1559_
timestamp 1623621585
transform 1 0 20332 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1623621585
transform 1 0 22080 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_208
timestamp 1623621585
transform 1 0 20240 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_218
timestamp 1623621585
transform 1 0 21160 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_226
timestamp 1623621585
transform 1 0 21896 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1209_
timestamp 1623621585
transform 1 0 23552 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_229
timestamp 1623621585
transform 1 0 22172 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_241
timestamp 1623621585
transform 1 0 23276 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_248
timestamp 1623621585
transform 1 0 23920 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1485_
timestamp 1623621585
transform 1 0 25208 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1493_
timestamp 1623621585
transform 1 0 24380 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1623621585
transform 1 0 25944 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_76_252
timestamp 1623621585
transform 1 0 24288 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_257
timestamp 1623621585
transform 1 0 24748 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_261
timestamp 1623621585
transform 1 0 25116 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_266
timestamp 1623621585
transform 1 0 25576 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_273
timestamp 1623621585
transform 1 0 26220 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1912_
timestamp 1623621585
transform 1 0 27876 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1914_
timestamp 1623621585
transform 1 0 26588 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1623621585
transform 1 0 27324 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_281
timestamp 1623621585
transform 1 0 26956 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_286
timestamp 1623621585
transform 1 0 27416 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_290
timestamp 1623621585
transform 1 0 27784 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_295
timestamp 1623621585
transform 1 0 28244 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1623621585
transform -1 0 28888 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1362_
timestamp 1623621585
transform 1 0 3036 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2024_
timestamp 1623621585
transform 1 0 1840 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1623621585
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_3
timestamp 1623621585
transform 1 0 1380 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_7
timestamp 1623621585
transform 1 0 1748 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_17
timestamp 1623621585
transform 1 0 2668 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1519_
timestamp 1623621585
transform 1 0 4784 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1623621585
transform 1 0 3772 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_24
timestamp 1623621585
transform 1 0 3312 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_28
timestamp 1623621585
transform 1 0 3680 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_30
timestamp 1623621585
transform 1 0 3864 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_38
timestamp 1623621585
transform 1 0 4600 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _2065_
timestamp 1623621585
transform 1 0 6440 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_77_49
timestamp 1623621585
transform 1 0 5612 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_57
timestamp 1623621585
transform 1 0 6348 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_67
timestamp 1623621585
transform 1 0 7268 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1413_
timestamp 1623621585
transform 1 0 7728 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1416_
timestamp 1623621585
transform 1 0 9476 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1623621585
transform 1 0 9016 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_71
timestamp 1623621585
transform 1 0 7636 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_76
timestamp 1623621585
transform 1 0 8096 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_84
timestamp 1623621585
transform 1 0 8832 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_87
timestamp 1623621585
transform 1 0 9108 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1411_
timestamp 1623621585
transform 1 0 10212 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_wb_clk_i
timestamp 1623621585
transform 1 0 11132 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_95
timestamp 1623621585
transform 1 0 9844 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_102
timestamp 1623621585
transform 1 0 10488 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_108
timestamp 1623621585
transform 1 0 11040 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_112
timestamp 1623621585
transform 1 0 11408 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _1377_
timestamp 1623621585
transform 1 0 13156 0 1 44064
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_77_124
timestamp 1623621585
transform 1 0 12512 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_130
timestamp 1623621585
transform 1 0 13064 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_136
timestamp 1623621585
transform 1 0 13616 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1623621585
transform 1 0 14260 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_142
timestamp 1623621585
transform 1 0 14168 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_144
timestamp 1623621585
transform 1 0 14352 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_156
timestamp 1623621585
transform 1 0 15456 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1455_
timestamp 1623621585
transform 1 0 16652 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1514_
timestamp 1623621585
transform 1 0 17848 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1700_
timestamp 1623621585
transform 1 0 16008 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_165
timestamp 1623621585
transform 1 0 16284 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_178
timestamp 1623621585
transform 1 0 17480 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1509_
timestamp 1623621585
transform 1 0 18768 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1623621585
transform 1 0 19504 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_wb_clk_i
timestamp 1623621585
transform 1 0 19964 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_188
timestamp 1623621585
transform 1 0 18400 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_196
timestamp 1623621585
transform 1 0 19136 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_201
timestamp 1623621585
transform 1 0 19596 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1556_
timestamp 1623621585
transform 1 0 21252 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_wb_clk_i
timestamp 1623621585
transform 1 0 21988 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_208
timestamp 1623621585
transform 1 0 20240 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_216
timestamp 1623621585
transform 1 0 20976 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_223
timestamp 1623621585
transform 1 0 21620 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1488_
timestamp 1623621585
transform 1 0 23368 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1490_
timestamp 1623621585
transform 1 0 24012 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_230
timestamp 1623621585
transform 1 0 22264 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_245
timestamp 1623621585
transform 1 0 23644 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _2194_
timestamp 1623621585
transform 1 0 25484 0 1 44064
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1623621585
transform 1 0 24748 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_253
timestamp 1623621585
transform 1 0 24380 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_258
timestamp 1623621585
transform 1 0 24840 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_264
timestamp 1623621585
transform 1 0 25392 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1913_
timestamp 1623621585
transform 1 0 27876 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_282
timestamp 1623621585
transform 1 0 27048 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_290
timestamp 1623621585
transform 1 0 27784 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_295
timestamp 1623621585
transform 1 0 28244 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1623621585
transform -1 0 28888 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2023_
timestamp 1623621585
transform 1 0 2484 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1623621585
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output276
timestamp 1623621585
transform 1 0 1748 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_3
timestamp 1623621585
transform 1 0 1380 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_11
timestamp 1623621585
transform 1 0 2116 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2028_
timestamp 1623621585
transform 1 0 3956 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_78_24
timestamp 1623621585
transform 1 0 3312 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_30
timestamp 1623621585
transform 1 0 3864 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_40
timestamp 1623621585
transform 1 0 4784 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1396_
timestamp 1623621585
transform 1 0 6808 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1714_
timestamp 1623621585
transform 1 0 5704 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1623621585
transform 1 0 6348 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_48
timestamp 1623621585
transform 1 0 5520 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_53
timestamp 1623621585
transform 1 0 5980 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_58
timestamp 1623621585
transform 1 0 6440 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_65
timestamp 1623621585
transform 1 0 7084 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1400_
timestamp 1623621585
transform 1 0 7544 0 -1 45152
box -38 -48 1326 592
use sky130_fd_sc_hd__o21bai_1  _1415_
timestamp 1623621585
transform 1 0 9200 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_69
timestamp 1623621585
transform 1 0 7452 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_84
timestamp 1623621585
transform 1 0 8832 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1623621585
transform 1 0 11592 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_94
timestamp 1623621585
transform 1 0 9752 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_106
timestamp 1623621585
transform 1 0 10856 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_2  _1438_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 12788 0 -1 45152
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_78_115
timestamp 1623621585
transform 1 0 11684 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_137
timestamp 1623621585
transform 1 0 13708 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2ai_2  _1440_
timestamp 1623621585
transform 1 0 14076 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _2071_
timestamp 1623621585
transform 1 0 15640 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_78_153
timestamp 1623621585
transform 1 0 15180 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_157
timestamp 1623621585
transform 1 0 15548 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__o31ai_4  _1515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 17664 0 -1 45152
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1623621585
transform 1 0 16836 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_167
timestamp 1623621585
transform 1 0 16468 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_172
timestamp 1623621585
transform 1 0 16928 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _2189_
timestamp 1623621585
transform 1 0 19596 0 -1 45152
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_78_197
timestamp 1623621585
transform 1 0 19228 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1623621585
transform 1 0 22080 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_218
timestamp 1623621585
transform 1 0 21160 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_226
timestamp 1623621585
transform 1 0 21896 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _1472_
timestamp 1623621585
transform 1 0 23276 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1491_
timestamp 1623621585
transform 1 0 24012 0 -1 45152
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1669_
timestamp 1623621585
transform 1 0 22632 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_229
timestamp 1623621585
transform 1 0 22172 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_233
timestamp 1623621585
transform 1 0 22540 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_237
timestamp 1623621585
transform 1 0 22908 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_244
timestamp 1623621585
transform 1 0 23552 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_248
timestamp 1623621585
transform 1 0 23920 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__o21bai_1  _1492_
timestamp 1623621585
transform 1 0 24840 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1623621585
transform 1 0 26036 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_254
timestamp 1623621585
transform 1 0 24472 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_264
timestamp 1623621585
transform 1 0 25392 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_270
timestamp 1623621585
transform 1 0 25944 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_274
timestamp 1623621585
transform 1 0 26312 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1915_
timestamp 1623621585
transform 1 0 27784 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1623621585
transform 1 0 27324 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1623621585
transform 1 0 26680 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_281
timestamp 1623621585
transform 1 0 26956 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_286
timestamp 1623621585
transform 1 0 27416 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_294
timestamp 1623621585
transform 1 0 28152 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1623621585
transform -1 0 28888 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_78_298
timestamp 1623621585
transform 1 0 28520 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_3
timestamp 1623621585
transform 1 0 1380 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_3
timestamp 1623621585
transform 1 0 1380 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output278
timestamp 1623621585
transform 1 0 1748 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1623621585
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1623621585
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1366_
timestamp 1623621585
transform 1 0 1564 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_80_19
timestamp 1623621585
transform 1 0 2852 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_11
timestamp 1623621585
transform 1 0 2116 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_79_14
timestamp 1623621585
transform 1 0 2392 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_20
timestamp 1623621585
transform 1 0 2944 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _2026_
timestamp 1623621585
transform 1 0 3036 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1771_
timestamp 1623621585
transform 1 0 3036 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2025_
timestamp 1623621585
transform 1 0 4232 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2027_
timestamp 1623621585
transform 1 0 4508 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1623621585
transform 1 0 3772 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_25
timestamp 1623621585
transform 1 0 3404 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_30
timestamp 1623621585
transform 1 0 3864 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_43
timestamp 1623621585
transform 1 0 5060 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_80_30
timestamp 1623621585
transform 1 0 3864 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_36
timestamp 1623621585
transform 1 0 4416 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1777_
timestamp 1623621585
transform 1 0 5704 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2066_
timestamp 1623621585
transform 1 0 5796 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1623621585
transform 1 0 6348 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_60
timestamp 1623621585
transform 1 0 6624 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_46
timestamp 1623621585
transform 1 0 5336 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_53
timestamp 1623621585
transform 1 0 5980 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_58
timestamp 1623621585
transform 1 0 6440 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_1  _1414_
timestamp 1623621585
transform 1 0 7912 0 1 45152
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1417_
timestamp 1623621585
transform 1 0 9476 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1623621585
transform 1 0 9016 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_72
timestamp 1623621585
transform 1 0 7728 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_79
timestamp 1623621585
transform 1 0 8372 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_85
timestamp 1623621585
transform 1 0 8924 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_87
timestamp 1623621585
transform 1 0 9108 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_70
timestamp 1623621585
transform 1 0 7544 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_82
timestamp 1623621585
transform 1 0 8648 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_1  _1428_
timestamp 1623621585
transform 1 0 10580 0 -1 46240
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1730_
timestamp 1623621585
transform 1 0 9936 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2207_
timestamp 1623621585
transform 1 0 11132 0 1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1623621585
transform 1 0 11592 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_95
timestamp 1623621585
transform 1 0 9844 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_107
timestamp 1623621585
transform 1 0 10948 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_94
timestamp 1623621585
transform 1 0 9752 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_99
timestamp 1623621585
transform 1 0 10212 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_110
timestamp 1623621585
transform 1 0 11224 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1380_
timestamp 1623621585
transform 1 0 12880 0 -1 46240
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1436_
timestamp 1623621585
transform 1 0 12236 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1437_
timestamp 1623621585
transform 1 0 13248 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_128
timestamp 1623621585
transform 1 0 12880 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_115
timestamp 1623621585
transform 1 0 11684 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_124
timestamp 1623621585
transform 1 0 12512 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_141
timestamp 1623621585
transform 1 0 14076 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_144
timestamp 1623621585
transform 1 0 14352 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_142
timestamp 1623621585
transform 1 0 14168 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_138
timestamp 1623621585
transform 1 0 13800 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1623621585
transform 1 0 14260 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1379_
timestamp 1623621585
transform 1 0 14444 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_80_154
timestamp 1623621585
transform 1 0 15272 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_148
timestamp 1623621585
transform 1 0 14720 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _2047_
timestamp 1623621585
transform 1 0 14812 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_79_158
timestamp 1623621585
transform 1 0 15640 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1744_
timestamp 1623621585
transform 1 0 15640 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1453_
timestamp 1623621585
transform 1 0 17296 0 -1 46240
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _1456_
timestamp 1623621585
transform 1 0 17572 0 1 45152
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _2072_
timestamp 1623621585
transform 1 0 16192 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1623621585
transform 1 0 16836 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_173
timestamp 1623621585
transform 1 0 17020 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_80_161
timestamp 1623621585
transform 1 0 15916 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_169
timestamp 1623621585
transform 1 0 16652 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_172
timestamp 1623621585
transform 1 0 16928 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_181
timestamp 1623621585
transform 1 0 17756 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1460_
timestamp 1623621585
transform 1 0 19688 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1513_
timestamp 1623621585
transform 1 0 18124 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1623621585
transform 1 0 19504 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_192
timestamp 1623621585
transform 1 0 18768 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_201
timestamp 1623621585
transform 1 0 19596 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_188
timestamp 1623621585
transform 1 0 18400 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_200
timestamp 1623621585
transform 1 0 19504 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2170_
timestamp 1623621585
transform 1 0 21160 0 1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1623621585
transform 1 0 22080 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_213
timestamp 1623621585
transform 1 0 20700 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_217
timestamp 1623621585
transform 1 0 21068 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_206
timestamp 1623621585
transform 1 0 20056 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_218
timestamp 1623621585
transform 1 0 21160 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_226
timestamp 1623621585
transform 1 0 21896 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__nand3_2  _1476_
timestamp 1623621585
transform 1 0 24196 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1558_
timestamp 1623621585
transform 1 0 23000 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2089_
timestamp 1623621585
transform 1 0 23000 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_79_234
timestamp 1623621585
transform 1 0 22632 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_247
timestamp 1623621585
transform 1 0 23828 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_80_229
timestamp 1623621585
transform 1 0 22172 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_237
timestamp 1623621585
transform 1 0 22908 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_247
timestamp 1623621585
transform 1 0 23828 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_259
timestamp 1623621585
transform 1 0 24932 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_258
timestamp 1623621585
transform 1 0 24840 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_255
timestamp 1623621585
transform 1 0 24564 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1623621585
transform 1 0 24748 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_267
timestamp 1623621585
transform 1 0 25668 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_263
timestamp 1623621585
transform 1 0 25300 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_265
timestamp 1623621585
transform 1 0 25484 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1623621585
transform 1 0 25392 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1473_
timestamp 1623621585
transform 1 0 25208 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_274
timestamp 1623621585
transform 1 0 26312 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_272
timestamp 1623621585
transform 1 0 26128 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1623621585
transform 1 0 26036 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1489_
timestamp 1623621585
transform 1 0 25852 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_281
timestamp 1623621585
transform 1 0 26956 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1623621585
transform 1 0 26680 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1623621585
transform 1 0 26864 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_286
timestamp 1623621585
transform 1 0 27416 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_291
timestamp 1623621585
transform 1 0 27876 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_283
timestamp 1623621585
transform 1 0 27140 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1623621585
transform 1 0 27324 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1917_
timestamp 1623621585
transform 1 0 27784 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1916_
timestamp 1623621585
transform 1 0 27508 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_294
timestamp 1623621585
transform 1 0 28152 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1623621585
transform -1 0 28888 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1623621585
transform -1 0 28888 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_298
timestamp 1623621585
transform 1 0 28520 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2217_
timestamp 1623621585
transform 1 0 1380 0 1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1623621585
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_19
timestamp 1623621585
transform 1 0 2852 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1772_
timestamp 1623621585
transform 1 0 4232 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1775_
timestamp 1623621585
transform 1 0 4876 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1623621585
transform 1 0 3772 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_27
timestamp 1623621585
transform 1 0 3588 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_30
timestamp 1623621585
transform 1 0 3864 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_37
timestamp 1623621585
transform 1 0 4508 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_44
timestamp 1623621585
transform 1 0 5152 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1717_
timestamp 1623621585
transform 1 0 5980 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_81_52
timestamp 1623621585
transform 1 0 5888 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_56
timestamp 1623621585
transform 1 0 6256 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_68
timestamp 1623621585
transform 1 0 7360 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1729_
timestamp 1623621585
transform 1 0 8372 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1623621585
transform 1 0 9016 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_76
timestamp 1623621585
transform 1 0 8096 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_82
timestamp 1623621585
transform 1 0 8648 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_87
timestamp 1623621585
transform 1 0 9108 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_91
timestamp 1623621585
transform 1 0 9476 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1429_
timestamp 1623621585
transform 1 0 11224 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2056_
timestamp 1623621585
transform 1 0 9568 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_81_101
timestamp 1623621585
transform 1 0 10396 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_109
timestamp 1623621585
transform 1 0 11132 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _2048_
timestamp 1623621585
transform 1 0 13064 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_81_119
timestamp 1623621585
transform 1 0 12052 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_127
timestamp 1623621585
transform 1 0 12788 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1525_
timestamp 1623621585
transform 1 0 14720 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1623621585
transform 1 0 14260 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_139
timestamp 1623621585
transform 1 0 13892 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_144
timestamp 1623621585
transform 1 0 14352 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_157
timestamp 1623621585
transform 1 0 15548 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1564_
timestamp 1623621585
transform 1 0 16192 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1701_
timestamp 1623621585
transform 1 0 17388 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_81_163
timestamp 1623621585
transform 1 0 16100 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_173
timestamp 1623621585
transform 1 0 17020 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_180
timestamp 1623621585
transform 1 0 17664 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _1462_
timestamp 1623621585
transform 1 0 19964 0 1 46240
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1623621585
transform 1 0 19504 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_192
timestamp 1623621585
transform 1 0 18768 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_201
timestamp 1623621585
transform 1 0 19596 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1463_
timestamp 1623621585
transform 1 0 20792 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_210
timestamp 1623621585
transform 1 0 20424 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_217
timestamp 1623621585
transform 1 0 21068 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _1477_
timestamp 1623621585
transform 1 0 23920 0 1 46240
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2090_
timestamp 1623621585
transform 1 0 22724 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_81_229
timestamp 1623621585
transform 1 0 22172 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_244
timestamp 1623621585
transform 1 0 23552 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1623621585
transform 1 0 24748 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1623621585
transform 1 0 25760 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_253
timestamp 1623621585
transform 1 0 24380 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_258
timestamp 1623621585
transform 1 0 24840 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_266
timestamp 1623621585
transform 1 0 25576 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_271
timestamp 1623621585
transform 1 0 26036 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1805_
timestamp 1623621585
transform 1 0 26404 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1918_
timestamp 1623621585
transform 1 0 27784 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1920_
timestamp 1623621585
transform 1 0 27048 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_278
timestamp 1623621585
transform 1 0 26680 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_286
timestamp 1623621585
transform 1 0 27416 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_294
timestamp 1623621585
transform 1 0 28152 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1623621585
transform -1 0 28888 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_81_298
timestamp 1623621585
transform 1 0 28520 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1623621585
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output279
timestamp 1623621585
transform 1 0 2484 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output280
timestamp 1623621585
transform 1 0 1748 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 1623621585
transform 1 0 1380 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_11
timestamp 1623621585
transform 1 0 2116 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_19
timestamp 1623621585
transform 1 0 2852 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output283
timestamp 1623621585
transform 1 0 3220 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output285
timestamp 1623621585
transform 1 0 3956 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output286
timestamp 1623621585
transform 1 0 4692 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_27
timestamp 1623621585
transform 1 0 3588 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1623621585
transform 1 0 4324 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_43
timestamp 1623621585
transform 1 0 5060 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1393_
timestamp 1623621585
transform 1 0 5520 0 -1 47328
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _1399_
timestamp 1623621585
transform 1 0 6808 0 -1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1623621585
transform 1 0 6348 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_47
timestamp 1623621585
transform 1 0 5428 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_53
timestamp 1623621585
transform 1 0 5980 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_58
timestamp 1623621585
transform 1 0 6440 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1384_
timestamp 1623621585
transform 1 0 8372 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2057_
timestamp 1623621585
transform 1 0 9016 0 -1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_82_71
timestamp 1623621585
transform 1 0 7636 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_82
timestamp 1623621585
transform 1 0 8648 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1387_
timestamp 1623621585
transform 1 0 10212 0 -1 47328
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1623621585
transform 1 0 11592 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_95
timestamp 1623621585
transform 1 0 9844 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_104
timestamp 1623621585
transform 1 0 10672 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_112
timestamp 1623621585
transform 1 0 11408 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  _1031_
timestamp 1623621585
transform 1 0 12512 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1743_
timestamp 1623621585
transform 1 0 13616 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_115
timestamp 1623621585
transform 1 0 11684 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_123
timestamp 1623621585
transform 1 0 12420 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_128
timestamp 1623621585
transform 1 0 12880 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2180_
timestamp 1623621585
transform 1 0 14352 0 -1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_82_139
timestamp 1623621585
transform 1 0 13892 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_143
timestamp 1623621585
transform 1 0 14260 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__o31ai_1  _1510_
timestamp 1623621585
transform 1 0 17848 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1623621585
transform 1 0 16836 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_160
timestamp 1623621585
transform 1 0 15824 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_168
timestamp 1623621585
transform 1 0 16560 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_172
timestamp 1623621585
transform 1 0 16928 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_180
timestamp 1623621585
transform 1 0 17664 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _1461_
timestamp 1623621585
transform 1 0 19136 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 19780 0 -1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_82_188
timestamp 1623621585
transform 1 0 18400 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_199
timestamp 1623621585
transform 1 0 19412 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1466_
timestamp 1623621585
transform 1 0 20792 0 -1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1623621585
transform 1 0 22080 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_210
timestamp 1623621585
transform 1 0 20424 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_221
timestamp 1623621585
transform 1 0 21436 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_227
timestamp 1623621585
transform 1 0 21988 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1478_
timestamp 1623621585
transform 1 0 24196 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1670_
timestamp 1623621585
transform 1 0 22908 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_229
timestamp 1623621585
transform 1 0 22172 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_240
timestamp 1623621585
transform 1 0 23184 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_248
timestamp 1623621585
transform 1 0 23920 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1504_
timestamp 1623621585
transform 1 0 25392 0 -1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_82_254
timestamp 1623621585
transform 1 0 24472 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_262
timestamp 1623621585
transform 1 0 25208 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_273
timestamp 1623621585
transform 1 0 26220 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1919_
timestamp 1623621585
transform 1 0 27784 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1921_
timestamp 1623621585
transform 1 0 26588 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1623621585
transform 1 0 27324 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_281
timestamp 1623621585
transform 1 0 26956 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_286
timestamp 1623621585
transform 1 0 27416 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_294
timestamp 1623621585
transform 1 0 28152 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1623621585
transform -1 0 28888 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_82_298
timestamp 1623621585
transform 1 0 28520 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1363_
timestamp 1623621585
transform 1 0 2576 0 1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1623621585
transform 1 0 1104 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output281
timestamp 1623621585
transform 1 0 1748 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_3
timestamp 1623621585
transform 1 0 1380 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_11
timestamp 1623621585
transform 1 0 2116 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_15
timestamp 1623621585
transform 1 0 2484 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__a211oi_4  _1398_
timestamp 1623621585
transform 1 0 5244 0 1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1773_
timestamp 1623621585
transform 1 0 4508 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1623621585
transform 1 0 3772 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_25
timestamp 1623621585
transform 1 0 3404 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_30
timestamp 1623621585
transform 1 0 3864 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_36
timestamp 1623621585
transform 1 0 4416 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_40
timestamp 1623621585
transform 1 0 4784 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_44
timestamp 1623621585
transform 1 0 5152 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1392_
timestamp 1623621585
transform 1 0 7084 0 1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_83_61
timestamp 1623621585
transform 1 0 6716 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1386_
timestamp 1623621585
transform 1 0 9476 0 1 47328
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1707_
timestamp 1623621585
transform 1 0 8280 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1623621585
transform 1 0 9016 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_74
timestamp 1623621585
transform 1 0 7912 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_82
timestamp 1623621585
transform 1 0 8648 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_87
timestamp 1623621585
transform 1 0 9108 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1385_
timestamp 1623621585
transform 1 0 10304 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1731_
timestamp 1623621585
transform 1 0 10948 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_96
timestamp 1623621585
transform 1 0 9936 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_103
timestamp 1623621585
transform 1 0 10580 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_110
timestamp 1623621585
transform 1 0 11224 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_122
timestamp 1623621585
transform 1 0 12328 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_134
timestamp 1623621585
transform 1 0 13432 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2164_
timestamp 1623621585
transform 1 0 15640 0 1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1623621585
transform 1 0 14260 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_83_142
timestamp 1623621585
transform 1 0 14168 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_144
timestamp 1623621585
transform 1 0 14352 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_156
timestamp 1623621585
transform 1 0 15456 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_83_174
timestamp 1623621585
transform 1 0 17112 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_182
timestamp 1623621585
transform 1 0 17848 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__o21bai_2  _1458_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 18032 0 1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1465_
timestamp 1623621585
transform 1 0 19964 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1623621585
transform 1 0 19504 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_193
timestamp 1623621585
transform 1 0 18860 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_199
timestamp 1623621585
transform 1 0 19412 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_201
timestamp 1623621585
transform 1 0 19596 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1503_
timestamp 1623621585
transform 1 0 21160 0 1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_83_209
timestamp 1623621585
transform 1 0 20332 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_217
timestamp 1623621585
transform 1 0 21068 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_225
timestamp 1623621585
transform 1 0 21804 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1801_
timestamp 1623621585
transform 1 0 24104 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_237
timestamp 1623621585
transform 1 0 22908 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_249
timestamp 1623621585
transform 1 0 24012 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2191_
timestamp 1623621585
transform 1 0 25576 0 1 47328
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1623621585
transform 1 0 24748 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_253
timestamp 1623621585
transform 1 0 24380 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_258
timestamp 1623621585
transform 1 0 24840 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1922_
timestamp 1623621585
transform 1 0 27692 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_285
timestamp 1623621585
transform 1 0 27324 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_293
timestamp 1623621585
transform 1 0 28060 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1623621585
transform -1 0 28888 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2219_
timestamp 1623621585
transform 1 0 2944 0 -1 48416
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1623621585
transform 1 0 1104 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output284
timestamp 1623621585
transform 1 0 1748 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_3
timestamp 1623621585
transform 1 0 1380 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_11
timestamp 1623621585
transform 1 0 2116 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_19
timestamp 1623621585
transform 1 0 2852 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1520_
timestamp 1623621585
transform 1 0 4784 0 -1 48416
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_84_36
timestamp 1623621585
transform 1 0 4416 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1394_
timestamp 1623621585
transform 1 0 6808 0 -1 48416
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1623621585
transform 1 0 6348 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_49
timestamp 1623621585
transform 1 0 5612 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_58
timestamp 1623621585
transform 1 0 6440 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2062_
timestamp 1623621585
transform 1 0 8004 0 -1 48416
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_84_71
timestamp 1623621585
transform 1 0 7636 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_84
timestamp 1623621585
transform 1 0 8832 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1389_
timestamp 1623621585
transform 1 0 9752 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1427_
timestamp 1623621585
transform 1 0 10856 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1623621585
transform 1 0 11592 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_92
timestamp 1623621585
transform 1 0 9568 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_84_98
timestamp 1623621585
transform 1 0 10120 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_110
timestamp 1623621585
transform 1 0 11224 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_115
timestamp 1623621585
transform 1 0 11684 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_127
timestamp 1623621585
transform 1 0 12788 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_139
timestamp 1623621585
transform 1 0 13892 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_151
timestamp 1623621585
transform 1 0 14996 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1457_
timestamp 1623621585
transform 1 0 17296 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1623621585
transform 1 0 16836 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_163
timestamp 1623621585
transform 1 0 16100 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_172
timestamp 1623621585
transform 1 0 16928 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_179
timestamp 1623621585
transform 1 0 17572 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1508_
timestamp 1623621585
transform 1 0 17940 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _1511_
timestamp 1623621585
transform 1 0 18860 0 -1 48416
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_84_189
timestamp 1623621585
transform 1 0 18492 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_198
timestamp 1623621585
transform 1 0 19320 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1501_
timestamp 1623621585
transform 1 0 20056 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1502_
timestamp 1623621585
transform 1 0 20700 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1623621585
transform 1 0 22080 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_209
timestamp 1623621585
transform 1 0 20332 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_217
timestamp 1623621585
transform 1 0 21068 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_225
timestamp 1623621585
transform 1 0 21804 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1480_
timestamp 1623621585
transform 1 0 23000 0 -1 48416
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _1802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 24012 0 -1 48416
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_84_229
timestamp 1623621585
transform 1 0 22172 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_237
timestamp 1623621585
transform 1 0 22908 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_243
timestamp 1623621585
transform 1 0 23460 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1623621585
transform 1 0 26036 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1623621585
transform 1 0 25392 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_84_256
timestamp 1623621585
transform 1 0 24656 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_267
timestamp 1623621585
transform 1 0 25668 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_274
timestamp 1623621585
transform 1 0 26312 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1923_
timestamp 1623621585
transform 1 0 27876 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1623621585
transform 1 0 27324 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1623621585
transform 1 0 26680 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_281
timestamp 1623621585
transform 1 0 26956 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_286
timestamp 1623621585
transform 1 0 27416 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_290
timestamp 1623621585
transform 1 0 27784 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_295
timestamp 1623621585
transform 1 0 28244 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1623621585
transform -1 0 28888 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_86_11
timestamp 1623621585
transform 1 0 2116 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_3
timestamp 1623621585
transform 1 0 1380 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_7
timestamp 1623621585
transform 1 0 1748 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_3
timestamp 1623621585
transform 1 0 1380 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output288
timestamp 1623621585
transform 1 0 1748 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1623621585
transform 1 0 1104 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1623621585
transform 1 0 1104 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_86_19
timestamp 1623621585
transform 1 0 2852 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output287
timestamp 1623621585
transform 1 0 2484 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2218_
timestamp 1623621585
transform 1 0 1840 0 1 48416
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _1361_
timestamp 1623621585
transform 1 0 4232 0 1 48416
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2185_
timestamp 1623621585
transform 1 0 3864 0 -1 49504
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1623621585
transform 1 0 3772 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_24
timestamp 1623621585
transform 1 0 3312 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_28
timestamp 1623621585
transform 1 0 3680 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_30
timestamp 1623621585
transform 1 0 3864 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_43
timestamp 1623621585
transform 1 0 5060 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_86_27
timestamp 1623621585
transform 1 0 3588 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_86_53
timestamp 1623621585
transform 1 0 5980 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_46
timestamp 1623621585
transform 1 0 5336 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1623621585
transform 1 0 5796 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_47
timestamp 1623621585
transform 1 0 5428 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1623621585
transform 1 0 6348 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _2063_
timestamp 1623621585
transform 1 0 6164 0 1 48416
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1723_
timestamp 1623621585
transform 1 0 5704 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1719_
timestamp 1623621585
transform 1 0 5520 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_85_64
timestamp 1623621585
transform 1 0 6992 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_58
timestamp 1623621585
transform 1 0 6440 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1522_
timestamp 1623621585
transform 1 0 7820 0 1 48416
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2183_
timestamp 1623621585
transform 1 0 7636 0 -1 49504
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1623621585
transform 1 0 9016 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_72
timestamp 1623621585
transform 1 0 7728 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_82
timestamp 1623621585
transform 1 0 8648 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_87
timestamp 1623621585
transform 1 0 9108 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_70
timestamp 1623621585
transform 1 0 7544 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_87
timestamp 1623621585
transform 1 0 9108 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_95
timestamp 1623621585
transform 1 0 9844 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_101
timestamp 1623621585
transform 1 0 10396 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_93
timestamp 1623621585
transform 1 0 9660 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_2  _1390_
timestamp 1623621585
transform 1 0 9752 0 1 48416
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1388_
timestamp 1623621585
transform 1 0 9936 0 -1 49504
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_86_110
timestamp 1623621585
transform 1 0 11224 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_103
timestamp 1623621585
transform 1 0 10580 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1623621585
transform 1 0 11592 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1426_
timestamp 1623621585
transform 1 0 10948 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1383_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 10764 0 1 48416
box -38 -48 1234 592
use sky130_fd_sc_hd__o21bai_2  _1382_
timestamp 1623621585
transform 1 0 12880 0 1 48416
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1430_
timestamp 1623621585
transform 1 0 12052 0 -1 49504
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1433_
timestamp 1623621585
transform 1 0 13340 0 -1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_85_118
timestamp 1623621585
transform 1 0 11960 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_126
timestamp 1623621585
transform 1 0 12696 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_85_137
timestamp 1623621585
transform 1 0 13708 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_115
timestamp 1623621585
transform 1 0 11684 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_126
timestamp 1623621585
transform 1 0 12696 0 -1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_132
timestamp 1623621585
transform 1 0 13248 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__o31ai_1  _1434_
timestamp 1623621585
transform 1 0 14260 0 -1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _1435_
timestamp 1623621585
transform 1 0 14720 0 1 48416
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1623621585
transform 1 0 14260 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_144
timestamp 1623621585
transform 1 0 14352 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_153
timestamp 1623621585
transform 1 0 15180 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_139
timestamp 1623621585
transform 1 0 13892 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_149
timestamp 1623621585
transform 1 0 14812 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_165
timestamp 1623621585
transform 1 0 16284 0 -1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_161
timestamp 1623621585
transform 1 0 15916 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_165
timestamp 1623621585
transform 1 0 16284 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1623621585
transform 1 0 16836 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1432_
timestamp 1623621585
transform 1 0 16008 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_86_172
timestamp 1623621585
transform 1 0 16928 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_85_173
timestamp 1623621585
transform 1 0 17020 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1452_
timestamp 1623621585
transform 1 0 17296 0 1 48416
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1013_
timestamp 1623621585
transform 1 0 17296 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_180
timestamp 1623621585
transform 1 0 17664 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_181
timestamp 1623621585
transform 1 0 17756 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__xor2_4  _1459_
timestamp 1623621585
transform 1 0 19596 0 -1 49504
box -38 -48 2062 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1623621585
transform 1 0 19504 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_85_193
timestamp 1623621585
transform 1 0 18860 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_199
timestamp 1623621585
transform 1 0 19412 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_201
timestamp 1623621585
transform 1 0 19596 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_192
timestamp 1623621585
transform 1 0 18768 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_200
timestamp 1623621585
transform 1 0 19504 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _1505_
timestamp 1623621585
transform 1 0 21160 0 1 48416
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1623621585
transform 1 0 22080 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_213
timestamp 1623621585
transform 1 0 20700 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_217
timestamp 1623621585
transform 1 0 21068 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_225
timestamp 1623621585
transform 1 0 21804 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_223
timestamp 1623621585
transform 1 0 21620 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_227
timestamp 1623621585
transform 1 0 21988 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_233
timestamp 1623621585
transform 1 0 22540 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_229
timestamp 1623621585
transform 1 0 22172 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_234
timestamp 1623621585
transform 1 0 22632 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_229
timestamp 1623621585
transform 1 0 22172 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _2093_
timestamp 1623621585
transform 1 0 22632 0 -1 49504
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1663_
timestamp 1623621585
transform 1 0 22264 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1479_
timestamp 1623621585
transform 1 0 23000 0 1 48416
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_86_243
timestamp 1623621585
transform 1 0 23460 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_85_243
timestamp 1623621585
transform 1 0 23460 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1482_
timestamp 1623621585
transform 1 0 23828 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1483_
timestamp 1623621585
transform 1 0 24196 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _1486_
timestamp 1623621585
transform 1 0 25208 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1506_
timestamp 1623621585
transform 1 0 25392 0 -1 49504
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1623621585
transform 1 0 24748 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_253
timestamp 1623621585
transform 1 0 24380 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_258
timestamp 1623621585
transform 1 0 24840 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_268
timestamp 1623621585
transform 1 0 25760 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_86_259
timestamp 1623621585
transform 1 0 24932 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_263
timestamp 1623621585
transform 1 0 25300 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_273
timestamp 1623621585
transform 1 0 26220 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_277
timestamp 1623621585
transform 1 0 26588 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1623621585
transform 1 0 26680 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1623621585
transform 1 0 26496 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_86_281
timestamp 1623621585
transform 1 0 26956 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_279
timestamp 1623621585
transform 1 0 26772 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1926_
timestamp 1623621585
transform 1 0 27140 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_286
timestamp 1623621585
transform 1 0 27416 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_287
timestamp 1623621585
transform 1 0 27508 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1623621585
transform 1 0 27324 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1925_
timestamp 1623621585
transform 1 0 27784 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1924_
timestamp 1623621585
transform 1 0 27876 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_294
timestamp 1623621585
transform 1 0 28152 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_295
timestamp 1623621585
transform 1 0 28244 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1623621585
transform -1 0 28888 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1623621585
transform -1 0 28888 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_86_298
timestamp 1623621585
transform 1 0 28520 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1623621585
transform 1 0 1104 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output289
timestamp 1623621585
transform 1 0 1748 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output290
timestamp 1623621585
transform 1 0 2484 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_3
timestamp 1623621585
transform 1 0 1380 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_11
timestamp 1623621585
transform 1 0 2116 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_19
timestamp 1623621585
transform 1 0 2852 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1623621585
transform 1 0 3772 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_27
timestamp 1623621585
transform 1 0 3588 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_30
timestamp 1623621585
transform 1 0 3864 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_42
timestamp 1623621585
transform 1 0 4968 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_54
timestamp 1623621585
transform 1 0 6072 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_66
timestamp 1623621585
transform 1 0 7176 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1718_
timestamp 1623621585
transform 1 0 7820 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1623621585
transform 1 0 9016 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_72
timestamp 1623621585
transform 1 0 7728 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_76
timestamp 1623621585
transform 1 0 8096 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_84
timestamp 1623621585
transform 1 0 8832 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_87
timestamp 1623621585
transform 1 0 9108 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_99
timestamp 1623621585
transform 1 0 10212 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_111
timestamp 1623621585
transform 1 0 11316 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1376_
timestamp 1623621585
transform 1 0 13432 0 1 49504
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1381_
timestamp 1623621585
transform 1 0 12788 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1735_
timestamp 1623621585
transform 1 0 11868 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_87_120
timestamp 1623621585
transform 1 0 12144 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_126
timestamp 1623621585
transform 1 0 12696 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_130
timestamp 1623621585
transform 1 0 13064 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2205_
timestamp 1623621585
transform 1 0 15088 0 1 49504
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1623621585
transform 1 0 14260 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_139
timestamp 1623621585
transform 1 0 13892 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_144
timestamp 1623621585
transform 1 0 14352 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2075_
timestamp 1623621585
transform 1 0 17204 0 1 49504
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_87_171
timestamp 1623621585
transform 1 0 16836 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1691_
timestamp 1623621585
transform 1 0 18400 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1692_
timestamp 1623621585
transform 1 0 19964 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1623621585
transform 1 0 19504 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_184
timestamp 1623621585
transform 1 0 18032 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_191
timestamp 1623621585
transform 1 0 18676 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_199
timestamp 1623621585
transform 1 0 19412 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_201
timestamp 1623621585
transform 1 0 19596 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1685_
timestamp 1623621585
transform 1 0 21068 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1686_
timestamp 1623621585
transform 1 0 21712 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_87_208
timestamp 1623621585
transform 1 0 20240 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_216
timestamp 1623621585
transform 1 0 20976 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_220
timestamp 1623621585
transform 1 0 21344 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_227
timestamp 1623621585
transform 1 0 21988 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1481_
timestamp 1623621585
transform 1 0 23920 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1664_
timestamp 1623621585
transform 1 0 22540 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_236
timestamp 1623621585
transform 1 0 22816 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_251
timestamp 1623621585
transform 1 0 24196 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2190_
timestamp 1623621585
transform 1 0 25484 0 1 49504
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1623621585
transform 1 0 24748 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_258
timestamp 1623621585
transform 1 0 24840 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_264
timestamp 1623621585
transform 1 0 25392 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1927_
timestamp 1623621585
transform 1 0 27784 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_284
timestamp 1623621585
transform 1 0 27232 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_87_294
timestamp 1623621585
transform 1 0 28152 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1623621585
transform -1 0 28888 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_87_298
timestamp 1623621585
transform 1 0 28520 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1623621585
transform 1 0 1104 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output291
timestamp 1623621585
transform 1 0 1748 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output292
timestamp 1623621585
transform 1 0 2484 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_3
timestamp 1623621585
transform 1 0 1380 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_11
timestamp 1623621585
transform 1 0 2116 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_19
timestamp 1623621585
transform 1 0 2852 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output306
timestamp 1623621585
transform 1 0 3220 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_27
timestamp 1623621585
transform 1 0 3588 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_39
timestamp 1623621585
transform 1 0 4692 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _1395_
timestamp 1623621585
transform 1 0 6992 0 -1 50592
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_1  _1418_
timestamp 1623621585
transform 1 0 5520 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1623621585
transform 1 0 6348 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_47
timestamp 1623621585
transform 1 0 5428 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_51
timestamp 1623621585
transform 1 0 5796 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_88_58
timestamp 1623621585
transform 1 0 6440 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _1423_
timestamp 1623621585
transform 1 0 9200 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_88_78
timestamp 1623621585
transform 1 0 8280 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_86
timestamp 1623621585
transform 1 0 9016 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1623621585
transform 1 0 11592 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_94
timestamp 1623621585
transform 1 0 9752 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_106
timestamp 1623621585
transform 1 0 10856 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _2054_
timestamp 1623621585
transform 1 0 12052 0 -1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_88_115
timestamp 1623621585
transform 1 0 11684 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_128
timestamp 1623621585
transform 1 0 12880 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_136
timestamp 1623621585
transform 1 0 13616 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _2051_
timestamp 1623621585
transform 1 0 13800 0 -1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_88_147
timestamp 1623621585
transform 1 0 14628 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_159
timestamp 1623621585
transform 1 0 15732 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1696_
timestamp 1623621585
transform 1 0 16192 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2074_
timestamp 1623621585
transform 1 0 17848 0 -1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1623621585
transform 1 0 16836 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_163
timestamp 1623621585
transform 1 0 16100 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_167
timestamp 1623621585
transform 1 0 16468 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_172
timestamp 1623621585
transform 1 0 16928 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_180
timestamp 1623621585
transform 1 0 17664 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_4  _2078_
timestamp 1623621585
transform 1 0 19044 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_191
timestamp 1623621585
transform 1 0 18676 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _2081_
timestamp 1623621585
transform 1 0 20700 0 -1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1623621585
transform 1 0 22080 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_207
timestamp 1623621585
transform 1 0 20148 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_88_222
timestamp 1623621585
transform 1 0 21528 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1487_
timestamp 1623621585
transform 1 0 23920 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1623621585
transform 1 0 23276 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input157
timestamp 1623621585
transform 1 0 22632 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_229
timestamp 1623621585
transform 1 0 22172 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_233
timestamp 1623621585
transform 1 0 22540 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_237
timestamp 1623621585
transform 1 0 22908 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_244
timestamp 1623621585
transform 1 0 23552 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1623621585
transform 1 0 26036 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1623621585
transform 1 0 25392 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1623621585
transform 1 0 24748 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_252
timestamp 1623621585
transform 1 0 24288 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_256
timestamp 1623621585
transform 1 0 24656 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_260
timestamp 1623621585
transform 1 0 25024 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_267
timestamp 1623621585
transform 1 0 25668 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_274
timestamp 1623621585
transform 1 0 26312 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1928_
timestamp 1623621585
transform 1 0 27876 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1623621585
transform 1 0 27324 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1623621585
transform 1 0 26680 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_281
timestamp 1623621585
transform 1 0 26956 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_286
timestamp 1623621585
transform 1 0 27416 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_290
timestamp 1623621585
transform 1 0 27784 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_295
timestamp 1623621585
transform 1 0 28244 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1623621585
transform -1 0 28888 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1623621585
transform 1 0 1104 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output294
timestamp 1623621585
transform 1 0 1748 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output305
timestamp 1623621585
transform 1 0 2484 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_3
timestamp 1623621585
transform 1 0 1380 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_11
timestamp 1623621585
transform 1 0 2116 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_19
timestamp 1623621585
transform 1 0 2852 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1623621585
transform 1 0 3772 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output307
timestamp 1623621585
transform 1 0 4232 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_27
timestamp 1623621585
transform 1 0 3588 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_30
timestamp 1623621585
transform 1 0 3864 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_38
timestamp 1623621585
transform 1 0 4600 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1420_
timestamp 1623621585
transform 1 0 7084 0 1 50592
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _2060_
timestamp 1623621585
transform 1 0 5520 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_46
timestamp 1623621585
transform 1 0 5336 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_60
timestamp 1623621585
transform 1 0 6624 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_64
timestamp 1623621585
transform 1 0 6992 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_1  _1419_
timestamp 1623621585
transform 1 0 8096 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1623621585
transform 1 0 9016 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_72
timestamp 1623621585
transform 1 0 7728 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_80
timestamp 1623621585
transform 1 0 8464 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_89_87
timestamp 1623621585
transform 1 0 9108 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1422_
timestamp 1623621585
transform 1 0 9752 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_93
timestamp 1623621585
transform 1 0 9660 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_100
timestamp 1623621585
transform 1 0 10304 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_112
timestamp 1623621585
transform 1 0 11408 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1736_
timestamp 1623621585
transform 1 0 12972 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1739_
timestamp 1623621585
transform 1 0 13616 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2053_
timestamp 1623621585
transform 1 0 11776 0 1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_89_125
timestamp 1623621585
transform 1 0 12604 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_132
timestamp 1623621585
transform 1 0 13248 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2050_
timestamp 1623621585
transform 1 0 14812 0 1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1623621585
transform 1 0 14260 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_139
timestamp 1623621585
transform 1 0 13892 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_144
timestamp 1623621585
transform 1 0 14352 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_148
timestamp 1623621585
transform 1 0 14720 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_158
timestamp 1623621585
transform 1 0 15640 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1563_
timestamp 1623621585
transform 1 0 16560 0 1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1697_
timestamp 1623621585
transform 1 0 17756 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_89_166
timestamp 1623621585
transform 1 0 16376 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_177
timestamp 1623621585
transform 1 0 17388 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2077_
timestamp 1623621585
transform 1 0 19964 0 1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1623621585
transform 1 0 19504 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_184
timestamp 1623621585
transform 1 0 18032 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_196
timestamp 1623621585
transform 1 0 19136 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_201
timestamp 1623621585
transform 1 0 19596 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2080_
timestamp 1623621585
transform 1 0 21160 0 1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_89_214
timestamp 1623621585
transform 1 0 20792 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_227
timestamp 1623621585
transform 1 0 21988 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2092_
timestamp 1623621585
transform 1 0 23000 0 1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1623621585
transform 1 0 22356 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_234
timestamp 1623621585
transform 1 0 22632 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_247
timestamp 1623621585
transform 1 0 23828 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1451_
timestamp 1623621585
transform 1 0 25208 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1623621585
transform 1 0 24748 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1623621585
transform 1 0 25852 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_89_255
timestamp 1623621585
transform 1 0 24564 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_258
timestamp 1623621585
transform 1 0 24840 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_265
timestamp 1623621585
transform 1 0 25484 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_272
timestamp 1623621585
transform 1 0 26128 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1929_
timestamp 1623621585
transform 1 0 27876 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1930_
timestamp 1623621585
transform 1 0 27140 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1623621585
transform 1 0 26496 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_279
timestamp 1623621585
transform 1 0 26772 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_287
timestamp 1623621585
transform 1 0 27508 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_295
timestamp 1623621585
transform 1 0 28244 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1623621585
transform -1 0 28888 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1623621585
transform 1 0 1104 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output295
timestamp 1623621585
transform 1 0 1748 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output297
timestamp 1623621585
transform 1 0 2484 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_3
timestamp 1623621585
transform 1 0 1380 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_11
timestamp 1623621585
transform 1 0 2116 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_19
timestamp 1623621585
transform 1 0 2852 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1521_
timestamp 1623621585
transform 1 0 4324 0 -1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output301
timestamp 1623621585
transform 1 0 3220 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_27
timestamp 1623621585
transform 1 0 3588 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_90_44
timestamp 1623621585
transform 1 0 5152 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2059_
timestamp 1623621585
transform 1 0 6808 0 -1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1623621585
transform 1 0 6348 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output308
timestamp 1623621585
transform 1 0 5520 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_52
timestamp 1623621585
transform 1 0 5888 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_56
timestamp 1623621585
transform 1 0 6256 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_58
timestamp 1623621585
transform 1 0 6440 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2208_
timestamp 1623621585
transform 1 0 8096 0 -1 51680
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_90_71
timestamp 1623621585
transform 1 0 7636 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_75
timestamp 1623621585
transform 1 0 8004 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1523_
timestamp 1623621585
transform 1 0 10396 0 -1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1623621585
transform 1 0 11592 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_95
timestamp 1623621585
transform 1 0 9844 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_90_110
timestamp 1623621585
transform 1 0 11224 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1431_
timestamp 1623621585
transform 1 0 12420 0 -1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1737_
timestamp 1623621585
transform 1 0 13616 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_90_115
timestamp 1623621585
transform 1 0 11684 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_90_132
timestamp 1623621585
transform 1 0 13248 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2181_
timestamp 1623621585
transform 1 0 14352 0 -1 51680
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_90_139
timestamp 1623621585
transform 1 0 13892 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_143
timestamp 1623621585
transform 1 0 14260 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1740_
timestamp 1623621585
transform 1 0 16192 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1623621585
transform 1 0 16836 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_160
timestamp 1623621585
transform 1 0 15824 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_167
timestamp 1623621585
transform 1 0 16468 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_172
timestamp 1623621585
transform 1 0 16928 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1562_
timestamp 1623621585
transform 1 0 18308 0 -1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1693_
timestamp 1623621585
transform 1 0 19504 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_90_184
timestamp 1623621585
transform 1 0 18032 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_90_196
timestamp 1623621585
transform 1 0 19136 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_203
timestamp 1623621585
transform 1 0 19780 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1561_
timestamp 1623621585
transform 1 0 20424 0 -1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1623621585
transform 1 0 22080 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_90_209
timestamp 1623621585
transform 1 0 20332 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_219
timestamp 1623621585
transform 1 0 21252 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_227
timestamp 1623621585
transform 1 0 21988 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1557_
timestamp 1623621585
transform 1 0 22540 0 -1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _2195_
timestamp 1623621585
transform 1 0 24104 0 -1 51680
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_90_229
timestamp 1623621585
transform 1 0 22172 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_242
timestamp 1623621585
transform 1 0 23368 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_90_267
timestamp 1623621585
transform 1 0 25668 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1931_
timestamp 1623621585
transform 1 0 27876 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1938_
timestamp 1623621585
transform 1 0 26588 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1623621585
transform 1 0 27324 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_275
timestamp 1623621585
transform 1 0 26404 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_281
timestamp 1623621585
transform 1 0 26956 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_286
timestamp 1623621585
transform 1 0 27416 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_290
timestamp 1623621585
transform 1 0 27784 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_295
timestamp 1623621585
transform 1 0 28244 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1623621585
transform -1 0 28888 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1623621585
transform 1 0 1104 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output296
timestamp 1623621585
transform 1 0 1748 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output299
timestamp 1623621585
transform 1 0 2484 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_3
timestamp 1623621585
transform 1 0 1380 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_11
timestamp 1623621585
transform 1 0 2116 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_91_19
timestamp 1623621585
transform 1 0 2852 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _1391_
timestamp 1623621585
transform 1 0 5060 0 1 51680
box -38 -48 2062 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1623621585
transform 1 0 3772 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output302
timestamp 1623621585
transform 1 0 4232 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_27
timestamp 1623621585
transform 1 0 3588 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_30
timestamp 1623621585
transform 1 0 3864 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_38
timestamp 1623621585
transform 1 0 4600 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_42
timestamp 1623621585
transform 1 0 4968 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_65
timestamp 1623621585
transform 1 0 7084 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1425_
timestamp 1623621585
transform 1 0 7820 0 1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _2209_
timestamp 1623621585
transform 1 0 9476 0 1 51680
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1623621585
transform 1 0 9016 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_82
timestamp 1623621585
transform 1 0 8648 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_87
timestamp 1623621585
transform 1 0 9108 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2182_
timestamp 1623621585
transform 1 0 11592 0 1 51680
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_91_110
timestamp 1623621585
transform 1 0 11224 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_130
timestamp 1623621585
transform 1 0 13064 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1524_
timestamp 1623621585
transform 1 0 14720 0 1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1623621585
transform 1 0 14260 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_91_142
timestamp 1623621585
transform 1 0 14168 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_144
timestamp 1623621585
transform 1 0 14352 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_91_157
timestamp 1623621585
transform 1 0 15548 0 1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2165_
timestamp 1623621585
transform 1 0 16100 0 1 51680
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_91_179
timestamp 1623621585
transform 1 0 17572 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2167_
timestamp 1623621585
transform 1 0 19964 0 1 51680
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1623621585
transform 1 0 19504 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_191
timestamp 1623621585
transform 1 0 18676 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_199
timestamp 1623621585
transform 1 0 19412 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_201
timestamp 1623621585
transform 1 0 19596 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2171_
timestamp 1623621585
transform 1 0 21804 0 1 51680
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_91_221
timestamp 1623621585
transform 1 0 21436 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1665_
timestamp 1623621585
transform 1 0 23644 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_241
timestamp 1623621585
transform 1 0 23276 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_91_248
timestamp 1623621585
transform 1 0 23920 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1939_
timestamp 1623621585
transform 1 0 25668 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1623621585
transform 1 0 24748 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_91_256
timestamp 1623621585
transform 1 0 24656 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_258
timestamp 1623621585
transform 1 0 24840 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_266
timestamp 1623621585
transform 1 0 25576 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_271
timestamp 1623621585
transform 1 0 26036 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1932_
timestamp 1623621585
transform 1 0 27876 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1933_
timestamp 1623621585
transform 1 0 27140 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1934_
timestamp 1623621585
transform 1 0 26404 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_279
timestamp 1623621585
transform 1 0 26772 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_287
timestamp 1623621585
transform 1 0 27508 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_295
timestamp 1623621585
transform 1 0 28244 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1623621585
transform -1 0 28888 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_3
timestamp 1623621585
transform 1 0 1380 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_3
timestamp 1623621585
transform 1 0 1380 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output298
timestamp 1623621585
transform 1 0 1748 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input159
timestamp 1623621585
transform 1 0 1748 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1623621585
transform 1 0 1104 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1623621585
transform 1 0 1104 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_13
timestamp 1623621585
transform 1 0 2300 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_11
timestamp 1623621585
transform 1 0 2116 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output300
timestamp 1623621585
transform 1 0 2484 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output160
timestamp 1623621585
transform 1 0 2668 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_93_21
timestamp 1623621585
transform 1 0 3036 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_92_19
timestamp 1623621585
transform 1 0 2852 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2184_
timestamp 1623621585
transform 1 0 3772 0 -1 52768
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1623621585
transform 1 0 3772 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output167
timestamp 1623621585
transform 1 0 4232 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output168
timestamp 1623621585
transform 1 0 4968 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_27
timestamp 1623621585
transform 1 0 3588 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_45
timestamp 1623621585
transform 1 0 5244 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_30
timestamp 1623621585
transform 1 0 3864 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_38
timestamp 1623621585
transform 1 0 4600 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_54
timestamp 1623621585
transform 1 0 6072 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_46
timestamp 1623621585
transform 1 0 5336 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_52
timestamp 1623621585
transform 1 0 5888 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output303
timestamp 1623621585
transform 1 0 5704 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1725_
timestamp 1623621585
transform 1 0 5612 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_59
timestamp 1623621585
transform 1 0 6532 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_58
timestamp 1623621585
transform 1 0 6440 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_56
timestamp 1623621585
transform 1 0 6256 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output169
timestamp 1623621585
transform 1 0 6900 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1623621585
transform 1 0 6440 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1623621585
transform 1 0 6348 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_93_67
timestamp 1623621585
transform 1 0 7268 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1424_
timestamp 1623621585
transform 1 0 7176 0 -1 52768
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1724_
timestamp 1623621585
transform 1 0 8188 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1623621585
transform 1 0 9108 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output170
timestamp 1623621585
transform 1 0 7820 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_73
timestamp 1623621585
transform 1 0 7820 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_80
timestamp 1623621585
transform 1 0 8464 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_77
timestamp 1623621585
transform 1 0 8188 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_85
timestamp 1623621585
transform 1 0 8924 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_88
timestamp 1623621585
transform 1 0 9200 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1623621585
transform 1 0 11592 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output171
timestamp 1623621585
transform 1 0 9568 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_92
timestamp 1623621585
transform 1 0 9568 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_104
timestamp 1623621585
transform 1 0 10672 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_112
timestamp 1623621585
transform 1 0 11408 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_96
timestamp 1623621585
transform 1 0 9936 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_108
timestamp 1623621585
transform 1 0 11040 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2206_
timestamp 1623621585
transform 1 0 12512 0 -1 52768
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1623621585
transform 1 0 11776 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output172
timestamp 1623621585
transform 1 0 12236 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output173
timestamp 1623621585
transform 1 0 13156 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_115
timestamp 1623621585
transform 1 0 11684 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_123
timestamp 1623621585
transform 1 0 12420 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_117
timestamp 1623621585
transform 1 0 11868 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_93_125
timestamp 1623621585
transform 1 0 12604 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_93_135
timestamp 1623621585
transform 1 0 13524 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1623621585
transform 1 0 14444 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output174
timestamp 1623621585
transform 1 0 14904 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_143
timestamp 1623621585
transform 1 0 14260 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_155
timestamp 1623621585
transform 1 0 15364 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_143
timestamp 1623621585
transform 1 0 14260 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_146
timestamp 1623621585
transform 1 0 14536 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_154
timestamp 1623621585
transform 1 0 15272 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1623621585
transform 1 0 16836 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1623621585
transform 1 0 17112 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output175
timestamp 1623621585
transform 1 0 16376 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_167
timestamp 1623621585
transform 1 0 16468 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_172
timestamp 1623621585
transform 1 0 16928 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_180
timestamp 1623621585
transform 1 0 17664 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_170
timestamp 1623621585
transform 1 0 16744 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_175
timestamp 1623621585
transform 1 0 17204 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_192
timestamp 1623621585
transform 1 0 18768 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_187
timestamp 1623621585
transform 1 0 18308 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output161
timestamp 1623621585
transform 1 0 18400 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_204
timestamp 1623621585
transform 1 0 19872 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_199
timestamp 1623621585
transform 1 0 19412 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_205
timestamp 1623621585
transform 1 0 19964 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_199
timestamp 1623621585
transform 1 0 19412 0 -1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1623621585
transform 1 0 19136 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1623621585
transform 1 0 19780 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2166_
timestamp 1623621585
transform 1 0 17940 0 -1 52768
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_92_209
timestamp 1623621585
transform 1 0 20332 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output162
timestamp 1623621585
transform 1 0 20240 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1623621585
transform 1 0 20056 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_212
timestamp 1623621585
transform 1 0 20608 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1623621585
transform 1 0 20700 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_220
timestamp 1623621585
transform 1 0 21344 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_216
timestamp 1623621585
transform 1 0 20976 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output166
timestamp 1623621585
transform 1 0 20976 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1687_
timestamp 1623621585
transform 1 0 21344 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_223
timestamp 1623621585
transform 1 0 21620 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output163
timestamp 1623621585
transform 1 0 21712 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_228
timestamp 1623621585
transform 1 0 22080 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_227
timestamp 1623621585
transform 1 0 21988 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1623621585
transform 1 0 22080 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_233
timestamp 1623621585
transform 1 0 22540 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_233
timestamp 1623621585
transform 1 0 22540 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_229
timestamp 1623621585
transform 1 0 22172 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1623621585
transform 1 0 22448 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_93_237
timestamp 1623621585
transform 1 0 22908 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_237
timestamp 1623621585
transform 1 0 22908 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output165
timestamp 1623621585
transform 1 0 23000 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1623621585
transform 1 0 22632 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_242
timestamp 1623621585
transform 1 0 23368 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1623621585
transform 1 0 23276 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_244
timestamp 1623621585
transform 1 0 23552 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output164
timestamp 1623621585
transform 1 0 23736 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_250
timestamp 1623621585
transform 1 0 24104 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_251
timestamp 1623621585
transform 1 0 24196 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1623621585
transform 1 0 23920 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1623621585
transform 1 0 24472 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1623621585
transform 1 0 24564 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_257
timestamp 1623621585
transform 1 0 24748 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_258
timestamp 1623621585
transform 1 0 24840 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_262
timestamp 1623621585
transform 1 0 25208 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_265
timestamp 1623621585
transform 1 0 25484 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1623621585
transform 1 0 25208 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1623621585
transform 1 0 25116 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_269
timestamp 1623621585
transform 1 0 25852 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1623621585
transform 1 0 25576 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1940_
timestamp 1623621585
transform 1 0 25852 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_273
timestamp 1623621585
transform 1 0 26220 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1941_
timestamp 1623621585
transform 1 0 26220 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_277
timestamp 1623621585
transform 1 0 26588 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_281
timestamp 1623621585
transform 1 0 26956 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1937_
timestamp 1623621585
transform 1 0 26956 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1936_
timestamp 1623621585
transform 1 0 26588 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_93_291
timestamp 1623621585
transform 1 0 27876 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_289
timestamp 1623621585
transform 1 0 27692 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_285
timestamp 1623621585
transform 1 0 27324 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_286
timestamp 1623621585
transform 1 0 27416 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1623621585
transform 1 0 27784 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1623621585
transform 1 0 27324 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1935_
timestamp 1623621585
transform 1 0 27784 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_294
timestamp 1623621585
transform 1 0 28152 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1623621585
transform -1 0 28888 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1623621585
transform -1 0 28888 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_92_298
timestamp 1623621585
transform 1 0 28520 0 -1 52768
box -38 -48 130 592
<< labels >>
rlabel metal2 s 6090 -800 6146 800 8 io_adr_i[0]
port 0 nsew signal input
rlabel metal2 s 7470 -800 7526 800 8 io_adr_i[1]
port 1 nsew signal input
rlabel metal2 s 3330 -800 3386 800 8 io_cs_i
port 2 nsew signal input
rlabel metal2 s 8758 -800 8814 800 8 io_dat_i[0]
port 3 nsew signal input
rlabel metal2 s 22466 -800 22522 800 8 io_dat_i[10]
port 4 nsew signal input
rlabel metal2 s 23754 -800 23810 800 8 io_dat_i[11]
port 5 nsew signal input
rlabel metal2 s 25134 -800 25190 800 8 io_dat_i[12]
port 6 nsew signal input
rlabel metal2 s 26514 -800 26570 800 8 io_dat_i[13]
port 7 nsew signal input
rlabel metal2 s 27894 -800 27950 800 8 io_dat_i[14]
port 8 nsew signal input
rlabel metal2 s 29274 -800 29330 800 8 io_dat_i[15]
port 9 nsew signal input
rlabel metal2 s 10138 -800 10194 800 8 io_dat_i[1]
port 10 nsew signal input
rlabel metal2 s 11518 -800 11574 800 8 io_dat_i[2]
port 11 nsew signal input
rlabel metal2 s 12898 -800 12954 800 8 io_dat_i[3]
port 12 nsew signal input
rlabel metal2 s 14278 -800 14334 800 8 io_dat_i[4]
port 13 nsew signal input
rlabel metal2 s 15658 -800 15714 800 8 io_dat_i[5]
port 14 nsew signal input
rlabel metal2 s 16946 -800 17002 800 8 io_dat_i[6]
port 15 nsew signal input
rlabel metal2 s 18326 -800 18382 800 8 io_dat_i[7]
port 16 nsew signal input
rlabel metal2 s 19706 -800 19762 800 8 io_dat_i[8]
port 17 nsew signal input
rlabel metal2 s 21086 -800 21142 800 8 io_dat_i[9]
port 18 nsew signal input
rlabel metal2 s 846 55200 902 56800 6 io_dat_o[0]
port 19 nsew signal tristate
rlabel metal2 s 18418 55200 18474 56800 6 io_dat_o[10]
port 20 nsew signal tristate
rlabel metal2 s 20166 55200 20222 56800 6 io_dat_o[11]
port 21 nsew signal tristate
rlabel metal2 s 22006 55200 22062 56800 6 io_dat_o[12]
port 22 nsew signal tristate
rlabel metal2 s 23754 55200 23810 56800 6 io_dat_o[13]
port 23 nsew signal tristate
rlabel metal2 s 25502 55200 25558 56800 6 io_dat_o[14]
port 24 nsew signal tristate
rlabel metal2 s 27250 55200 27306 56800 6 io_dat_o[15]
port 25 nsew signal tristate
rlabel metal2 s 2594 55200 2650 56800 6 io_dat_o[1]
port 26 nsew signal tristate
rlabel metal2 s 4342 55200 4398 56800 6 io_dat_o[2]
port 27 nsew signal tristate
rlabel metal2 s 6090 55200 6146 56800 6 io_dat_o[3]
port 28 nsew signal tristate
rlabel metal2 s 7838 55200 7894 56800 6 io_dat_o[4]
port 29 nsew signal tristate
rlabel metal2 s 9586 55200 9642 56800 6 io_dat_o[5]
port 30 nsew signal tristate
rlabel metal2 s 11426 55200 11482 56800 6 io_dat_o[6]
port 31 nsew signal tristate
rlabel metal2 s 13174 55200 13230 56800 6 io_dat_o[7]
port 32 nsew signal tristate
rlabel metal2 s 14922 55200 14978 56800 6 io_dat_o[8]
port 33 nsew signal tristate
rlabel metal2 s 16670 55200 16726 56800 6 io_dat_o[9]
port 34 nsew signal tristate
rlabel metal3 s 29200 29520 30800 29640 6 io_eo[0]
port 35 nsew signal input
rlabel metal3 s 29200 33600 30800 33720 6 io_eo[10]
port 36 nsew signal input
rlabel metal3 s 29200 34008 30800 34128 6 io_eo[11]
port 37 nsew signal input
rlabel metal3 s 29200 34416 30800 34536 6 io_eo[12]
port 38 nsew signal input
rlabel metal3 s 29200 34824 30800 34944 6 io_eo[13]
port 39 nsew signal input
rlabel metal3 s 29200 35232 30800 35352 6 io_eo[14]
port 40 nsew signal input
rlabel metal3 s 29200 35640 30800 35760 6 io_eo[15]
port 41 nsew signal input
rlabel metal3 s 29200 36048 30800 36168 6 io_eo[16]
port 42 nsew signal input
rlabel metal3 s 29200 36456 30800 36576 6 io_eo[17]
port 43 nsew signal input
rlabel metal3 s 29200 36864 30800 36984 6 io_eo[18]
port 44 nsew signal input
rlabel metal3 s 29200 37272 30800 37392 6 io_eo[19]
port 45 nsew signal input
rlabel metal3 s 29200 29928 30800 30048 6 io_eo[1]
port 46 nsew signal input
rlabel metal3 s 29200 37680 30800 37800 6 io_eo[20]
port 47 nsew signal input
rlabel metal3 s 29200 38088 30800 38208 6 io_eo[21]
port 48 nsew signal input
rlabel metal3 s 29200 38496 30800 38616 6 io_eo[22]
port 49 nsew signal input
rlabel metal3 s 29200 38904 30800 39024 6 io_eo[23]
port 50 nsew signal input
rlabel metal3 s 29200 39312 30800 39432 6 io_eo[24]
port 51 nsew signal input
rlabel metal3 s 29200 39720 30800 39840 6 io_eo[25]
port 52 nsew signal input
rlabel metal3 s 29200 40128 30800 40248 6 io_eo[26]
port 53 nsew signal input
rlabel metal3 s 29200 40536 30800 40656 6 io_eo[27]
port 54 nsew signal input
rlabel metal3 s 29200 40944 30800 41064 6 io_eo[28]
port 55 nsew signal input
rlabel metal3 s 29200 41352 30800 41472 6 io_eo[29]
port 56 nsew signal input
rlabel metal3 s 29200 30336 30800 30456 6 io_eo[2]
port 57 nsew signal input
rlabel metal3 s 29200 41760 30800 41880 6 io_eo[30]
port 58 nsew signal input
rlabel metal3 s 29200 42168 30800 42288 6 io_eo[31]
port 59 nsew signal input
rlabel metal3 s 29200 42576 30800 42696 6 io_eo[32]
port 60 nsew signal input
rlabel metal3 s 29200 42984 30800 43104 6 io_eo[33]
port 61 nsew signal input
rlabel metal3 s 29200 43392 30800 43512 6 io_eo[34]
port 62 nsew signal input
rlabel metal3 s 29200 43800 30800 43920 6 io_eo[35]
port 63 nsew signal input
rlabel metal3 s 29200 44208 30800 44328 6 io_eo[36]
port 64 nsew signal input
rlabel metal3 s 29200 44616 30800 44736 6 io_eo[37]
port 65 nsew signal input
rlabel metal3 s 29200 45024 30800 45144 6 io_eo[38]
port 66 nsew signal input
rlabel metal3 s 29200 45432 30800 45552 6 io_eo[39]
port 67 nsew signal input
rlabel metal3 s 29200 30744 30800 30864 6 io_eo[3]
port 68 nsew signal input
rlabel metal3 s 29200 45840 30800 45960 6 io_eo[40]
port 69 nsew signal input
rlabel metal3 s 29200 46248 30800 46368 6 io_eo[41]
port 70 nsew signal input
rlabel metal3 s 29200 46656 30800 46776 6 io_eo[42]
port 71 nsew signal input
rlabel metal3 s 29200 47064 30800 47184 6 io_eo[43]
port 72 nsew signal input
rlabel metal3 s 29200 47472 30800 47592 6 io_eo[44]
port 73 nsew signal input
rlabel metal3 s 29200 47880 30800 48000 6 io_eo[45]
port 74 nsew signal input
rlabel metal3 s 29200 48288 30800 48408 6 io_eo[46]
port 75 nsew signal input
rlabel metal3 s 29200 48696 30800 48816 6 io_eo[47]
port 76 nsew signal input
rlabel metal3 s 29200 49104 30800 49224 6 io_eo[48]
port 77 nsew signal input
rlabel metal3 s 29200 49512 30800 49632 6 io_eo[49]
port 78 nsew signal input
rlabel metal3 s 29200 31152 30800 31272 6 io_eo[4]
port 79 nsew signal input
rlabel metal3 s 29200 49920 30800 50040 6 io_eo[50]
port 80 nsew signal input
rlabel metal3 s 29200 50328 30800 50448 6 io_eo[51]
port 81 nsew signal input
rlabel metal3 s 29200 50736 30800 50856 6 io_eo[52]
port 82 nsew signal input
rlabel metal3 s 29200 51144 30800 51264 6 io_eo[53]
port 83 nsew signal input
rlabel metal3 s 29200 51552 30800 51672 6 io_eo[54]
port 84 nsew signal input
rlabel metal3 s 29200 51960 30800 52080 6 io_eo[55]
port 85 nsew signal input
rlabel metal3 s 29200 52368 30800 52488 6 io_eo[56]
port 86 nsew signal input
rlabel metal3 s 29200 52776 30800 52896 6 io_eo[57]
port 87 nsew signal input
rlabel metal3 s 29200 53184 30800 53304 6 io_eo[58]
port 88 nsew signal input
rlabel metal3 s 29200 53592 30800 53712 6 io_eo[59]
port 89 nsew signal input
rlabel metal3 s 29200 31560 30800 31680 6 io_eo[5]
port 90 nsew signal input
rlabel metal3 s 29200 54000 30800 54120 6 io_eo[60]
port 91 nsew signal input
rlabel metal3 s 29200 54408 30800 54528 6 io_eo[61]
port 92 nsew signal input
rlabel metal3 s 29200 54816 30800 54936 6 io_eo[62]
port 93 nsew signal input
rlabel metal3 s 29200 55224 30800 55344 6 io_eo[63]
port 94 nsew signal input
rlabel metal3 s 29200 31968 30800 32088 6 io_eo[6]
port 95 nsew signal input
rlabel metal3 s 29200 32376 30800 32496 6 io_eo[7]
port 96 nsew signal input
rlabel metal3 s 29200 32784 30800 32904 6 io_eo[8]
port 97 nsew signal input
rlabel metal3 s 29200 33192 30800 33312 6 io_eo[9]
port 98 nsew signal input
rlabel metal3 s -800 144 800 264 4 io_i_0_ci
port 99 nsew signal input
rlabel metal3 s -800 3408 800 3528 4 io_i_0_in1[0]
port 100 nsew signal input
rlabel metal3 s -800 6672 800 6792 4 io_i_0_in1[1]
port 101 nsew signal input
rlabel metal3 s -800 9936 800 10056 4 io_i_0_in1[2]
port 102 nsew signal input
rlabel metal3 s -800 13200 800 13320 4 io_i_0_in1[3]
port 103 nsew signal input
rlabel metal3 s -800 16464 800 16584 4 io_i_0_in1[4]
port 104 nsew signal input
rlabel metal3 s -800 19728 800 19848 4 io_i_0_in1[5]
port 105 nsew signal input
rlabel metal3 s -800 22992 800 23112 4 io_i_0_in1[6]
port 106 nsew signal input
rlabel metal3 s -800 26256 800 26376 4 io_i_0_in1[7]
port 107 nsew signal input
rlabel metal3 s -800 552 800 672 4 io_i_1_ci
port 108 nsew signal input
rlabel metal3 s -800 3816 800 3936 4 io_i_1_in1[0]
port 109 nsew signal input
rlabel metal3 s -800 7080 800 7200 4 io_i_1_in1[1]
port 110 nsew signal input
rlabel metal3 s -800 10344 800 10464 4 io_i_1_in1[2]
port 111 nsew signal input
rlabel metal3 s -800 13608 800 13728 4 io_i_1_in1[3]
port 112 nsew signal input
rlabel metal3 s -800 16872 800 16992 4 io_i_1_in1[4]
port 113 nsew signal input
rlabel metal3 s -800 20136 800 20256 4 io_i_1_in1[5]
port 114 nsew signal input
rlabel metal3 s -800 23400 800 23520 4 io_i_1_in1[6]
port 115 nsew signal input
rlabel metal3 s -800 26664 800 26784 4 io_i_1_in1[7]
port 116 nsew signal input
rlabel metal3 s -800 960 800 1080 4 io_i_2_ci
port 117 nsew signal input
rlabel metal3 s -800 4224 800 4344 4 io_i_2_in1[0]
port 118 nsew signal input
rlabel metal3 s -800 7488 800 7608 4 io_i_2_in1[1]
port 119 nsew signal input
rlabel metal3 s -800 10752 800 10872 4 io_i_2_in1[2]
port 120 nsew signal input
rlabel metal3 s -800 14016 800 14136 4 io_i_2_in1[3]
port 121 nsew signal input
rlabel metal3 s -800 17280 800 17400 4 io_i_2_in1[4]
port 122 nsew signal input
rlabel metal3 s -800 20544 800 20664 4 io_i_2_in1[5]
port 123 nsew signal input
rlabel metal3 s -800 23808 800 23928 4 io_i_2_in1[6]
port 124 nsew signal input
rlabel metal3 s -800 27072 800 27192 4 io_i_2_in1[7]
port 125 nsew signal input
rlabel metal3 s -800 1368 800 1488 4 io_i_3_ci
port 126 nsew signal input
rlabel metal3 s -800 4632 800 4752 4 io_i_3_in1[0]
port 127 nsew signal input
rlabel metal3 s -800 7896 800 8016 4 io_i_3_in1[1]
port 128 nsew signal input
rlabel metal3 s -800 11160 800 11280 4 io_i_3_in1[2]
port 129 nsew signal input
rlabel metal3 s -800 14424 800 14544 4 io_i_3_in1[3]
port 130 nsew signal input
rlabel metal3 s -800 17688 800 17808 4 io_i_3_in1[4]
port 131 nsew signal input
rlabel metal3 s -800 20952 800 21072 4 io_i_3_in1[5]
port 132 nsew signal input
rlabel metal3 s -800 24216 800 24336 4 io_i_3_in1[6]
port 133 nsew signal input
rlabel metal3 s -800 27480 800 27600 4 io_i_3_in1[7]
port 134 nsew signal input
rlabel metal3 s -800 1776 800 1896 4 io_i_4_ci
port 135 nsew signal input
rlabel metal3 s -800 5040 800 5160 4 io_i_4_in1[0]
port 136 nsew signal input
rlabel metal3 s -800 8304 800 8424 4 io_i_4_in1[1]
port 137 nsew signal input
rlabel metal3 s -800 11568 800 11688 4 io_i_4_in1[2]
port 138 nsew signal input
rlabel metal3 s -800 14832 800 14952 4 io_i_4_in1[3]
port 139 nsew signal input
rlabel metal3 s -800 18096 800 18216 4 io_i_4_in1[4]
port 140 nsew signal input
rlabel metal3 s -800 21360 800 21480 4 io_i_4_in1[5]
port 141 nsew signal input
rlabel metal3 s -800 24624 800 24744 4 io_i_4_in1[6]
port 142 nsew signal input
rlabel metal3 s -800 27888 800 28008 4 io_i_4_in1[7]
port 143 nsew signal input
rlabel metal3 s -800 2184 800 2304 4 io_i_5_ci
port 144 nsew signal input
rlabel metal3 s -800 5448 800 5568 4 io_i_5_in1[0]
port 145 nsew signal input
rlabel metal3 s -800 8712 800 8832 4 io_i_5_in1[1]
port 146 nsew signal input
rlabel metal3 s -800 11976 800 12096 4 io_i_5_in1[2]
port 147 nsew signal input
rlabel metal3 s -800 15240 800 15360 4 io_i_5_in1[3]
port 148 nsew signal input
rlabel metal3 s -800 18504 800 18624 4 io_i_5_in1[4]
port 149 nsew signal input
rlabel metal3 s -800 21768 800 21888 4 io_i_5_in1[5]
port 150 nsew signal input
rlabel metal3 s -800 25032 800 25152 4 io_i_5_in1[6]
port 151 nsew signal input
rlabel metal3 s -800 28296 800 28416 4 io_i_5_in1[7]
port 152 nsew signal input
rlabel metal3 s -800 2592 800 2712 4 io_i_6_ci
port 153 nsew signal input
rlabel metal3 s -800 5856 800 5976 4 io_i_6_in1[0]
port 154 nsew signal input
rlabel metal3 s -800 9120 800 9240 4 io_i_6_in1[1]
port 155 nsew signal input
rlabel metal3 s -800 12384 800 12504 4 io_i_6_in1[2]
port 156 nsew signal input
rlabel metal3 s -800 15648 800 15768 4 io_i_6_in1[3]
port 157 nsew signal input
rlabel metal3 s -800 18912 800 19032 4 io_i_6_in1[4]
port 158 nsew signal input
rlabel metal3 s -800 22176 800 22296 4 io_i_6_in1[5]
port 159 nsew signal input
rlabel metal3 s -800 25440 800 25560 4 io_i_6_in1[6]
port 160 nsew signal input
rlabel metal3 s -800 28704 800 28824 4 io_i_6_in1[7]
port 161 nsew signal input
rlabel metal3 s -800 3000 800 3120 4 io_i_7_ci
port 162 nsew signal input
rlabel metal3 s -800 6264 800 6384 4 io_i_7_in1[0]
port 163 nsew signal input
rlabel metal3 s -800 9528 800 9648 4 io_i_7_in1[1]
port 164 nsew signal input
rlabel metal3 s -800 12792 800 12912 4 io_i_7_in1[2]
port 165 nsew signal input
rlabel metal3 s -800 16056 800 16176 4 io_i_7_in1[3]
port 166 nsew signal input
rlabel metal3 s -800 19320 800 19440 4 io_i_7_in1[4]
port 167 nsew signal input
rlabel metal3 s -800 22584 800 22704 4 io_i_7_in1[5]
port 168 nsew signal input
rlabel metal3 s -800 25848 800 25968 4 io_i_7_in1[6]
port 169 nsew signal input
rlabel metal3 s -800 29112 800 29232 4 io_i_7_in1[7]
port 170 nsew signal input
rlabel metal3 s 29200 144 30800 264 6 io_o_0_co
port 171 nsew signal tristate
rlabel metal3 s 29200 3408 30800 3528 6 io_o_0_out[0]
port 172 nsew signal tristate
rlabel metal3 s 29200 6672 30800 6792 6 io_o_0_out[1]
port 173 nsew signal tristate
rlabel metal3 s 29200 9936 30800 10056 6 io_o_0_out[2]
port 174 nsew signal tristate
rlabel metal3 s 29200 13200 30800 13320 6 io_o_0_out[3]
port 175 nsew signal tristate
rlabel metal3 s 29200 16464 30800 16584 6 io_o_0_out[4]
port 176 nsew signal tristate
rlabel metal3 s 29200 19728 30800 19848 6 io_o_0_out[5]
port 177 nsew signal tristate
rlabel metal3 s 29200 22992 30800 23112 6 io_o_0_out[6]
port 178 nsew signal tristate
rlabel metal3 s 29200 26256 30800 26376 6 io_o_0_out[7]
port 179 nsew signal tristate
rlabel metal3 s 29200 552 30800 672 6 io_o_1_co
port 180 nsew signal tristate
rlabel metal3 s 29200 3816 30800 3936 6 io_o_1_out[0]
port 181 nsew signal tristate
rlabel metal3 s 29200 7080 30800 7200 6 io_o_1_out[1]
port 182 nsew signal tristate
rlabel metal3 s 29200 10344 30800 10464 6 io_o_1_out[2]
port 183 nsew signal tristate
rlabel metal3 s 29200 13608 30800 13728 6 io_o_1_out[3]
port 184 nsew signal tristate
rlabel metal3 s 29200 16872 30800 16992 6 io_o_1_out[4]
port 185 nsew signal tristate
rlabel metal3 s 29200 20136 30800 20256 6 io_o_1_out[5]
port 186 nsew signal tristate
rlabel metal3 s 29200 23400 30800 23520 6 io_o_1_out[6]
port 187 nsew signal tristate
rlabel metal3 s 29200 26664 30800 26784 6 io_o_1_out[7]
port 188 nsew signal tristate
rlabel metal3 s 29200 960 30800 1080 6 io_o_2_co
port 189 nsew signal tristate
rlabel metal3 s 29200 4224 30800 4344 6 io_o_2_out[0]
port 190 nsew signal tristate
rlabel metal3 s 29200 7488 30800 7608 6 io_o_2_out[1]
port 191 nsew signal tristate
rlabel metal3 s 29200 10752 30800 10872 6 io_o_2_out[2]
port 192 nsew signal tristate
rlabel metal3 s 29200 14016 30800 14136 6 io_o_2_out[3]
port 193 nsew signal tristate
rlabel metal3 s 29200 17280 30800 17400 6 io_o_2_out[4]
port 194 nsew signal tristate
rlabel metal3 s 29200 20544 30800 20664 6 io_o_2_out[5]
port 195 nsew signal tristate
rlabel metal3 s 29200 23808 30800 23928 6 io_o_2_out[6]
port 196 nsew signal tristate
rlabel metal3 s 29200 27072 30800 27192 6 io_o_2_out[7]
port 197 nsew signal tristate
rlabel metal3 s 29200 1368 30800 1488 6 io_o_3_co
port 198 nsew signal tristate
rlabel metal3 s 29200 4632 30800 4752 6 io_o_3_out[0]
port 199 nsew signal tristate
rlabel metal3 s 29200 7896 30800 8016 6 io_o_3_out[1]
port 200 nsew signal tristate
rlabel metal3 s 29200 11160 30800 11280 6 io_o_3_out[2]
port 201 nsew signal tristate
rlabel metal3 s 29200 14424 30800 14544 6 io_o_3_out[3]
port 202 nsew signal tristate
rlabel metal3 s 29200 17688 30800 17808 6 io_o_3_out[4]
port 203 nsew signal tristate
rlabel metal3 s 29200 20952 30800 21072 6 io_o_3_out[5]
port 204 nsew signal tristate
rlabel metal3 s 29200 24216 30800 24336 6 io_o_3_out[6]
port 205 nsew signal tristate
rlabel metal3 s 29200 27480 30800 27600 6 io_o_3_out[7]
port 206 nsew signal tristate
rlabel metal3 s 29200 1776 30800 1896 6 io_o_4_co
port 207 nsew signal tristate
rlabel metal3 s 29200 5040 30800 5160 6 io_o_4_out[0]
port 208 nsew signal tristate
rlabel metal3 s 29200 8304 30800 8424 6 io_o_4_out[1]
port 209 nsew signal tristate
rlabel metal3 s 29200 11568 30800 11688 6 io_o_4_out[2]
port 210 nsew signal tristate
rlabel metal3 s 29200 14832 30800 14952 6 io_o_4_out[3]
port 211 nsew signal tristate
rlabel metal3 s 29200 18096 30800 18216 6 io_o_4_out[4]
port 212 nsew signal tristate
rlabel metal3 s 29200 21360 30800 21480 6 io_o_4_out[5]
port 213 nsew signal tristate
rlabel metal3 s 29200 24624 30800 24744 6 io_o_4_out[6]
port 214 nsew signal tristate
rlabel metal3 s 29200 27888 30800 28008 6 io_o_4_out[7]
port 215 nsew signal tristate
rlabel metal3 s 29200 2184 30800 2304 6 io_o_5_co
port 216 nsew signal tristate
rlabel metal3 s 29200 5448 30800 5568 6 io_o_5_out[0]
port 217 nsew signal tristate
rlabel metal3 s 29200 8712 30800 8832 6 io_o_5_out[1]
port 218 nsew signal tristate
rlabel metal3 s 29200 11976 30800 12096 6 io_o_5_out[2]
port 219 nsew signal tristate
rlabel metal3 s 29200 15240 30800 15360 6 io_o_5_out[3]
port 220 nsew signal tristate
rlabel metal3 s 29200 18504 30800 18624 6 io_o_5_out[4]
port 221 nsew signal tristate
rlabel metal3 s 29200 21768 30800 21888 6 io_o_5_out[5]
port 222 nsew signal tristate
rlabel metal3 s 29200 25032 30800 25152 6 io_o_5_out[6]
port 223 nsew signal tristate
rlabel metal3 s 29200 28296 30800 28416 6 io_o_5_out[7]
port 224 nsew signal tristate
rlabel metal3 s 29200 2592 30800 2712 6 io_o_6_co
port 225 nsew signal tristate
rlabel metal3 s 29200 5856 30800 5976 6 io_o_6_out[0]
port 226 nsew signal tristate
rlabel metal3 s 29200 9120 30800 9240 6 io_o_6_out[1]
port 227 nsew signal tristate
rlabel metal3 s 29200 12384 30800 12504 6 io_o_6_out[2]
port 228 nsew signal tristate
rlabel metal3 s 29200 15648 30800 15768 6 io_o_6_out[3]
port 229 nsew signal tristate
rlabel metal3 s 29200 18912 30800 19032 6 io_o_6_out[4]
port 230 nsew signal tristate
rlabel metal3 s 29200 22176 30800 22296 6 io_o_6_out[5]
port 231 nsew signal tristate
rlabel metal3 s 29200 25440 30800 25560 6 io_o_6_out[6]
port 232 nsew signal tristate
rlabel metal3 s 29200 28704 30800 28824 6 io_o_6_out[7]
port 233 nsew signal tristate
rlabel metal3 s 29200 3000 30800 3120 6 io_o_7_co
port 234 nsew signal tristate
rlabel metal3 s 29200 6264 30800 6384 6 io_o_7_out[0]
port 235 nsew signal tristate
rlabel metal3 s 29200 9528 30800 9648 6 io_o_7_out[1]
port 236 nsew signal tristate
rlabel metal3 s 29200 12792 30800 12912 6 io_o_7_out[2]
port 237 nsew signal tristate
rlabel metal3 s 29200 16056 30800 16176 6 io_o_7_out[3]
port 238 nsew signal tristate
rlabel metal3 s 29200 19320 30800 19440 6 io_o_7_out[4]
port 239 nsew signal tristate
rlabel metal3 s 29200 22584 30800 22704 6 io_o_7_out[5]
port 240 nsew signal tristate
rlabel metal3 s 29200 25848 30800 25968 6 io_o_7_out[6]
port 241 nsew signal tristate
rlabel metal3 s 29200 29112 30800 29232 6 io_o_7_out[7]
port 242 nsew signal tristate
rlabel metal2 s 662 -800 718 800 8 io_vci
port 243 nsew signal input
rlabel metal2 s 1950 -800 2006 800 8 io_vco
port 244 nsew signal tristate
rlabel metal2 s 28998 55200 29054 56800 6 io_vi
port 245 nsew signal input
rlabel metal2 s 4710 -800 4766 800 8 io_we_i
port 246 nsew signal input
rlabel metal3 s -800 29520 800 29640 4 io_wo[0]
port 247 nsew signal tristate
rlabel metal3 s -800 33600 800 33720 4 io_wo[10]
port 248 nsew signal tristate
rlabel metal3 s -800 34008 800 34128 4 io_wo[11]
port 249 nsew signal tristate
rlabel metal3 s -800 34416 800 34536 4 io_wo[12]
port 250 nsew signal tristate
rlabel metal3 s -800 34824 800 34944 4 io_wo[13]
port 251 nsew signal tristate
rlabel metal3 s -800 35232 800 35352 4 io_wo[14]
port 252 nsew signal tristate
rlabel metal3 s -800 35640 800 35760 4 io_wo[15]
port 253 nsew signal tristate
rlabel metal3 s -800 36048 800 36168 4 io_wo[16]
port 254 nsew signal tristate
rlabel metal3 s -800 36456 800 36576 4 io_wo[17]
port 255 nsew signal tristate
rlabel metal3 s -800 36864 800 36984 4 io_wo[18]
port 256 nsew signal tristate
rlabel metal3 s -800 37272 800 37392 4 io_wo[19]
port 257 nsew signal tristate
rlabel metal3 s -800 29928 800 30048 4 io_wo[1]
port 258 nsew signal tristate
rlabel metal3 s -800 37680 800 37800 4 io_wo[20]
port 259 nsew signal tristate
rlabel metal3 s -800 38088 800 38208 4 io_wo[21]
port 260 nsew signal tristate
rlabel metal3 s -800 38496 800 38616 4 io_wo[22]
port 261 nsew signal tristate
rlabel metal3 s -800 38904 800 39024 4 io_wo[23]
port 262 nsew signal tristate
rlabel metal3 s -800 39312 800 39432 4 io_wo[24]
port 263 nsew signal tristate
rlabel metal3 s -800 39720 800 39840 4 io_wo[25]
port 264 nsew signal tristate
rlabel metal3 s -800 40128 800 40248 4 io_wo[26]
port 265 nsew signal tristate
rlabel metal3 s -800 40536 800 40656 4 io_wo[27]
port 266 nsew signal tristate
rlabel metal3 s -800 40944 800 41064 4 io_wo[28]
port 267 nsew signal tristate
rlabel metal3 s -800 41352 800 41472 4 io_wo[29]
port 268 nsew signal tristate
rlabel metal3 s -800 30336 800 30456 4 io_wo[2]
port 269 nsew signal tristate
rlabel metal3 s -800 41760 800 41880 4 io_wo[30]
port 270 nsew signal tristate
rlabel metal3 s -800 42168 800 42288 4 io_wo[31]
port 271 nsew signal tristate
rlabel metal3 s -800 42576 800 42696 4 io_wo[32]
port 272 nsew signal tristate
rlabel metal3 s -800 42984 800 43104 4 io_wo[33]
port 273 nsew signal tristate
rlabel metal3 s -800 43392 800 43512 4 io_wo[34]
port 274 nsew signal tristate
rlabel metal3 s -800 43800 800 43920 4 io_wo[35]
port 275 nsew signal tristate
rlabel metal3 s -800 44208 800 44328 4 io_wo[36]
port 276 nsew signal tristate
rlabel metal3 s -800 44616 800 44736 4 io_wo[37]
port 277 nsew signal tristate
rlabel metal3 s -800 45024 800 45144 4 io_wo[38]
port 278 nsew signal tristate
rlabel metal3 s -800 45432 800 45552 4 io_wo[39]
port 279 nsew signal tristate
rlabel metal3 s -800 30744 800 30864 4 io_wo[3]
port 280 nsew signal tristate
rlabel metal3 s -800 45840 800 45960 4 io_wo[40]
port 281 nsew signal tristate
rlabel metal3 s -800 46248 800 46368 4 io_wo[41]
port 282 nsew signal tristate
rlabel metal3 s -800 46656 800 46776 4 io_wo[42]
port 283 nsew signal tristate
rlabel metal3 s -800 47064 800 47184 4 io_wo[43]
port 284 nsew signal tristate
rlabel metal3 s -800 47472 800 47592 4 io_wo[44]
port 285 nsew signal tristate
rlabel metal3 s -800 47880 800 48000 4 io_wo[45]
port 286 nsew signal tristate
rlabel metal3 s -800 48288 800 48408 4 io_wo[46]
port 287 nsew signal tristate
rlabel metal3 s -800 48696 800 48816 4 io_wo[47]
port 288 nsew signal tristate
rlabel metal3 s -800 49104 800 49224 4 io_wo[48]
port 289 nsew signal tristate
rlabel metal3 s -800 49512 800 49632 4 io_wo[49]
port 290 nsew signal tristate
rlabel metal3 s -800 31152 800 31272 4 io_wo[4]
port 291 nsew signal tristate
rlabel metal3 s -800 49920 800 50040 4 io_wo[50]
port 292 nsew signal tristate
rlabel metal3 s -800 50328 800 50448 4 io_wo[51]
port 293 nsew signal tristate
rlabel metal3 s -800 50736 800 50856 4 io_wo[52]
port 294 nsew signal tristate
rlabel metal3 s -800 51144 800 51264 4 io_wo[53]
port 295 nsew signal tristate
rlabel metal3 s -800 51552 800 51672 4 io_wo[54]
port 296 nsew signal tristate
rlabel metal3 s -800 51960 800 52080 4 io_wo[55]
port 297 nsew signal tristate
rlabel metal3 s -800 52368 800 52488 4 io_wo[56]
port 298 nsew signal tristate
rlabel metal3 s -800 52776 800 52896 4 io_wo[57]
port 299 nsew signal tristate
rlabel metal3 s -800 53184 800 53304 4 io_wo[58]
port 300 nsew signal tristate
rlabel metal3 s -800 53592 800 53712 4 io_wo[59]
port 301 nsew signal tristate
rlabel metal3 s -800 31560 800 31680 4 io_wo[5]
port 302 nsew signal tristate
rlabel metal3 s -800 54000 800 54120 4 io_wo[60]
port 303 nsew signal tristate
rlabel metal3 s -800 54408 800 54528 4 io_wo[61]
port 304 nsew signal tristate
rlabel metal3 s -800 54816 800 54936 4 io_wo[62]
port 305 nsew signal tristate
rlabel metal3 s -800 55224 800 55344 4 io_wo[63]
port 306 nsew signal tristate
rlabel metal3 s -800 31968 800 32088 4 io_wo[6]
port 307 nsew signal tristate
rlabel metal3 s -800 32376 800 32496 4 io_wo[7]
port 308 nsew signal tristate
rlabel metal3 s -800 32784 800 32904 4 io_wo[8]
port 309 nsew signal tristate
rlabel metal3 s -800 33192 800 33312 4 io_wo[9]
port 310 nsew signal tristate
rlabel metal3 s 29200 55632 30800 55752 6 wb_clk_i
port 311 nsew signal input
rlabel metal3 s -800 55632 800 55752 4 wb_rst_i
port 312 nsew signal input
rlabel metal4 s 24104 2128 24424 53360 6 vccd1
port 313 nsew power bidirectional
rlabel metal4 s 14840 2128 15160 53360 6 vccd1
port 314 nsew power bidirectional
rlabel metal4 s 5576 2128 5896 53360 6 vccd1
port 315 nsew power bidirectional
rlabel metal4 s 19472 2128 19792 53360 6 vssd1
port 316 nsew ground bidirectional
rlabel metal4 s 10208 2128 10528 53360 6 vssd1
port 317 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 56000
<< end >>
