* NGSPICE file created from cic_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

.subckt cic_block io_adr_i[0] io_adr_i[1] io_cs_i io_dat_i[0] io_dat_i[10] io_dat_i[11]
+ io_dat_i[12] io_dat_i[13] io_dat_i[14] io_dat_i[15] io_dat_i[1] io_dat_i[2] io_dat_i[3]
+ io_dat_i[4] io_dat_i[5] io_dat_i[6] io_dat_i[7] io_dat_i[8] io_dat_i[9] io_dat_o[0]
+ io_dat_o[10] io_dat_o[11] io_dat_o[12] io_dat_o[13] io_dat_o[14] io_dat_o[15] io_dat_o[1]
+ io_dat_o[2] io_dat_o[3] io_dat_o[4] io_dat_o[5] io_dat_o[6] io_dat_o[7] io_dat_o[8]
+ io_dat_o[9] io_eo[0] io_eo[10] io_eo[11] io_eo[12] io_eo[13] io_eo[14] io_eo[15]
+ io_eo[16] io_eo[17] io_eo[18] io_eo[19] io_eo[1] io_eo[20] io_eo[21] io_eo[22] io_eo[23]
+ io_eo[24] io_eo[25] io_eo[26] io_eo[27] io_eo[28] io_eo[29] io_eo[2] io_eo[30] io_eo[31]
+ io_eo[32] io_eo[33] io_eo[34] io_eo[35] io_eo[36] io_eo[37] io_eo[38] io_eo[39]
+ io_eo[3] io_eo[40] io_eo[41] io_eo[42] io_eo[43] io_eo[44] io_eo[45] io_eo[46] io_eo[47]
+ io_eo[48] io_eo[49] io_eo[4] io_eo[50] io_eo[51] io_eo[52] io_eo[53] io_eo[54] io_eo[55]
+ io_eo[56] io_eo[57] io_eo[58] io_eo[59] io_eo[5] io_eo[60] io_eo[61] io_eo[62] io_eo[63]
+ io_eo[6] io_eo[7] io_eo[8] io_eo[9] io_i_0_ci io_i_0_in1[0] io_i_0_in1[1] io_i_0_in1[2]
+ io_i_0_in1[3] io_i_0_in1[4] io_i_0_in1[5] io_i_0_in1[6] io_i_0_in1[7] io_i_1_ci
+ io_i_1_in1[0] io_i_1_in1[1] io_i_1_in1[2] io_i_1_in1[3] io_i_1_in1[4] io_i_1_in1[5]
+ io_i_1_in1[6] io_i_1_in1[7] io_i_2_ci io_i_2_in1[0] io_i_2_in1[1] io_i_2_in1[2]
+ io_i_2_in1[3] io_i_2_in1[4] io_i_2_in1[5] io_i_2_in1[6] io_i_2_in1[7] io_i_3_ci
+ io_i_3_in1[0] io_i_3_in1[1] io_i_3_in1[2] io_i_3_in1[3] io_i_3_in1[4] io_i_3_in1[5]
+ io_i_3_in1[6] io_i_3_in1[7] io_i_4_ci io_i_4_in1[0] io_i_4_in1[1] io_i_4_in1[2]
+ io_i_4_in1[3] io_i_4_in1[4] io_i_4_in1[5] io_i_4_in1[6] io_i_4_in1[7] io_i_5_ci
+ io_i_5_in1[0] io_i_5_in1[1] io_i_5_in1[2] io_i_5_in1[3] io_i_5_in1[4] io_i_5_in1[5]
+ io_i_5_in1[6] io_i_5_in1[7] io_i_6_ci io_i_6_in1[0] io_i_6_in1[1] io_i_6_in1[2]
+ io_i_6_in1[3] io_i_6_in1[4] io_i_6_in1[5] io_i_6_in1[6] io_i_6_in1[7] io_i_7_ci
+ io_i_7_in1[0] io_i_7_in1[1] io_i_7_in1[2] io_i_7_in1[3] io_i_7_in1[4] io_i_7_in1[5]
+ io_i_7_in1[6] io_i_7_in1[7] io_o_0_co io_o_0_out[0] io_o_0_out[1] io_o_0_out[2]
+ io_o_0_out[3] io_o_0_out[4] io_o_0_out[5] io_o_0_out[6] io_o_0_out[7] io_o_1_co
+ io_o_1_out[0] io_o_1_out[1] io_o_1_out[2] io_o_1_out[3] io_o_1_out[4] io_o_1_out[5]
+ io_o_1_out[6] io_o_1_out[7] io_o_2_co io_o_2_out[0] io_o_2_out[1] io_o_2_out[2]
+ io_o_2_out[3] io_o_2_out[4] io_o_2_out[5] io_o_2_out[6] io_o_2_out[7] io_o_3_co
+ io_o_3_out[0] io_o_3_out[1] io_o_3_out[2] io_o_3_out[3] io_o_3_out[4] io_o_3_out[5]
+ io_o_3_out[6] io_o_3_out[7] io_o_4_co io_o_4_out[0] io_o_4_out[1] io_o_4_out[2]
+ io_o_4_out[3] io_o_4_out[4] io_o_4_out[5] io_o_4_out[6] io_o_4_out[7] io_o_5_co
+ io_o_5_out[0] io_o_5_out[1] io_o_5_out[2] io_o_5_out[3] io_o_5_out[4] io_o_5_out[5]
+ io_o_5_out[6] io_o_5_out[7] io_o_6_co io_o_6_out[0] io_o_6_out[1] io_o_6_out[2]
+ io_o_6_out[3] io_o_6_out[4] io_o_6_out[5] io_o_6_out[6] io_o_6_out[7] io_o_7_co
+ io_o_7_out[0] io_o_7_out[1] io_o_7_out[2] io_o_7_out[3] io_o_7_out[4] io_o_7_out[5]
+ io_o_7_out[6] io_o_7_out[7] io_vci io_vco io_vi io_we_i io_wo[0] io_wo[10] io_wo[11]
+ io_wo[12] io_wo[13] io_wo[14] io_wo[15] io_wo[16] io_wo[17] io_wo[18] io_wo[19]
+ io_wo[1] io_wo[20] io_wo[21] io_wo[22] io_wo[23] io_wo[24] io_wo[25] io_wo[26] io_wo[27]
+ io_wo[28] io_wo[29] io_wo[2] io_wo[30] io_wo[31] io_wo[32] io_wo[33] io_wo[34] io_wo[35]
+ io_wo[36] io_wo[37] io_wo[38] io_wo[39] io_wo[3] io_wo[40] io_wo[41] io_wo[42] io_wo[43]
+ io_wo[44] io_wo[45] io_wo[46] io_wo[47] io_wo[48] io_wo[49] io_wo[4] io_wo[50] io_wo[51]
+ io_wo[52] io_wo[53] io_wo[54] io_wo[55] io_wo[56] io_wo[57] io_wo[58] io_wo[59]
+ io_wo[5] io_wo[60] io_wo[61] io_wo[62] io_wo[63] io_wo[6] io_wo[7] io_wo[8] io_wo[9]
+ wb_clk_i wb_rst_i vccd1 vssd1
XFILLER_54_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2106_ input86/X _1695_/A _1658_/A _2119_/A0 _2244_/Q _2245_/Q vssd1 vssd1 vccd1
+ vccd1 _2106_/X sky130_fd_sc_hd__mux4_2
X_2037_ _1759_/Y _1684_/Y _2294_/Q vssd1 vssd1 vccd1 vccd1 _2037_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1270_ _1268_/Y _1269_/Y _1258_/A vssd1 vssd1 vccd1 vccd1 _1270_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1606_ _1607_/A _2137_/X _2138_/X _2139_/X vssd1 vssd1 vccd1 vccd1 _1606_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_86_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1399_ _1399_/A _1399_/B vssd1 vssd1 vccd1 vccd1 _1414_/B sky130_fd_sc_hd__nor2_4
X_1468_ _1963_/X _2087_/X vssd1 vssd1 vccd1 vccd1 _1475_/A sky130_fd_sc_hd__nor2_2
X_1537_ _1536_/X _2178_/Q _1546_/S vssd1 vssd1 vccd1 vccd1 _2178_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1253_ _1248_/B _1253_/B _1253_/C vssd1 vssd1 vccd1 vccd1 _1254_/B sky130_fd_sc_hd__nand3b_1
X_1322_ _2116_/X vssd1 vssd1 vccd1 vccd1 _1752_/A sky130_fd_sc_hd__inv_2
X_1184_ _1172_/X _1876_/C _1187_/C vssd1 vssd1 vccd1 vccd1 _1184_/Y sky130_fd_sc_hd__nand3b_1
Xoutput286 _1921_/X vssd1 vssd1 vccd1 vccd1 io_wo[43] sky130_fd_sc_hd__clkbuf_2
Xoutput275 _1911_/X vssd1 vssd1 vccd1 vccd1 io_wo[33] sky130_fd_sc_hd__clkbuf_2
Xoutput264 _1901_/X vssd1 vssd1 vccd1 vccd1 io_wo[23] sky130_fd_sc_hd__clkbuf_2
Xoutput253 _1891_/X vssd1 vssd1 vccd1 vccd1 io_wo[13] sky130_fd_sc_hd__clkbuf_2
Xoutput220 _2179_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput231 _2148_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput242 _2142_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput297 _1931_/X vssd1 vssd1 vccd1 vccd1 io_wo[53] sky130_fd_sc_hd__clkbuf_2
XFILLER_74_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1940_ _1940_/A vssd1 vssd1 vccd1 vccd1 _1940_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1871_ _1871_/A _2282_/Q vssd1 vssd1 vccd1 vccd1 _1871_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2285_ _2299_/CLK _2285_/D vssd1 vssd1 vccd1 vccd1 _2285_/Q sky130_fd_sc_hd__dfxtp_1
X_1236_ _1236_/A _1236_/B _1236_/C vssd1 vssd1 vccd1 vccd1 _1269_/B sky130_fd_sc_hd__nand3_4
XFILLER_49_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1305_ _2113_/X _1304_/Y _1758_/A _2038_/X vssd1 vssd1 vccd1 vccd1 _1305_/Y sky130_fd_sc_hd__o2bb2ai_2
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1098_ _2281_/Q _1095_/X _1088_/X _1097_/Y vssd1 vssd1 vccd1 vccd1 _2281_/D sky130_fd_sc_hd__o211a_1
X_1167_ _2258_/Q _1159_/X _1165_/X _1166_/Y vssd1 vssd1 vccd1 vccd1 _2258_/D sky130_fd_sc_hd__o211a_1
XFILLER_60_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2070_ _2070_/A0 _2227_/Q _2248_/Q vssd1 vssd1 vccd1 vccd1 _2070_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1021_ _1219_/A vssd1 vssd1 vccd1 vccd1 _1193_/A sky130_fd_sc_hd__inv_2
XFILLER_61_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1923_ _1923_/A vssd1 vssd1 vccd1 vccd1 _1923_/X sky130_fd_sc_hd__clkbuf_2
X_1854_ _2269_/Q _1849_/X _1850_/X _1853_/X vssd1 vssd1 vccd1 vccd1 _1854_/X sky130_fd_sc_hd__a31o_1
X_1785_ _2213_/Q vssd1 vssd1 vccd1 vccd1 _1785_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1219_ _1219_/A _1949_/X vssd1 vssd1 vccd1 vccd1 _2236_/D sky130_fd_sc_hd__nor2b_1
XFILLER_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2268_ _2268_/CLK _2268_/D vssd1 vssd1 vccd1 vccd1 _2268_/Q sky130_fd_sc_hd__dfxtp_2
X_2199_ _2231_/CLK _2199_/D vssd1 vssd1 vccd1 vccd1 _2199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ _1569_/Y _2129_/X _2127_/X _2128_/X vssd1 vssd1 vccd1 vccd1 _1583_/B sky130_fd_sc_hd__and4b_1
XFILLER_6_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2053_ _1737_/Y _1736_/Y _2296_/Q vssd1 vssd1 vccd1 vccd1 _2053_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2122_ _2122_/A0 _2192_/Q _2208_/Q _2232_/Q _2252_/Q _2253_/Q vssd1 vssd1 vccd1 vccd1
+ _2122_/X sky130_fd_sc_hd__mux4_2
XFILLER_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1906_ _1906_/A vssd1 vssd1 vccd1 vccd1 _1906_/X sky130_fd_sc_hd__clkbuf_2
X_1837_ _1745_/Y _1814_/Y _1836_/Y vssd1 vssd1 vccd1 vccd1 _1837_/Y sky130_fd_sc_hd__o21ai_1
X_1768_ _2196_/Q vssd1 vssd1 vccd1 vccd1 _1768_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1699_ _1699_/A vssd1 vssd1 vccd1 vccd1 _1699_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput153 io_i_7_in1[5] vssd1 vssd1 vccd1 vccd1 _1672_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput120 io_i_4_ci vssd1 vssd1 vccd1 vccd1 _2003_/A0 sky130_fd_sc_hd__buf_1
Xinput131 io_i_5_in1[1] vssd1 vssd1 vccd1 vccd1 _1754_/A sky130_fd_sc_hd__clkbuf_1
Xinput142 io_i_6_in1[3] vssd1 vssd1 vccd1 vccd1 _1727_/A sky130_fd_sc_hd__clkbuf_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1622_ _2134_/X _1622_/B vssd1 vssd1 vccd1 vccd1 _1622_/Y sky130_fd_sc_hd__xnor2_1
X_1484_ _1951_/X vssd1 vssd1 vccd1 vccd1 _1485_/A sky130_fd_sc_hd__inv_2
XFILLER_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1553_ _1949_/X _1550_/Y _1552_/Y vssd1 vssd1 vccd1 vccd1 _2173_/D sky130_fd_sc_hd__o21ai_1
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2105_ input85/X _1699_/A _1742_/A _1803_/A _2244_/Q _2245_/Q vssd1 vssd1 vccd1 vccd1
+ _2105_/X sky130_fd_sc_hd__mux4_2
X_2036_ _1760_/Y _2035_/X _2295_/Q vssd1 vssd1 vccd1 vccd1 _2036_/X sky130_fd_sc_hd__mux2_2
XFILLER_62_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1536_ _1536_/A _1541_/B vssd1 vssd1 vccd1 vccd1 _1536_/X sky130_fd_sc_hd__xor2_1
X_1605_ _1618_/A _1618_/B vssd1 vssd1 vccd1 vccd1 _1607_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1398_ _1981_/X _2063_/X _1979_/X _2060_/X vssd1 vssd1 vccd1 vccd1 _1399_/B sky130_fd_sc_hd__a211oi_4
X_1467_ _1961_/X _2084_/X vssd1 vssd1 vccd1 vccd1 _1499_/A sky130_fd_sc_hd__xor2_4
X_2019_ _1781_/Y _1728_/Y _2292_/Q vssd1 vssd1 vccd1 vccd1 _2019_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1252_ _1262_/A _1252_/B _1262_/B vssd1 vssd1 vccd1 vccd1 _1253_/B sky130_fd_sc_hd__nand3_4
Xclkbuf_4_12_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2299_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1321_ _1350_/B _1350_/A _1348_/A _1305_/Y vssd1 vssd1 vccd1 vccd1 _1344_/B sky130_fd_sc_hd__a31oi_4
X_1183_ _2252_/Q _1175_/X _1179_/X _1182_/Y vssd1 vssd1 vccd1 vccd1 _2252_/D sky130_fd_sc_hd__o211a_1
XFILLER_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput298 _1932_/X vssd1 vssd1 vccd1 vccd1 io_wo[54] sky130_fd_sc_hd__clkbuf_2
Xoutput287 _1922_/X vssd1 vssd1 vccd1 vccd1 io_wo[44] sky130_fd_sc_hd__clkbuf_2
Xoutput276 _1912_/X vssd1 vssd1 vccd1 vccd1 io_wo[34] sky130_fd_sc_hd__clkbuf_2
X_1519_ _2186_/Q _1983_/X _1522_/S vssd1 vssd1 vccd1 vccd1 _2186_/D sky130_fd_sc_hd__mux2_1
Xoutput265 _1902_/X vssd1 vssd1 vccd1 vccd1 io_wo[24] sky130_fd_sc_hd__clkbuf_2
Xoutput254 _1892_/X vssd1 vssd1 vccd1 vccd1 io_wo[14] sky130_fd_sc_hd__clkbuf_2
Xoutput210 _2194_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput243 _2143_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput221 _1572_/X vssd1 vssd1 vccd1 vccd1 io_o_5_co sky130_fd_sc_hd__clkbuf_2
Xoutput232 _2149_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1870_ _1871_/A _2284_/Q vssd1 vssd1 vccd1 vccd1 _1870_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2284_ _2299_/CLK _2284_/D vssd1 vssd1 vccd1 vccd1 _2284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1166_ _1110_/X _1166_/B _1173_/C vssd1 vssd1 vccd1 vccd1 _1166_/Y sky130_fd_sc_hd__nand3b_1
X_1235_ _1235_/A vssd1 vssd1 vccd1 vccd1 _1236_/C sky130_fd_sc_hd__inv_2
X_1304_ _1758_/A _2038_/X _2036_/X vssd1 vssd1 vccd1 vccd1 _1304_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1097_ _1096_/X _1105_/B _1191_/B vssd1 vssd1 vccd1 vccd1 _1097_/Y sky130_fd_sc_hd__nand3b_1
X_1999_ _1999_/A0 _1572_/X _2272_/Q vssd1 vssd1 vccd1 vccd1 _1999_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1020_ _1032_/A vssd1 vssd1 vccd1 vccd1 _1020_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1922_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1922_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1853_ _2253_/Q _1203_/C _1111_/B _2285_/Q vssd1 vssd1 vccd1 vccd1 _1853_/X sky130_fd_sc_hd__a22o_1
X_1784_ _1784_/A _1821_/A vssd1 vssd1 vccd1 vccd1 _1784_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1218_ _1219_/A _1992_/A0 vssd1 vssd1 vccd1 vccd1 _2237_/D sky130_fd_sc_hd__nor2b_1
XFILLER_37_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2267_ _2268_/CLK _2267_/D vssd1 vssd1 vccd1 vccd1 _2267_/Q sky130_fd_sc_hd__dfxtp_2
X_2198_ _2231_/CLK _2198_/D vssd1 vssd1 vccd1 vccd1 _2198_/Q sky130_fd_sc_hd__dfxtp_1
X_1149_ _1151_/A _1196_/B vssd1 vssd1 vccd1 vccd1 _1149_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2052_ _2052_/A0 _2221_/Q _2248_/Q vssd1 vssd1 vccd1 vccd1 _2052_/X sky130_fd_sc_hd__mux2_1
X_2121_ _2121_/A0 _2191_/Q _2207_/Q _2231_/Q _2252_/Q _2253_/Q vssd1 vssd1 vccd1 vccd1
+ _2121_/X sky130_fd_sc_hd__mux4_2
X_1905_ _1905_/A vssd1 vssd1 vccd1 vccd1 _1905_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1836_ _1849_/A _1845_/B _2248_/Q vssd1 vssd1 vccd1 vccd1 _1836_/Y sky130_fd_sc_hd__nand3_1
X_1767_ _1767_/A _1989_/X vssd1 vssd1 vccd1 vccd1 _1767_/Y sky130_fd_sc_hd__nand2_1
X_1698_ _2073_/X vssd1 vssd1 vccd1 vccd1 _1698_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput110 io_i_2_in1[7] vssd1 vssd1 vccd1 vccd1 _2070_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput154 io_i_7_in1[6] vssd1 vssd1 vccd1 vccd1 _1667_/A sky130_fd_sc_hd__clkbuf_2
Xinput143 io_i_6_in1[4] vssd1 vssd1 vccd1 vccd1 _1721_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput121 io_i_4_in1[0] vssd1 vssd1 vccd1 vccd1 _1803_/A sky130_fd_sc_hd__buf_1
Xinput132 io_i_5_in1[2] vssd1 vssd1 vccd1 vccd1 _2127_/A0 sky130_fd_sc_hd__buf_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1552_ _1552_/A _1949_/X _1552_/C vssd1 vssd1 vccd1 vccd1 _1552_/Y sky130_fd_sc_hd__nand3_1
X_1621_ _1620_/X _2151_/Q _1628_/S vssd1 vssd1 vccd1 vccd1 _2151_/D sky130_fd_sc_hd__mux2_1
X_1483_ _1801_/A _1481_/A _1478_/Y _1476_/Y vssd1 vssd1 vccd1 vccd1 _1483_/X sky130_fd_sc_hd__o211a_1
XFILLER_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2104_ _1803_/Y _1512_/Y _1439_/Y _1291_/Y _2252_/Q _2253_/Q vssd1 vssd1 vccd1 vccd1
+ _2104_/X sky130_fd_sc_hd__mux4_2
X_2035_ _1761_/Y _1690_/Y _2294_/Q vssd1 vssd1 vccd1 vccd1 _2035_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1819_ _1850_/A _2276_/Q _1839_/A vssd1 vssd1 vccd1 vccd1 _1819_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_93_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1535_ _1546_/S _2179_/Q _1532_/Y _1534_/Y vssd1 vssd1 vccd1 vccd1 _2179_/D sky130_fd_sc_hd__o2bb2ai_1
X_1604_ _1622_/B _2134_/X _2135_/X vssd1 vssd1 vccd1 vccd1 _1618_/B sky130_fd_sc_hd__nand3b_2
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1466_ _1505_/B _1505_/A _1503_/A _1465_/Y vssd1 vssd1 vccd1 vccd1 _1499_/B sky130_fd_sc_hd__a31o_1
X_1397_ _1412_/A vssd1 vssd1 vccd1 vccd1 _1400_/B sky130_fd_sc_hd__inv_2
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2018_ _1782_/Y _2017_/X _2293_/Q vssd1 vssd1 vccd1 vccd1 _2018_/X sky130_fd_sc_hd__mux2_2
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1320_ _1320_/A vssd1 vssd1 vccd1 vccd1 _1344_/A sky130_fd_sc_hd__inv_2
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1251_ _1245_/C _1239_/A _1239_/B vssd1 vssd1 vccd1 vccd1 _1262_/B sky130_fd_sc_hd__a21oi_4
X_1182_ _1172_/X _1182_/B _1187_/C vssd1 vssd1 vccd1 vccd1 _1182_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_91_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput200 _2209_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[5] sky130_fd_sc_hd__clkbuf_2
Xoutput299 _1933_/X vssd1 vssd1 vccd1 vccd1 io_wo[55] sky130_fd_sc_hd__clkbuf_2
Xoutput288 _1923_/X vssd1 vssd1 vccd1 vccd1 io_wo[45] sky130_fd_sc_hd__clkbuf_2
Xoutput277 _1913_/X vssd1 vssd1 vccd1 vccd1 io_wo[35] sky130_fd_sc_hd__clkbuf_2
X_1518_ _2187_/Q _1985_/X _1522_/S vssd1 vssd1 vccd1 vccd1 _2187_/D sky130_fd_sc_hd__mux2_1
Xoutput266 _1903_/X vssd1 vssd1 vccd1 vccd1 io_wo[25] sky130_fd_sc_hd__clkbuf_2
Xoutput255 _1893_/X vssd1 vssd1 vccd1 vccd1 io_wo[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput211 _2195_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput244 _2144_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput222 _2156_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[0] sky130_fd_sc_hd__clkbuf_2
X_1449_ _2197_/Q _1991_/X _1450_/S vssd1 vssd1 vccd1 vccd1 _2197_/D sky130_fd_sc_hd__mux2_1
Xoutput233 _2150_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2283_ _2299_/CLK _2283_/D vssd1 vssd1 vccd1 vccd1 _2283_/Q sky130_fd_sc_hd__dfxtp_1
X_1303_ _2114_/X vssd1 vssd1 vccd1 vccd1 _1758_/A sky130_fd_sc_hd__inv_2
X_1096_ _1110_/A vssd1 vssd1 vccd1 vccd1 _1096_/X sky130_fd_sc_hd__buf_1
X_1234_ _2108_/X _2020_/X vssd1 vssd1 vccd1 vccd1 _1235_/A sky130_fd_sc_hd__and2b_1
X_1165_ _1165_/A vssd1 vssd1 vccd1 vccd1 _1165_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1998_ _2274_/Q _1997_/X _2275_/Q vssd1 vssd1 vccd1 vccd1 _1998_/X sky130_fd_sc_hd__mux2_2
XFILLER_85_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1921_ _1921_/A vssd1 vssd1 vccd1 vccd1 _1921_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1852_ _2268_/Q _1849_/X _1850_/X _1851_/X vssd1 vssd1 vccd1 vccd1 _1852_/X sky130_fd_sc_hd__a31o_1
XFILLER_6_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1783_ _2214_/Q vssd1 vssd1 vccd1 vccd1 _1783_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2266_ _2268_/CLK _2266_/D vssd1 vssd1 vccd1 vccd1 _2266_/Q sky130_fd_sc_hd__dfxtp_1
X_1217_ _1219_/A _1216_/X vssd1 vssd1 vccd1 vccd1 _2238_/D sky130_fd_sc_hd__nor2b_1
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1079_ input5/X vssd1 vssd1 vccd1 vccd1 _1177_/B sky130_fd_sc_hd__inv_2
X_2197_ _2231_/CLK _2197_/D vssd1 vssd1 vccd1 vccd1 _2197_/Q sky130_fd_sc_hd__dfxtp_1
X_1148_ _1165_/A vssd1 vssd1 vccd1 vccd1 _1148_/X sky130_fd_sc_hd__buf_2
XFILLER_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2120_ _2120_/A0 _2190_/Q _2206_/Q _2230_/Q _2252_/Q _2253_/Q vssd1 vssd1 vccd1 vccd1
+ _2120_/X sky130_fd_sc_hd__mux4_2
X_2051_ _1739_/Y _2050_/X _2297_/Q vssd1 vssd1 vccd1 vccd1 _2051_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1904_ _1904_/A vssd1 vssd1 vccd1 vccd1 _1904_/X sky130_fd_sc_hd__clkbuf_2
X_1835_ _2295_/Q _1824_/X _2279_/Q _1825_/X _1834_/X vssd1 vssd1 vccd1 vccd1 _1835_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1697_ _2165_/Q vssd1 vssd1 vccd1 vccd1 _1697_/Y sky130_fd_sc_hd__inv_2
X_1766_ _1766_/A vssd1 vssd1 vccd1 vccd1 _1766_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2249_ _2254_/CLK _2249_/D vssd1 vssd1 vccd1 vccd1 _2249_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput100 io_i_1_in1[6] vssd1 vssd1 vccd1 vccd1 _2117_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput144 io_i_6_in1[5] vssd1 vssd1 vccd1 vccd1 _1716_/A sky130_fd_sc_hd__clkbuf_2
Xinput133 io_i_5_in1[3] vssd1 vssd1 vccd1 vccd1 _2128_/A0 sky130_fd_sc_hd__buf_1
Xinput111 io_i_3_ci vssd1 vssd1 vccd1 vccd1 _1703_/A sky130_fd_sc_hd__clkbuf_1
Xinput122 io_i_4_in1[1] vssd1 vssd1 vccd1 vccd1 _2119_/A0 sky130_fd_sc_hd__buf_1
Xinput155 io_i_7_in1[7] vssd1 vssd1 vccd1 vccd1 _1661_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1482_ _1476_/Y _1478_/Y _1481_/Y vssd1 vssd1 vccd1 vccd1 _1482_/Y sky130_fd_sc_hd__a21boi_1
X_1620_ _2135_/X _1620_/B vssd1 vssd1 vccd1 vccd1 _1620_/X sky130_fd_sc_hd__xor2_1
X_1551_ _1539_/A _2004_/X _2119_/X vssd1 vssd1 vccd1 vccd1 _1552_/A sky130_fd_sc_hd__a21o_1
XFILLER_54_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2103_ _1766_/Y _1804_/Y _1512_/Y _1354_/Y _2254_/Q _2255_/Q vssd1 vssd1 vccd1 vccd1
+ _2103_/X sky130_fd_sc_hd__mux4_2
X_2034_ input95/X _2229_/Q _2246_/Q vssd1 vssd1 vccd1 vccd1 _2034_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1818_ _1823_/B vssd1 vssd1 vccd1 vccd1 _1850_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1749_ _2203_/Q vssd1 vssd1 vccd1 vccd1 _1749_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1465_ _1685_/B _2081_/X _1464_/X vssd1 vssd1 vccd1 vccd1 _1465_/Y sky130_fd_sc_hd__o21ai_1
X_1534_ _2125_/X _1533_/Y _1555_/S vssd1 vssd1 vccd1 vccd1 _1534_/Y sky130_fd_sc_hd__o21bai_1
X_1603_ _2133_/X _1611_/B _2000_/X vssd1 vssd1 vccd1 vccd1 _1622_/B sky130_fd_sc_hd__nand3b_4
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1396_ _1983_/X _2066_/X vssd1 vssd1 vccd1 vccd1 _1412_/A sky130_fd_sc_hd__nor2_1
X_2017_ _1783_/Y _1734_/Y _2292_/Q vssd1 vssd1 vccd1 vccd1 _2017_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1250_ _2108_/X _1229_/Y _1236_/B _1269_/C _1236_/A vssd1 vssd1 vccd1 vccd1 _1262_/A
+ sky130_fd_sc_hd__o2111ai_4
X_1181_ _2253_/Q _1175_/X _1179_/X _1180_/Y vssd1 vssd1 vccd1 vccd1 _2253_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput201 _2210_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput212 _1532_/Y vssd1 vssd1 vccd1 vccd1 io_o_4_co sky130_fd_sc_hd__clkbuf_2
Xoutput223 _2157_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput234 _2151_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput289 _1924_/X vssd1 vssd1 vccd1 vccd1 io_wo[46] sky130_fd_sc_hd__clkbuf_2
Xoutput278 _1914_/X vssd1 vssd1 vccd1 vccd1 io_wo[36] sky130_fd_sc_hd__clkbuf_2
X_1517_ _1969_/X vssd1 vssd1 vccd1 vccd1 _1522_/S sky130_fd_sc_hd__buf_2
Xoutput267 _1904_/X vssd1 vssd1 vccd1 vccd1 io_wo[26] sky130_fd_sc_hd__clkbuf_2
Xoutput256 _1894_/X vssd1 vssd1 vccd1 vccd1 io_wo[16] sky130_fd_sc_hd__clkbuf_2
Xoutput245 _2145_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_4_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1448_ _2198_/Q _1760_/A _1450_/S vssd1 vssd1 vccd1 vccd1 _2198_/D sky130_fd_sc_hd__mux2_1
X_1379_ _1971_/X _2048_/X vssd1 vssd1 vccd1 vccd1 _1436_/A sky130_fd_sc_hd__nor2_4
XFILLER_74_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2282_ _2298_/CLK _2282_/D vssd1 vssd1 vccd1 vccd1 _2282_/Q sky130_fd_sc_hd__dfxtp_1
X_1233_ _2109_/X _2022_/X vssd1 vssd1 vccd1 vccd1 _1236_/B sky130_fd_sc_hd__xnor2_4
XFILLER_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1302_ _2114_/X _2038_/X vssd1 vssd1 vccd1 vccd1 _1348_/A sky130_fd_sc_hd__xnor2_4
X_1095_ _1095_/A vssd1 vssd1 vccd1 vccd1 _1095_/X sky130_fd_sc_hd__clkbuf_2
X_1164_ _2259_/Q _1159_/X _1148_/X _1163_/Y vssd1 vssd1 vccd1 vccd1 _2259_/D sky130_fd_sc_hd__o211a_1
X_1997_ _1789_/A _1608_/X _2274_/Q vssd1 vssd1 vccd1 vccd1 _1997_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1920_ _1920_/A vssd1 vssd1 vccd1 vccd1 _1920_/X sky130_fd_sc_hd__clkbuf_2
X_1851_ _2252_/Q _1203_/C _1111_/B _2284_/Q vssd1 vssd1 vccd1 vccd1 _1851_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1782_ _1782_/A _1821_/A vssd1 vssd1 vccd1 vccd1 _1782_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1216_ _1374_/S vssd1 vssd1 vccd1 vccd1 _1216_/X sky130_fd_sc_hd__buf_2
X_2196_ _2231_/CLK _2196_/D vssd1 vssd1 vccd1 vccd1 _2196_/Q sky130_fd_sc_hd__dfxtp_1
X_2265_ _2268_/CLK _2265_/D vssd1 vssd1 vccd1 vccd1 _2265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1078_ _1110_/A vssd1 vssd1 vccd1 vccd1 _1078_/X sky130_fd_sc_hd__buf_1
XFILLER_37_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1147_ _2264_/Q _1143_/X _1135_/X _1146_/Y vssd1 vssd1 vccd1 vccd1 _2264_/D sky130_fd_sc_hd__o211a_1
XFILLER_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2050_ _1740_/Y _1432_/Y _2296_/Q vssd1 vssd1 vccd1 vccd1 _2050_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1903_ _1903_/A vssd1 vssd1 vccd1 vccd1 _1903_/X sky130_fd_sc_hd__clkbuf_2
X_1834_ _2247_/Q _1203_/C _1833_/Y vssd1 vssd1 vccd1 vccd1 _1834_/X sky130_fd_sc_hd__a21bo_1
X_1765_ _2031_/X vssd1 vssd1 vccd1 vccd1 _1765_/Y sky130_fd_sc_hd__inv_2
X_1696_ _1700_/A _1955_/X vssd1 vssd1 vccd1 vccd1 _1696_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2179_ _2254_/CLK _2179_/D vssd1 vssd1 vccd1 vccd1 _2179_/Q sky130_fd_sc_hd__dfxtp_1
X_2248_ _2251_/CLK _2248_/D vssd1 vssd1 vccd1 vccd1 _2248_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_40_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput101 io_i_1_in1[7] vssd1 vssd1 vccd1 vccd1 _2118_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput145 io_i_6_in1[6] vssd1 vssd1 vccd1 vccd1 _1711_/A sky130_fd_sc_hd__clkbuf_2
Xinput134 io_i_5_in1[4] vssd1 vssd1 vccd1 vccd1 _2129_/A0 sky130_fd_sc_hd__buf_1
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput156 io_vci vssd1 vssd1 vccd1 vccd1 _1992_/A0 sky130_fd_sc_hd__clkbuf_2
Xinput112 io_i_3_in1[0] vssd1 vssd1 vccd1 vccd1 _2073_/A0 sky130_fd_sc_hd__buf_1
Xinput123 io_i_4_in1[2] vssd1 vssd1 vccd1 vccd1 _2120_/A0 sky130_fd_sc_hd__buf_1
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1481_ _1481_/A _1801_/A vssd1 vssd1 vccd1 vccd1 _1481_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_4_9_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2295_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1550_ _2173_/Q vssd1 vssd1 vccd1 vccd1 _1550_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2102_ _1742_/Y _1808_/Y _1804_/Y _1439_/Y _2256_/Q _2257_/Q vssd1 vssd1 vccd1 vccd1
+ _2102_/X sky130_fd_sc_hd__mux4_2
X_2033_ _1763_/Y _2032_/X _2295_/Q vssd1 vssd1 vccd1 vccd1 _2033_/X sky130_fd_sc_hd__mux2_2
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1748_ _1748_/A _1767_/A vssd1 vssd1 vccd1 vccd1 _1748_/Y sky130_fd_sc_hd__nand2_1
X_1817_ _1817_/A _1845_/B _2244_/Q vssd1 vssd1 vccd1 vccd1 _1817_/Y sky130_fd_sc_hd__nand3_2
XFILLER_30_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1679_ _1685_/A _1961_/X vssd1 vssd1 vccd1 vccd1 _1679_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1602_ _2102_/X vssd1 vssd1 vccd1 vccd1 _1611_/B sky130_fd_sc_hd__inv_2
X_1395_ _1424_/B _1424_/A _1420_/A vssd1 vssd1 vccd1 vccd1 _1414_/A sky130_fd_sc_hd__nand3_4
X_1464_ _1685_/B _2081_/X _1957_/X _2078_/X vssd1 vssd1 vccd1 vccd1 _1464_/X sky130_fd_sc_hd__a211o_1
XFILLER_79_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1533_ _1536_/A _1541_/B vssd1 vssd1 vccd1 vccd1 _1533_/Y sky130_fd_sc_hd__nor2_1
X_2016_ _1784_/Y _2015_/X _2293_/Q vssd1 vssd1 vccd1 vccd1 _2016_/X sky130_fd_sc_hd__mux2_2
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1180_ _1172_/X _1180_/B _1187_/C vssd1 vssd1 vccd1 vccd1 _1180_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_17_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1516_ _1209_/X _1512_/Y _1514_/X _1515_/Y vssd1 vssd1 vccd1 vccd1 _2188_/D sky130_fd_sc_hd__o22ai_4
Xoutput268 _1905_/X vssd1 vssd1 vccd1 vccd1 io_wo[27] sky130_fd_sc_hd__clkbuf_2
Xoutput257 _1895_/X vssd1 vssd1 vccd1 vccd1 io_wo[17] sky130_fd_sc_hd__clkbuf_2
Xoutput202 _2211_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput246 _2146_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput235 _2152_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput213 _2172_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput224 _2158_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput279 _1915_/X vssd1 vssd1 vccd1 vccd1 io_wo[37] sky130_fd_sc_hd__clkbuf_2
X_1378_ _2008_/X vssd1 vssd1 vccd1 vccd1 _1378_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1447_ _2113_/X vssd1 vssd1 vccd1 vccd1 _1760_/A sky130_fd_sc_hd__inv_2
XFILLER_90_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2281_ _2295_/CLK _2281_/D vssd1 vssd1 vccd1 vccd1 _2281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1301_ _2113_/X _2036_/X vssd1 vssd1 vccd1 vccd1 _1350_/A sky130_fd_sc_hd__xnor2_4
X_1232_ _1280_/A _1280_/B _1231_/Y vssd1 vssd1 vccd1 vccd1 _1236_/A sky130_fd_sc_hd__o21bai_4
X_1094_ _2282_/Q _1077_/X _1088_/X _1093_/Y vssd1 vssd1 vccd1 vccd1 _2282_/D sky130_fd_sc_hd__o211a_1
XFILLER_64_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1163_ _1110_/X _1163_/B _1173_/C vssd1 vssd1 vccd1 vccd1 _1163_/Y sky130_fd_sc_hd__nand3b_1
X_1996_ _1695_/A _2149_/Q _2258_/Q vssd1 vssd1 vccd1 vccd1 _1996_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_11_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2297_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1850_ _1850_/A vssd1 vssd1 vccd1 vccd1 _1850_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1781_ _2215_/Q vssd1 vssd1 vccd1 vccd1 _1781_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2195_ _2195_/CLK _2195_/D vssd1 vssd1 vccd1 vccd1 _2195_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1215_ _1993_/X vssd1 vssd1 vccd1 vccd1 _1374_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_1_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1146_ _1151_/A _1194_/B vssd1 vssd1 vccd1 vccd1 _1146_/Y sky130_fd_sc_hd__nand2_1
X_2264_ _2268_/CLK _2264_/D vssd1 vssd1 vccd1 vccd1 _2264_/Q sky130_fd_sc_hd__dfxtp_1
X_1077_ _1095_/A vssd1 vssd1 vccd1 vccd1 _1077_/X sky130_fd_sc_hd__clkbuf_2
X_1979_ _1720_/Y _1978_/X _2249_/Q vssd1 vssd1 vccd1 vccd1 _1979_/X sky130_fd_sc_hd__mux2_8
XFILLER_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1902_ _1902_/A vssd1 vssd1 vccd1 vccd1 _1902_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1833_ _1823_/A _2263_/Q _1833_/C vssd1 vssd1 vccd1 vccd1 _1833_/Y sky130_fd_sc_hd__nand3b_1
X_1764_ _2197_/Q vssd1 vssd1 vccd1 vccd1 _1764_/Y sky130_fd_sc_hd__inv_2
X_1695_ _1695_/A vssd1 vssd1 vccd1 vccd1 _1695_/Y sky130_fd_sc_hd__inv_2
X_2178_ _2254_/CLK _2178_/D vssd1 vssd1 vccd1 vccd1 _2178_/Q sky130_fd_sc_hd__dfxtp_1
X_2247_ _2251_/CLK _2247_/D vssd1 vssd1 vccd1 vccd1 _2247_/Q sky130_fd_sc_hd__dfxtp_4
X_1129_ _2271_/Q _1116_/X _1122_/X _1128_/Y vssd1 vssd1 vccd1 vccd1 _2271_/D sky130_fd_sc_hd__o211a_1
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput157 io_vi vssd1 vssd1 vccd1 vccd1 _1805_/A sky130_fd_sc_hd__buf_1
XFILLER_56_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput146 io_i_6_in1[7] vssd1 vssd1 vccd1 vccd1 _1705_/A sky130_fd_sc_hd__clkbuf_2
Xinput135 io_i_5_in1[5] vssd1 vssd1 vccd1 vccd1 _2130_/A0 sky130_fd_sc_hd__buf_1
Xinput102 io_i_2_ci vssd1 vssd1 vccd1 vccd1 _1746_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput113 io_i_3_in1[1] vssd1 vssd1 vccd1 vccd1 _2076_/A0 sky130_fd_sc_hd__buf_1
Xinput124 io_i_4_in1[3] vssd1 vssd1 vccd1 vccd1 _2121_/A0 sky130_fd_sc_hd__buf_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ _1967_/X _2093_/X vssd1 vssd1 vccd1 vccd1 _1801_/A sky130_fd_sc_hd__and2_1
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2101_ _1699_/Y _1869_/Y _1808_/Y _1512_/Y _2258_/Q _2259_/Q vssd1 vssd1 vccd1 vccd1
+ _2101_/X sky130_fd_sc_hd__mux4_2
X_2032_ _1764_/Y _1757_/Y _2294_/Q vssd1 vssd1 vccd1 vccd1 _2032_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1678_ _2224_/Q vssd1 vssd1 vccd1 vccd1 _1678_/Y sky130_fd_sc_hd__inv_2
X_1816_ _1816_/A vssd1 vssd1 vccd1 vccd1 _1845_/B sky130_fd_sc_hd__buf_2
X_1747_ _2294_/Q vssd1 vssd1 vccd1 vccd1 _1767_/A sky130_fd_sc_hd__buf_2
XFILLER_26_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1532_ _1536_/A _1541_/B _2125_/X vssd1 vssd1 vccd1 vccd1 _1532_/Y sky130_fd_sc_hd__nor3b_4
X_1601_ _2136_/X vssd1 vssd1 vccd1 vccd1 _1618_/A sky130_fd_sc_hd__inv_2
X_1394_ _1399_/A _1394_/B vssd1 vssd1 vccd1 vccd1 _1420_/A sky130_fd_sc_hd__nor2_4
X_1463_ _1463_/A _1463_/B vssd1 vssd1 vccd1 vccd1 _1503_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2015_ _1785_/Y _1285_/Y _2292_/Q vssd1 vssd1 vccd1 vccd1 _2015_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1515_ _2006_/X _1455_/Y _1513_/Y _1564_/S vssd1 vssd1 vccd1 vccd1 _1515_/Y sky130_fd_sc_hd__o31ai_4
Xoutput269 _1906_/X vssd1 vssd1 vccd1 vccd1 io_wo[28] sky130_fd_sc_hd__clkbuf_2
Xoutput258 _1896_/X vssd1 vssd1 vccd1 vccd1 io_wo[18] sky130_fd_sc_hd__clkbuf_2
Xoutput247 _2147_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput236 _2153_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[5] sky130_fd_sc_hd__clkbuf_2
Xoutput225 _2159_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput203 _1802_/X vssd1 vssd1 vccd1 vccd1 io_o_3_co sky130_fd_sc_hd__clkbuf_2
Xoutput214 _2173_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[1] sky130_fd_sc_hd__clkbuf_2
X_1377_ _1971_/X _2048_/X vssd1 vssd1 vccd1 vccd1 _1377_/Y sky130_fd_sc_hd__nand2_2
XFILLER_67_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1446_ _2199_/Q _1758_/A _1450_/S vssd1 vssd1 vccd1 vccd1 _2199_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2280_ _2297_/CLK _2280_/D vssd1 vssd1 vccd1 vccd1 _2280_/Q sky130_fd_sc_hd__dfxtp_1
X_1162_ _1855_/A vssd1 vssd1 vccd1 vccd1 _1173_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_36_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1300_ _1352_/A _1352_/B _1299_/Y vssd1 vssd1 vccd1 vccd1 _1350_/B sky130_fd_sc_hd__o21bai_4
X_1231_ _2108_/X _1229_/Y _2018_/X _1782_/A vssd1 vssd1 vccd1 vccd1 _1231_/Y sky130_fd_sc_hd__o2bb2ai_1
X_1093_ _1078_/X _1105_/B _1187_/B vssd1 vssd1 vccd1 vccd1 _1093_/Y sky130_fd_sc_hd__nand3b_1
X_1995_ _1872_/Y _1994_/X _2259_/Q vssd1 vssd1 vccd1 vccd1 _1995_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1429_ _1428_/Y _2207_/Q _1431_/S vssd1 vssd1 vccd1 vccd1 _2207_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1780_ _1780_/A _1780_/B vssd1 vssd1 vccd1 vccd1 _1780_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2194_ _2195_/CLK _2194_/D vssd1 vssd1 vccd1 vccd1 _2194_/Q sky130_fd_sc_hd__dfxtp_2
X_1214_ _1214_/A _1342_/B vssd1 vssd1 vccd1 vccd1 _2239_/D sky130_fd_sc_hd__nor2b_1
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1145_ _2265_/Q _1143_/X _1135_/X _1144_/Y vssd1 vssd1 vccd1 vccd1 _2265_/D sky130_fd_sc_hd__o211a_1
X_2263_ _2268_/CLK _2263_/D vssd1 vssd1 vccd1 vccd1 _2263_/Q sky130_fd_sc_hd__dfxtp_1
X_1076_ _2287_/Q _1055_/X _1069_/X _1075_/Y vssd1 vssd1 vccd1 vccd1 _2287_/D sky130_fd_sc_hd__o211a_1
XFILLER_52_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1978_ _1722_/Y _1721_/Y _2248_/Q vssd1 vssd1 vccd1 vccd1 _1978_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1901_ _1901_/A vssd1 vssd1 vccd1 vccd1 _1901_/X sky130_fd_sc_hd__clkbuf_2
X_1832_ _1760_/B _1824_/X _2278_/Q _1825_/X _1831_/Y vssd1 vssd1 vccd1 vccd1 _1832_/X
+ sky130_fd_sc_hd__a221o_2
X_1763_ _1767_/A _1991_/X vssd1 vssd1 vccd1 vccd1 _1763_/Y sky130_fd_sc_hd__nand2_1
X_1694_ _2076_/X vssd1 vssd1 vccd1 vccd1 _1694_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2246_ _2251_/CLK _2246_/D vssd1 vssd1 vccd1 vccd1 _2246_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_65_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1059_ _1825_/A vssd1 vssd1 vccd1 vccd1 _1071_/B sky130_fd_sc_hd__clkbuf_2
X_2177_ _2254_/CLK _2177_/D vssd1 vssd1 vccd1 vccd1 _2177_/Q sky130_fd_sc_hd__dfxtp_1
X_1128_ _1138_/A _1173_/B vssd1 vssd1 vccd1 vccd1 _1128_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput136 io_i_5_in1[6] vssd1 vssd1 vccd1 vccd1 _2131_/A0 sky130_fd_sc_hd__buf_1
Xinput125 io_i_4_in1[4] vssd1 vssd1 vccd1 vccd1 _2122_/A0 sky130_fd_sc_hd__buf_1
Xinput158 io_we_i vssd1 vssd1 vccd1 vccd1 _1017_/A sky130_fd_sc_hd__buf_1
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput147 io_i_7_ci vssd1 vssd1 vccd1 vccd1 _1789_/A sky130_fd_sc_hd__clkbuf_2
Xinput103 io_i_2_in1[0] vssd1 vssd1 vccd1 vccd1 _2049_/A0 sky130_fd_sc_hd__buf_1
Xinput114 io_i_3_in1[2] vssd1 vssd1 vccd1 vccd1 _2079_/A0 sky130_fd_sc_hd__clkbuf_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2100_ _1689_/A _2150_/Q _2158_/Q _2190_/Q _2258_/Q _2259_/Q vssd1 vssd1 vccd1 vccd1
+ _2100_/X sky130_fd_sc_hd__mux4_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2031_ input94/X _2228_/Q _2246_/Q vssd1 vssd1 vccd1 vccd1 _2031_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1815_ _1829_/A vssd1 vssd1 vccd1 vccd1 _1817_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1677_ _1677_/A vssd1 vssd1 vccd1 vccd1 _1677_/Y sky130_fd_sc_hd__inv_2
X_1746_ _1746_/A vssd1 vssd1 vccd1 vccd1 _1746_/Y sky130_fd_sc_hd__inv_2
X_2229_ _2231_/CLK _2229_/D vssd1 vssd1 vccd1 vccd1 _2229_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1462_ _1959_/X _2081_/X vssd1 vssd1 vccd1 vccd1 _1463_/B sky130_fd_sc_hd__and2_1
X_1600_ _1628_/S vssd1 vssd1 vccd1 vccd1 _1616_/A sky130_fd_sc_hd__clkbuf_2
X_1531_ _1543_/B _2122_/X _2123_/X vssd1 vssd1 vccd1 vccd1 _1541_/B sky130_fd_sc_hd__nand3_4
X_1393_ _1981_/X _2063_/X vssd1 vssd1 vccd1 vccd1 _1394_/B sky130_fd_sc_hd__and2_1
X_2014_ _1786_/Y _2013_/X _2293_/Q vssd1 vssd1 vccd1 vccd1 _2014_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1729_ _1729_/A _1729_/B vssd1 vssd1 vccd1 vccd1 _1729_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1514_ _1455_/Y _1513_/Y _2006_/X vssd1 vssd1 vccd1 vccd1 _1514_/X sky130_fd_sc_hd__o21a_1
Xoutput259 _1897_/X vssd1 vssd1 vccd1 vccd1 io_wo[19] sky130_fd_sc_hd__clkbuf_2
Xoutput237 _2154_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput226 _2160_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[4] sky130_fd_sc_hd__clkbuf_2
X_1445_ _2200_/Q _1755_/A _1445_/S vssd1 vssd1 vccd1 vccd1 _2200_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput248 _1943_/X vssd1 vssd1 vccd1 vccd1 io_vco sky130_fd_sc_hd__clkbuf_2
Xoutput204 _2188_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput215 _2174_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[2] sky130_fd_sc_hd__clkbuf_2
X_1376_ _1973_/X _2051_/X vssd1 vssd1 vccd1 vccd1 _1376_/X sky130_fd_sc_hd__and2_1
XFILLER_82_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
X_1092_ _1825_/A vssd1 vssd1 vccd1 vccd1 _1105_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1161_ _1202_/A vssd1 vssd1 vccd1 vccd1 _1855_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1230_ _2107_/X vssd1 vssd1 vccd1 vccd1 _1782_/A sky130_fd_sc_hd__inv_2
X_1994_ _1659_/Y _1507_/Y _2258_/Q vssd1 vssd1 vccd1 vccd1 _1994_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1428_ _1428_/A _1428_/B vssd1 vssd1 vccd1 vccd1 _1428_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_70_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1359_ _1342_/B _1354_/Y _1356_/X _1358_/Y vssd1 vssd1 vccd1 vccd1 _2220_/D sky130_fd_sc_hd__o22ai_1
XFILLER_18_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1213_ _1987_/X vssd1 vssd1 vccd1 vccd1 _1342_/B sky130_fd_sc_hd__buf_2
X_2262_ _2268_/CLK _2262_/D vssd1 vssd1 vccd1 vccd1 _2262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2193_ _2195_/CLK _2193_/D vssd1 vssd1 vccd1 vccd1 _2193_/Q sky130_fd_sc_hd__dfxtp_2
X_1075_ _1056_/X _1090_/B _1173_/B vssd1 vssd1 vccd1 vccd1 _1075_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1144_ _1151_/A _1191_/B vssd1 vssd1 vccd1 vccd1 _1144_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1977_ _1726_/Y _1976_/X _2249_/Q vssd1 vssd1 vccd1 vccd1 _1977_/X sky130_fd_sc_hd__mux2_2
XFILLER_20_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1900_ _1900_/A vssd1 vssd1 vccd1 vccd1 _1900_/X sky130_fd_sc_hd__clkbuf_2
X_1831_ _1769_/Y _1814_/Y _1830_/Y vssd1 vssd1 vccd1 vccd1 _1831_/Y sky130_fd_sc_hd__o21ai_1
X_1693_ _2166_/Q vssd1 vssd1 vccd1 vccd1 _1693_/Y sky130_fd_sc_hd__inv_2
X_1762_ _2034_/X vssd1 vssd1 vccd1 vccd1 _1762_/Y sky130_fd_sc_hd__inv_2
X_2245_ _2251_/CLK _2245_/D vssd1 vssd1 vccd1 vccd1 _2245_/Q sky130_fd_sc_hd__dfxtp_4
X_2176_ _2254_/CLK _2176_/D vssd1 vssd1 vccd1 vccd1 _2176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1058_ _1858_/A vssd1 vssd1 vccd1 vccd1 _1825_/A sky130_fd_sc_hd__buf_1
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1127_ _1140_/A vssd1 vssd1 vccd1 vccd1 _1138_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput126 io_i_4_in1[5] vssd1 vssd1 vccd1 vccd1 _2123_/A0 sky130_fd_sc_hd__buf_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput104 io_i_2_in1[1] vssd1 vssd1 vccd1 vccd1 _2052_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput115 io_i_3_in1[3] vssd1 vssd1 vccd1 vccd1 _2082_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput159 wb_rst_i vssd1 vssd1 vccd1 vccd1 _1219_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput137 io_i_5_in1[7] vssd1 vssd1 vccd1 vccd1 _2132_/A0 sky130_fd_sc_hd__buf_1
Xinput148 io_i_7_in1[0] vssd1 vssd1 vccd1 vccd1 _1699_/A sky130_fd_sc_hd__buf_1
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2030_ _1767_/Y _2029_/X _2295_/Q vssd1 vssd1 vccd1 vccd1 _2030_/X sky130_fd_sc_hd__mux2_2
XFILLER_62_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1814_ _1829_/A _1833_/C vssd1 vssd1 vccd1 vccd1 _1814_/Y sky130_fd_sc_hd__nand2_2
XFILLER_30_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1745_ _2264_/Q vssd1 vssd1 vccd1 vccd1 _1745_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1676_ _2085_/X vssd1 vssd1 vccd1 vccd1 _1676_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2228_ _2231_/CLK _2228_/D vssd1 vssd1 vccd1 vccd1 _2228_/Q sky130_fd_sc_hd__dfxtp_2
X_2159_ _2272_/CLK _2159_/D vssd1 vssd1 vccd1 vccd1 _2159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1392_ _1981_/X _2063_/X vssd1 vssd1 vccd1 vccd1 _1399_/A sky130_fd_sc_hd__nor2_4
X_1461_ _1685_/B _2081_/X vssd1 vssd1 vccd1 vccd1 _1463_/A sky130_fd_sc_hd__nor2_1
X_1530_ _1530_/A _2120_/X _2121_/X _2119_/X vssd1 vssd1 vccd1 vccd1 _1543_/B sky130_fd_sc_hd__and4_2
XFILLER_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2013_ _1787_/Y _1291_/Y _2292_/Q vssd1 vssd1 vccd1 vccd1 _2013_/X sky130_fd_sc_hd__mux2_1
X_1728_ _2231_/Q vssd1 vssd1 vccd1 vccd1 _1728_/Y sky130_fd_sc_hd__inv_2
X_1659_ _2157_/Q vssd1 vssd1 vccd1 vccd1 _1659_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_8_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2292_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput205 _2189_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput216 _2175_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[3] sky130_fd_sc_hd__clkbuf_2
X_1513_ _1513_/A vssd1 vssd1 vccd1 vccd1 _1513_/Y sky130_fd_sc_hd__inv_2
X_1375_ _2211_/Q vssd1 vssd1 vccd1 vccd1 _1375_/Y sky130_fd_sc_hd__inv_2
Xoutput249 _1878_/X vssd1 vssd1 vccd1 vccd1 io_wo[0] sky130_fd_sc_hd__clkbuf_2
Xoutput238 _2155_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput227 _2161_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[5] sky130_fd_sc_hd__clkbuf_2
X_1444_ _2201_/Q _1752_/A _1445_/S vssd1 vssd1 vccd1 vccd1 _2201_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1091_ _2283_/Q _1077_/X _1088_/X _1090_/Y vssd1 vssd1 vccd1 vccd1 _2283_/D sky130_fd_sc_hd__o211a_1
XFILLER_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1160_ input2/X input1/X vssd1 vssd1 vccd1 vccd1 _1202_/A sky130_fd_sc_hd__nor2_1
X_1993_ _1807_/Y _1992_/X _2277_/Q vssd1 vssd1 vccd1 vccd1 _1993_/X sky130_fd_sc_hd__mux2_2
XFILLER_87_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1427_ _1430_/B _1430_/A _1426_/Y vssd1 vssd1 vccd1 vccd1 _1428_/B sky130_fd_sc_hd__a21oi_1
XFILLER_55_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1358_ _2010_/X _1296_/Y _1355_/Y _1450_/S vssd1 vssd1 vccd1 vccd1 _1358_/Y sky130_fd_sc_hd__o31ai_1
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1289_ _1287_/Y _1223_/X _1288_/Y vssd1 vssd1 vccd1 vccd1 _1289_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1212_ _1214_/A _1211_/X vssd1 vssd1 vccd1 vccd1 _2240_/D sky130_fd_sc_hd__nor2b_1
X_2192_ _2291_/CLK _2192_/D vssd1 vssd1 vccd1 vccd1 _2192_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2261_ _2268_/CLK _2261_/D vssd1 vssd1 vccd1 vccd1 _2261_/Q sky130_fd_sc_hd__dfxtp_1
X_1074_ input6/X vssd1 vssd1 vccd1 vccd1 _1173_/B sky130_fd_sc_hd__inv_2
XFILLER_1_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1143_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1143_/X sky130_fd_sc_hd__clkbuf_2
X_1976_ _1728_/Y _1727_/Y _2248_/Q vssd1 vssd1 vccd1 vccd1 _1976_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1830_ _1849_/A _1845_/B _2246_/Q vssd1 vssd1 vccd1 vccd1 _1830_/Y sky130_fd_sc_hd__nand3_1
X_1761_ _2198_/Q vssd1 vssd1 vccd1 vccd1 _1761_/Y sky130_fd_sc_hd__inv_2
X_1692_ _2190_/Q vssd1 vssd1 vccd1 vccd1 _1692_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_10_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2219_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2244_ _2251_/CLK _2244_/D vssd1 vssd1 vccd1 vccd1 _2244_/Q sky130_fd_sc_hd__dfxtp_4
X_2175_ _2272_/CLK _2175_/D vssd1 vssd1 vccd1 vccd1 _2175_/Q sky130_fd_sc_hd__dfxtp_1
X_1126_ _2272_/Q _1116_/X _1122_/X _1125_/Y vssd1 vssd1 vccd1 vccd1 _2272_/D sky130_fd_sc_hd__o211a_1
X_1057_ _1823_/B input2/X vssd1 vssd1 vccd1 vccd1 _1858_/A sky130_fd_sc_hd__and2b_1
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1959_ _1682_/Y _1958_/X _2251_/Q vssd1 vssd1 vccd1 vccd1 _1959_/X sky130_fd_sc_hd__mux2_2
Xinput127 io_i_4_in1[6] vssd1 vssd1 vccd1 vccd1 _2124_/A0 sky130_fd_sc_hd__buf_1
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput138 io_i_6_ci vssd1 vssd1 vccd1 vccd1 _1999_/A0 sky130_fd_sc_hd__buf_1
Xinput149 io_i_7_in1[1] vssd1 vssd1 vccd1 vccd1 _1695_/A sky130_fd_sc_hd__clkbuf_2
Xinput105 io_i_2_in1[2] vssd1 vssd1 vccd1 vccd1 _2055_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput116 io_i_3_in1[4] vssd1 vssd1 vccd1 vccd1 _2085_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_72_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1744_ _2180_/Q vssd1 vssd1 vccd1 vccd1 _1744_/Y sky130_fd_sc_hd__inv_2
X_1813_ _1813_/A vssd1 vssd1 vccd1 vccd1 _1813_/Y sky130_fd_sc_hd__inv_2
X_1675_ _2169_/Q vssd1 vssd1 vccd1 vccd1 _1675_/Y sky130_fd_sc_hd__inv_2
X_2089_ _1670_/Y _1488_/Y _2298_/Q vssd1 vssd1 vccd1 vccd1 _2089_/X sky130_fd_sc_hd__mux2_1
X_1109_ _2277_/Q _1095_/X _1104_/X _1108_/Y vssd1 vssd1 vccd1 vccd1 _2277_/D sky130_fd_sc_hd__o211a_1
X_2227_ _2292_/CLK _2227_/D vssd1 vssd1 vccd1 vccd1 _2227_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2158_ _2275_/CLK _2158_/D vssd1 vssd1 vccd1 vccd1 _2158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1391_ _1979_/X _2060_/X vssd1 vssd1 vccd1 vccd1 _1424_/A sky130_fd_sc_hd__xor2_4
X_1460_ _1959_/X vssd1 vssd1 vccd1 vccd1 _1685_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2012_ _1788_/Y _2011_/X _2261_/Q vssd1 vssd1 vccd1 vccd1 _2012_/X sky130_fd_sc_hd__mux2_2
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1727_ _1727_/A vssd1 vssd1 vccd1 vccd1 _1727_/Y sky130_fd_sc_hd__inv_2
X_1658_ _1658_/A vssd1 vssd1 vccd1 vccd1 _1658_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1589_ _1207_/X _2159_/Q vssd1 vssd1 vccd1 vccd1 _1589_/X sky130_fd_sc_hd__and2b_1
XFILLER_85_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput228 _2162_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput217 _2176_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput239 _1637_/X vssd1 vssd1 vccd1 vccd1 io_o_7_co sky130_fd_sc_hd__clkbuf_2
X_1512_ _2188_/Q vssd1 vssd1 vccd1 vccd1 _1512_/Y sky130_fd_sc_hd__clkinv_4
Xoutput206 _2190_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_67_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1443_ _2202_/Q _1750_/A _1445_/S vssd1 vssd1 vccd1 vccd1 _2202_/D sky130_fd_sc_hd__mux2_1
X_1374_ _2212_/Q _1786_/A _1374_/S vssd1 vssd1 vccd1 vccd1 _2212_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1090_ _1078_/X _1090_/B _1876_/C vssd1 vssd1 vccd1 vccd1 _1090_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1992_ _1992_/A0 _2237_/Q _2276_/Q vssd1 vssd1 vccd1 vccd1 _1992_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1426_ _1975_/X _2054_/X vssd1 vssd1 vccd1 vccd1 _1426_/Y sky130_fd_sc_hd__nor2_1
X_1357_ _1987_/X vssd1 vssd1 vccd1 vccd1 _1450_/S sky130_fd_sc_hd__buf_2
X_1288_ _2012_/X vssd1 vssd1 vccd1 vccd1 _1288_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2191_ _2195_/CLK _2191_/D vssd1 vssd1 vccd1 vccd1 _2191_/Q sky130_fd_sc_hd__dfxtp_4
X_1211_ _1969_/X vssd1 vssd1 vccd1 vccd1 _1211_/X sky130_fd_sc_hd__clkbuf_2
X_1142_ _2266_/Q _1130_/X _1135_/X _1141_/Y vssd1 vssd1 vccd1 vccd1 _2266_/D sky130_fd_sc_hd__o211a_1
X_2260_ _2268_/CLK _2260_/D vssd1 vssd1 vccd1 vccd1 _2260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1073_ _1825_/A vssd1 vssd1 vccd1 vccd1 _1090_/B sky130_fd_sc_hd__buf_1
XFILLER_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1975_ _1732_/Y _1974_/X _2249_/Q vssd1 vssd1 vccd1 vccd1 _1975_/X sky130_fd_sc_hd__mux2_4
X_1409_ _1406_/Y _1407_/X _1417_/A vssd1 vssd1 vccd1 vccd1 _1409_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1691_ _1700_/A _1957_/X vssd1 vssd1 vccd1 vccd1 _1691_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1760_ _1760_/A _1760_/B vssd1 vssd1 vccd1 vccd1 _1760_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2243_ _2291_/CLK _2243_/D vssd1 vssd1 vccd1 vccd1 _2243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1125_ _1125_/A _1170_/B vssd1 vssd1 vccd1 vccd1 _1125_/Y sky130_fd_sc_hd__nand2_1
X_2174_ _2272_/CLK _2174_/D vssd1 vssd1 vccd1 vccd1 _2174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1056_ _1110_/A vssd1 vssd1 vccd1 vccd1 _1056_/X sky130_fd_sc_hd__buf_1
X_1889_ _1889_/A vssd1 vssd1 vccd1 vccd1 _1889_/X sky130_fd_sc_hd__clkbuf_2
X_1958_ _1684_/Y _1683_/Y _2250_/Q vssd1 vssd1 vccd1 vccd1 _1958_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput128 io_i_4_in1[7] vssd1 vssd1 vccd1 vccd1 _2125_/A0 sky130_fd_sc_hd__buf_1
Xinput117 io_i_3_in1[5] vssd1 vssd1 vccd1 vccd1 _2088_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput139 io_i_6_in1[0] vssd1 vssd1 vccd1 vccd1 _1742_/A sky130_fd_sc_hd__buf_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput106 io_i_2_in1[3] vssd1 vssd1 vccd1 vccd1 _2058_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1743_ _1743_/A _1971_/X vssd1 vssd1 vccd1 vccd1 _1743_/Y sky130_fd_sc_hd__nand2_1
X_1674_ _2193_/Q vssd1 vssd1 vccd1 vccd1 _1674_/Y sky130_fd_sc_hd__inv_2
X_1812_ _1812_/A vssd1 vssd1 vccd1 vccd1 _1812_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2226_ _2226_/CLK _2226_/D vssd1 vssd1 vccd1 vccd1 _2226_/Q sky130_fd_sc_hd__dfxtp_2
X_1039_ _2294_/Q vssd1 vssd1 vccd1 vccd1 _1760_/B sky130_fd_sc_hd__buf_2
X_1108_ _1096_/X _1111_/B _1200_/B vssd1 vssd1 vccd1 vccd1 _1108_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2088_ _2088_/A0 _2209_/Q _2250_/Q vssd1 vssd1 vccd1 vccd1 _2088_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2157_ _2275_/CLK _2157_/D vssd1 vssd1 vccd1 vccd1 _2157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1390_ _1430_/B _1430_/A _1428_/A _1389_/Y vssd1 vssd1 vccd1 vccd1 _1424_/B sky130_fd_sc_hd__a31o_2
XFILLER_79_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2011_ _1790_/Y _1789_/Y _2260_/Q vssd1 vssd1 vccd1 vccd1 _2011_/X sky130_fd_sc_hd__mux2_1
X_1726_ _2058_/X vssd1 vssd1 vccd1 vccd1 _1726_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1657_ _1656_/Y _2140_/Q _1657_/S vssd1 vssd1 vccd1 vccd1 _2140_/D sky130_fd_sc_hd__mux2_1
X_1588_ _1579_/A _1579_/B _2127_/X _1597_/B _2128_/X vssd1 vssd1 vccd1 vccd1 _1588_/X
+ sky130_fd_sc_hd__a41o_1
X_2209_ _2219_/CLK _2209_/D vssd1 vssd1 vccd1 vccd1 _2209_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1511_ _1209_/X _1507_/Y _1508_/X _1510_/Y vssd1 vssd1 vccd1 vccd1 _2189_/D sky130_fd_sc_hd__o22ai_1
X_1442_ _2203_/Q _1748_/A _1445_/S vssd1 vssd1 vccd1 vccd1 _2203_/D sky130_fd_sc_hd__mux2_1
Xoutput229 _2163_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput218 _2177_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_4_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput207 _2191_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1373_ _2105_/X vssd1 vssd1 vccd1 vccd1 _1786_/A sky130_fd_sc_hd__inv_2
XFILLER_4_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1709_ _2187_/Q vssd1 vssd1 vccd1 vccd1 _1709_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1991_ _1762_/Y _1990_/X _2247_/Q vssd1 vssd1 vccd1 vccd1 _1991_/X sky130_fd_sc_hd__mux2_2
XFILLER_13_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1425_ _1424_/X _2208_/Q _1431_/S vssd1 vssd1 vccd1 vccd1 _2208_/D sky130_fd_sc_hd__mux2_1
X_1356_ _1296_/Y _1355_/Y _2010_/X vssd1 vssd1 vccd1 vccd1 _1356_/X sky130_fd_sc_hd__o21a_1
X_1287_ _1287_/A vssd1 vssd1 vccd1 vccd1 _1287_/Y sky130_fd_sc_hd__inv_2
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2190_ _2195_/CLK _2190_/D vssd1 vssd1 vccd1 vccd1 _2190_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_77_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1210_ _1214_/A _1209_/X vssd1 vssd1 vccd1 vccd1 _2241_/D sky130_fd_sc_hd__nor2b_1
X_1072_ _2288_/Q _1055_/X _1069_/X _1071_/Y vssd1 vssd1 vccd1 vccd1 _2288_/D sky130_fd_sc_hd__o211a_1
XFILLER_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1141_ _1151_/A _1187_/B vssd1 vssd1 vccd1 vccd1 _1141_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1974_ _1734_/Y _1733_/Y _2248_/Q vssd1 vssd1 vccd1 vccd1 _1974_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1408_ _1969_/X vssd1 vssd1 vccd1 vccd1 _1417_/A sky130_fd_sc_hd__inv_2
XFILLER_29_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1339_ _2225_/Q vssd1 vssd1 vccd1 vccd1 _1339_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1690_ _2222_/Q vssd1 vssd1 vccd1 vccd1 _1690_/Y sky130_fd_sc_hd__inv_2
X_2242_ _2299_/CLK _2242_/D vssd1 vssd1 vccd1 vccd1 _2242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1055_ _1095_/A vssd1 vssd1 vccd1 vccd1 _1055_/X sky130_fd_sc_hd__clkbuf_2
X_1124_ _2273_/Q _1116_/X _1122_/X _1123_/Y vssd1 vssd1 vccd1 vccd1 _2273_/D sky130_fd_sc_hd__o211a_1
X_2173_ _2272_/CLK _2173_/D vssd1 vssd1 vccd1 vccd1 _2173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1957_ _1688_/Y _1956_/X _2251_/Q vssd1 vssd1 vccd1 vccd1 _1957_/X sky130_fd_sc_hd__mux2_8
X_1888_ _1888_/A vssd1 vssd1 vccd1 vccd1 _1888_/X sky130_fd_sc_hd__clkbuf_2
Xinput118 io_i_3_in1[6] vssd1 vssd1 vccd1 vccd1 _2091_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput129 io_i_5_ci vssd1 vssd1 vccd1 vccd1 _2001_/A0 sky130_fd_sc_hd__buf_1
Xinput107 io_i_2_in1[4] vssd1 vssd1 vccd1 vccd1 _2061_/A0 sky130_fd_sc_hd__clkbuf_1
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1811_ _1811_/A vssd1 vssd1 vccd1 vccd1 _1811_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1673_ _1685_/A _1963_/X vssd1 vssd1 vccd1 vccd1 _1673_/Y sky130_fd_sc_hd__nand2_1
X_1742_ _1742_/A vssd1 vssd1 vccd1 vccd1 _1742_/Y sky130_fd_sc_hd__inv_2
X_2225_ _2226_/CLK _2225_/D vssd1 vssd1 vccd1 vccd1 _2225_/Q sky130_fd_sc_hd__dfxtp_2
X_2087_ _1673_/Y _2086_/X _2299_/Q vssd1 vssd1 vccd1 vccd1 _2087_/X sky130_fd_sc_hd__mux2_2
X_1038_ _2295_/Q _1020_/X _1023_/X _1037_/Y vssd1 vssd1 vccd1 vccd1 _2295_/D sky130_fd_sc_hd__o211a_1
X_1107_ _1858_/A vssd1 vssd1 vccd1 vccd1 _1111_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_53_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2156_ _2275_/CLK _2156_/D vssd1 vssd1 vccd1 vccd1 _2156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2010_ _1769_/Y _2009_/X _2263_/Q vssd1 vssd1 vccd1 vccd1 _2010_/X sky130_fd_sc_hd__mux2_2
X_1725_ _2184_/Q vssd1 vssd1 vccd1 vccd1 _1725_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1587_ _1581_/A _1585_/Y _1583_/B _1586_/Y vssd1 vssd1 vccd1 vccd1 _2160_/D sky130_fd_sc_hd__o31ai_1
X_1656_ _2101_/X _1998_/X vssd1 vssd1 vccd1 vccd1 _1656_/Y sky130_fd_sc_hd__xnor2_1
X_2208_ _2219_/CLK _2208_/D vssd1 vssd1 vccd1 vccd1 _2208_/Q sky130_fd_sc_hd__dfxtp_4
X_2139_ _1705_/A _2163_/Q _2179_/Q _2211_/Q _2256_/Q _2257_/Q vssd1 vssd1 vccd1 vccd1
+ _2139_/X sky130_fd_sc_hd__mux4_2
XFILLER_34_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1510_ _1457_/Y _1452_/X _1456_/Y _1564_/S vssd1 vssd1 vccd1 vccd1 _1510_/Y sky130_fd_sc_hd__o31ai_1
X_1441_ _2118_/X vssd1 vssd1 vccd1 vccd1 _1748_/A sky130_fd_sc_hd__inv_2
Xoutput219 _2178_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput208 _2192_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1372_ _2213_/Q _1784_/A _1372_/S vssd1 vssd1 vccd1 vccd1 _2213_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1708_ _1729_/A _1985_/X vssd1 vssd1 vccd1 vccd1 _1708_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1639_ _2095_/X _1638_/X _1657_/S vssd1 vssd1 vccd1 vccd1 _1639_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_64_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1990_ _1695_/Y _1754_/Y _2246_/Q vssd1 vssd1 vccd1 vccd1 _1990_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1424_ _1424_/A _1424_/B vssd1 vssd1 vccd1 vccd1 _1424_/X sky130_fd_sc_hd__xor2_1
XFILLER_87_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_7_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2163_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1355_ _1355_/A vssd1 vssd1 vccd1 vccd1 _1355_/Y sky130_fd_sc_hd__inv_2
X_1286_ _1283_/X _1284_/Y _1216_/X _1285_/Y vssd1 vssd1 vccd1 vccd1 _2229_/D sky130_fd_sc_hd__o2bb2ai_1
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1071_ _1056_/X _1071_/B _1170_/B vssd1 vssd1 vccd1 vccd1 _1071_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_52_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1140_ _1140_/A vssd1 vssd1 vccd1 vccd1 _1151_/A sky130_fd_sc_hd__clkbuf_2
X_1973_ _1738_/Y _1972_/X _2249_/Q vssd1 vssd1 vccd1 vccd1 _1973_/X sky130_fd_sc_hd__mux2_4
X_1407_ _1799_/A _1405_/A _1402_/Y _1400_/Y vssd1 vssd1 vccd1 vccd1 _1407_/X sky130_fd_sc_hd__o211a_1
X_1338_ _1335_/X _1342_/B _1337_/Y vssd1 vssd1 vccd1 vccd1 _2226_/D sky130_fd_sc_hd__a21oi_1
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1269_ _1239_/A _1269_/B _1269_/C vssd1 vssd1 vccd1 vccd1 _1269_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2241_ _2298_/CLK _2241_/D vssd1 vssd1 vccd1 vccd1 _2241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2172_ _2272_/CLK _2172_/D vssd1 vssd1 vccd1 vccd1 _2172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1054_ _1833_/C _1829_/A _1158_/C vssd1 vssd1 vccd1 vccd1 _1095_/A sky130_fd_sc_hd__nor3_4
X_1123_ _1125_/A _1168_/B vssd1 vssd1 vccd1 vccd1 _1123_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1887_ _1887_/A vssd1 vssd1 vccd1 vccd1 _1887_/X sky130_fd_sc_hd__clkbuf_2
X_1956_ _1690_/Y _1689_/Y _2250_/Q vssd1 vssd1 vccd1 vccd1 _1956_/X sky130_fd_sc_hd__mux2_1
Xinput108 io_i_2_in1[5] vssd1 vssd1 vccd1 vccd1 _2064_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput119 io_i_3_in1[7] vssd1 vssd1 vccd1 vccd1 _2094_/A0 sky130_fd_sc_hd__clkbuf_1
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1810_ _1871_/A _2278_/Q vssd1 vssd1 vccd1 vccd1 _1810_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1741_ _2049_/X vssd1 vssd1 vccd1 vccd1 _1741_/Y sky130_fd_sc_hd__inv_2
X_1672_ _1672_/A vssd1 vssd1 vccd1 vccd1 _1672_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1106_ _2278_/Q _1095_/X _1104_/X _1105_/Y vssd1 vssd1 vccd1 vccd1 _2278_/D sky130_fd_sc_hd__o211a_1
X_2155_ _2163_/CLK _2155_/D vssd1 vssd1 vccd1 vccd1 _2155_/Q sky130_fd_sc_hd__dfxtp_1
X_2224_ _2226_/CLK _2224_/D vssd1 vssd1 vccd1 vccd1 _2224_/Q sky130_fd_sc_hd__dfxtp_2
X_2086_ _1675_/Y _1674_/Y _2298_/Q vssd1 vssd1 vccd1 vccd1 _2086_/X sky130_fd_sc_hd__mux2_1
X_1037_ _1049_/A _1196_/B vssd1 vssd1 vccd1 vccd1 _1037_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1939_ _1939_/A vssd1 vssd1 vccd1 vccd1 _1939_/X sky130_fd_sc_hd__clkbuf_2
Xinput90 io_i_0_in1[5] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1724_ _2208_/Q vssd1 vssd1 vccd1 vccd1 _1724_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1586_ _1598_/S _2160_/Q vssd1 vssd1 vccd1 vccd1 _1586_/Y sky130_fd_sc_hd__nand2_1
X_1655_ _1647_/S _2141_/Q _1654_/Y vssd1 vssd1 vccd1 vccd1 _2141_/D sky130_fd_sc_hd__a21bo_1
X_2207_ _2297_/CLK _2207_/D vssd1 vssd1 vccd1 vccd1 _2207_/Q sky130_fd_sc_hd__dfxtp_4
X_2069_ _1708_/Y _2068_/X _2297_/Q vssd1 vssd1 vccd1 vccd1 _2069_/X sky130_fd_sc_hd__mux2_2
XFILLER_53_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2138_ _1711_/A _2162_/Q _2178_/Q _2210_/Q _2256_/Q _2257_/Q vssd1 vssd1 vccd1 vccd1
+ _2138_/X sky130_fd_sc_hd__mux4_2
XFILLER_78_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1440_ _1437_/X _1438_/Y _1211_/X _1439_/Y vssd1 vssd1 vccd1 vccd1 _2204_/D sky130_fd_sc_hd__o2bb2ai_2
XFILLER_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput209 _2193_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[5] sky130_fd_sc_hd__clkbuf_2
X_1371_ _2214_/Q _1782_/A _1372_/S vssd1 vssd1 vccd1 vccd1 _2214_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1707_ _2296_/Q vssd1 vssd1 vccd1 vccd1 _1729_/A sky130_fd_sc_hd__clkbuf_2
X_1638_ _1644_/B _2097_/X _2096_/X vssd1 vssd1 vccd1 vccd1 _1638_/X sky130_fd_sc_hd__and3_1
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1569_ _1579_/A _1579_/B _2002_/X vssd1 vssd1 vccd1 vccd1 _1569_/Y sky130_fd_sc_hd__nand3_2
XFILLER_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1423_ _1431_/S _1420_/X _1422_/X vssd1 vssd1 vccd1 vccd1 _2209_/D sky130_fd_sc_hd__o21bai_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1354_ _2220_/Q vssd1 vssd1 vccd1 vccd1 _1354_/Y sky130_fd_sc_hd__inv_2
X_1285_ _2229_/Q vssd1 vssd1 vccd1 vccd1 _1285_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1070_ input7/X vssd1 vssd1 vccd1 vccd1 _1170_/B sky130_fd_sc_hd__inv_2
XFILLER_81_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1972_ _1285_/Y _1658_/Y _2248_/Q vssd1 vssd1 vccd1 vccd1 _1972_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1406_ _1400_/Y _1402_/Y _1405_/Y vssd1 vssd1 vccd1 vccd1 _1406_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1268_ _1239_/A _1267_/Y _1269_/C vssd1 vssd1 vccd1 vccd1 _1268_/Y sky130_fd_sc_hd__o21bai_1
X_1337_ _1445_/S _2226_/Q vssd1 vssd1 vccd1 vccd1 _1337_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1199_ _2246_/Q _1189_/X _1193_/X _1198_/Y vssd1 vssd1 vccd1 vccd1 _2246_/D sky130_fd_sc_hd__o211a_1
XPHY_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2171_ _2195_/CLK _2171_/D vssd1 vssd1 vccd1 vccd1 _2171_/Q sky130_fd_sc_hd__dfxtp_1
X_2240_ _2298_/CLK _2240_/D vssd1 vssd1 vccd1 vccd1 _2240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1122_ _1165_/A vssd1 vssd1 vccd1 vccd1 _1122_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1053_ _1186_/A vssd1 vssd1 vccd1 vccd1 _1158_/C sky130_fd_sc_hd__buf_2
XFILLER_18_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1886_ _1886_/A vssd1 vssd1 vccd1 vccd1 _1886_/X sky130_fd_sc_hd__clkbuf_2
X_1955_ _1694_/Y _1954_/X _2251_/Q vssd1 vssd1 vccd1 vccd1 _1955_/X sky130_fd_sc_hd__mux2_4
Xinput109 io_i_2_in1[6] vssd1 vssd1 vccd1 vccd1 _2067_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_71_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1740_ _2181_/Q vssd1 vssd1 vccd1 vccd1 _1740_/Y sky130_fd_sc_hd__inv_2
X_1671_ _2088_/X vssd1 vssd1 vccd1 vccd1 _1671_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1105_ _1096_/X _1105_/B _1198_/B vssd1 vssd1 vccd1 vccd1 _1105_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2154_ _2163_/CLK _2154_/D vssd1 vssd1 vccd1 vccd1 _2154_/Q sky130_fd_sc_hd__dfxtp_1
X_2085_ _2085_/A0 _2208_/Q _2250_/Q vssd1 vssd1 vccd1 vccd1 _2085_/X sky130_fd_sc_hd__mux2_1
X_2223_ _2231_/CLK _2223_/D vssd1 vssd1 vccd1 vccd1 _2223_/Q sky130_fd_sc_hd__dfxtp_2
X_1036_ _1036_/A vssd1 vssd1 vccd1 vccd1 _1196_/B sky130_fd_sc_hd__inv_2
XFILLER_21_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1938_ _1938_/A vssd1 vssd1 vccd1 vccd1 _1938_/X sky130_fd_sc_hd__clkbuf_2
Xinput80 io_eo[6] vssd1 vssd1 vccd1 vccd1 _1884_/A sky130_fd_sc_hd__clkbuf_1
Xinput91 io_i_0_in1[6] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__clkbuf_1
X_1869_ _2148_/Q vssd1 vssd1 vccd1 vccd1 _1869_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1723_ _1729_/A _1979_/X vssd1 vssd1 vccd1 vccd1 _1723_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1654_ _1654_/A _1943_/X _1654_/C vssd1 vssd1 vccd1 vccd1 _1654_/Y sky130_fd_sc_hd__nand3_1
X_2206_ _2297_/CLK _2206_/D vssd1 vssd1 vccd1 vccd1 _2206_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1585_ _1579_/X _2128_/X _2129_/X vssd1 vssd1 vccd1 vccd1 _1585_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2068_ _1709_/Y _1375_/Y _2296_/Q vssd1 vssd1 vccd1 vccd1 _2068_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_1019_ _1019_/A _1110_/A vssd1 vssd1 vccd1 vccd1 _1032_/A sky130_fd_sc_hd__nor2_1
X_2137_ _1716_/A _2161_/Q _2177_/Q _2209_/Q _2256_/Q _2257_/Q vssd1 vssd1 vccd1 vccd1
+ _2137_/X sky130_fd_sc_hd__mux4_2
XFILLER_34_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1370_ _2215_/Q _1780_/A _1372_/S vssd1 vssd1 vccd1 vccd1 _2215_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1706_ _2235_/Q vssd1 vssd1 vccd1 vccd1 _1706_/Y sky130_fd_sc_hd__inv_2
X_1637_ _1637_/A vssd1 vssd1 vccd1 vccd1 _1637_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1499_ _1499_/A _1499_/B vssd1 vssd1 vccd1 vccd1 _1499_/X sky130_fd_sc_hd__xor2_1
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1568_ _2126_/X vssd1 vssd1 vccd1 vccd1 _1579_/B sky130_fd_sc_hd__inv_2
XFILLER_81_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1422_ _1525_/S _2209_/Q vssd1 vssd1 vccd1 vccd1 _1422_/X sky130_fd_sc_hd__and2b_1
X_1353_ _1352_/X _2221_/Q _1353_/S vssd1 vssd1 vccd1 vccd1 _2221_/D sky130_fd_sc_hd__mux2_1
X_1284_ _1224_/Y _1282_/Y _1226_/Y _1281_/S vssd1 vssd1 vccd1 vccd1 _1284_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1971_ _1741_/Y _1970_/X _2249_/Q vssd1 vssd1 vccd1 vccd1 _1971_/X sky130_fd_sc_hd__mux2_4
X_1405_ _1405_/A _1799_/A vssd1 vssd1 vccd1 vccd1 _1405_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1267_ _1269_/B vssd1 vssd1 vccd1 vccd1 _1267_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1198_ _1186_/X _1198_/B _1200_/C vssd1 vssd1 vccd1 vccd1 _1198_/Y sky130_fd_sc_hd__nand3b_1
X_1336_ _1987_/X vssd1 vssd1 vccd1 vccd1 _1445_/S sky130_fd_sc_hd__buf_2
Xinput1 io_adr_i[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
XFILLER_61_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE3_0 _1913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2170_ _2195_/CLK _2170_/D vssd1 vssd1 vccd1 vccd1 _2170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1052_ input2/X vssd1 vssd1 vccd1 vccd1 _1829_/A sky130_fd_sc_hd__inv_2
X_1121_ _2274_/Q _1116_/X _1104_/X _1120_/Y vssd1 vssd1 vccd1 vccd1 _2274_/D sky130_fd_sc_hd__o211a_1
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1954_ _1757_/Y _1695_/Y _2250_/Q vssd1 vssd1 vccd1 vccd1 _1954_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1885_ _1885_/A vssd1 vssd1 vccd1 vccd1 _1885_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2299_ _2299_/CLK _2299_/D vssd1 vssd1 vccd1 vccd1 _2299_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1319_ _1327_/B _1319_/B _1333_/B vssd1 vssd1 vccd1 vccd1 _1319_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_24_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput190 _2224_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[4] sky130_fd_sc_hd__clkbuf_2
XPHY_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1670_ _2170_/Q vssd1 vssd1 vccd1 vccd1 _1670_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_2222_ _2231_/CLK _2222_/D vssd1 vssd1 vccd1 vccd1 _2222_/Q sky130_fd_sc_hd__dfxtp_2
X_2084_ _1679_/Y _2083_/X _2299_/Q vssd1 vssd1 vccd1 vccd1 _2084_/X sky130_fd_sc_hd__mux2_4
X_1035_ _1743_/A _1020_/X _1023_/X _1034_/Y vssd1 vssd1 vccd1 vccd1 _2296_/D sky130_fd_sc_hd__o211a_1
XFILLER_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2153_ _2163_/CLK _2153_/D vssd1 vssd1 vccd1 vccd1 _2153_/Q sky130_fd_sc_hd__dfxtp_1
X_1104_ _1165_/A vssd1 vssd1 vccd1 vccd1 _1104_/X sky130_fd_sc_hd__clkbuf_4
X_1937_ _1937_/A vssd1 vssd1 vccd1 vccd1 _1937_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput70 io_eo[55] vssd1 vssd1 vccd1 vccd1 _1933_/A sky130_fd_sc_hd__clkbuf_1
X_1799_ _1799_/A vssd1 vssd1 vccd1 vccd1 _1799_/Y sky130_fd_sc_hd__inv_2
X_1868_ _2275_/Q _1817_/A _1821_/C _1867_/X vssd1 vssd1 vccd1 vccd1 _1868_/X sky130_fd_sc_hd__a31o_1
Xinput81 io_eo[7] vssd1 vssd1 vccd1 vccd1 _1885_/A sky130_fd_sc_hd__clkbuf_1
Xinput92 io_i_0_in1[7] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1722_ _2232_/Q vssd1 vssd1 vccd1 vccd1 _1722_/Y sky130_fd_sc_hd__inv_2
X_1584_ _1583_/X _2161_/Q _1598_/S vssd1 vssd1 vccd1 vccd1 _2161_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1653_ _1633_/B _1998_/X _1995_/X vssd1 vssd1 vccd1 vccd1 _1654_/A sky130_fd_sc_hd__a21bo_1
X_2205_ _2298_/CLK _2205_/D vssd1 vssd1 vccd1 vccd1 _2205_/Q sky130_fd_sc_hd__dfxtp_4
X_1018_ _1186_/A vssd1 vssd1 vccd1 vccd1 _1110_/A sky130_fd_sc_hd__clkbuf_2
X_2067_ _2067_/A0 _2226_/Q _2248_/Q vssd1 vssd1 vccd1 vccd1 _2067_/X sky130_fd_sc_hd__mux2_1
X_2136_ _1721_/A _2160_/Q _2176_/Q _2208_/Q _2256_/Q _2257_/Q vssd1 vssd1 vccd1 vccd1
+ _2136_/X sky130_fd_sc_hd__mux4_2
XFILLER_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1705_ _1705_/A vssd1 vssd1 vccd1 vccd1 _1705_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1636_ _1644_/B _2097_/X _2096_/X _2095_/X vssd1 vssd1 vccd1 vccd1 _1637_/A sky130_fd_sc_hd__and4_1
X_1567_ _2103_/X vssd1 vssd1 vccd1 vccd1 _1579_/A sky130_fd_sc_hd__inv_2
X_1498_ _1506_/S _1496_/X _1497_/X vssd1 vssd1 vccd1 vccd1 _2193_/D sky130_fd_sc_hd__o21bai_1
XFILLER_73_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2119_ _2119_/A0 _2189_/Q _2205_/Q _2229_/Q _2252_/Q _2253_/Q vssd1 vssd1 vccd1 vccd1
+ _2119_/X sky130_fd_sc_hd__mux4_2
XFILLER_81_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1421_ _1969_/X vssd1 vssd1 vccd1 vccd1 _1525_/S sky130_fd_sc_hd__clkbuf_2
X_1352_ _1352_/A _1352_/B vssd1 vssd1 vccd1 vccd1 _1352_/X sky130_fd_sc_hd__xor2_1
X_1283_ _1282_/Y _1226_/Y _1224_/Y vssd1 vssd1 vccd1 vccd1 _1283_/X sky130_fd_sc_hd__a21o_1
XFILLER_63_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1619_ _1618_/X _2152_/Q _1628_/S vssd1 vssd1 vccd1 vccd1 _2152_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1970_ _1291_/Y _1742_/Y _2248_/Q vssd1 vssd1 vccd1 vccd1 _1970_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1404_ _1985_/X _2069_/X vssd1 vssd1 vccd1 vccd1 _1799_/A sky130_fd_sc_hd__and2_1
X_1335_ _1335_/A _1335_/B vssd1 vssd1 vccd1 vccd1 _1335_/X sky130_fd_sc_hd__xor2_1
XFILLER_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1266_ _2233_/Q vssd1 vssd1 vccd1 vccd1 _1266_/Y sky130_fd_sc_hd__inv_2
X_1197_ _2247_/Q _1189_/X _1193_/X _1196_/Y vssd1 vssd1 vccd1 vccd1 _2247_/D sky130_fd_sc_hd__o211a_1
XFILLER_28_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput2 io_adr_i[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_51_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2254_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1051_ _1823_/B vssd1 vssd1 vccd1 vccd1 _1833_/C sky130_fd_sc_hd__clkbuf_4
X_1120_ _1125_/A _1166_/B vssd1 vssd1 vccd1 vccd1 _1120_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1884_ _1884_/A vssd1 vssd1 vccd1 vccd1 _1884_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1953_ _1698_/Y _1952_/X _2251_/Q vssd1 vssd1 vccd1 vccd1 _1953_/X sky130_fd_sc_hd__mux2_4
X_2298_ _2298_/CLK _2298_/D vssd1 vssd1 vccd1 vccd1 _2298_/Q sky130_fd_sc_hd__dfxtp_4
X_1318_ _1750_/A _2044_/X vssd1 vssd1 vccd1 vccd1 _1333_/B sky130_fd_sc_hd__nand2_2
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1249_ _2110_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _1269_/C sky130_fd_sc_hd__xnor2_2
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput191 _2225_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[5] sky130_fd_sc_hd__clkbuf_2
Xoutput180 _2231_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2152_ _2163_/CLK _2152_/D vssd1 vssd1 vccd1 vccd1 _2152_/Q sky130_fd_sc_hd__dfxtp_1
X_2221_ _2231_/CLK _2221_/D vssd1 vssd1 vccd1 vccd1 _2221_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2083_ _1681_/Y _1680_/Y _2298_/Q vssd1 vssd1 vccd1 vccd1 _2083_/X sky130_fd_sc_hd__mux2_1
X_1034_ _1049_/A _1194_/B vssd1 vssd1 vccd1 vccd1 _1034_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1103_ _1193_/A vssd1 vssd1 vccd1 vccd1 _1165_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1936_ _1936_/A vssd1 vssd1 vccd1 vccd1 _1936_/X sky130_fd_sc_hd__clkbuf_2
X_1867_ _2259_/Q _1855_/A _1858_/X _2291_/Q vssd1 vssd1 vccd1 vccd1 _1867_/X sky130_fd_sc_hd__a22o_1
Xinput71 io_eo[56] vssd1 vssd1 vccd1 vccd1 _1934_/A sky130_fd_sc_hd__clkbuf_1
Xinput60 io_eo[46] vssd1 vssd1 vccd1 vccd1 _1924_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput82 io_eo[8] vssd1 vssd1 vccd1 vccd1 _1886_/A sky130_fd_sc_hd__clkbuf_1
X_1798_ _1319_/B _1796_/Y _1333_/B _1797_/X vssd1 vssd1 vccd1 vccd1 _1812_/A sky130_fd_sc_hd__a31oi_4
Xinput93 io_i_1_ci vssd1 vssd1 vccd1 vccd1 _1770_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _1721_/A vssd1 vssd1 vccd1 vccd1 _1721_/Y sky130_fd_sc_hd__inv_2
X_1583_ _2130_/X _1583_/B vssd1 vssd1 vccd1 vccd1 _1583_/X sky130_fd_sc_hd__xor2_1
X_1652_ _1651_/Y _2142_/Q _1657_/S vssd1 vssd1 vccd1 vccd1 _2142_/D sky130_fd_sc_hd__mux2_1
X_2204_ _2251_/CLK _2204_/D vssd1 vssd1 vccd1 vccd1 _2204_/Q sky130_fd_sc_hd__dfxtp_2
X_2135_ _1727_/A _2159_/Q _2175_/Q _2207_/Q _2256_/Q _2257_/Q vssd1 vssd1 vccd1 vccd1
+ _2135_/X sky130_fd_sc_hd__mux4_2
X_2066_ _1713_/Y _2065_/X _2297_/Q vssd1 vssd1 vccd1 vccd1 _2066_/X sky130_fd_sc_hd__mux2_1
X_1017_ _1017_/A input3/X vssd1 vssd1 vccd1 vccd1 _1186_/A sky130_fd_sc_hd__nand2_4
XFILLER_19_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1919_ _1919_/A vssd1 vssd1 vccd1 vccd1 _1919_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1704_ _2070_/X vssd1 vssd1 vccd1 vccd1 _1704_/Y sky130_fd_sc_hd__inv_2
X_1497_ _1951_/X _2193_/Q vssd1 vssd1 vccd1 vccd1 _1497_/X sky130_fd_sc_hd__and2b_1
XFILLER_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1566_ _1575_/A vssd1 vssd1 vccd1 vccd1 _1581_/A sky130_fd_sc_hd__clkbuf_2
X_1635_ _1646_/A _1646_/B vssd1 vssd1 vccd1 vccd1 _1644_/B sky130_fd_sc_hd__nor2_2
XFILLER_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2118_ _2118_/A0 _2235_/Q _1661_/A _2132_/A0 _2246_/Q _2247_/Q vssd1 vssd1 vccd1
+ vccd1 _2118_/X sky130_fd_sc_hd__mux4_2
X_2049_ _2049_/A0 _2220_/Q _2248_/Q vssd1 vssd1 vccd1 vccd1 _2049_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1420_ _1420_/A _1420_/B vssd1 vssd1 vccd1 vccd1 _1420_/X sky130_fd_sc_hd__xor2_1
XFILLER_79_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1351_ _1350_/X _2222_/Q _1353_/S vssd1 vssd1 vccd1 vccd1 _2222_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1282_ _1282_/A vssd1 vssd1 vccd1 vccd1 _1282_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1618_ _1618_/A _1618_/B vssd1 vssd1 vccd1 vccd1 _1618_/X sky130_fd_sc_hd__xor2_1
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1549_ _1548_/Y _2174_/Q _1555_/S vssd1 vssd1 vccd1 vccd1 _2174_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1403_ _1985_/X _2069_/X vssd1 vssd1 vccd1 vccd1 _1405_/A sky130_fd_sc_hd__nor2_4
X_1265_ _1263_/Y _1216_/X _1264_/Y vssd1 vssd1 vccd1 vccd1 _2234_/D sky130_fd_sc_hd__a21oi_1
X_1334_ _1334_/A _1334_/B vssd1 vssd1 vccd1 vccd1 _1335_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1196_ _1186_/X _1196_/B _1200_/C vssd1 vssd1 vccd1 vccd1 _1196_/Y sky130_fd_sc_hd__nand3b_1
Xinput3 io_cs_i vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_1
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1050_ _1821_/A _1029_/A _1043_/X _1049_/Y vssd1 vssd1 vccd1 vccd1 _2292_/D sky130_fd_sc_hd__o211a_1
X_1883_ _1883_/A vssd1 vssd1 vccd1 vccd1 _1883_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1952_ _1354_/Y _1699_/Y _2250_/Q vssd1 vssd1 vccd1 vccd1 _1952_/X sky130_fd_sc_hd__mux2_1
X_2297_ _2297_/CLK _2297_/D vssd1 vssd1 vccd1 vccd1 _2297_/Q sky130_fd_sc_hd__dfxtp_4
X_1248_ _1248_/A _1248_/B _1252_/B vssd1 vssd1 vccd1 vccd1 _1254_/A sky130_fd_sc_hd__nand3_1
XFILLER_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1317_ _2117_/X vssd1 vssd1 vccd1 vccd1 _1750_/A sky130_fd_sc_hd__inv_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1179_ _1193_/A vssd1 vssd1 vccd1 vccd1 _1179_/X sky130_fd_sc_hd__clkbuf_2
Xoutput170 _1838_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[4] sky130_fd_sc_hd__clkbuf_2
Xoutput192 _2226_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput181 _2232_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1102_ _2279_/Q _1095_/X _1088_/X _1101_/Y vssd1 vssd1 vccd1 vccd1 _2279_/D sky130_fd_sc_hd__o211a_1
X_2151_ _2275_/CLK _2151_/D vssd1 vssd1 vccd1 vccd1 _2151_/Q sky130_fd_sc_hd__dfxtp_1
X_2220_ _2268_/CLK _2220_/D vssd1 vssd1 vccd1 vccd1 _2220_/Q sky130_fd_sc_hd__dfxtp_1
X_2082_ _2082_/A0 _2207_/Q _2250_/Q vssd1 vssd1 vccd1 vccd1 _2082_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1033_ _1033_/A vssd1 vssd1 vccd1 vccd1 _1194_/B sky130_fd_sc_hd__inv_2
X_1935_ _1935_/A vssd1 vssd1 vccd1 vccd1 _1935_/X sky130_fd_sc_hd__clkbuf_2
Xinput72 io_eo[57] vssd1 vssd1 vccd1 vccd1 _1935_/A sky130_fd_sc_hd__clkbuf_1
Xinput61 io_eo[47] vssd1 vssd1 vccd1 vccd1 _1925_/A sky130_fd_sc_hd__clkbuf_1
Xinput50 io_eo[37] vssd1 vssd1 vccd1 vccd1 _1915_/A sky130_fd_sc_hd__clkbuf_1
X_1866_ _2274_/Q _1817_/A _1821_/C _1865_/X vssd1 vssd1 vccd1 vccd1 _1866_/X sky130_fd_sc_hd__a31o_1
X_1797_ _2046_/X _2118_/X vssd1 vssd1 vccd1 vccd1 _1797_/X sky130_fd_sc_hd__and2b_1
XFILLER_88_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput83 io_eo[9] vssd1 vssd1 vccd1 vccd1 _1887_/A sky130_fd_sc_hd__clkbuf_1
Xinput94 io_i_1_in1[0] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1720_ _2061_/X vssd1 vssd1 vccd1 vccd1 _1720_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1651_ _2100_/X _1654_/C vssd1 vssd1 vccd1 vccd1 _1651_/Y sky130_fd_sc_hd__xnor2_1
X_1582_ _1581_/A _1580_/Y _1574_/X _1581_/Y vssd1 vssd1 vccd1 vccd1 _2162_/D sky130_fd_sc_hd__o31ai_1
XFILLER_85_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2065_ _1714_/Y _1411_/Y _2296_/Q vssd1 vssd1 vccd1 vccd1 _2065_/X sky130_fd_sc_hd__mux2_1
X_2203_ _2292_/CLK _2203_/D vssd1 vssd1 vccd1 vccd1 _2203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2134_ _1733_/A _2158_/Q _2174_/Q _2206_/Q _2256_/Q _2257_/Q vssd1 vssd1 vccd1 vccd1
+ _2134_/X sky130_fd_sc_hd__mux4_2
X_1016_ _1823_/A _1823_/B vssd1 vssd1 vccd1 vccd1 _1019_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1918_ _1918_/A vssd1 vssd1 vccd1 vccd1 _1918_/X sky130_fd_sc_hd__clkbuf_2
X_1849_ _1849_/A vssd1 vssd1 vccd1 vccd1 _1849_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1703_ _1703_/A vssd1 vssd1 vccd1 vccd1 _1703_/Y sky130_fd_sc_hd__inv_2
XPHY_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1634_ _1654_/C _2100_/X _2099_/X vssd1 vssd1 vccd1 vccd1 _1646_/B sky130_fd_sc_hd__nand3b_4
X_1496_ _1496_/A _1496_/B vssd1 vssd1 vccd1 vccd1 _1496_/X sky130_fd_sc_hd__xor2_1
X_1565_ _1947_/X vssd1 vssd1 vccd1 vccd1 _1575_/A sky130_fd_sc_hd__inv_2
X_2048_ _1743_/Y _2047_/X _2297_/Q vssd1 vssd1 vccd1 vccd1 _2048_/X sky130_fd_sc_hd__mux2_2
X_2117_ _2117_/A0 _2234_/Q _1667_/A _2131_/A0 _2246_/Q _2247_/Q vssd1 vssd1 vccd1
+ vccd1 _2117_/X sky130_fd_sc_hd__mux4_2
XFILLER_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_1350_ _1350_/A _1350_/B vssd1 vssd1 vccd1 vccd1 _1350_/X sky130_fd_sc_hd__xor2_1
X_1281_ _1280_/X _2230_/Q _1281_/S vssd1 vssd1 vccd1 vccd1 _2230_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1617_ _1616_/A _1615_/Y _1613_/B _1616_/Y vssd1 vssd1 vccd1 vccd1 _2153_/D sky130_fd_sc_hd__o31ai_1
XFILLER_5_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1479_ _1967_/X _2093_/X vssd1 vssd1 vccd1 vccd1 _1481_/A sky130_fd_sc_hd__nor2_2
XFILLER_75_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1548_ _2120_/X _1552_/C vssd1 vssd1 vccd1 vccd1 _1548_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1402_ _1412_/B vssd1 vssd1 vccd1 vccd1 _1402_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1264_ _1363_/S _2234_/Q vssd1 vssd1 vccd1 vccd1 _1264_/Y sky130_fd_sc_hd__nor2_1
X_1333_ _1333_/A _1333_/B vssd1 vssd1 vccd1 vccd1 _1335_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 io_dat_i[0] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1195_ _2248_/Q _1189_/X _1193_/X _1194_/Y vssd1 vssd1 vccd1 vccd1 _2248_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1951_ _1871_/Y _1950_/X _2283_/Q vssd1 vssd1 vccd1 vccd1 _1951_/X sky130_fd_sc_hd__mux2_2
X_1882_ _1882_/A vssd1 vssd1 vccd1 vccd1 _1882_/X sky130_fd_sc_hd__clkbuf_2
X_2296_ _2297_/CLK _2296_/D vssd1 vssd1 vccd1 vccd1 _2296_/Q sky130_fd_sc_hd__dfxtp_4
X_1247_ _2026_/X _2111_/X vssd1 vssd1 vccd1 vccd1 _1252_/B sky130_fd_sc_hd__or2b_2
XFILLER_56_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1316_ _1334_/A _1333_/A _1334_/B vssd1 vssd1 vccd1 vccd1 _1319_/B sky130_fd_sc_hd__nand3_4
X_1178_ _2254_/Q _1175_/X _1165_/X _1177_/Y vssd1 vssd1 vccd1 vccd1 _2254_/D sky130_fd_sc_hd__o211a_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput171 _1841_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[5] sky130_fd_sc_hd__clkbuf_2
Xoutput160 _1822_/Y vssd1 vssd1 vccd1 vccd1 io_dat_o[0] sky130_fd_sc_hd__clkbuf_2
Xoutput193 _2227_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput182 _2233_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[5] sky130_fd_sc_hd__clkbuf_2
XPHY_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2081_ _1685_/Y _2080_/X _2299_/Q vssd1 vssd1 vccd1 vccd1 _2081_/X sky130_fd_sc_hd__mux2_2
XFILLER_87_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1101_ _1096_/X _1105_/B _1196_/B vssd1 vssd1 vccd1 vccd1 _1101_/Y sky130_fd_sc_hd__nand3b_1
X_1032_ _1032_/A vssd1 vssd1 vccd1 vccd1 _1049_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2150_ _2275_/CLK _2150_/D vssd1 vssd1 vccd1 vccd1 _2150_/Q sky130_fd_sc_hd__dfxtp_1
X_1934_ _1934_/A vssd1 vssd1 vccd1 vccd1 _1934_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput73 io_eo[58] vssd1 vssd1 vccd1 vccd1 _1936_/A sky130_fd_sc_hd__clkbuf_1
Xinput62 io_eo[48] vssd1 vssd1 vccd1 vccd1 _1926_/A sky130_fd_sc_hd__clkbuf_1
Xinput51 io_eo[38] vssd1 vssd1 vccd1 vccd1 _1916_/A sky130_fd_sc_hd__clkbuf_1
Xinput40 io_eo[28] vssd1 vssd1 vccd1 vccd1 _1906_/A sky130_fd_sc_hd__clkbuf_1
X_1865_ _2258_/Q _1855_/X _1858_/X _2290_/Q vssd1 vssd1 vccd1 vccd1 _1865_/X sky130_fd_sc_hd__a22o_1
X_1796_ _1796_/A vssd1 vssd1 vccd1 vccd1 _1796_/Y sky130_fd_sc_hd__inv_2
Xinput84 io_i_0_ci vssd1 vssd1 vccd1 vccd1 _1790_/A sky130_fd_sc_hd__clkbuf_1
Xinput95 io_i_1_in1[1] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_1
X_2279_ _2297_/CLK _2279_/D vssd1 vssd1 vccd1 vccd1 _2279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1581_ _1581_/A _2162_/Q vssd1 vssd1 vccd1 vccd1 _1581_/Y sky130_fd_sc_hd__nand2_1
X_1650_ _1649_/X _2143_/Q _1657_/S vssd1 vssd1 vccd1 vccd1 _2143_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2202_ _2292_/CLK _2202_/D vssd1 vssd1 vccd1 vccd1 _2202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1015_ input1/X vssd1 vssd1 vccd1 vccd1 _1823_/B sky130_fd_sc_hd__buf_1
X_2064_ _2064_/A0 _2225_/Q _2248_/Q vssd1 vssd1 vccd1 vccd1 _2064_/X sky130_fd_sc_hd__mux2_1
X_2133_ _1658_/Y _1659_/Y _1550_/Y _1432_/Y _2256_/Q _2257_/Q vssd1 vssd1 vccd1 vccd1
+ _2133_/X sky130_fd_sc_hd__mux4_2
X_1917_ _1917_/A vssd1 vssd1 vccd1 vccd1 _1917_/X sky130_fd_sc_hd__clkbuf_2
X_1779_ _2216_/Q vssd1 vssd1 vccd1 vccd1 _1779_/Y sky130_fd_sc_hd__inv_2
X_1848_ _2299_/Q _1876_/B _2283_/Q _1071_/B _1847_/Y vssd1 vssd1 vccd1 vccd1 _1848_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1564_ _2164_/Q _1953_/X _1564_/S vssd1 vssd1 vccd1 vccd1 _2164_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1702_ _2266_/Q vssd1 vssd1 vccd1 vccd1 _1702_/Y sky130_fd_sc_hd__inv_2
X_1633_ _1995_/X _1633_/B _1998_/X vssd1 vssd1 vccd1 vccd1 _1654_/C sky130_fd_sc_hd__nand3b_4
X_1495_ _1499_/B _1499_/A _1494_/Y vssd1 vssd1 vccd1 vccd1 _1496_/B sky130_fd_sc_hd__a21oi_1
XFILLER_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2047_ _1744_/Y _1439_/Y _2296_/Q vssd1 vssd1 vccd1 vccd1 _2047_/X sky130_fd_sc_hd__mux2_1
X_2116_ input99/X _2233_/Q _1672_/A _2130_/A0 _2246_/Q _2247_/Q vssd1 vssd1 vccd1
+ vccd1 _2116_/X sky130_fd_sc_hd__mux4_2
XFILLER_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1280_ _1280_/A _1280_/B vssd1 vssd1 vccd1 vccd1 _1280_/X sky130_fd_sc_hd__xor2_1
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1616_ _1616_/A _2153_/Q vssd1 vssd1 vccd1 vccd1 _1616_/Y sky130_fd_sc_hd__nand2_1
X_1547_ _2104_/X _2004_/X _2119_/X vssd1 vssd1 vccd1 vccd1 _1552_/C sky130_fd_sc_hd__nand3b_2
X_1478_ _1489_/B vssd1 vssd1 vccd1 vccd1 _1478_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1401_ _1983_/X _2066_/X vssd1 vssd1 vccd1 vccd1 _1412_/B sky130_fd_sc_hd__and2_1
XFILLER_5_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1263_ _1263_/A _1263_/B vssd1 vssd1 vccd1 vccd1 _1263_/Y sky130_fd_sc_hd__xnor2_1
X_1332_ _1332_/A _1332_/B vssd1 vssd1 vccd1 vccd1 _2227_/D sky130_fd_sc_hd__nand2_1
X_1194_ _1186_/X _1194_/B _1200_/C vssd1 vssd1 vccd1 vccd1 _1194_/Y sky130_fd_sc_hd__nand3b_1
Xinput5 io_dat_i[10] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1950_ _1969_/X _2240_/Q _2282_/Q vssd1 vssd1 vccd1 vccd1 _1950_/X sky130_fd_sc_hd__mux2_1
X_1881_ _1881_/A vssd1 vssd1 vccd1 vccd1 _1881_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1315_ _1326_/C _1313_/X _1314_/X vssd1 vssd1 vccd1 vccd1 _1334_/B sky130_fd_sc_hd__a21oi_4
X_1246_ _2112_/X _2028_/X vssd1 vssd1 vccd1 vccd1 _1248_/B sky130_fd_sc_hd__xnor2_1
XFILLER_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2295_ _2295_/CLK _2295_/D vssd1 vssd1 vccd1 vccd1 _2295_/Q sky130_fd_sc_hd__dfxtp_4
X_1177_ _1172_/X _1177_/B _1187_/C vssd1 vssd1 vccd1 vccd1 _1177_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_2_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput161 _1857_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[10] sky130_fd_sc_hd__clkbuf_2
Xoutput172 _1844_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[6] sky130_fd_sc_hd__clkbuf_2
Xoutput183 _2234_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput194 _1811_/Y vssd1 vssd1 vccd1 vccd1 io_o_2_co sky130_fd_sc_hd__clkbuf_2
XPHY_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2080_ _1687_/Y _1686_/Y _2298_/Q vssd1 vssd1 vccd1 vccd1 _2080_/X sky130_fd_sc_hd__mux2_1
X_1031_ _2296_/Q vssd1 vssd1 vccd1 vccd1 _1743_/A sky130_fd_sc_hd__clkbuf_2
X_1100_ _2280_/Q _1095_/X _1088_/X _1099_/Y vssd1 vssd1 vccd1 vccd1 _2280_/D sky130_fd_sc_hd__o211a_1
X_1933_ _1933_/A vssd1 vssd1 vccd1 vccd1 _1933_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput74 io_eo[59] vssd1 vssd1 vccd1 vccd1 _1937_/A sky130_fd_sc_hd__clkbuf_1
Xinput63 io_eo[49] vssd1 vssd1 vccd1 vccd1 _1927_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput52 io_eo[39] vssd1 vssd1 vccd1 vccd1 _1917_/A sky130_fd_sc_hd__clkbuf_1
Xinput41 io_eo[29] vssd1 vssd1 vccd1 vccd1 _1907_/A sky130_fd_sc_hd__clkbuf_1
Xinput30 io_eo[19] vssd1 vssd1 vccd1 vccd1 _1897_/A sky130_fd_sc_hd__clkbuf_1
X_1864_ _2273_/Q _1817_/A _1821_/C _1863_/X vssd1 vssd1 vccd1 vccd1 _1864_/X sky130_fd_sc_hd__a31o_1
X_1795_ _2118_/X _2046_/X vssd1 vssd1 vccd1 vccd1 _1796_/A sky130_fd_sc_hd__and2b_1
Xinput85 io_i_0_in1[0] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__clkbuf_1
Xinput96 io_i_1_in1[2] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_5_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2275_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2278_ _2295_/CLK _2278_/D vssd1 vssd1 vccd1 vccd1 _2278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1229_ _2020_/X vssd1 vssd1 vccd1 vccd1 _1229_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1580_ _2129_/X _1579_/X _2130_/X _2128_/X _2131_/X vssd1 vssd1 vccd1 vccd1 _1580_/Y
+ sky130_fd_sc_hd__a41oi_2
XFILLER_11_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2132_ _2132_/A0 _2179_/Q _2195_/Q _2227_/Q _2254_/Q _2255_/Q vssd1 vssd1 vccd1 vccd1
+ _2132_/X sky130_fd_sc_hd__mux4_2
X_2201_ _2226_/CLK _2201_/D vssd1 vssd1 vccd1 vccd1 _2201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2063_ _1717_/Y _2062_/X _2297_/Q vssd1 vssd1 vccd1 vccd1 _2063_/X sky130_fd_sc_hd__mux2_2
X_1014_ input2/X vssd1 vssd1 vccd1 vccd1 _1823_/A sky130_fd_sc_hd__buf_1
XFILLER_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1916_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1916_/X sky130_fd_sc_hd__clkbuf_2
X_1847_ _1847_/A _1847_/B vssd1 vssd1 vccd1 vccd1 _1847_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1778_ _1778_/A _1780_/B vssd1 vssd1 vccd1 vccd1 _1778_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1701_ _2164_/Q vssd1 vssd1 vccd1 vccd1 _1701_/Y sky130_fd_sc_hd__inv_2
XPHY_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1563_ _2165_/Q _1955_/X _1564_/S vssd1 vssd1 vccd1 vccd1 _2165_/D sky130_fd_sc_hd__mux2_1
X_1494_ _1961_/X _2084_/X vssd1 vssd1 vccd1 vccd1 _1494_/Y sky130_fd_sc_hd__nor2_1
X_1632_ _2101_/X vssd1 vssd1 vccd1 vccd1 _1633_/B sky130_fd_sc_hd__inv_2
XFILLER_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2115_ input98/X _2232_/Q _1677_/A _2129_/A0 _2246_/Q _2247_/Q vssd1 vssd1 vccd1
+ vccd1 _2115_/X sky130_fd_sc_hd__mux4_2
X_2046_ _1748_/Y _2045_/X _2295_/Q vssd1 vssd1 vccd1 vccd1 _2046_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1477_ _1965_/X _2090_/X vssd1 vssd1 vccd1 vccd1 _1489_/B sky130_fd_sc_hd__and2_1
X_1615_ _1620_/B _2135_/X _2136_/X _2137_/X vssd1 vssd1 vccd1 vccd1 _1615_/Y sky130_fd_sc_hd__a31oi_1
X_1546_ _1545_/X _2175_/Q _1546_/S vssd1 vssd1 vccd1 vccd1 _2175_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2029_ _1768_/Y _1354_/Y _2294_/Q vssd1 vssd1 vccd1 vccd1 _2029_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1400_ _1414_/A _1400_/B _1414_/B vssd1 vssd1 vccd1 vccd1 _1400_/Y sky130_fd_sc_hd__nand3_4
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1331_ _1353_/S _2227_/Q vssd1 vssd1 vccd1 vccd1 _1332_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1262_ _1262_/A _1262_/B vssd1 vssd1 vccd1 vccd1 _1263_/B sky130_fd_sc_hd__nand2_1
X_1193_ _1193_/A vssd1 vssd1 vccd1 vccd1 _1193_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 io_dat_i[11] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput310 _1885_/X vssd1 vssd1 vccd1 vccd1 io_wo[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_10_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1529_ _2104_/X _2004_/X vssd1 vssd1 vccd1 vccd1 _1530_/A sky130_fd_sc_hd__and2b_1
XFILLER_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1880_ _1880_/A vssd1 vssd1 vccd1 vccd1 _1880_/X sky130_fd_sc_hd__clkbuf_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2294_ _2295_/CLK _2294_/D vssd1 vssd1 vccd1 vccd1 _2294_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1314_ _2042_/X _2116_/X vssd1 vssd1 vccd1 vccd1 _1314_/X sky130_fd_sc_hd__and2b_1
X_1245_ _1245_/A _1253_/C _1245_/C vssd1 vssd1 vccd1 vccd1 _1248_/A sky130_fd_sc_hd__nand3_1
XFILLER_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1176_ _1855_/A vssd1 vssd1 vccd1 vccd1 _1187_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput162 _1860_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[11] sky130_fd_sc_hd__clkbuf_2
Xoutput173 _1848_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[7] sky130_fd_sc_hd__clkbuf_2
Xoutput184 _2235_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput195 _2204_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_21_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1030_ _2297_/Q _1020_/X _1023_/X _1029_/Y vssd1 vssd1 vccd1 vccd1 _2297_/D sky130_fd_sc_hd__o211a_1
XFILLER_46_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1932_ _1932_/A vssd1 vssd1 vccd1 vccd1 _1932_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1863_ _2257_/Q _1855_/X _1858_/X _2289_/Q vssd1 vssd1 vccd1 vccd1 _1863_/X sky130_fd_sc_hd__a22o_1
Xinput20 io_eo[0] vssd1 vssd1 vccd1 vccd1 _1878_/A sky130_fd_sc_hd__clkbuf_1
Xinput31 io_eo[1] vssd1 vssd1 vccd1 vccd1 _1879_/A sky130_fd_sc_hd__clkbuf_1
X_1794_ _1253_/B _1792_/Y _1253_/C _1793_/X vssd1 vssd1 vccd1 vccd1 _1813_/A sky130_fd_sc_hd__a31oi_4
Xinput53 io_eo[3] vssd1 vssd1 vccd1 vccd1 _1881_/A sky130_fd_sc_hd__clkbuf_1
Xinput75 io_eo[5] vssd1 vssd1 vccd1 vccd1 _1883_/A sky130_fd_sc_hd__clkbuf_1
Xinput42 io_eo[2] vssd1 vssd1 vccd1 vccd1 _1880_/A sky130_fd_sc_hd__clkbuf_1
Xinput64 io_eo[4] vssd1 vssd1 vccd1 vccd1 _1882_/A sky130_fd_sc_hd__clkbuf_1
Xinput86 io_i_0_in1[1] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__clkbuf_1
Xinput97 io_i_1_in1[3] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_1
X_2277_ _2295_/CLK _2277_/D vssd1 vssd1 vccd1 vccd1 _2277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1228_ _1224_/Y _1226_/Y _1282_/A vssd1 vssd1 vccd1 vccd1 _1280_/B sky130_fd_sc_hd__a21oi_4
X_1159_ _1189_/A vssd1 vssd1 vccd1 vccd1 _1159_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2062_ _1719_/Y _1718_/Y _2296_/Q vssd1 vssd1 vccd1 vccd1 _2062_/X sky130_fd_sc_hd__mux2_1
X_2131_ _2131_/A0 _2178_/Q _2194_/Q _2226_/Q _2254_/Q _2255_/Q vssd1 vssd1 vccd1 vccd1
+ _2131_/X sky130_fd_sc_hd__mux4_2
X_2200_ _2226_/CLK _2200_/D vssd1 vssd1 vccd1 vccd1 _2200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1013_ _2298_/Q vssd1 vssd1 vccd1 vccd1 _1700_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1777_ _2217_/Q vssd1 vssd1 vccd1 vccd1 _1777_/Y sky130_fd_sc_hd__inv_2
X_1915_ _1915_/A vssd1 vssd1 vccd1 vccd1 _1915_/X sky130_fd_sc_hd__clkbuf_2
X_1846_ _1839_/A _2267_/Q _1850_/A vssd1 vssd1 vccd1 vccd1 _1847_/B sky130_fd_sc_hd__nand3b_1
XFILLER_84_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1700_ _1700_/A _1953_/X vssd1 vssd1 vccd1 vccd1 _1700_/Y sky130_fd_sc_hd__nand2_1
X_1631_ _2098_/X vssd1 vssd1 vccd1 vccd1 _1646_/A sky130_fd_sc_hd__inv_2
XPHY_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1562_ _2166_/Q _1957_/X _1564_/S vssd1 vssd1 vccd1 vccd1 _2166_/D sky130_fd_sc_hd__mux2_1
X_1493_ _1209_/X _1488_/Y _1492_/Y vssd1 vssd1 vccd1 vccd1 _2194_/D sky130_fd_sc_hd__o21ai_1
XFILLER_66_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2045_ _1749_/Y _1662_/Y _2294_/Q vssd1 vssd1 vccd1 vccd1 _2045_/X sky130_fd_sc_hd__mux2_1
X_2114_ input97/X _2231_/Q _1683_/A _2128_/A0 _2246_/Q _2247_/Q vssd1 vssd1 vccd1
+ vccd1 _2114_/X sky130_fd_sc_hd__mux4_2
XFILLER_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1829_ _1829_/A vssd1 vssd1 vccd1 vccd1 _1849_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1614_ _1613_/X _2154_/Q _1616_/A vssd1 vssd1 vccd1 vccd1 _2154_/D sky130_fd_sc_hd__mux2_1
XFILLER_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1476_ _1491_/A _1476_/B _1491_/B vssd1 vssd1 vccd1 vccd1 _1476_/Y sky130_fd_sc_hd__nand3_2
X_1545_ _2121_/X _1545_/B vssd1 vssd1 vccd1 vccd1 _1545_/X sky130_fd_sc_hd__xor2_1
X_2028_ _1772_/Y _2027_/X _2293_/Q vssd1 vssd1 vccd1 vccd1 _2028_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1261_ _2111_/X _2026_/X vssd1 vssd1 vccd1 vccd1 _1263_/A sky130_fd_sc_hd__xnor2_1
XFILLER_68_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1330_ _1330_/A vssd1 vssd1 vccd1 vccd1 _1353_/S sky130_fd_sc_hd__buf_2
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1192_ _2249_/Q _1189_/X _1179_/X _1191_/Y vssd1 vssd1 vccd1 vccd1 _2249_/D sky130_fd_sc_hd__o211a_1
Xinput7 io_dat_i[12] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput300 _1934_/X vssd1 vssd1 vccd1 vccd1 io_wo[56] sky130_fd_sc_hd__clkbuf_2
Xoutput311 _1886_/X vssd1 vssd1 vccd1 vccd1 io_wo[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_10_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1459_ _1957_/X _2078_/X vssd1 vssd1 vccd1 vccd1 _1505_/A sky130_fd_sc_hd__xor2_4
X_1528_ _2124_/X vssd1 vssd1 vccd1 vccd1 _1536_/A sky130_fd_sc_hd__inv_2
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1244_ _1244_/A vssd1 vssd1 vccd1 vccd1 _1245_/C sky130_fd_sc_hd__inv_2
X_2293_ _2295_/CLK _2293_/D vssd1 vssd1 vccd1 vccd1 _2293_/Q sky130_fd_sc_hd__dfxtp_4
X_1313_ _2040_/X _2115_/X vssd1 vssd1 vccd1 vccd1 _1313_/X sky130_fd_sc_hd__and2b_1
XFILLER_2_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1175_ _1189_/A vssd1 vssd1 vccd1 vccd1 _1175_/X sky130_fd_sc_hd__clkbuf_2
Xoutput163 _1862_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[12] sky130_fd_sc_hd__clkbuf_2
Xoutput174 _1852_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[8] sky130_fd_sc_hd__clkbuf_2
Xoutput185 _1812_/Y vssd1 vssd1 vccd1 vccd1 io_o_1_co sky130_fd_sc_hd__clkbuf_2
Xoutput196 _2205_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1931_ _1931_/A vssd1 vssd1 vccd1 vccd1 _1931_/X sky130_fd_sc_hd__clkbuf_2
Xinput54 io_eo[40] vssd1 vssd1 vccd1 vccd1 _1918_/A sky130_fd_sc_hd__clkbuf_1
Xinput43 io_eo[30] vssd1 vssd1 vccd1 vccd1 _1908_/A sky130_fd_sc_hd__clkbuf_1
X_1793_ _2028_/X _2112_/X vssd1 vssd1 vccd1 vccd1 _1793_/X sky130_fd_sc_hd__and2b_1
Xinput32 io_eo[20] vssd1 vssd1 vccd1 vccd1 _1898_/A sky130_fd_sc_hd__clkbuf_1
Xinput21 io_eo[10] vssd1 vssd1 vccd1 vccd1 _1888_/A sky130_fd_sc_hd__clkbuf_1
X_1862_ _2272_/Q _1849_/X _1850_/X _1861_/X vssd1 vssd1 vccd1 vccd1 _1862_/X sky130_fd_sc_hd__a31o_1
Xinput10 io_dat_i[15] vssd1 vssd1 vccd1 vccd1 _1060_/A sky130_fd_sc_hd__clkbuf_1
Xinput76 io_eo[60] vssd1 vssd1 vccd1 vccd1 _1938_/A sky130_fd_sc_hd__clkbuf_1
Xinput65 io_eo[50] vssd1 vssd1 vccd1 vccd1 _1928_/A sky130_fd_sc_hd__clkbuf_1
Xinput87 io_i_0_in1[2] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_1
Xinput98 io_i_1_in1[4] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_1
X_2276_ _2299_/CLK _2276_/D vssd1 vssd1 vccd1 vccd1 _2276_/Q sky130_fd_sc_hd__dfxtp_2
X_1158_ _1839_/A _1833_/C _1158_/C vssd1 vssd1 vccd1 vccd1 _1189_/A sky130_fd_sc_hd__nor3_4
XFILLER_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1227_ _2016_/X _2106_/X vssd1 vssd1 vccd1 vccd1 _1282_/A sky130_fd_sc_hd__and2b_1
XFILLER_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1089_ _1089_/A vssd1 vssd1 vccd1 vccd1 _1876_/C sky130_fd_sc_hd__inv_2
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2130_ _2130_/A0 _2177_/Q _2193_/Q _2225_/Q _2254_/Q _2255_/Q vssd1 vssd1 vccd1 vccd1
+ _2130_/X sky130_fd_sc_hd__mux4_2
X_2061_ _2061_/A0 _2224_/Q _2248_/Q vssd1 vssd1 vccd1 vccd1 _2061_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1914_ _1914_/A vssd1 vssd1 vccd1 vccd1 _1914_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1776_ _1776_/A _1780_/B vssd1 vssd1 vccd1 vccd1 _1776_/Y sky130_fd_sc_hd__nand2_1
X_1845_ _1849_/A _1845_/B _2251_/Q vssd1 vssd1 vccd1 vccd1 _1847_/A sky130_fd_sc_hd__nand3_1
X_2259_ _2291_/CLK _2259_/D vssd1 vssd1 vccd1 vccd1 _2259_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1630_ _1657_/S vssd1 vssd1 vccd1 vccd1 _1647_/S sky130_fd_sc_hd__buf_2
XPHY_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1561_ _2167_/Q _1685_/B _1561_/S vssd1 vssd1 vccd1 vccd1 _2167_/D sky130_fd_sc_hd__mux2_1
X_1492_ _1490_/Y _1491_/X _1485_/A vssd1 vssd1 vccd1 vccd1 _1492_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_66_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2044_ _1750_/Y _2043_/X _2295_/Q vssd1 vssd1 vccd1 vccd1 _2044_/X sky130_fd_sc_hd__mux2_1
X_2113_ input96/X _2230_/Q _1689_/A _2127_/A0 _2246_/Q _2247_/Q vssd1 vssd1 vccd1
+ vccd1 _2113_/X sky130_fd_sc_hd__mux4_2
XFILLER_30_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1828_ _2293_/Q _1824_/X _2277_/Q _1825_/X _1827_/X vssd1 vssd1 vccd1 vccd1 _1828_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1759_ _2199_/Q vssd1 vssd1 vccd1 vccd1 _1759_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1613_ _2138_/X _1613_/B vssd1 vssd1 vccd1 vccd1 _1613_/X sky130_fd_sc_hd__xor2_1
X_1544_ _1543_/X _2176_/Q _1546_/S vssd1 vssd1 vccd1 vccd1 _2176_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1475_ _1475_/A _1475_/B vssd1 vssd1 vccd1 vccd1 _1491_/B sky130_fd_sc_hd__nor2_2
XFILLER_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2027_ _1773_/Y _1706_/Y _2292_/Q vssd1 vssd1 vccd1 vccd1 _2027_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1260_ _1260_/A _1260_/B vssd1 vssd1 vccd1 vccd1 _2235_/D sky130_fd_sc_hd__nand2_1
X_1191_ _1186_/X _1191_/B _1200_/C vssd1 vssd1 vccd1 vccd1 _1191_/Y sky130_fd_sc_hd__nand3b_1
Xinput8 io_dat_i[13] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput301 _1935_/X vssd1 vssd1 vccd1 vccd1 io_wo[57] sky130_fd_sc_hd__clkbuf_2
Xoutput312 _1887_/X vssd1 vssd1 vccd1 vccd1 io_wo[9] sky130_fd_sc_hd__clkbuf_2
X_1527_ _1555_/S vssd1 vssd1 vccd1 vccd1 _1546_/S sky130_fd_sc_hd__clkbuf_2
X_1389_ _1729_/B _2057_/X _1388_/X vssd1 vssd1 vccd1 vccd1 _1389_/Y sky130_fd_sc_hd__o21ai_1
X_1458_ _1452_/X _1456_/Y _1457_/Y vssd1 vssd1 vccd1 vccd1 _1505_/B sky130_fd_sc_hd__o21bai_2
XFILLER_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1243_ _2110_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _1244_/A sky130_fd_sc_hd__and2b_1
X_2292_ _2292_/CLK _2292_/D vssd1 vssd1 vccd1 vccd1 _2292_/Q sky130_fd_sc_hd__dfxtp_4
X_1174_ _2255_/Q _1159_/X _1165_/X _1173_/Y vssd1 vssd1 vccd1 vccd1 _2255_/D sky130_fd_sc_hd__o211a_1
X_1312_ _1312_/A vssd1 vssd1 vccd1 vccd1 _1326_/C sky130_fd_sc_hd__inv_2
XFILLER_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput164 _1864_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[13] sky130_fd_sc_hd__clkbuf_2
Xoutput175 _1854_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[9] sky130_fd_sc_hd__clkbuf_2
Xoutput186 _2220_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput197 _2206_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[2] sky130_fd_sc_hd__clkbuf_2
XPHY_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1930_ _1930_/A vssd1 vssd1 vccd1 vccd1 _1930_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput77 io_eo[61] vssd1 vssd1 vccd1 vccd1 _1939_/A sky130_fd_sc_hd__clkbuf_1
Xinput66 io_eo[51] vssd1 vssd1 vccd1 vccd1 _1929_/A sky130_fd_sc_hd__clkbuf_1
Xinput55 io_eo[41] vssd1 vssd1 vccd1 vccd1 _1919_/A sky130_fd_sc_hd__clkbuf_1
Xinput44 io_eo[31] vssd1 vssd1 vccd1 vccd1 _1909_/A sky130_fd_sc_hd__clkbuf_1
Xinput33 io_eo[21] vssd1 vssd1 vccd1 vccd1 _1899_/A sky130_fd_sc_hd__clkbuf_1
X_1792_ _1792_/A vssd1 vssd1 vccd1 vccd1 _1792_/Y sky130_fd_sc_hd__inv_2
Xinput22 io_eo[11] vssd1 vssd1 vccd1 vccd1 _1889_/A sky130_fd_sc_hd__clkbuf_1
X_1861_ _2256_/Q _1855_/X _1858_/X _2288_/Q vssd1 vssd1 vccd1 vccd1 _1861_/X sky130_fd_sc_hd__a22o_1
Xinput11 io_dat_i[1] vssd1 vssd1 vccd1 vccd1 _1044_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput88 io_i_0_in1[3] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__clkbuf_1
Xinput99 io_i_1_in1[5] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1157_ _1823_/A vssd1 vssd1 vccd1 vccd1 _1839_/A sky130_fd_sc_hd__buf_2
XFILLER_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2275_ _2275_/CLK _2275_/D vssd1 vssd1 vccd1 vccd1 _2275_/Q sky130_fd_sc_hd__dfxtp_2
X_1226_ _1784_/A _2016_/X vssd1 vssd1 vccd1 vccd1 _1226_/Y sky130_fd_sc_hd__nand2_2
XFILLER_16_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1088_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1088_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2060_ _1723_/Y _2059_/X _2297_/Q vssd1 vssd1 vccd1 vccd1 _2060_/X sky130_fd_sc_hd__mux2_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1913_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1913_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1775_ _2218_/Q vssd1 vssd1 vccd1 vccd1 _1775_/Y sky130_fd_sc_hd__inv_2
X_1844_ _1700_/A _1824_/X _2282_/Q _1825_/X _1843_/Y vssd1 vssd1 vccd1 vccd1 _1844_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2258_ _2291_/CLK _2258_/D vssd1 vssd1 vccd1 vccd1 _2258_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2189_ _2195_/CLK _2189_/D vssd1 vssd1 vccd1 vccd1 _2189_/Q sky130_fd_sc_hd__dfxtp_2
X_1209_ _1951_/X vssd1 vssd1 vccd1 vccd1 _1209_/X sky130_fd_sc_hd__buf_2
XFILLER_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_4_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2272_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1560_ _2168_/Q _1961_/X _1561_/S vssd1 vssd1 vccd1 vccd1 _2168_/D sky130_fd_sc_hd__mux2_1
X_1491_ _1491_/A _1491_/B _1491_/C vssd1 vssd1 vccd1 vccd1 _1491_/X sky130_fd_sc_hd__and3_1
X_2112_ input92/X _1661_/A _1705_/A _2125_/A0 _2244_/Q _2245_/Q vssd1 vssd1 vccd1
+ vccd1 _2112_/X sky130_fd_sc_hd__mux4_2
XFILLER_3_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2043_ _1751_/Y _1668_/Y _2294_/Q vssd1 vssd1 vccd1 vccd1 _2043_/X sky130_fd_sc_hd__mux2_1
X_1827_ _2245_/Q _1203_/C _1826_/Y vssd1 vssd1 vccd1 vccd1 _1827_/X sky130_fd_sc_hd__a21bo_1
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1689_ _1689_/A vssd1 vssd1 vccd1 vccd1 _1689_/Y sky130_fd_sc_hd__inv_2
X_1758_ _1758_/A _1760_/B vssd1 vssd1 vccd1 vccd1 _1758_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1474_ _1963_/X _2087_/X _1961_/X _2084_/X vssd1 vssd1 vccd1 vccd1 _1475_/B sky130_fd_sc_hd__a211oi_4
X_1612_ _1620_/B _2135_/X _2136_/X _2137_/X vssd1 vssd1 vccd1 vccd1 _1613_/B sky130_fd_sc_hd__and4_1
X_1543_ _2122_/X _1543_/B vssd1 vssd1 vccd1 vccd1 _1543_/X sky130_fd_sc_hd__xor2_1
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2026_ _1774_/Y _2025_/X _2293_/Q vssd1 vssd1 vccd1 vccd1 _2026_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1190_ _1855_/A vssd1 vssd1 vccd1 vccd1 _1200_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 io_dat_i[14] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput302 _1936_/X vssd1 vssd1 vccd1 vccd1 io_wo[58] sky130_fd_sc_hd__clkbuf_2
X_1457_ _1955_/X _2075_/X vssd1 vssd1 vccd1 vccd1 _1457_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1526_ _1949_/X vssd1 vssd1 vccd1 vccd1 _1555_/S sky130_fd_sc_hd__inv_2
X_1388_ _1729_/B _2057_/X _1975_/X _2054_/X vssd1 vssd1 vccd1 vccd1 _1388_/X sky130_fd_sc_hd__a211o_1
XFILLER_82_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2009_ _1770_/Y _1813_/A _2262_/Q vssd1 vssd1 vccd1 vccd1 _2009_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2291_ _2291_/CLK _2291_/D vssd1 vssd1 vccd1 vccd1 _2291_/Q sky130_fd_sc_hd__dfxtp_1
X_1311_ _2116_/X _2042_/X vssd1 vssd1 vccd1 vccd1 _1312_/A sky130_fd_sc_hd__and2b_1
X_1242_ _1242_/A vssd1 vssd1 vccd1 vccd1 _1253_/C sky130_fd_sc_hd__inv_2
X_1173_ _1172_/X _1173_/B _1173_/C vssd1 vssd1 vccd1 vccd1 _1173_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput165 _1866_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[14] sky130_fd_sc_hd__clkbuf_2
X_1509_ _1951_/X vssd1 vssd1 vccd1 vccd1 _1564_/S sky130_fd_sc_hd__buf_2
Xoutput176 _1813_/Y vssd1 vssd1 vccd1 vccd1 io_o_0_co sky130_fd_sc_hd__clkbuf_2
Xoutput187 _2221_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput198 _2207_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[3] sky130_fd_sc_hd__clkbuf_2
XPHY_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1860_ _2271_/Q _1849_/X _1850_/X _1859_/X vssd1 vssd1 vccd1 vccd1 _1860_/X sky130_fd_sc_hd__a31o_1
XFILLER_14_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput67 io_eo[52] vssd1 vssd1 vccd1 vccd1 _1930_/A sky130_fd_sc_hd__clkbuf_1
Xinput78 io_eo[62] vssd1 vssd1 vccd1 vccd1 _1940_/A sky130_fd_sc_hd__clkbuf_1
Xinput56 io_eo[42] vssd1 vssd1 vccd1 vccd1 _1920_/A sky130_fd_sc_hd__clkbuf_1
Xinput45 io_eo[32] vssd1 vssd1 vccd1 vccd1 _1910_/A sky130_fd_sc_hd__clkbuf_1
X_1791_ _2112_/X _2028_/X vssd1 vssd1 vccd1 vccd1 _1792_/A sky130_fd_sc_hd__and2b_1
Xinput34 io_eo[22] vssd1 vssd1 vccd1 vccd1 _1900_/A sky130_fd_sc_hd__clkbuf_1
Xinput23 io_eo[12] vssd1 vssd1 vccd1 vccd1 _1890_/A sky130_fd_sc_hd__clkbuf_1
Xinput12 io_dat_i[2] vssd1 vssd1 vccd1 vccd1 _1040_/A sky130_fd_sc_hd__clkbuf_1
Xinput89 io_i_0_in1[4] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2274_ _2275_/CLK _2274_/D vssd1 vssd1 vccd1 vccd1 _2274_/Q sky130_fd_sc_hd__dfxtp_2
X_1087_ _2284_/Q _1077_/X _1069_/X _1086_/Y vssd1 vssd1 vccd1 vccd1 _2284_/D sky130_fd_sc_hd__o211a_1
XFILLER_52_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1156_ _2260_/Q _1125_/A _1148_/X _1155_/Y vssd1 vssd1 vccd1 vccd1 _2260_/D sky130_fd_sc_hd__o211a_1
X_1225_ _2106_/X vssd1 vssd1 vccd1 vccd1 _1784_/A sky130_fd_sc_hd__inv_2
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1989_ _1765_/Y _1988_/X _2247_/Q vssd1 vssd1 vccd1 vccd1 _1989_/X sky130_fd_sc_hd__mux2_2
XFILLER_57_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1912_ _1912_/A vssd1 vssd1 vccd1 vccd1 _1912_/X sky130_fd_sc_hd__clkbuf_2
X_1843_ _1702_/Y _1814_/Y _1842_/Y vssd1 vssd1 vccd1 vccd1 _1843_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1774_ _1774_/A _1780_/B vssd1 vssd1 vccd1 vccd1 _1774_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1208_ _1214_/A _1207_/X vssd1 vssd1 vccd1 vccd1 _2242_/D sky130_fd_sc_hd__nor2b_1
X_2257_ _2291_/CLK _2257_/D vssd1 vssd1 vccd1 vccd1 _2257_/Q sky130_fd_sc_hd__dfxtp_4
X_2188_ _2272_/CLK _2188_/D vssd1 vssd1 vccd1 vccd1 _2188_/Q sky130_fd_sc_hd__dfxtp_1
X_1139_ _2267_/Q _1130_/X _1135_/X _1138_/Y vssd1 vssd1 vccd1 vccd1 _2267_/D sky130_fd_sc_hd__o211a_1
XFILLER_25_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1490_ _1491_/A _1491_/B _1491_/C vssd1 vssd1 vccd1 vccd1 _1490_/Y sky130_fd_sc_hd__a21oi_1
X_2111_ input91/X _1667_/A _1711_/A _2124_/A0 _2244_/Q _2245_/Q vssd1 vssd1 vccd1
+ vccd1 _2111_/X sky130_fd_sc_hd__mux4_2
X_2042_ _1752_/Y _2041_/X _2295_/Q vssd1 vssd1 vccd1 vccd1 _2042_/X sky130_fd_sc_hd__mux2_2
XFILLER_81_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1826_ _1823_/A _2261_/Q _1833_/C vssd1 vssd1 vccd1 vccd1 _1826_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_89_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1757_ _2221_/Q vssd1 vssd1 vccd1 vccd1 _1757_/Y sky130_fd_sc_hd__inv_2
X_1688_ _2079_/X vssd1 vssd1 vccd1 vccd1 _1688_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1611_ _2133_/X _1611_/B _2134_/X _2000_/X vssd1 vssd1 vccd1 vccd1 _1620_/B sky130_fd_sc_hd__and4b_1
X_1473_ _1489_/A vssd1 vssd1 vccd1 vccd1 _1476_/B sky130_fd_sc_hd__inv_2
X_1542_ _1546_/S _2177_/Q _1541_/Y vssd1 vssd1 vccd1 vccd1 _2177_/D sky130_fd_sc_hd__a21bo_1
XFILLER_5_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2025_ _1775_/Y _1712_/Y _2292_/Q vssd1 vssd1 vccd1 vccd1 _2025_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1809_ _1871_/A _2280_/Q vssd1 vssd1 vccd1 vccd1 _1809_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput303 _1937_/X vssd1 vssd1 vccd1 vccd1 io_wo[59] sky130_fd_sc_hd__clkbuf_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1387_ _1387_/A _1387_/B vssd1 vssd1 vccd1 vccd1 _1428_/A sky130_fd_sc_hd__nor2_2
X_1525_ _2180_/Q _1971_/X _1525_/S vssd1 vssd1 vccd1 vccd1 _2180_/D sky130_fd_sc_hd__mux2_1
X_1456_ _1513_/A _1454_/Y _1455_/Y vssd1 vssd1 vccd1 vccd1 _1456_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_19_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2008_ _1745_/Y _2007_/X _2265_/Q vssd1 vssd1 vccd1 vccd1 _2008_/X sky130_fd_sc_hd__mux2_2
XFILLER_51_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1241_ _2111_/X _2026_/X vssd1 vssd1 vccd1 vccd1 _1242_/A sky130_fd_sc_hd__and2b_1
X_2290_ _2291_/CLK _2290_/D vssd1 vssd1 vccd1 vccd1 _2290_/Q sky130_fd_sc_hd__dfxtp_1
X_1310_ _2044_/X _2117_/X vssd1 vssd1 vccd1 vccd1 _1333_/A sky130_fd_sc_hd__or2b_2
XFILLER_66_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1172_ _1186_/A vssd1 vssd1 vccd1 vccd1 _1172_/X sky130_fd_sc_hd__buf_1
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput166 _1868_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[15] sky130_fd_sc_hd__clkbuf_2
Xoutput177 _2228_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[0] sky130_fd_sc_hd__clkbuf_2
X_1508_ _1457_/Y _1452_/X _1456_/Y vssd1 vssd1 vccd1 vccd1 _1508_/X sky130_fd_sc_hd__o21a_1
Xoutput199 _2208_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput188 _2222_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[2] sky130_fd_sc_hd__clkbuf_2
X_1439_ _2204_/Q vssd1 vssd1 vccd1 vccd1 _1439_/Y sky130_fd_sc_hd__inv_2
XPHY_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1790_ _1790_/A vssd1 vssd1 vccd1 vccd1 _1790_/Y sky130_fd_sc_hd__inv_2
Xinput13 io_dat_i[3] vssd1 vssd1 vccd1 vccd1 _1036_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput68 io_eo[53] vssd1 vssd1 vccd1 vccd1 _1931_/A sky130_fd_sc_hd__clkbuf_1
Xinput79 io_eo[63] vssd1 vssd1 vccd1 vccd1 _1941_/A sky130_fd_sc_hd__clkbuf_1
Xinput57 io_eo[43] vssd1 vssd1 vccd1 vccd1 _1921_/A sky130_fd_sc_hd__clkbuf_1
Xinput46 io_eo[33] vssd1 vssd1 vccd1 vccd1 _1911_/A sky130_fd_sc_hd__clkbuf_1
Xinput35 io_eo[23] vssd1 vssd1 vccd1 vccd1 _1901_/A sky130_fd_sc_hd__clkbuf_1
Xinput24 io_eo[13] vssd1 vssd1 vccd1 vccd1 _1891_/A sky130_fd_sc_hd__clkbuf_1
X_2273_ _2275_/CLK _2273_/D vssd1 vssd1 vccd1 vccd1 _2273_/Q sky130_fd_sc_hd__dfxtp_2
X_1224_ _2012_/X _1287_/A _1223_/X vssd1 vssd1 vccd1 vccd1 _1224_/Y sky130_fd_sc_hd__o21ai_4
X_1086_ _1078_/X _1090_/B _1182_/B vssd1 vssd1 vccd1 vccd1 _1086_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_37_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1155_ _1155_/A _1203_/B vssd1 vssd1 vccd1 vccd1 _1155_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1988_ _1699_/Y _1766_/Y _2246_/Q vssd1 vssd1 vccd1 vccd1 _1988_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1773_ _2219_/Q vssd1 vssd1 vccd1 vccd1 _1773_/Y sky130_fd_sc_hd__inv_2
X_1911_ _1911_/A vssd1 vssd1 vccd1 vccd1 _1911_/X sky130_fd_sc_hd__clkbuf_2
X_1842_ _1849_/A _1845_/B _2250_/Q vssd1 vssd1 vccd1 vccd1 _1842_/Y sky130_fd_sc_hd__nand3_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2187_ _2219_/CLK _2187_/D vssd1 vssd1 vccd1 vccd1 _2187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1207_ _1947_/X vssd1 vssd1 vccd1 vccd1 _1207_/X sky130_fd_sc_hd__clkbuf_2
X_2256_ _2291_/CLK _2256_/D vssd1 vssd1 vccd1 vccd1 _2256_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1069_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1138_ _1138_/A _1876_/C vssd1 vssd1 vccd1 vccd1 _1138_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2041_ _1753_/Y _1339_/Y _2294_/Q vssd1 vssd1 vccd1 vccd1 _2041_/X sky130_fd_sc_hd__mux2_1
X_2110_ input90/X _1672_/A _1716_/A _2123_/A0 _2244_/Q _2245_/Q vssd1 vssd1 vccd1
+ vccd1 _2110_/X sky130_fd_sc_hd__mux4_2
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1825_ _1825_/A vssd1 vssd1 vccd1 vccd1 _1825_/X sky130_fd_sc_hd__clkbuf_2
X_1756_ _2200_/Q vssd1 vssd1 vccd1 vccd1 _1756_/Y sky130_fd_sc_hd__inv_2
X_1687_ _2167_/Q vssd1 vssd1 vccd1 vccd1 _1687_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2239_ _2297_/CLK _2239_/D vssd1 vssd1 vccd1 vccd1 _2239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1610_ _1616_/A _1606_/Y _1608_/X _1609_/Y vssd1 vssd1 vccd1 vccd1 _2155_/D sky130_fd_sc_hd__o31ai_1
XFILLER_5_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1472_ _1965_/X _2090_/X vssd1 vssd1 vccd1 vccd1 _1489_/A sky130_fd_sc_hd__nor2_1
X_1541_ _1541_/A _1541_/B _1949_/X vssd1 vssd1 vccd1 vccd1 _1541_/Y sky130_fd_sc_hd__nand3_1
XFILLER_5_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2024_ _1776_/Y _2023_/X _2293_/Q vssd1 vssd1 vccd1 vccd1 _2024_/X sky130_fd_sc_hd__mux2_2
XFILLER_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1739_ _1743_/A _1973_/X vssd1 vssd1 vccd1 vccd1 _1739_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1808_ _2156_/Q vssd1 vssd1 vccd1 vccd1 _1808_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1524_ _2181_/Q _1973_/X _1525_/S vssd1 vssd1 vccd1 vccd1 _2181_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput304 _1883_/X vssd1 vssd1 vccd1 vccd1 io_wo[5] sky130_fd_sc_hd__clkbuf_2
X_1386_ _1977_/X _2057_/X vssd1 vssd1 vccd1 vccd1 _1387_/B sky130_fd_sc_hd__and2_1
X_1455_ _1953_/X _2072_/X vssd1 vssd1 vccd1 vccd1 _1455_/Y sky130_fd_sc_hd__nor2_4
XFILLER_4_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2007_ _1746_/Y _1812_/A _2264_/Q vssd1 vssd1 vccd1 vccd1 _2007_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1240_ _1269_/B _1240_/B vssd1 vssd1 vccd1 vccd1 _1245_/A sky130_fd_sc_hd__nand2_1
X_1171_ _2256_/Q _1159_/X _1165_/X _1170_/Y vssd1 vssd1 vccd1 vccd1 _2256_/D sky130_fd_sc_hd__o211a_1
XFILLER_1_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput167 _1828_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[1] sky130_fd_sc_hd__clkbuf_2
Xoutput178 _2229_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[1] sky130_fd_sc_hd__clkbuf_2
X_1507_ _2189_/Q vssd1 vssd1 vccd1 vccd1 _1507_/Y sky130_fd_sc_hd__inv_2
Xoutput189 _2223_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[3] sky130_fd_sc_hd__clkbuf_2
X_1438_ _1436_/Y _1378_/Y _1377_/Y _1431_/S vssd1 vssd1 vccd1 vccd1 _1438_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1369_ _2108_/X vssd1 vssd1 vccd1 vccd1 _1780_/A sky130_fd_sc_hd__inv_2
XPHY_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput36 io_eo[24] vssd1 vssd1 vccd1 vccd1 _1902_/A sky130_fd_sc_hd__clkbuf_1
Xinput25 io_eo[14] vssd1 vssd1 vccd1 vccd1 _1892_/A sky130_fd_sc_hd__clkbuf_1
Xinput14 io_dat_i[4] vssd1 vssd1 vccd1 vccd1 _1033_/A sky130_fd_sc_hd__clkbuf_1
Xinput69 io_eo[54] vssd1 vssd1 vccd1 vccd1 _1932_/A sky130_fd_sc_hd__clkbuf_1
Xinput58 io_eo[44] vssd1 vssd1 vccd1 vccd1 _1922_/A sky130_fd_sc_hd__clkbuf_1
Xinput47 io_eo[34] vssd1 vssd1 vccd1 vccd1 _1912_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_37_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2272_ _2272_/CLK _2272_/D vssd1 vssd1 vccd1 vccd1 _2272_/Q sky130_fd_sc_hd__dfxtp_2
X_1154_ _2261_/Q _1143_/X _1148_/X _1153_/Y vssd1 vssd1 vccd1 vccd1 _2261_/D sky130_fd_sc_hd__o211a_1
X_1223_ _2014_/X _2105_/X vssd1 vssd1 vccd1 vccd1 _1223_/X sky130_fd_sc_hd__or2b_2
XFILLER_52_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1085_ _1085_/A vssd1 vssd1 vccd1 vccd1 _1182_/B sky130_fd_sc_hd__inv_2
XFILLER_20_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1987_ _1810_/Y _1986_/X _2279_/Q vssd1 vssd1 vccd1 vccd1 _1987_/X sky130_fd_sc_hd__mux2_4
XFILLER_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1910_ _1910_/A vssd1 vssd1 vccd1 vccd1 _1910_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1772_ _1772_/A _1780_/B vssd1 vssd1 vccd1 vccd1 _1772_/Y sky130_fd_sc_hd__nand2_1
X_1841_ _2265_/Q _1817_/A _1821_/C _1839_/Y _1840_/X vssd1 vssd1 vccd1 vccd1 _1841_/X
+ sky130_fd_sc_hd__a311o_2
XFILLER_8_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2186_ _2219_/CLK _2186_/D vssd1 vssd1 vccd1 vccd1 _2186_/Q sky130_fd_sc_hd__dfxtp_1
X_1206_ _1214_/A _1945_/X vssd1 vssd1 vccd1 vccd1 _2243_/D sky130_fd_sc_hd__nor2b_1
X_2255_ _2291_/CLK _2255_/D vssd1 vssd1 vccd1 vccd1 _2255_/Q sky130_fd_sc_hd__dfxtp_4
X_1137_ _2268_/Q _1130_/X _1135_/X _1136_/Y vssd1 vssd1 vccd1 vccd1 _2268_/D sky130_fd_sc_hd__o211a_1
X_1068_ _2289_/Q _1055_/X _1043_/X _1067_/Y vssd1 vssd1 vccd1 vccd1 _2289_/D sky130_fd_sc_hd__o211a_1
XFILLER_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2040_ _1755_/Y _2039_/X _2295_/Q vssd1 vssd1 vccd1 vccd1 _2040_/X sky130_fd_sc_hd__mux2_2
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1686_ _2191_/Q vssd1 vssd1 vccd1 vccd1 _1686_/Y sky130_fd_sc_hd__inv_2
X_1824_ _1876_/B vssd1 vssd1 vccd1 vccd1 _1824_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1755_ _1755_/A _1760_/B vssd1 vssd1 vccd1 vccd1 _1755_/Y sky130_fd_sc_hd__nand2_1
X_2238_ _2292_/CLK _2238_/D vssd1 vssd1 vccd1 vccd1 _2238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2169_ _2195_/CLK _2169_/D vssd1 vssd1 vccd1 vccd1 _2169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1540_ _1545_/B _2122_/X _2121_/X _2123_/X vssd1 vssd1 vccd1 vccd1 _1541_/A sky130_fd_sc_hd__a31o_1
XFILLER_12_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1471_ _1499_/B _1499_/A _1496_/A vssd1 vssd1 vccd1 vccd1 _1491_/A sky130_fd_sc_hd__nand3_2
XFILLER_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2023_ _1777_/Y _1266_/Y _2292_/Q vssd1 vssd1 vccd1 vccd1 _2023_/X sky130_fd_sc_hd__mux2_1
X_1807_ _1871_/A _2276_/Q vssd1 vssd1 vccd1 vccd1 _1807_/Y sky130_fd_sc_hd__nand2_1
X_1669_ _1685_/A _1965_/X vssd1 vssd1 vccd1 vccd1 _1669_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_4_3_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2251_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1738_ _2052_/X vssd1 vssd1 vccd1 vccd1 _1738_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1523_ _2182_/Q _1975_/X _1525_/S vssd1 vssd1 vccd1 vccd1 _2182_/D sky130_fd_sc_hd__mux2_1
Xoutput305 _1938_/X vssd1 vssd1 vccd1 vccd1 io_wo[60] sky130_fd_sc_hd__clkbuf_2
X_1454_ _2006_/X vssd1 vssd1 vccd1 vccd1 _1454_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1385_ _1729_/B _2057_/X vssd1 vssd1 vccd1 vccd1 _1387_/A sky130_fd_sc_hd__nor2_1
XFILLER_67_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2006_ _1702_/Y _2005_/X _2267_/Q vssd1 vssd1 vccd1 vccd1 _2006_/X sky130_fd_sc_hd__mux2_4
XFILLER_58_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1170_ _1110_/X _1170_/B _1173_/C vssd1 vssd1 vccd1 vccd1 _1170_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput168 _1832_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[2] sky130_fd_sc_hd__clkbuf_2
X_1506_ _1505_/X _2190_/Q _1506_/S vssd1 vssd1 vccd1 vccd1 _2190_/D sky130_fd_sc_hd__mux2_1
X_1437_ _1436_/Y _1377_/Y _1378_/Y vssd1 vssd1 vccd1 vccd1 _1437_/X sky130_fd_sc_hd__a21o_1
Xoutput179 _2230_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[2] sky130_fd_sc_hd__clkbuf_2
X_1368_ _2216_/Q _1778_/A _1372_/S vssd1 vssd1 vccd1 vccd1 _2216_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1299_ _1991_/X _2033_/X vssd1 vssd1 vccd1 vccd1 _1299_/Y sky130_fd_sc_hd__nor2_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput59 io_eo[45] vssd1 vssd1 vccd1 vccd1 _1923_/A sky130_fd_sc_hd__clkbuf_1
Xinput48 io_eo[35] vssd1 vssd1 vccd1 vccd1 _1913_/A sky130_fd_sc_hd__clkbuf_1
Xinput37 io_eo[25] vssd1 vssd1 vccd1 vccd1 _1903_/A sky130_fd_sc_hd__clkbuf_1
Xinput26 io_eo[15] vssd1 vssd1 vccd1 vccd1 _1893_/A sky130_fd_sc_hd__clkbuf_1
Xinput15 io_dat_i[5] vssd1 vssd1 vccd1 vccd1 _1028_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2271_ _2272_/CLK _2271_/D vssd1 vssd1 vccd1 vccd1 _2271_/Q sky130_fd_sc_hd__dfxtp_2
X_1084_ _2285_/Q _1077_/X _1069_/X _1083_/Y vssd1 vssd1 vccd1 vccd1 _2285_/D sky130_fd_sc_hd__o211a_1
XFILLER_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1153_ _1155_/A _1200_/B vssd1 vssd1 vccd1 vccd1 _1153_/Y sky130_fd_sc_hd__nand2_1
X_1222_ _2105_/X _2014_/X vssd1 vssd1 vccd1 vccd1 _1287_/A sky130_fd_sc_hd__and2b_1
X_1986_ _1993_/X _2238_/Q _2278_/Q vssd1 vssd1 vccd1 vccd1 _1986_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1840_ _1876_/B _2297_/Q _2281_/Q _1825_/A vssd1 vssd1 vccd1 vccd1 _1840_/X sky130_fd_sc_hd__a22o_1
X_1771_ _2292_/Q vssd1 vssd1 vccd1 vccd1 _1780_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2254_ _2254_/CLK _2254_/D vssd1 vssd1 vccd1 vccd1 _2254_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2185_ _2219_/CLK _2185_/D vssd1 vssd1 vccd1 vccd1 _2185_/Q sky130_fd_sc_hd__dfxtp_1
X_1205_ _1219_/A vssd1 vssd1 vccd1 vccd1 _1214_/A sky130_fd_sc_hd__clkbuf_2
X_1067_ _1056_/X _1071_/B _1168_/B vssd1 vssd1 vccd1 vccd1 _1067_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1136_ _1138_/A _1182_/B vssd1 vssd1 vccd1 vccd1 _1136_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1969_ _1809_/Y _1968_/X _2281_/Q vssd1 vssd1 vccd1 vccd1 _1969_/X sky130_fd_sc_hd__mux2_2
XFILLER_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1823_ _1823_/A _1823_/B vssd1 vssd1 vccd1 vccd1 _1876_/B sky130_fd_sc_hd__and2_1
X_1685_ _1685_/A _1685_/B vssd1 vssd1 vccd1 vccd1 _1685_/Y sky130_fd_sc_hd__nand2_1
X_1754_ _1754_/A vssd1 vssd1 vccd1 vccd1 _1754_/Y sky130_fd_sc_hd__inv_2
X_2237_ _2292_/CLK _2237_/D vssd1 vssd1 vccd1 vccd1 _2237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2168_ _2195_/CLK _2168_/D vssd1 vssd1 vccd1 vccd1 _2168_/Q sky130_fd_sc_hd__dfxtp_1
X_1119_ _2275_/Q _1116_/X _1104_/X _1118_/Y vssd1 vssd1 vccd1 vccd1 _2275_/D sky130_fd_sc_hd__o211a_1
X_2099_ _1683_/A _2151_/Q _2159_/Q _2191_/Q _2258_/Q _2259_/Q vssd1 vssd1 vccd1 vccd1
+ _2099_/X sky130_fd_sc_hd__mux4_2
XFILLER_88_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1470_ _1475_/A _1470_/B vssd1 vssd1 vccd1 vccd1 _1496_/A sky130_fd_sc_hd__nor2_2
XFILLER_5_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2022_ _1778_/Y _2021_/X _2293_/Q vssd1 vssd1 vccd1 vccd1 _2022_/X sky130_fd_sc_hd__mux2_2
XFILLER_62_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1806_ _1875_/A vssd1 vssd1 vccd1 vccd1 _1871_/A sky130_fd_sc_hd__clkbuf_2
X_1737_ _2182_/Q vssd1 vssd1 vccd1 vccd1 _1737_/Y sky130_fd_sc_hd__inv_2
X_1668_ _2226_/Q vssd1 vssd1 vccd1 vccd1 _1668_/Y sky130_fd_sc_hd__inv_2
X_1599_ _1945_/X vssd1 vssd1 vccd1 vccd1 _1628_/S sky130_fd_sc_hd__inv_2
XFILLER_53_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput306 _1939_/X vssd1 vssd1 vccd1 vccd1 io_wo[61] sky130_fd_sc_hd__clkbuf_2
X_1522_ _2183_/Q _1729_/B _1522_/S vssd1 vssd1 vccd1 vccd1 _2183_/D sky130_fd_sc_hd__mux2_1
X_1453_ _1953_/X _2072_/X vssd1 vssd1 vccd1 vccd1 _1513_/A sky130_fd_sc_hd__nand2_2
XFILLER_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1384_ _1977_/X vssd1 vssd1 vccd1 vccd1 _1729_/B sky130_fd_sc_hd__buf_1
XFILLER_67_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2005_ _1703_/Y _1811_/A _2266_/Q vssd1 vssd1 vccd1 vccd1 _2005_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput169 _1835_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[3] sky130_fd_sc_hd__clkbuf_2
X_1505_ _1505_/A _1505_/B vssd1 vssd1 vccd1 vccd1 _1505_/X sky130_fd_sc_hd__xor2_1
X_1436_ _1436_/A vssd1 vssd1 vccd1 vccd1 _1436_/Y sky130_fd_sc_hd__inv_2
X_1367_ _2109_/X vssd1 vssd1 vccd1 vccd1 _1778_/A sky130_fd_sc_hd__inv_2
XPHY_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1298_ _1991_/X _2033_/X vssd1 vssd1 vccd1 vccd1 _1352_/B sky130_fd_sc_hd__xnor2_2
XFILLER_23_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput49 io_eo[36] vssd1 vssd1 vccd1 vccd1 _1914_/A sky130_fd_sc_hd__clkbuf_1
Xinput38 io_eo[26] vssd1 vssd1 vccd1 vccd1 _1904_/A sky130_fd_sc_hd__clkbuf_1
Xinput27 io_eo[16] vssd1 vssd1 vccd1 vccd1 _1894_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput16 io_dat_i[6] vssd1 vssd1 vccd1 vccd1 _1025_/A sky130_fd_sc_hd__clkbuf_1
X_2270_ _2272_/CLK _2270_/D vssd1 vssd1 vccd1 vccd1 _2270_/Q sky130_fd_sc_hd__dfxtp_2
X_1221_ _1221_/A vssd1 vssd1 vccd1 vccd1 _1280_/A sky130_fd_sc_hd__inv_2
X_1083_ _1078_/X _1090_/B _1180_/B vssd1 vssd1 vccd1 vccd1 _1083_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_45_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1152_ _2262_/Q _1143_/X _1148_/X _1151_/Y vssd1 vssd1 vccd1 vccd1 _2262_/D sky130_fd_sc_hd__o211a_1
X_1985_ _1704_/Y _1984_/X _2249_/Q vssd1 vssd1 vccd1 vccd1 _1985_/X sky130_fd_sc_hd__mux2_2
XFILLER_9_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1419_ _1424_/B _1424_/A _1418_/Y vssd1 vssd1 vccd1 vccd1 _1420_/B sky130_fd_sc_hd__a21oi_1
XFILLER_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1770_ _1770_/A vssd1 vssd1 vccd1 vccd1 _1770_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2184_ _2219_/CLK _2184_/D vssd1 vssd1 vccd1 vccd1 _2184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1204_ _2244_/Q _1189_/A _1193_/X _1203_/Y vssd1 vssd1 vccd1 vccd1 _2244_/D sky130_fd_sc_hd__o211a_1
X_2253_ _2254_/CLK _2253_/D vssd1 vssd1 vccd1 vccd1 _2253_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_1066_ input8/X vssd1 vssd1 vccd1 vccd1 _1168_/B sky130_fd_sc_hd__inv_2
X_1135_ _1165_/A vssd1 vssd1 vccd1 vccd1 _1135_/X sky130_fd_sc_hd__clkbuf_2
X_1968_ _1987_/X _2239_/Q _2280_/Q vssd1 vssd1 vccd1 vccd1 _1968_/X sky130_fd_sc_hd__mux2_1
X_1899_ _1899_/A vssd1 vssd1 vccd1 vccd1 _1899_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1822_ _1788_/Y _1814_/Y _1817_/Y _1819_/Y _1821_/Y vssd1 vssd1 vccd1 vccd1 _1822_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_1753_ _2201_/Q vssd1 vssd1 vccd1 vccd1 _1753_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1684_ _2223_/Q vssd1 vssd1 vccd1 vccd1 _1684_/Y sky130_fd_sc_hd__inv_2
X_2167_ _2195_/CLK _2167_/D vssd1 vssd1 vccd1 vccd1 _2167_/Q sky130_fd_sc_hd__dfxtp_1
X_2236_ _2299_/CLK _2236_/D vssd1 vssd1 vccd1 vccd1 _2236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1049_ _1049_/A _1203_/B vssd1 vssd1 vccd1 vccd1 _1049_/Y sky130_fd_sc_hd__nand2_1
X_2098_ _1677_/A _2152_/Q _2160_/Q _2192_/Q _2258_/Q _2259_/Q vssd1 vssd1 vccd1 vccd1
+ _2098_/X sky130_fd_sc_hd__mux4_2
X_1118_ _1125_/A _1163_/B vssd1 vssd1 vccd1 vccd1 _1118_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2021_ _1779_/Y _1722_/Y _2292_/Q vssd1 vssd1 vccd1 vccd1 _2021_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1736_ _2206_/Q vssd1 vssd1 vccd1 vccd1 _1736_/Y sky130_fd_sc_hd__inv_2
X_1805_ _1805_/A vssd1 vssd1 vccd1 vccd1 _1875_/A sky130_fd_sc_hd__inv_2
XFILLER_85_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1667_ _1667_/A vssd1 vssd1 vccd1 vccd1 _1667_/Y sky130_fd_sc_hd__inv_2
X_1598_ _1597_/Y _2156_/Q _1598_/S vssd1 vssd1 vccd1 vccd1 _2156_/D sky130_fd_sc_hd__mux2_1
X_2219_ _2219_/CLK _2219_/D vssd1 vssd1 vccd1 vccd1 _2219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput307 _1940_/X vssd1 vssd1 vccd1 vccd1 io_wo[62] sky130_fd_sc_hd__clkbuf_2
X_1521_ _2184_/Q _1979_/X _1522_/S vssd1 vssd1 vccd1 vccd1 _2184_/D sky130_fd_sc_hd__mux2_1
X_1452_ _1955_/X _2075_/X vssd1 vssd1 vccd1 vccd1 _1452_/X sky130_fd_sc_hd__and2_1
X_1383_ _1975_/X _2054_/X vssd1 vssd1 vccd1 vccd1 _1430_/A sky130_fd_sc_hd__xor2_2
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2004_ _2268_/Q _2003_/X _2269_/Q vssd1 vssd1 vccd1 vccd1 _2004_/X sky130_fd_sc_hd__mux2_2
XFILLER_90_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1719_ _2185_/Q vssd1 vssd1 vccd1 vccd1 _1719_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1504_ _1503_/Y _2191_/Q _1506_/S vssd1 vssd1 vccd1 vccd1 _2191_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1435_ _1211_/X _1432_/Y _1433_/X _1434_/Y vssd1 vssd1 vccd1 vccd1 _2205_/D sky130_fd_sc_hd__o22ai_1
X_1366_ _2217_/Q _1776_/A _1372_/S vssd1 vssd1 vccd1 vccd1 _2217_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1297_ _1355_/A _1295_/Y _1296_/Y vssd1 vssd1 vccd1 vccd1 _1352_/A sky130_fd_sc_hd__a21oi_4
XFILLER_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput39 io_eo[27] vssd1 vssd1 vccd1 vccd1 _1905_/A sky130_fd_sc_hd__clkbuf_1
Xinput28 io_eo[17] vssd1 vssd1 vccd1 vccd1 _1895_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput17 io_dat_i[7] vssd1 vssd1 vccd1 vccd1 _1089_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_77_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1220_ _2107_/X _2018_/X vssd1 vssd1 vccd1 vccd1 _1221_/A sky130_fd_sc_hd__xnor2_1
X_1151_ _1151_/A _1198_/B vssd1 vssd1 vccd1 vccd1 _1151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1082_ _1082_/A vssd1 vssd1 vccd1 vccd1 _1180_/B sky130_fd_sc_hd__inv_2
XFILLER_60_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1984_ _1706_/Y _1705_/Y _2248_/Q vssd1 vssd1 vccd1 vccd1 _1984_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_1418_ _1979_/X _2060_/X vssd1 vssd1 vccd1 vccd1 _1418_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1349_ _1348_/Y _2223_/Q _1353_/S vssd1 vssd1 vccd1 vccd1 _2223_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2183_ _2219_/CLK _2183_/D vssd1 vssd1 vccd1 vccd1 _2183_/Q sky130_fd_sc_hd__dfxtp_1
X_2252_ _2254_/CLK _2252_/D vssd1 vssd1 vccd1 vccd1 _2252_/Q sky130_fd_sc_hd__dfxtp_4
X_1203_ _1158_/C _1203_/B _1203_/C vssd1 vssd1 vccd1 vccd1 _1203_/Y sky130_fd_sc_hd__nand3b_1
X_1134_ _2269_/Q _1130_/X _1122_/X _1133_/Y vssd1 vssd1 vccd1 vccd1 _2269_/D sky130_fd_sc_hd__o211a_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1065_ _2290_/Q _1055_/X _1043_/X _1064_/Y vssd1 vssd1 vccd1 vccd1 _2290_/D sky130_fd_sc_hd__o211a_1
XFILLER_33_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1898_ _1898_/A vssd1 vssd1 vccd1 vccd1 _1898_/X sky130_fd_sc_hd__clkbuf_2
X_1967_ _1660_/Y _1966_/X _2251_/Q vssd1 vssd1 vccd1 vccd1 _1967_/X sky130_fd_sc_hd__mux2_4
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1821_ _1821_/A _1839_/A _1821_/C vssd1 vssd1 vccd1 vccd1 _1821_/Y sky130_fd_sc_hd__nand3_2
X_1752_ _1752_/A _1767_/A vssd1 vssd1 vccd1 vccd1 _1752_/Y sky130_fd_sc_hd__nand2_1
X_1683_ _1683_/A vssd1 vssd1 vccd1 vccd1 _1683_/Y sky130_fd_sc_hd__inv_2
X_2166_ _2298_/CLK _2166_/D vssd1 vssd1 vccd1 vccd1 _2166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2235_ _2292_/CLK _2235_/D vssd1 vssd1 vccd1 vccd1 _2235_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2097_ _1672_/A _2153_/Q _2161_/Q _2193_/Q _2258_/Q _2259_/Q vssd1 vssd1 vccd1 vccd1
+ _2097_/X sky130_fd_sc_hd__mux4_2
X_1117_ _1140_/A vssd1 vssd1 vccd1 vccd1 _1125_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1048_ input4/X vssd1 vssd1 vccd1 vccd1 _1203_/B sky130_fd_sc_hd__inv_2
XFILLER_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2020_ _1780_/Y _2019_/X _2293_/Q vssd1 vssd1 vccd1 vccd1 _2020_/X sky130_fd_sc_hd__mux2_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1735_ _1743_/A _1975_/X vssd1 vssd1 vccd1 vccd1 _1735_/Y sky130_fd_sc_hd__nand2_1
X_1666_ _2091_/X vssd1 vssd1 vccd1 vccd1 _1666_/Y sky130_fd_sc_hd__inv_2
X_1804_ _2172_/Q vssd1 vssd1 vccd1 vccd1 _1804_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1597_ _2103_/X _1597_/B vssd1 vssd1 vccd1 vccd1 _1597_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2218_ _2219_/CLK _2218_/D vssd1 vssd1 vccd1 vccd1 _2218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2149_ _2275_/CLK _2149_/D vssd1 vssd1 vccd1 vccd1 _2149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput308 _1941_/X vssd1 vssd1 vccd1 vccd1 io_wo[63] sky130_fd_sc_hd__clkbuf_2
X_1520_ _2185_/Q _1981_/X _1522_/S vssd1 vssd1 vccd1 vccd1 _2185_/D sky130_fd_sc_hd__mux2_1
X_1451_ _2195_/Q vssd1 vssd1 vccd1 vccd1 _1451_/Y sky130_fd_sc_hd__inv_2
X_1382_ _1376_/X _1380_/Y _1381_/Y vssd1 vssd1 vccd1 vccd1 _1430_/B sky130_fd_sc_hd__o21bai_2
XFILLER_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2003_ _2003_/A0 _1802_/X _2268_/Q vssd1 vssd1 vccd1 vccd1 _2003_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1718_ _2209_/Q vssd1 vssd1 vccd1 vccd1 _1718_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1649_ _2099_/X _1649_/B vssd1 vssd1 vccd1 vccd1 _1649_/X sky130_fd_sc_hd__xor2_1
XFILLER_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2226_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1503_ _1503_/A _1503_/B vssd1 vssd1 vccd1 vccd1 _1503_/Y sky130_fd_sc_hd__xnor2_1
X_1434_ _1381_/Y _1376_/X _1380_/Y _1525_/S vssd1 vssd1 vccd1 vccd1 _1434_/Y sky130_fd_sc_hd__o31ai_1
X_1365_ _1374_/S vssd1 vssd1 vccd1 vccd1 _1372_/S sky130_fd_sc_hd__buf_2
X_1296_ _1989_/X _2030_/X vssd1 vssd1 vccd1 vccd1 _1296_/Y sky130_fd_sc_hd__nor2_4
XPHY_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 io_dat_i[8] vssd1 vssd1 vccd1 vccd1 _1085_/A sky130_fd_sc_hd__clkbuf_1
Xinput29 io_eo[18] vssd1 vssd1 vccd1 vccd1 _1896_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_37_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1150_ _2263_/Q _1143_/X _1148_/X _1149_/Y vssd1 vssd1 vccd1 vccd1 _2263_/D sky130_fd_sc_hd__o211a_1
X_1081_ _2286_/Q _1077_/X _1069_/X _1080_/Y vssd1 vssd1 vccd1 vccd1 _2286_/D sky130_fd_sc_hd__o211a_1
XFILLER_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1983_ _1710_/Y _1982_/X _2249_/Q vssd1 vssd1 vccd1 vccd1 _1983_/X sky130_fd_sc_hd__mux2_2
X_1417_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1431_/S sky130_fd_sc_hd__buf_2
XFILLER_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1279_ _1278_/X _2231_/Q _1281_/S vssd1 vssd1 vccd1 vccd1 _2231_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1348_ _1348_/A _1348_/B vssd1 vssd1 vccd1 vccd1 _1348_/Y sky130_fd_sc_hd__xnor2_1
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2251_ _2251_/CLK _2251_/D vssd1 vssd1 vccd1 vccd1 _2251_/Q sky130_fd_sc_hd__dfxtp_4
X_2182_ _2297_/CLK _2182_/D vssd1 vssd1 vccd1 vccd1 _2182_/Q sky130_fd_sc_hd__dfxtp_1
X_1064_ _1056_/X _1071_/B _1166_/B vssd1 vssd1 vccd1 vccd1 _1064_/Y sky130_fd_sc_hd__nand3b_1
X_1202_ _1202_/A vssd1 vssd1 vccd1 vccd1 _1203_/C sky130_fd_sc_hd__clkbuf_2
X_1133_ _1138_/A _1180_/B vssd1 vssd1 vccd1 vccd1 _1133_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1966_ _1662_/Y _1661_/Y _2250_/Q vssd1 vssd1 vccd1 vccd1 _1966_/X sky130_fd_sc_hd__mux2_1
X_1897_ _1897_/A vssd1 vssd1 vccd1 vccd1 _1897_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1820_ _1850_/A vssd1 vssd1 vccd1 vccd1 _1821_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_15_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1751_ _2202_/Q vssd1 vssd1 vccd1 vccd1 _1751_/Y sky130_fd_sc_hd__inv_2
X_1682_ _2082_/X vssd1 vssd1 vccd1 vccd1 _1682_/Y sky130_fd_sc_hd__inv_2
X_2234_ _2292_/CLK _2234_/D vssd1 vssd1 vccd1 vccd1 _2234_/Q sky130_fd_sc_hd__dfxtp_2
X_2165_ _2298_/CLK _2165_/D vssd1 vssd1 vccd1 vccd1 _2165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1047_ _2292_/Q vssd1 vssd1 vccd1 vccd1 _1821_/A sky130_fd_sc_hd__buf_2
X_2096_ _1667_/A _2154_/Q _2162_/Q _2194_/Q _2258_/Q _2259_/Q vssd1 vssd1 vccd1 vccd1
+ _2096_/X sky130_fd_sc_hd__mux4_2
X_1116_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1116_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_15_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2195_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1949_ _1870_/Y _1948_/X _2285_/Q vssd1 vssd1 vccd1 vccd1 _1949_/X sky130_fd_sc_hd__mux2_4
XFILLER_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1803_ _1803_/A vssd1 vssd1 vccd1 vccd1 _1803_/Y sky130_fd_sc_hd__inv_2
X_1665_ _2171_/Q vssd1 vssd1 vccd1 vccd1 _1665_/Y sky130_fd_sc_hd__inv_2
X_1596_ _1594_/X _1207_/X _1569_/Y _1595_/X vssd1 vssd1 vccd1 vccd1 _2157_/D sky130_fd_sc_hd__a31o_1
X_1734_ _2230_/Q vssd1 vssd1 vccd1 vccd1 _1734_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2217_ _2219_/CLK _2217_/D vssd1 vssd1 vccd1 vccd1 _2217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2148_ _2275_/CLK _2148_/D vssd1 vssd1 vccd1 vccd1 _2148_/Q sky130_fd_sc_hd__dfxtp_1
X_2079_ _2079_/A0 _2206_/Q _2250_/Q vssd1 vssd1 vccd1 vccd1 _2079_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput309 _1884_/X vssd1 vssd1 vccd1 vccd1 io_wo[6] sky130_fd_sc_hd__clkbuf_2
X_1450_ _2196_/Q _1989_/X _1450_/S vssd1 vssd1 vccd1 vccd1 _2196_/D sky130_fd_sc_hd__mux2_1
X_1381_ _1973_/X _2051_/X vssd1 vssd1 vccd1 vccd1 _1381_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2002_ _2270_/Q _2001_/X _2271_/Q vssd1 vssd1 vccd1 vccd1 _2002_/X sky130_fd_sc_hd__mux2_1
X_1717_ _1729_/A _1981_/X vssd1 vssd1 vccd1 vccd1 _1717_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1579_ _1579_/A _1579_/B _2127_/X _1597_/B vssd1 vssd1 vccd1 vccd1 _1579_/X sky130_fd_sc_hd__and4_1
X_1648_ _1654_/C _2100_/X vssd1 vssd1 vccd1 vccd1 _1649_/B sky130_fd_sc_hd__and2b_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1433_ _1381_/Y _1376_/X _1380_/Y vssd1 vssd1 vccd1 vccd1 _1433_/X sky130_fd_sc_hd__o21a_1
X_1502_ _1505_/B _1505_/A _1501_/Y vssd1 vssd1 vccd1 vccd1 _1503_/B sky130_fd_sc_hd__a21oi_1
X_1364_ _2110_/X vssd1 vssd1 vccd1 vccd1 _1776_/A sky130_fd_sc_hd__inv_2
XFILLER_48_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1295_ _2010_/X vssd1 vssd1 vccd1 vccd1 _1295_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput19 io_dat_i[9] vssd1 vssd1 vccd1 vccd1 _1082_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_77_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1080_ _1078_/X _1090_/B _1177_/B vssd1 vssd1 vccd1 vccd1 _1080_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1982_ _1712_/Y _1711_/Y _2248_/Q vssd1 vssd1 vccd1 vccd1 _1982_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1416_ _1211_/X _1411_/Y _1415_/Y vssd1 vssd1 vccd1 vccd1 _2210_/D sky130_fd_sc_hd__o21ai_1
X_1347_ _1350_/B _1350_/A _1346_/X vssd1 vssd1 vccd1 vccd1 _1348_/B sky130_fd_sc_hd__a21oi_1
XPHY_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1278_ _1278_/A _1278_/B vssd1 vssd1 vccd1 vccd1 _1278_/X sky130_fd_sc_hd__xor2_1
XFILLER_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1201_ _2245_/Q _1189_/X _1193_/X _1200_/Y vssd1 vssd1 vccd1 vccd1 _2245_/D sky130_fd_sc_hd__o211a_1
X_2250_ _2254_/CLK _2250_/D vssd1 vssd1 vccd1 vccd1 _2250_/Q sky130_fd_sc_hd__dfxtp_4
X_2181_ _2297_/CLK _2181_/D vssd1 vssd1 vccd1 vccd1 _2181_/Q sky130_fd_sc_hd__dfxtp_1
X_1132_ _2270_/Q _1130_/X _1122_/X _1131_/Y vssd1 vssd1 vccd1 vccd1 _2270_/D sky130_fd_sc_hd__o211a_1
X_1063_ input9/X vssd1 vssd1 vccd1 vccd1 _1166_/B sky130_fd_sc_hd__inv_2
X_1965_ _1666_/Y _1964_/X _2251_/Q vssd1 vssd1 vccd1 vccd1 _1965_/X sky130_fd_sc_hd__mux2_2
X_1896_ _1896_/A vssd1 vssd1 vccd1 vccd1 _1896_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1750_ _1750_/A _1767_/A vssd1 vssd1 vccd1 vccd1 _1750_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1681_ _2168_/Q vssd1 vssd1 vccd1 vccd1 _1681_/Y sky130_fd_sc_hd__inv_2
X_2164_ _2298_/CLK _2164_/D vssd1 vssd1 vccd1 vccd1 _2164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2233_ _2292_/CLK _2233_/D vssd1 vssd1 vccd1 vccd1 _2233_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1046_ _2293_/Q _1029_/A _1043_/X _1045_/Y vssd1 vssd1 vccd1 vccd1 _2293_/D sky130_fd_sc_hd__o211a_1
X_2095_ _1661_/A _2155_/Q _2163_/Q _2195_/Q _2258_/Q _2259_/Q vssd1 vssd1 vccd1 vccd1
+ _2095_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1115_ _1140_/A vssd1 vssd1 vccd1 vccd1 _1155_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1948_ _1951_/X _2241_/Q _2284_/Q vssd1 vssd1 vccd1 vccd1 _1948_/X sky130_fd_sc_hd__mux2_1
X_1879_ _1879_/A vssd1 vssd1 vccd1 vccd1 _1879_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1802_ _1476_/Y _1801_/Y _1478_/Y _1481_/A vssd1 vssd1 vccd1 vccd1 _1802_/X sky130_fd_sc_hd__a31o_2
XPHY_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1733_ _1733_/A vssd1 vssd1 vccd1 vccd1 _1733_/Y sky130_fd_sc_hd__inv_2
X_1664_ _1685_/A _1967_/X vssd1 vssd1 vccd1 vccd1 _1664_/Y sky130_fd_sc_hd__nand2_1
X_1595_ _1207_/X _2157_/Q vssd1 vssd1 vccd1 vccd1 _1595_/X sky130_fd_sc_hd__and2b_1
X_2216_ _2219_/CLK _2216_/D vssd1 vssd1 vccd1 vccd1 _2216_/Q sky130_fd_sc_hd__dfxtp_1
X_2147_ _2291_/CLK _2147_/D vssd1 vssd1 vccd1 vccd1 _2147_/Q sky130_fd_sc_hd__dfxtp_1
X_2078_ _1691_/Y _2077_/X _2299_/Q vssd1 vssd1 vccd1 vccd1 _2078_/X sky130_fd_sc_hd__mux2_4
X_1029_ _1029_/A _1191_/B vssd1 vssd1 vccd1 vccd1 _1029_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1380_ _1377_/Y _1378_/Y _1436_/A vssd1 vssd1 vccd1 vccd1 _1380_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_4_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2001_ _2001_/A0 _1532_/Y _2270_/Q vssd1 vssd1 vccd1 vccd1 _2001_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1716_ _1716_/A vssd1 vssd1 vccd1 vccd1 _1716_/Y sky130_fd_sc_hd__inv_2
X_1647_ _1646_/X _2144_/Q _1647_/S vssd1 vssd1 vccd1 vccd1 _2144_/D sky130_fd_sc_hd__mux2_1
X_1578_ _2002_/X vssd1 vssd1 vccd1 vccd1 _1597_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_92_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1432_ _2205_/Q vssd1 vssd1 vccd1 vccd1 _1432_/Y sky130_fd_sc_hd__inv_2
X_1501_ _1957_/X _2078_/X vssd1 vssd1 vccd1 vccd1 _1501_/Y sky130_fd_sc_hd__nor2_1
X_1363_ _2218_/Q _1774_/A _1363_/S vssd1 vssd1 vccd1 vccd1 _2218_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1294_ _1989_/X _2030_/X vssd1 vssd1 vccd1 vccd1 _1355_/A sky130_fd_sc_hd__nand2_2
XFILLER_63_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1981_ _1715_/Y _1980_/X _2249_/Q vssd1 vssd1 vccd1 vccd1 _1981_/X sky130_fd_sc_hd__mux2_4
XFILLER_13_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1415_ _1413_/Y _1414_/X _1417_/A vssd1 vssd1 vccd1 vccd1 _1415_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1346_ _2036_/X _2113_/X vssd1 vssd1 vccd1 vccd1 _1346_/X sky130_fd_sc_hd__and2b_1
XPHY_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1277_ _1280_/A _1280_/B _1276_/X vssd1 vssd1 vccd1 vccd1 _1278_/B sky130_fd_sc_hd__o21bai_1
XFILLER_22_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2180_ _2297_/CLK _2180_/D vssd1 vssd1 vccd1 vccd1 _2180_/Q sky130_fd_sc_hd__dfxtp_1
X_1200_ _1158_/C _1200_/B _1200_/C vssd1 vssd1 vccd1 vccd1 _1200_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_92_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1062_ _2291_/Q _1055_/X _1043_/X _1061_/Y vssd1 vssd1 vccd1 vccd1 _2291_/D sky130_fd_sc_hd__o211a_1
X_1131_ _1138_/A _1177_/B vssd1 vssd1 vccd1 vccd1 _1131_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1895_ _1895_/A vssd1 vssd1 vccd1 vccd1 _1895_/X sky130_fd_sc_hd__clkbuf_2
X_1964_ _1668_/Y _1667_/Y _2250_/Q vssd1 vssd1 vccd1 vccd1 _1964_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1329_ _1319_/Y _1327_/Y _1330_/A vssd1 vssd1 vccd1 vccd1 _1332_/A sky130_fd_sc_hd__a21o_1
XPHY_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput290 _1925_/X vssd1 vssd1 vccd1 vccd1 io_wo[47] sky130_fd_sc_hd__clkbuf_2
XFILLER_58_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1680_ _2192_/Q vssd1 vssd1 vccd1 vccd1 _1680_/Y sky130_fd_sc_hd__inv_2
X_2232_ _2292_/CLK _2232_/D vssd1 vssd1 vccd1 vccd1 _2232_/Q sky130_fd_sc_hd__dfxtp_2
X_2163_ _2163_/CLK _2163_/D vssd1 vssd1 vccd1 vccd1 _2163_/Q sky130_fd_sc_hd__dfxtp_1
X_1114_ input2/X _1816_/A _1186_/A vssd1 vssd1 vccd1 vccd1 _1140_/A sky130_fd_sc_hd__nor3_4
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1045_ _1049_/A _1200_/B vssd1 vssd1 vccd1 vccd1 _1045_/Y sky130_fd_sc_hd__nand2_1
X_2094_ _2094_/A0 _2211_/Q _2250_/Q vssd1 vssd1 vccd1 vccd1 _2094_/X sky130_fd_sc_hd__mux2_1
X_1947_ _1874_/Y _1946_/X _2287_/Q vssd1 vssd1 vccd1 vccd1 _1947_/X sky130_fd_sc_hd__mux2_1
X_1878_ _1878_/A vssd1 vssd1 vccd1 vccd1 _1878_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1663_ _2298_/Q vssd1 vssd1 vccd1 vccd1 _1685_/A sky130_fd_sc_hd__clkbuf_2
X_1801_ _1801_/A vssd1 vssd1 vccd1 vccd1 _1801_/Y sky130_fd_sc_hd__inv_2
XPHY_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1732_ _2055_/X vssd1 vssd1 vccd1 vccd1 _1732_/Y sky130_fd_sc_hd__inv_2
X_1594_ _1579_/A _1597_/B _1579_/B vssd1 vssd1 vccd1 vccd1 _1594_/X sky130_fd_sc_hd__a21o_1
X_2077_ _1693_/Y _1692_/Y _2298_/Q vssd1 vssd1 vccd1 vccd1 _2077_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2215_ _2292_/CLK _2215_/D vssd1 vssd1 vccd1 vccd1 _2215_/Q sky130_fd_sc_hd__dfxtp_1
X_2146_ _2163_/CLK _2146_/D vssd1 vssd1 vccd1 vccd1 _2146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1028_ _1028_/A vssd1 vssd1 vccd1 vccd1 _1191_/B sky130_fd_sc_hd__inv_2
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2000_ _2272_/Q _1999_/X _2273_/Q vssd1 vssd1 vccd1 vccd1 _2000_/X sky130_fd_sc_hd__mux2_2
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1715_ _2064_/X vssd1 vssd1 vccd1 vccd1 _1715_/Y sky130_fd_sc_hd__inv_2
X_1646_ _1646_/A _1646_/B vssd1 vssd1 vccd1 vccd1 _1646_/X sky130_fd_sc_hd__xor2_1
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1577_ _1581_/A _2163_/Q _1572_/X _1576_/Y vssd1 vssd1 vccd1 vccd1 _2163_/D sky130_fd_sc_hd__o2bb2ai_1
XFILLER_41_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2129_ _2129_/A0 _2176_/Q _2192_/Q _2224_/Q _2254_/Q _2255_/Q vssd1 vssd1 vccd1 vccd1
+ _2129_/X sky130_fd_sc_hd__mux4_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1500_ _1499_/X _2192_/Q _1506_/S vssd1 vssd1 vccd1 vccd1 _2192_/D sky130_fd_sc_hd__mux2_1
X_1431_ _1430_/X _2206_/Q _1431_/S vssd1 vssd1 vccd1 vccd1 _2206_/D sky130_fd_sc_hd__mux2_1
X_1362_ _2111_/X vssd1 vssd1 vccd1 vccd1 _1774_/A sky130_fd_sc_hd__inv_2
X_1293_ _2118_/X _2046_/X vssd1 vssd1 vccd1 vccd1 _1327_/B sky130_fd_sc_hd__xnor2_1
XFILLER_48_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1629_ _1943_/X vssd1 vssd1 vccd1 vccd1 _1657_/S sky130_fd_sc_hd__inv_2
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1980_ _1266_/Y _1716_/Y _2248_/Q vssd1 vssd1 vccd1 vccd1 _1980_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1414_ _1414_/A _1414_/B _1414_/C vssd1 vssd1 vccd1 vccd1 _1414_/X sky130_fd_sc_hd__and3_1
X_1345_ _1344_/X _2224_/Q _1353_/S vssd1 vssd1 vccd1 vccd1 _2224_/D sky130_fd_sc_hd__mux2_1
X_1276_ _2018_/X _2107_/X vssd1 vssd1 vccd1 vccd1 _1276_/X sky130_fd_sc_hd__and2b_1
XPHY_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_1_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2268_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1130_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1130_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1061_ _1056_/X _1071_/B _1163_/B vssd1 vssd1 vccd1 vccd1 _1061_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1894_ _1894_/A vssd1 vssd1 vccd1 vccd1 _1894_/X sky130_fd_sc_hd__clkbuf_2
X_1963_ _1671_/Y _1962_/X _2251_/Q vssd1 vssd1 vccd1 vccd1 _1963_/X sky130_fd_sc_hd__mux2_4
XFILLER_83_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1259_ _1281_/S _2235_/Q vssd1 vssd1 vccd1 vccd1 _1260_/B sky130_fd_sc_hd__nand2_1
X_1328_ _1987_/X vssd1 vssd1 vccd1 vccd1 _1330_/A sky130_fd_sc_hd__inv_2
XFILLER_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput291 _1926_/X vssd1 vssd1 vccd1 vccd1 io_wo[48] sky130_fd_sc_hd__clkbuf_2
Xoutput280 _1916_/X vssd1 vssd1 vccd1 vccd1 io_wo[38] sky130_fd_sc_hd__clkbuf_2
XFILLER_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2231_ _2231_/CLK _2231_/D vssd1 vssd1 vccd1 vccd1 _2231_/Q sky130_fd_sc_hd__dfxtp_2
X_2093_ _1664_/Y _2092_/X _2299_/Q vssd1 vssd1 vccd1 vccd1 _2093_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2162_ _2254_/CLK _2162_/D vssd1 vssd1 vccd1 vccd1 _2162_/Q sky130_fd_sc_hd__dfxtp_1
X_1044_ _1044_/A vssd1 vssd1 vccd1 vccd1 _1200_/B sky130_fd_sc_hd__inv_2
X_1113_ input1/X vssd1 vssd1 vccd1 vccd1 _1816_/A sky130_fd_sc_hd__inv_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1946_ _1949_/X _2236_/Q _2286_/Q vssd1 vssd1 vccd1 vccd1 _1946_/X sky130_fd_sc_hd__mux2_1
X_1877_ _2299_/Q _1029_/A _1088_/A _1876_/Y vssd1 vssd1 vccd1 vccd1 _2299_/D sky130_fd_sc_hd__o211a_1
XFILLER_9_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1800_ _1400_/Y _1799_/Y _1402_/Y _1405_/A vssd1 vssd1 vccd1 vccd1 _1811_/A sky130_fd_sc_hd__a31oi_4
XFILLER_62_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1731_ _2183_/Q vssd1 vssd1 vccd1 vccd1 _1731_/Y sky130_fd_sc_hd__inv_2
XPHY_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1662_ _2227_/Q vssd1 vssd1 vccd1 vccd1 _1662_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2214_ _2226_/CLK _2214_/D vssd1 vssd1 vccd1 vccd1 _2214_/Q sky130_fd_sc_hd__dfxtp_1
X_1593_ _1581_/A _1591_/Y _1579_/X _1592_/Y vssd1 vssd1 vccd1 vccd1 _2158_/D sky130_fd_sc_hd__o31ai_1
XFILLER_93_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1027_ _1700_/A _1020_/X _1023_/X _1026_/Y vssd1 vssd1 vccd1 vccd1 _2298_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2145_ _2163_/CLK _2145_/D vssd1 vssd1 vccd1 vccd1 _2145_/Q sky130_fd_sc_hd__dfxtp_1
X_2076_ _2076_/A0 _2205_/Q _2250_/Q vssd1 vssd1 vccd1 vccd1 _2076_/X sky130_fd_sc_hd__mux2_1
X_1929_ _1929_/A vssd1 vssd1 vccd1 vccd1 _1929_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_14_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2298_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1714_ _2186_/Q vssd1 vssd1 vccd1 vccd1 _1714_/Y sky130_fd_sc_hd__inv_2
X_1576_ _2132_/X _1574_/X _1598_/S vssd1 vssd1 vccd1 vccd1 _1576_/Y sky130_fd_sc_hd__o21bai_1
X_1645_ _1644_/X _2145_/Q _1647_/S vssd1 vssd1 vccd1 vccd1 _2145_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2059_ _1725_/Y _1724_/Y _2296_/Q vssd1 vssd1 vccd1 vccd1 _2059_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2128_ _2128_/A0 _2175_/Q _2191_/Q _2223_/Q _2254_/Q _2255_/Q vssd1 vssd1 vccd1 vccd1
+ _2128_/X sky130_fd_sc_hd__mux4_2
XFILLER_41_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1430_ _1430_/A _1430_/B vssd1 vssd1 vccd1 vccd1 _1430_/X sky130_fd_sc_hd__xor2_1
X_1361_ _2219_/Q _1772_/A _1363_/S vssd1 vssd1 vccd1 vccd1 _2219_/D sky130_fd_sc_hd__mux2_1
X_1292_ _1289_/X _1290_/Y _1216_/X _1291_/Y vssd1 vssd1 vccd1 vccd1 _2228_/D sky130_fd_sc_hd__o2bb2ai_1
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1559_ _2169_/Q _1963_/X _1561_/S vssd1 vssd1 vccd1 vccd1 _2169_/D sky130_fd_sc_hd__mux2_1
X_1628_ _1627_/Y _2148_/Q _1628_/S vssd1 vssd1 vccd1 vccd1 _2148_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1413_ _1414_/A _1414_/B _1414_/C vssd1 vssd1 vccd1 vccd1 _1413_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1275_ _2108_/X _2020_/X vssd1 vssd1 vccd1 vccd1 _1278_/A sky130_fd_sc_hd__xnor2_2
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1344_ _1344_/A _1344_/B vssd1 vssd1 vccd1 vccd1 _1344_/X sky130_fd_sc_hd__xor2_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1060_ _1060_/A vssd1 vssd1 vccd1 vccd1 _1163_/B sky130_fd_sc_hd__inv_2
X_1962_ _1339_/Y _1672_/Y _2250_/Q vssd1 vssd1 vccd1 vccd1 _1962_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1893_ _1893_/A vssd1 vssd1 vccd1 vccd1 _1893_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1258_ _1258_/A vssd1 vssd1 vccd1 vccd1 _1281_/S sky130_fd_sc_hd__buf_2
X_1327_ _1327_/A _1327_/B _1333_/A vssd1 vssd1 vccd1 vccd1 _1327_/Y sky130_fd_sc_hd__nand3_1
X_1189_ _1189_/A vssd1 vssd1 vccd1 vccd1 _1189_/X sky130_fd_sc_hd__clkbuf_2
XPHY_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput270 _1907_/X vssd1 vssd1 vccd1 vccd1 io_wo[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_3_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput292 _1927_/X vssd1 vssd1 vccd1 vccd1 io_wo[49] sky130_fd_sc_hd__clkbuf_2
Xoutput281 _1917_/X vssd1 vssd1 vccd1 vccd1 io_wo[39] sky130_fd_sc_hd__clkbuf_2
XFILLER_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2230_ _2231_/CLK _2230_/D vssd1 vssd1 vccd1 vccd1 _2230_/Q sky130_fd_sc_hd__dfxtp_2
X_2092_ _1665_/Y _1451_/Y _2298_/Q vssd1 vssd1 vccd1 vccd1 _2092_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1043_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1043_/X sky130_fd_sc_hd__clkbuf_2
X_1112_ _2276_/Q _1095_/A _1104_/X _1111_/Y vssd1 vssd1 vccd1 vccd1 _2276_/D sky130_fd_sc_hd__o211a_1
X_2161_ _2163_/CLK _2161_/D vssd1 vssd1 vccd1 vccd1 _2161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1945_ _1873_/Y _1944_/X _2289_/Q vssd1 vssd1 vccd1 vccd1 _1945_/X sky130_fd_sc_hd__mux2_4
XFILLER_9_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1876_ _1158_/C _1876_/B _1876_/C vssd1 vssd1 vccd1 vccd1 _1876_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1730_ _2207_/Q vssd1 vssd1 vccd1 vccd1 _1730_/Y sky130_fd_sc_hd__inv_2
X_1661_ _1661_/A vssd1 vssd1 vccd1 vccd1 _1661_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1592_ _1598_/S _2158_/Q vssd1 vssd1 vccd1 vccd1 _1592_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2213_ _2226_/CLK _2213_/D vssd1 vssd1 vccd1 vccd1 _2213_/Q sky130_fd_sc_hd__dfxtp_1
X_2144_ _2163_/CLK _2144_/D vssd1 vssd1 vccd1 vccd1 _2144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2075_ _1696_/Y _2074_/X _2299_/Q vssd1 vssd1 vccd1 vccd1 _2075_/X sky130_fd_sc_hd__mux2_1
X_1026_ _1029_/A _1187_/B vssd1 vssd1 vccd1 vccd1 _1026_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1928_ _1928_/A vssd1 vssd1 vccd1 vccd1 _1928_/X sky130_fd_sc_hd__clkbuf_2
X_1859_ _2255_/Q _1855_/X _1858_/X _2287_/Q vssd1 vssd1 vccd1 vccd1 _1859_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1713_ _1729_/A _1983_/X vssd1 vssd1 vccd1 vccd1 _1713_/Y sky130_fd_sc_hd__nand2_1
XPHY_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1575_ _1575_/A vssd1 vssd1 vccd1 vccd1 _1598_/S sky130_fd_sc_hd__clkbuf_2
X_1644_ _2097_/X _1644_/B vssd1 vssd1 vccd1 vccd1 _1644_/X sky130_fd_sc_hd__xor2_1
XFILLER_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2127_ _2127_/A0 _2174_/Q _2190_/Q _2222_/Q _2254_/Q _2255_/Q vssd1 vssd1 vccd1 vccd1
+ _2127_/X sky130_fd_sc_hd__mux4_2
XFILLER_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2058_ _2058_/A0 _2223_/Q _2248_/Q vssd1 vssd1 vccd1 vccd1 _2058_/X sky130_fd_sc_hd__mux2_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1360_ _2112_/X vssd1 vssd1 vccd1 vccd1 _1772_/A sky130_fd_sc_hd__inv_2
XFILLER_48_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1291_ _2228_/Q vssd1 vssd1 vccd1 vccd1 _1291_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1489_ _1489_/A _1489_/B vssd1 vssd1 vccd1 vccd1 _1491_/C sky130_fd_sc_hd__nor2_1
X_1558_ _2170_/Q _1965_/X _1561_/S vssd1 vssd1 vccd1 vccd1 _2170_/D sky130_fd_sc_hd__mux2_1
X_1627_ _2102_/X _2000_/X vssd1 vssd1 vccd1 vccd1 _1627_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1412_ _1412_/A _1412_/B vssd1 vssd1 vccd1 vccd1 _1414_/C sky130_fd_sc_hd__nor2_1
X_1343_ _1342_/B _1339_/Y _1342_/Y vssd1 vssd1 vccd1 vccd1 _2225_/D sky130_fd_sc_hd__o21ai_1
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1274_ _1272_/X _1363_/S _1269_/B _1273_/X vssd1 vssd1 vccd1 vccd1 _2232_/D sky130_fd_sc_hd__a31o_1
XFILLER_51_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1892_ _1892_/A vssd1 vssd1 vccd1 vccd1 _1892_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1961_ _1676_/Y _1960_/X _2251_/Q vssd1 vssd1 vccd1 vccd1 _1961_/X sky130_fd_sc_hd__mux2_8
XFILLER_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1326_ _1326_/A _1333_/B _1326_/C vssd1 vssd1 vccd1 vccd1 _1327_/A sky130_fd_sc_hd__nand3_1
X_1257_ _1993_/X vssd1 vssd1 vccd1 vccd1 _1258_/A sky130_fd_sc_hd__inv_2
X_1188_ _2250_/Q _1175_/X _1179_/X _1187_/Y vssd1 vssd1 vccd1 vccd1 _2250_/D sky130_fd_sc_hd__o211a_1
XPHY_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput293 _1882_/X vssd1 vssd1 vccd1 vccd1 io_wo[4] sky130_fd_sc_hd__clkbuf_2
Xoutput282 _1881_/X vssd1 vssd1 vccd1 vccd1 io_wo[3] sky130_fd_sc_hd__clkbuf_2
Xoutput260 _1879_/X vssd1 vssd1 vccd1 vccd1 io_wo[1] sky130_fd_sc_hd__clkbuf_2
Xoutput271 _1880_/X vssd1 vssd1 vccd1 vccd1 io_wo[2] sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_0 _2001_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2160_ _2163_/CLK _2160_/D vssd1 vssd1 vccd1 vccd1 _2160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1042_ _1760_/B _1020_/X _1023_/X _1041_/Y vssd1 vssd1 vccd1 vccd1 _2294_/D sky130_fd_sc_hd__o211a_1
X_1111_ _1110_/X _1111_/B _1203_/B vssd1 vssd1 vccd1 vccd1 _1111_/Y sky130_fd_sc_hd__nand3b_1
X_2091_ _2091_/A0 _2210_/Q _2250_/Q vssd1 vssd1 vccd1 vccd1 _2091_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1944_ _1947_/X _2242_/Q _2288_/Q vssd1 vssd1 vccd1 vccd1 _1944_/X sky130_fd_sc_hd__mux2_1
X_1875_ _1875_/A _2290_/Q vssd1 vssd1 vccd1 vccd1 _1875_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2289_ _2291_/CLK _2289_/D vssd1 vssd1 vccd1 vccd1 _2289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1309_ _1309_/A _1320_/A _1341_/A vssd1 vssd1 vccd1 vccd1 _1334_/A sky130_fd_sc_hd__nand3_4
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1660_ _2094_/X vssd1 vssd1 vccd1 vccd1 _1660_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1591_ _1579_/A _1579_/B _1597_/B _2127_/X vssd1 vssd1 vccd1 vccd1 _1591_/Y sky130_fd_sc_hd__a31oi_1
X_2212_ _2226_/CLK _2212_/D vssd1 vssd1 vccd1 vccd1 _2212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2143_ _2275_/CLK _2143_/D vssd1 vssd1 vccd1 vccd1 _2143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2074_ _1697_/Y _1507_/Y _2298_/Q vssd1 vssd1 vccd1 vccd1 _2074_/X sky130_fd_sc_hd__mux2_1
X_1025_ _1025_/A vssd1 vssd1 vccd1 vccd1 _1187_/B sky130_fd_sc_hd__inv_2
X_1927_ _1927_/A vssd1 vssd1 vccd1 vccd1 _1927_/X sky130_fd_sc_hd__clkbuf_2
X_1858_ _1858_/A vssd1 vssd1 vccd1 vccd1 _1858_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1789_ _1789_/A vssd1 vssd1 vccd1 vccd1 _1789_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1712_ _2234_/Q vssd1 vssd1 vccd1 vccd1 _1712_/Y sky130_fd_sc_hd__inv_2
X_1643_ _1642_/X _2146_/Q _1647_/S vssd1 vssd1 vccd1 vccd1 _2146_/D sky130_fd_sc_hd__mux2_1
XPHY_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1574_ _1573_/Y _2131_/X _2129_/X _2130_/X vssd1 vssd1 vccd1 vccd1 _1574_/X sky130_fd_sc_hd__and4b_1
X_2057_ _1729_/Y _2056_/X _2297_/Q vssd1 vssd1 vccd1 vccd1 _2057_/X sky130_fd_sc_hd__mux2_2
XFILLER_81_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2126_ _1754_/Y _1550_/Y _1507_/Y _1757_/Y _2254_/Q _2255_/Q vssd1 vssd1 vccd1 vccd1
+ _2126_/X sky130_fd_sc_hd__mux4_2
XFILLER_25_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1290_ _1287_/Y _1288_/Y _1223_/X _1281_/S vssd1 vssd1 vccd1 vccd1 _1290_/Y sky130_fd_sc_hd__a31oi_1
X_1626_ _1624_/X _1945_/X _1622_/B _1625_/X vssd1 vssd1 vccd1 vccd1 _2149_/D sky130_fd_sc_hd__a31o_1
X_1557_ _2171_/Q _1967_/X _1561_/S vssd1 vssd1 vccd1 vccd1 _2171_/D sky130_fd_sc_hd__mux2_1
X_1488_ _2194_/Q vssd1 vssd1 vccd1 vccd1 _1488_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2109_ input89/X _1677_/A _1721_/A _2122_/A0 _2244_/Q _2245_/Q vssd1 vssd1 vccd1
+ vccd1 _2109_/X sky130_fd_sc_hd__mux4_2
XFILLER_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1411_ _2210_/Q vssd1 vssd1 vccd1 vccd1 _1411_/Y sky130_fd_sc_hd__inv_2
X_1273_ _1374_/S _2232_/Q vssd1 vssd1 vccd1 vccd1 _1273_/X sky130_fd_sc_hd__and2b_1
X_1342_ _1342_/A _1342_/B vssd1 vssd1 vccd1 vccd1 _1342_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1609_ _1616_/A _2155_/Q vssd1 vssd1 vccd1 vccd1 _1609_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1891_ _1891_/A vssd1 vssd1 vccd1 vccd1 _1891_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1960_ _1678_/Y _1677_/Y _2250_/Q vssd1 vssd1 vccd1 vccd1 _1960_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1256_ _1256_/A _1363_/S vssd1 vssd1 vccd1 vccd1 _1260_/A sky130_fd_sc_hd__nand2_1
X_1325_ _1344_/A _1344_/B _1324_/Y vssd1 vssd1 vccd1 vccd1 _1326_/A sky130_fd_sc_hd__o21bai_1
XFILLER_91_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1187_ _1186_/X _1187_/B _1187_/C vssd1 vssd1 vccd1 vccd1 _1187_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput294 _1928_/X vssd1 vssd1 vccd1 vccd1 io_wo[50] sky130_fd_sc_hd__clkbuf_2
Xoutput283 _1918_/X vssd1 vssd1 vccd1 vccd1 io_wo[40] sky130_fd_sc_hd__clkbuf_2
Xoutput272 _1908_/X vssd1 vssd1 vccd1 vccd1 io_wo[30] sky130_fd_sc_hd__clkbuf_2
Xoutput261 _1898_/X vssd1 vssd1 vccd1 vccd1 io_wo[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput250 _1888_/X vssd1 vssd1 vccd1 vccd1 io_wo[10] sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_1 _1999_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2090_ _1669_/Y _2089_/X _2299_/Q vssd1 vssd1 vccd1 vccd1 _2090_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1110_ _1110_/A vssd1 vssd1 vccd1 vccd1 _1110_/X sky130_fd_sc_hd__buf_1
X_1041_ _1049_/A _1198_/B vssd1 vssd1 vccd1 vccd1 _1041_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2231_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1874_ _1875_/A _2286_/Q vssd1 vssd1 vccd1 vccd1 _1874_/Y sky130_fd_sc_hd__nand2_1
X_1943_ _1875_/Y _1942_/X _2291_/Q vssd1 vssd1 vccd1 vccd1 _1943_/X sky130_fd_sc_hd__mux2_4
XFILLER_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1239_ _1239_/A _1239_/B vssd1 vssd1 vccd1 vccd1 _1240_/B sky130_fd_sc_hd__nor2_1
X_2288_ _2299_/CLK _2288_/D vssd1 vssd1 vccd1 vccd1 _2288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1308_ _2116_/X _2042_/X vssd1 vssd1 vccd1 vccd1 _1341_/A sky130_fd_sc_hd__xnor2_2
XFILLER_28_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1590_ _1573_/Y _1588_/X _1207_/X _1589_/X vssd1 vssd1 vccd1 vccd1 _2159_/D sky130_fd_sc_hd__a31o_1
XFILLER_93_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2211_ _2219_/CLK _2211_/D vssd1 vssd1 vccd1 vccd1 _2211_/Q sky130_fd_sc_hd__dfxtp_2
X_1024_ _1032_/A vssd1 vssd1 vccd1 vccd1 _1029_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2073_ _2073_/A0 _2204_/Q _2250_/Q vssd1 vssd1 vccd1 vccd1 _2073_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2142_ _2275_/CLK _2142_/D vssd1 vssd1 vccd1 vccd1 _2142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1926_ _1926_/A vssd1 vssd1 vccd1 vccd1 _1926_/X sky130_fd_sc_hd__clkbuf_2
X_1857_ _2270_/Q _1849_/X _1850_/X _1856_/X vssd1 vssd1 vccd1 vccd1 _1857_/X sky130_fd_sc_hd__a31o_1
X_1788_ _2260_/Q vssd1 vssd1 vccd1 vccd1 _1788_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1711_ _1711_/A vssd1 vssd1 vccd1 vccd1 _1711_/Y sky130_fd_sc_hd__inv_2
X_1642_ _2096_/X _1642_/B vssd1 vssd1 vccd1 vccd1 _1642_/X sky130_fd_sc_hd__xor2_1
XPHY_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ _1569_/Y _2127_/X _2128_/X vssd1 vssd1 vccd1 vccd1 _1573_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2056_ _1731_/Y _1730_/Y _2296_/Q vssd1 vssd1 vccd1 vccd1 _2056_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2125_ _2125_/A0 _2195_/Q _2211_/Q _2235_/Q _2252_/Q _2253_/Q vssd1 vssd1 vccd1 vccd1
+ _2125_/X sky130_fd_sc_hd__mux4_2
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1909_ _1909_/A vssd1 vssd1 vccd1 vccd1 _1909_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput150 io_i_7_in1[2] vssd1 vssd1 vccd1 vccd1 _1689_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1556_ _1951_/X vssd1 vssd1 vccd1 vccd1 _1561_/S sky130_fd_sc_hd__buf_2
X_1625_ _1945_/X _2149_/Q vssd1 vssd1 vccd1 vccd1 _1625_/X sky130_fd_sc_hd__and2b_1
X_1487_ _1209_/X _1451_/Y _1486_/Y vssd1 vssd1 vccd1 vccd1 _2195_/D sky130_fd_sc_hd__o21ai_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2039_ _1756_/Y _1678_/Y _2294_/Q vssd1 vssd1 vccd1 vccd1 _2039_/X sky130_fd_sc_hd__mux2_1
X_2108_ input88/X _1683_/A _1727_/A _2121_/A0 _2244_/Q _2245_/Q vssd1 vssd1 vccd1
+ vccd1 _2108_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_4_13_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2291_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1410_ _1211_/X _1375_/Y _1409_/Y vssd1 vssd1 vccd1 vccd1 _2211_/D sky130_fd_sc_hd__o21ai_1
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1272_ _1236_/A _1236_/C _1236_/B vssd1 vssd1 vccd1 vccd1 _1272_/X sky130_fd_sc_hd__a21o_1
X_1341_ _1341_/A _1341_/B vssd1 vssd1 vccd1 vccd1 _1342_/A sky130_fd_sc_hd__xor2_1
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1608_ _1608_/A vssd1 vssd1 vccd1 vccd1 _1608_/X sky130_fd_sc_hd__clkbuf_2
X_1539_ _1539_/A _2120_/X _2004_/X _2119_/X vssd1 vssd1 vccd1 vccd1 _1545_/B sky130_fd_sc_hd__and4_1
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1890_ _1890_/A vssd1 vssd1 vccd1 vccd1 _1890_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1255_ _1374_/S vssd1 vssd1 vccd1 vccd1 _1363_/S sky130_fd_sc_hd__clkbuf_2
X_1324_ _2042_/X _1752_/A _1755_/A _2040_/X vssd1 vssd1 vccd1 vccd1 _1324_/Y sky130_fd_sc_hd__o22ai_1
X_1186_ _1186_/A vssd1 vssd1 vccd1 vccd1 _1186_/X sky130_fd_sc_hd__buf_1
XFILLER_33_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput295 _1929_/X vssd1 vssd1 vccd1 vccd1 io_wo[51] sky130_fd_sc_hd__clkbuf_2
Xoutput284 _1919_/X vssd1 vssd1 vccd1 vccd1 io_wo[41] sky130_fd_sc_hd__clkbuf_2
Xoutput273 _1909_/X vssd1 vssd1 vccd1 vccd1 io_wo[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_74_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput262 _1899_/X vssd1 vssd1 vccd1 vccd1 io_wo[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput251 _1889_/X vssd1 vssd1 vccd1 vccd1 io_wo[11] sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_2 _2235_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput240 _2140_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1040_ _1040_/A vssd1 vssd1 vccd1 vccd1 _1198_/B sky130_fd_sc_hd__inv_2
XFILLER_73_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1942_ _1945_/X _2243_/Q _2290_/Q vssd1 vssd1 vccd1 vccd1 _1942_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1873_ _1875_/A _2288_/Q vssd1 vssd1 vccd1 vccd1 _1873_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1238_ _2024_/X _2110_/X vssd1 vssd1 vccd1 vccd1 _1239_/B sky130_fd_sc_hd__and2b_1
XFILLER_64_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2287_ _2291_/CLK _2287_/D vssd1 vssd1 vccd1 vccd1 _2287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1169_ _2257_/Q _1159_/X _1165_/X _1168_/Y vssd1 vssd1 vccd1 vccd1 _2257_/D sky130_fd_sc_hd__o211a_1
XFILLER_44_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1307_ _2115_/X _2040_/X vssd1 vssd1 vccd1 vccd1 _1320_/A sky130_fd_sc_hd__xnor2_2
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2210_ _2219_/CLK _2210_/D vssd1 vssd1 vccd1 vccd1 _2210_/Q sky130_fd_sc_hd__dfxtp_2
X_2072_ _1700_/Y _2071_/X _2299_/Q vssd1 vssd1 vccd1 vccd1 _2072_/X sky130_fd_sc_hd__mux2_2
X_1023_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1023_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2141_ _2275_/CLK _2141_/D vssd1 vssd1 vccd1 vccd1 _2141_/Q sky130_fd_sc_hd__dfxtp_1
X_1925_ _1925_/A vssd1 vssd1 vccd1 vccd1 _1925_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1856_ _2254_/Q _1855_/X _1111_/B _2286_/Q vssd1 vssd1 vccd1 vccd1 _1856_/X sky130_fd_sc_hd__a22o_1
X_1787_ _2212_/Q vssd1 vssd1 vccd1 vccd1 _1787_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1710_ _2067_/X vssd1 vssd1 vccd1 vccd1 _1710_/Y sky130_fd_sc_hd__inv_2
X_1641_ _1646_/A _1646_/B _2097_/X vssd1 vssd1 vccd1 vccd1 _1642_/B sky130_fd_sc_hd__nor3b_4
X_1572_ _1572_/A vssd1 vssd1 vccd1 vccd1 _1572_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2124_ _2124_/A0 _2194_/Q _2210_/Q _2234_/Q _2252_/Q _2253_/Q vssd1 vssd1 vccd1 vccd1
+ _2124_/X sky130_fd_sc_hd__mux4_2
XFILLER_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2055_ _2055_/A0 _2222_/Q _2248_/Q vssd1 vssd1 vccd1 vccd1 _2055_/X sky130_fd_sc_hd__mux2_1
X_1908_ _1908_/A vssd1 vssd1 vccd1 vccd1 _1908_/X sky130_fd_sc_hd__clkbuf_2
X_1839_ _1839_/A _1850_/A _2249_/Q vssd1 vssd1 vccd1 vccd1 _1839_/Y sky130_fd_sc_hd__nor3b_2
XFILLER_72_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput140 io_i_6_in1[1] vssd1 vssd1 vccd1 vccd1 _1658_/A sky130_fd_sc_hd__buf_1
Xinput151 io_i_7_in1[3] vssd1 vssd1 vccd1 vccd1 _1683_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1555_ _1554_/Y _2172_/Q _1555_/S vssd1 vssd1 vccd1 vccd1 _2172_/D sky130_fd_sc_hd__mux2_1
X_1624_ _1611_/B _2000_/X _2133_/X vssd1 vssd1 vccd1 vccd1 _1624_/X sky130_fd_sc_hd__a21bo_1
X_1486_ _1482_/Y _1483_/X _1506_/S vssd1 vssd1 vccd1 vccd1 _1486_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_54_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2107_ input87/X _1689_/A _1733_/A _2120_/A0 _2244_/Q _2245_/Q vssd1 vssd1 vccd1
+ vccd1 _2107_/X sky130_fd_sc_hd__mux4_2
XFILLER_62_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2038_ _1758_/Y _2037_/X _2295_/Q vssd1 vssd1 vccd1 vccd1 _2038_/X sky130_fd_sc_hd__mux2_4
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1340_ _1344_/A _1344_/B _1313_/X vssd1 vssd1 vccd1 vccd1 _1341_/B sky130_fd_sc_hd__o21bai_1
X_1271_ _1216_/X _1266_/Y _1270_/X vssd1 vssd1 vccd1 vccd1 _2233_/D sky130_fd_sc_hd__o21ai_1
XFILLER_36_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1469_ _1963_/X _2087_/X vssd1 vssd1 vccd1 vccd1 _1470_/B sky130_fd_sc_hd__and2_1
X_1607_ _1607_/A _2137_/X _2138_/X _2139_/X vssd1 vssd1 vccd1 vccd1 _1608_/A sky130_fd_sc_hd__and4_1
X_1538_ _2104_/X vssd1 vssd1 vccd1 vccd1 _1539_/A sky130_fd_sc_hd__inv_2
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1323_ _2115_/X vssd1 vssd1 vccd1 vccd1 _1755_/A sky130_fd_sc_hd__inv_2
X_1254_ _1254_/A _1254_/B vssd1 vssd1 vccd1 vccd1 _1256_/A sky130_fd_sc_hd__nand2_1
X_1185_ _2251_/Q _1175_/X _1179_/X _1184_/Y vssd1 vssd1 vccd1 vccd1 _2251_/D sky130_fd_sc_hd__o211a_1
Xoutput252 _1890_/X vssd1 vssd1 vccd1 vccd1 io_wo[12] sky130_fd_sc_hd__clkbuf_2
Xoutput230 _1608_/X vssd1 vssd1 vccd1 vccd1 io_o_6_co sky130_fd_sc_hd__clkbuf_2
Xoutput241 _2141_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput296 _1930_/X vssd1 vssd1 vccd1 vccd1 io_wo[52] sky130_fd_sc_hd__clkbuf_2
Xoutput285 _1920_/X vssd1 vssd1 vccd1 vccd1 io_wo[42] sky130_fd_sc_hd__clkbuf_2
Xoutput274 _1910_/X vssd1 vssd1 vccd1 vccd1 io_wo[32] sky130_fd_sc_hd__clkbuf_2
Xoutput263 _1900_/X vssd1 vssd1 vccd1 vccd1 io_wo[22] sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_3 _1890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1941_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1941_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1872_ _1996_/X vssd1 vssd1 vccd1 vccd1 _1872_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2286_ _2299_/CLK _2286_/D vssd1 vssd1 vccd1 vccd1 _2286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1306_ _1350_/B _1350_/A _1348_/A _1305_/Y vssd1 vssd1 vccd1 vccd1 _1309_/A sky130_fd_sc_hd__a31o_1
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1237_ _2022_/X _2109_/X vssd1 vssd1 vccd1 vccd1 _1239_/A sky130_fd_sc_hd__and2b_2
X_1099_ _1096_/X _1105_/B _1194_/B vssd1 vssd1 vccd1 vccd1 _1099_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1168_ _1110_/X _1168_/B _1173_/C vssd1 vssd1 vccd1 vccd1 _1168_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2140_ _2275_/CLK _2140_/D vssd1 vssd1 vccd1 vccd1 _2140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2071_ _1701_/Y _1512_/Y _2298_/Q vssd1 vssd1 vccd1 vccd1 _2071_/X sky130_fd_sc_hd__mux2_1
X_1022_ _1193_/A vssd1 vssd1 vccd1 vccd1 _1088_/A sky130_fd_sc_hd__buf_1
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1924_ _1924_/A vssd1 vssd1 vccd1 vccd1 _1924_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1855_ _1855_/A vssd1 vssd1 vccd1 vccd1 _1855_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1786_ _1786_/A _1821_/A vssd1 vssd1 vccd1 vccd1 _1786_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2269_ _2272_/CLK _2269_/D vssd1 vssd1 vccd1 vccd1 _2269_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1640_ _2147_/Q _1647_/S _1637_/X _1639_/Y vssd1 vssd1 vccd1 vccd1 _2147_/D sky130_fd_sc_hd__o2bb2ai_1
X_1571_ _1583_/B _2131_/X _2132_/X _2130_/X vssd1 vssd1 vccd1 vccd1 _1572_/A sky130_fd_sc_hd__and4_1
XFILLER_6_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2123_ _2123_/A0 _2193_/Q _2209_/Q _2233_/Q _2252_/Q _2253_/Q vssd1 vssd1 vccd1 vccd1
+ _2123_/X sky130_fd_sc_hd__mux4_2
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2054_ _1735_/Y _2053_/X _2297_/Q vssd1 vssd1 vccd1 vccd1 _2054_/X sky130_fd_sc_hd__mux2_2
XFILLER_81_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1907_ _1907_/A vssd1 vssd1 vccd1 vccd1 _1907_/X sky130_fd_sc_hd__clkbuf_2
X_1838_ _1743_/A _1824_/X _2280_/Q _1825_/X _1837_/Y vssd1 vssd1 vccd1 vccd1 _1838_/X
+ sky130_fd_sc_hd__a221o_1
X_1769_ _2262_/Q vssd1 vssd1 vccd1 vccd1 _1769_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput152 io_i_7_in1[4] vssd1 vssd1 vccd1 vccd1 _1677_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput130 io_i_5_in1[0] vssd1 vssd1 vccd1 vccd1 _1766_/A sky130_fd_sc_hd__clkbuf_1
Xinput141 io_i_6_in1[2] vssd1 vssd1 vccd1 vccd1 _1733_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1485_ _1485_/A vssd1 vssd1 vccd1 vccd1 _1506_/S sky130_fd_sc_hd__clkbuf_2
X_1554_ _2104_/X _2004_/X vssd1 vssd1 vccd1 vccd1 _1554_/Y sky130_fd_sc_hd__xnor2_1
X_1623_ _1622_/Y _2150_/Q _1628_/S vssd1 vssd1 vccd1 vccd1 _2150_/D sky130_fd_sc_hd__mux2_1
.ends

