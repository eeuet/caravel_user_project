* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for cic_block abstract view
.subckt cic_block io_adr_i[0] io_adr_i[1] io_cs_i io_dat_i[0] io_dat_i[10] io_dat_i[11]
+ io_dat_i[12] io_dat_i[13] io_dat_i[14] io_dat_i[15] io_dat_i[1] io_dat_i[2] io_dat_i[3]
+ io_dat_i[4] io_dat_i[5] io_dat_i[6] io_dat_i[7] io_dat_i[8] io_dat_i[9] io_dat_o[0]
+ io_dat_o[10] io_dat_o[11] io_dat_o[12] io_dat_o[13] io_dat_o[14] io_dat_o[15] io_dat_o[1]
+ io_dat_o[2] io_dat_o[3] io_dat_o[4] io_dat_o[5] io_dat_o[6] io_dat_o[7] io_dat_o[8]
+ io_dat_o[9] io_eo[0] io_eo[10] io_eo[11] io_eo[12] io_eo[13] io_eo[14] io_eo[15]
+ io_eo[16] io_eo[17] io_eo[18] io_eo[19] io_eo[1] io_eo[20] io_eo[21] io_eo[22] io_eo[23]
+ io_eo[24] io_eo[25] io_eo[26] io_eo[27] io_eo[28] io_eo[29] io_eo[2] io_eo[30] io_eo[31]
+ io_eo[32] io_eo[33] io_eo[34] io_eo[35] io_eo[36] io_eo[37] io_eo[38] io_eo[39]
+ io_eo[3] io_eo[40] io_eo[41] io_eo[42] io_eo[43] io_eo[44] io_eo[45] io_eo[46] io_eo[47]
+ io_eo[48] io_eo[49] io_eo[4] io_eo[50] io_eo[51] io_eo[52] io_eo[53] io_eo[54] io_eo[55]
+ io_eo[56] io_eo[57] io_eo[58] io_eo[59] io_eo[5] io_eo[60] io_eo[61] io_eo[62] io_eo[63]
+ io_eo[6] io_eo[7] io_eo[8] io_eo[9] io_i_0_ci io_i_0_in1[0] io_i_0_in1[1] io_i_0_in1[2]
+ io_i_0_in1[3] io_i_0_in1[4] io_i_0_in1[5] io_i_0_in1[6] io_i_0_in1[7] io_i_1_ci
+ io_i_1_in1[0] io_i_1_in1[1] io_i_1_in1[2] io_i_1_in1[3] io_i_1_in1[4] io_i_1_in1[5]
+ io_i_1_in1[6] io_i_1_in1[7] io_i_2_ci io_i_2_in1[0] io_i_2_in1[1] io_i_2_in1[2]
+ io_i_2_in1[3] io_i_2_in1[4] io_i_2_in1[5] io_i_2_in1[6] io_i_2_in1[7] io_i_3_ci
+ io_i_3_in1[0] io_i_3_in1[1] io_i_3_in1[2] io_i_3_in1[3] io_i_3_in1[4] io_i_3_in1[5]
+ io_i_3_in1[6] io_i_3_in1[7] io_i_4_ci io_i_4_in1[0] io_i_4_in1[1] io_i_4_in1[2]
+ io_i_4_in1[3] io_i_4_in1[4] io_i_4_in1[5] io_i_4_in1[6] io_i_4_in1[7] io_i_5_ci
+ io_i_5_in1[0] io_i_5_in1[1] io_i_5_in1[2] io_i_5_in1[3] io_i_5_in1[4] io_i_5_in1[5]
+ io_i_5_in1[6] io_i_5_in1[7] io_i_6_ci io_i_6_in1[0] io_i_6_in1[1] io_i_6_in1[2]
+ io_i_6_in1[3] io_i_6_in1[4] io_i_6_in1[5] io_i_6_in1[6] io_i_6_in1[7] io_i_7_ci
+ io_i_7_in1[0] io_i_7_in1[1] io_i_7_in1[2] io_i_7_in1[3] io_i_7_in1[4] io_i_7_in1[5]
+ io_i_7_in1[6] io_i_7_in1[7] io_o_0_co io_o_0_out[0] io_o_0_out[1] io_o_0_out[2]
+ io_o_0_out[3] io_o_0_out[4] io_o_0_out[5] io_o_0_out[6] io_o_0_out[7] io_o_1_co
+ io_o_1_out[0] io_o_1_out[1] io_o_1_out[2] io_o_1_out[3] io_o_1_out[4] io_o_1_out[5]
+ io_o_1_out[6] io_o_1_out[7] io_o_2_co io_o_2_out[0] io_o_2_out[1] io_o_2_out[2]
+ io_o_2_out[3] io_o_2_out[4] io_o_2_out[5] io_o_2_out[6] io_o_2_out[7] io_o_3_co
+ io_o_3_out[0] io_o_3_out[1] io_o_3_out[2] io_o_3_out[3] io_o_3_out[4] io_o_3_out[5]
+ io_o_3_out[6] io_o_3_out[7] io_o_4_co io_o_4_out[0] io_o_4_out[1] io_o_4_out[2]
+ io_o_4_out[3] io_o_4_out[4] io_o_4_out[5] io_o_4_out[6] io_o_4_out[7] io_o_5_co
+ io_o_5_out[0] io_o_5_out[1] io_o_5_out[2] io_o_5_out[3] io_o_5_out[4] io_o_5_out[5]
+ io_o_5_out[6] io_o_5_out[7] io_o_6_co io_o_6_out[0] io_o_6_out[1] io_o_6_out[2]
+ io_o_6_out[3] io_o_6_out[4] io_o_6_out[5] io_o_6_out[6] io_o_6_out[7] io_o_7_co
+ io_o_7_out[0] io_o_7_out[1] io_o_7_out[2] io_o_7_out[3] io_o_7_out[4] io_o_7_out[5]
+ io_o_7_out[6] io_o_7_out[7] io_vci io_vco io_vi io_we_i io_wo[0] io_wo[10] io_wo[11]
+ io_wo[12] io_wo[13] io_wo[14] io_wo[15] io_wo[16] io_wo[17] io_wo[18] io_wo[19]
+ io_wo[1] io_wo[20] io_wo[21] io_wo[22] io_wo[23] io_wo[24] io_wo[25] io_wo[26] io_wo[27]
+ io_wo[28] io_wo[29] io_wo[2] io_wo[30] io_wo[31] io_wo[32] io_wo[33] io_wo[34] io_wo[35]
+ io_wo[36] io_wo[37] io_wo[38] io_wo[39] io_wo[3] io_wo[40] io_wo[41] io_wo[42] io_wo[43]
+ io_wo[44] io_wo[45] io_wo[46] io_wo[47] io_wo[48] io_wo[49] io_wo[4] io_wo[50] io_wo[51]
+ io_wo[52] io_wo[53] io_wo[54] io_wo[55] io_wo[56] io_wo[57] io_wo[58] io_wo[59]
+ io_wo[5] io_wo[60] io_wo[61] io_wo[62] io_wo[63] io_wo[6] io_wo[7] io_wo[8] io_wo[9]
+ wb_clk_i wb_rst_i vccd1 vssd1
.ends

* Black-box entry subcircuit for motor_top abstract view
.subckt motor_top clock io_QEI_ChA io_QEI_ChB io_irq io_pwm_h io_pwm_l io_wb_ack_o
+ io_wb_adr_i[0] io_wb_adr_i[10] io_wb_adr_i[11] io_wb_adr_i[1] io_wb_adr_i[2] io_wb_adr_i[3]
+ io_wb_adr_i[4] io_wb_adr_i[5] io_wb_adr_i[6] io_wb_adr_i[7] io_wb_adr_i[8] io_wb_adr_i[9]
+ io_wb_cs_i io_wb_dat_i[0] io_wb_dat_i[10] io_wb_dat_i[11] io_wb_dat_i[12] io_wb_dat_i[13]
+ io_wb_dat_i[14] io_wb_dat_i[15] io_wb_dat_i[16] io_wb_dat_i[17] io_wb_dat_i[18]
+ io_wb_dat_i[19] io_wb_dat_i[1] io_wb_dat_i[20] io_wb_dat_i[21] io_wb_dat_i[22] io_wb_dat_i[23]
+ io_wb_dat_i[24] io_wb_dat_i[25] io_wb_dat_i[26] io_wb_dat_i[27] io_wb_dat_i[28]
+ io_wb_dat_i[29] io_wb_dat_i[2] io_wb_dat_i[30] io_wb_dat_i[31] io_wb_dat_i[3] io_wb_dat_i[4]
+ io_wb_dat_i[5] io_wb_dat_i[6] io_wb_dat_i[7] io_wb_dat_i[8] io_wb_dat_i[9] io_wb_dat_o[0]
+ io_wb_dat_o[10] io_wb_dat_o[11] io_wb_dat_o[12] io_wb_dat_o[13] io_wb_dat_o[14]
+ io_wb_dat_o[15] io_wb_dat_o[16] io_wb_dat_o[17] io_wb_dat_o[18] io_wb_dat_o[19]
+ io_wb_dat_o[1] io_wb_dat_o[20] io_wb_dat_o[21] io_wb_dat_o[22] io_wb_dat_o[23] io_wb_dat_o[24]
+ io_wb_dat_o[25] io_wb_dat_o[26] io_wb_dat_o[27] io_wb_dat_o[28] io_wb_dat_o[29]
+ io_wb_dat_o[2] io_wb_dat_o[30] io_wb_dat_o[31] io_wb_dat_o[3] io_wb_dat_o[4] io_wb_dat_o[5]
+ io_wb_dat_o[6] io_wb_dat_o[7] io_wb_dat_o[8] io_wb_dat_o[9] io_wb_we_i reset vccd1
+ vssd1
.ends

* Black-box entry subcircuit for sin3 abstract view
.subckt sin3 ao_reg[0] ao_reg[10] ao_reg[11] ao_reg[12] ao_reg[13] ao_reg[14] ao_reg[15]
+ ao_reg[16] ao_reg[17] ao_reg[18] ao_reg[19] ao_reg[1] ao_reg[20] ao_reg[21] ao_reg[22]
+ ao_reg[23] ao_reg[24] ao_reg[25] ao_reg[26] ao_reg[27] ao_reg[28] ao_reg[29] ao_reg[2]
+ ao_reg[30] ao_reg[31] ao_reg[3] ao_reg[4] ao_reg[5] ao_reg[6] ao_reg[7] ao_reg[8]
+ ao_reg[9] asel bo_reg[0] bo_reg[10] bo_reg[11] bo_reg[12] bo_reg[13] bo_reg[14]
+ bo_reg[15] bo_reg[16] bo_reg[17] bo_reg[18] bo_reg[19] bo_reg[1] bo_reg[20] bo_reg[21]
+ bo_reg[22] bo_reg[23] bo_reg[24] bo_reg[25] bo_reg[26] bo_reg[27] bo_reg[28] bo_reg[29]
+ bo_reg[2] bo_reg[30] bo_reg[31] bo_reg[3] bo_reg[4] bo_reg[5] bo_reg[6] bo_reg[7]
+ bo_reg[8] bo_reg[9] clk e_i[0] e_i[10] e_i[11] e_i[12] e_i[13] e_i[14] e_i[15] e_i[16]
+ e_i[17] e_i[18] e_i[19] e_i[1] e_i[20] e_i[21] e_i[22] e_i[23] e_i[24] e_i[25] e_i[26]
+ e_i[27] e_i[28] e_i[29] e_i[2] e_i[30] e_i[31] e_i[3] e_i[4] e_i[5] e_i[6] e_i[7]
+ e_i[8] e_i[9] e_o[0] e_o[10] e_o[11] e_o[12] e_o[13] e_o[14] e_o[15] e_o[16] e_o[17]
+ e_o[18] e_o[19] e_o[1] e_o[20] e_o[21] e_o[22] e_o[23] e_o[24] e_o[25] e_o[26] e_o[27]
+ e_o[28] e_o[29] e_o[2] e_o[30] e_o[31] e_o[3] e_o[4] e_o[5] e_o[6] e_o[7] e_o[8]
+ e_o[9] se_i[0] se_i[10] se_i[11] se_i[12] se_i[13] se_i[14] se_i[15] se_i[16] se_i[17]
+ se_i[18] se_i[19] se_i[1] se_i[20] se_i[21] se_i[22] se_i[23] se_i[24] se_i[25]
+ se_i[26] se_i[27] se_i[28] se_i[29] se_i[2] se_i[30] se_i[31] se_i[3] se_i[4] se_i[5]
+ se_i[6] se_i[7] se_i[8] se_i[9] se_o[0] se_o[10] se_o[11] se_o[12] se_o[13] se_o[14]
+ se_o[15] se_o[16] se_o[17] se_o[18] se_o[19] se_o[1] se_o[20] se_o[21] se_o[22]
+ se_o[23] se_o[24] se_o[25] se_o[26] se_o[27] se_o[28] se_o[29] se_o[2] se_o[30]
+ se_o[31] se_o[3] se_o[4] se_o[5] se_o[6] se_o[7] se_o[8] se_o[9] sw_i[0] sw_i[10]
+ sw_i[11] sw_i[12] sw_i[13] sw_i[14] sw_i[15] sw_i[16] sw_i[17] sw_i[18] sw_i[19]
+ sw_i[1] sw_i[20] sw_i[21] sw_i[22] sw_i[23] sw_i[24] sw_i[25] sw_i[26] sw_i[27]
+ sw_i[28] sw_i[29] sw_i[2] sw_i[30] sw_i[31] sw_i[3] sw_i[4] sw_i[5] sw_i[6] sw_i[7]
+ sw_i[8] sw_i[9] sw_o[0] sw_o[10] sw_o[11] sw_o[12] sw_o[13] sw_o[14] sw_o[15] sw_o[16]
+ sw_o[17] sw_o[18] sw_o[19] sw_o[1] sw_o[20] sw_o[21] sw_o[22] sw_o[23] sw_o[24]
+ sw_o[25] sw_o[26] sw_o[27] sw_o[28] sw_o[29] sw_o[2] sw_o[30] sw_o[31] sw_o[3] sw_o[4]
+ sw_o[5] sw_o[6] sw_o[7] sw_o[8] sw_o[9] w_i[0] w_i[10] w_i[11] w_i[12] w_i[13] w_i[14]
+ w_i[15] w_i[16] w_i[17] w_i[18] w_i[19] w_i[1] w_i[20] w_i[21] w_i[22] w_i[23] w_i[24]
+ w_i[25] w_i[26] w_i[27] w_i[28] w_i[29] w_i[2] w_i[30] w_i[31] w_i[3] w_i[4] w_i[5]
+ w_i[6] w_i[7] w_i[8] w_i[9] w_o[0] w_o[10] w_o[11] w_o[12] w_o[13] w_o[14] w_o[15]
+ w_o[16] w_o[17] w_o[18] w_o[19] w_o[1] w_o[20] w_o[21] w_o[22] w_o[23] w_o[24] w_o[25]
+ w_o[26] w_o[27] w_o[28] w_o[29] w_o[2] w_o[30] w_o[31] w_o[3] w_o[4] w_o[5] w_o[6]
+ w_o[7] w_o[8] w_o[9] vccd1 vssd1
.ends

* Black-box entry subcircuit for cic_con abstract view
.subckt cic_con io_ack_o io_adr_i[0] io_adr_i[10] io_adr_i[11] io_adr_i[1] io_adr_i[2]
+ io_adr_i[3] io_adr_i[4] io_adr_i[5] io_adr_i[6] io_adr_i[7] io_adr_i[8] io_adr_i[9]
+ io_b_adr_i[0] io_b_adr_i[1] io_b_cs_i_0 io_b_cs_i_1 io_b_cs_i_10 io_b_cs_i_2 io_b_cs_i_3
+ io_b_cs_i_4 io_b_cs_i_5 io_b_cs_i_6 io_b_cs_i_7 io_b_cs_i_8 io_b_cs_i_9 io_b_dat_i[0]
+ io_b_dat_i[10] io_b_dat_i[11] io_b_dat_i[12] io_b_dat_i[13] io_b_dat_i[14] io_b_dat_i[15]
+ io_b_dat_i[1] io_b_dat_i[2] io_b_dat_i[3] io_b_dat_i[4] io_b_dat_i[5] io_b_dat_i[6]
+ io_b_dat_i[7] io_b_dat_i[8] io_b_dat_i[9] io_b_dat_o_0[0] io_b_dat_o_0[10] io_b_dat_o_0[11]
+ io_b_dat_o_0[12] io_b_dat_o_0[13] io_b_dat_o_0[14] io_b_dat_o_0[15] io_b_dat_o_0[1]
+ io_b_dat_o_0[2] io_b_dat_o_0[3] io_b_dat_o_0[4] io_b_dat_o_0[5] io_b_dat_o_0[6]
+ io_b_dat_o_0[7] io_b_dat_o_0[8] io_b_dat_o_0[9] io_b_dat_o_10[0] io_b_dat_o_10[10]
+ io_b_dat_o_10[11] io_b_dat_o_10[12] io_b_dat_o_10[13] io_b_dat_o_10[14] io_b_dat_o_10[15]
+ io_b_dat_o_10[1] io_b_dat_o_10[2] io_b_dat_o_10[3] io_b_dat_o_10[4] io_b_dat_o_10[5]
+ io_b_dat_o_10[6] io_b_dat_o_10[7] io_b_dat_o_10[8] io_b_dat_o_10[9] io_b_dat_o_1[0]
+ io_b_dat_o_1[10] io_b_dat_o_1[11] io_b_dat_o_1[12] io_b_dat_o_1[13] io_b_dat_o_1[14]
+ io_b_dat_o_1[15] io_b_dat_o_1[1] io_b_dat_o_1[2] io_b_dat_o_1[3] io_b_dat_o_1[4]
+ io_b_dat_o_1[5] io_b_dat_o_1[6] io_b_dat_o_1[7] io_b_dat_o_1[8] io_b_dat_o_1[9]
+ io_b_dat_o_2[0] io_b_dat_o_2[10] io_b_dat_o_2[11] io_b_dat_o_2[12] io_b_dat_o_2[13]
+ io_b_dat_o_2[14] io_b_dat_o_2[15] io_b_dat_o_2[1] io_b_dat_o_2[2] io_b_dat_o_2[3]
+ io_b_dat_o_2[4] io_b_dat_o_2[5] io_b_dat_o_2[6] io_b_dat_o_2[7] io_b_dat_o_2[8]
+ io_b_dat_o_2[9] io_b_dat_o_3[0] io_b_dat_o_3[10] io_b_dat_o_3[11] io_b_dat_o_3[12]
+ io_b_dat_o_3[13] io_b_dat_o_3[14] io_b_dat_o_3[15] io_b_dat_o_3[1] io_b_dat_o_3[2]
+ io_b_dat_o_3[3] io_b_dat_o_3[4] io_b_dat_o_3[5] io_b_dat_o_3[6] io_b_dat_o_3[7]
+ io_b_dat_o_3[8] io_b_dat_o_3[9] io_b_dat_o_4[0] io_b_dat_o_4[10] io_b_dat_o_4[11]
+ io_b_dat_o_4[12] io_b_dat_o_4[13] io_b_dat_o_4[14] io_b_dat_o_4[15] io_b_dat_o_4[1]
+ io_b_dat_o_4[2] io_b_dat_o_4[3] io_b_dat_o_4[4] io_b_dat_o_4[5] io_b_dat_o_4[6]
+ io_b_dat_o_4[7] io_b_dat_o_4[8] io_b_dat_o_4[9] io_b_dat_o_5[0] io_b_dat_o_5[10]
+ io_b_dat_o_5[11] io_b_dat_o_5[12] io_b_dat_o_5[13] io_b_dat_o_5[14] io_b_dat_o_5[15]
+ io_b_dat_o_5[1] io_b_dat_o_5[2] io_b_dat_o_5[3] io_b_dat_o_5[4] io_b_dat_o_5[5]
+ io_b_dat_o_5[6] io_b_dat_o_5[7] io_b_dat_o_5[8] io_b_dat_o_5[9] io_b_dat_o_6[0]
+ io_b_dat_o_6[10] io_b_dat_o_6[11] io_b_dat_o_6[12] io_b_dat_o_6[13] io_b_dat_o_6[14]
+ io_b_dat_o_6[15] io_b_dat_o_6[1] io_b_dat_o_6[2] io_b_dat_o_6[3] io_b_dat_o_6[4]
+ io_b_dat_o_6[5] io_b_dat_o_6[6] io_b_dat_o_6[7] io_b_dat_o_6[8] io_b_dat_o_6[9]
+ io_b_dat_o_7[0] io_b_dat_o_7[10] io_b_dat_o_7[11] io_b_dat_o_7[12] io_b_dat_o_7[13]
+ io_b_dat_o_7[14] io_b_dat_o_7[15] io_b_dat_o_7[1] io_b_dat_o_7[2] io_b_dat_o_7[3]
+ io_b_dat_o_7[4] io_b_dat_o_7[5] io_b_dat_o_7[6] io_b_dat_o_7[7] io_b_dat_o_7[8]
+ io_b_dat_o_7[9] io_b_dat_o_8[0] io_b_dat_o_8[10] io_b_dat_o_8[11] io_b_dat_o_8[12]
+ io_b_dat_o_8[13] io_b_dat_o_8[14] io_b_dat_o_8[15] io_b_dat_o_8[1] io_b_dat_o_8[2]
+ io_b_dat_o_8[3] io_b_dat_o_8[4] io_b_dat_o_8[5] io_b_dat_o_8[6] io_b_dat_o_8[7]
+ io_b_dat_o_8[8] io_b_dat_o_8[9] io_b_dat_o_9[0] io_b_dat_o_9[10] io_b_dat_o_9[11]
+ io_b_dat_o_9[12] io_b_dat_o_9[13] io_b_dat_o_9[14] io_b_dat_o_9[15] io_b_dat_o_9[1]
+ io_b_dat_o_9[2] io_b_dat_o_9[3] io_b_dat_o_9[4] io_b_dat_o_9[5] io_b_dat_o_9[6]
+ io_b_dat_o_9[7] io_b_dat_o_9[8] io_b_dat_o_9[9] io_b_we_i io_cs_i io_dat_i[0] io_dat_i[10]
+ io_dat_i[11] io_dat_i[12] io_dat_i[13] io_dat_i[14] io_dat_i[15] io_dat_i[16] io_dat_i[17]
+ io_dat_i[18] io_dat_i[19] io_dat_i[1] io_dat_i[20] io_dat_i[21] io_dat_i[22] io_dat_i[23]
+ io_dat_i[24] io_dat_i[25] io_dat_i[26] io_dat_i[27] io_dat_i[28] io_dat_i[29] io_dat_i[2]
+ io_dat_i[30] io_dat_i[31] io_dat_i[3] io_dat_i[4] io_dat_i[5] io_dat_i[6] io_dat_i[7]
+ io_dat_i[8] io_dat_i[9] io_dat_o[0] io_dat_o[10] io_dat_o[11] io_dat_o[12] io_dat_o[13]
+ io_dat_o[14] io_dat_o[15] io_dat_o[16] io_dat_o[17] io_dat_o[18] io_dat_o[19] io_dat_o[1]
+ io_dat_o[20] io_dat_o[21] io_dat_o[22] io_dat_o[23] io_dat_o[24] io_dat_o[25] io_dat_o[26]
+ io_dat_o[27] io_dat_o[28] io_dat_o[29] io_dat_o[2] io_dat_o[30] io_dat_o[31] io_dat_o[3]
+ io_dat_o[4] io_dat_o[5] io_dat_o[6] io_dat_o[7] io_dat_o[8] io_dat_o[9] io_dataLastBlock[0]
+ io_dataLastBlock[10] io_dataLastBlock[11] io_dataLastBlock[12] io_dataLastBlock[13]
+ io_dataLastBlock[14] io_dataLastBlock[15] io_dataLastBlock[16] io_dataLastBlock[17]
+ io_dataLastBlock[18] io_dataLastBlock[19] io_dataLastBlock[1] io_dataLastBlock[20]
+ io_dataLastBlock[21] io_dataLastBlock[22] io_dataLastBlock[23] io_dataLastBlock[24]
+ io_dataLastBlock[25] io_dataLastBlock[26] io_dataLastBlock[27] io_dataLastBlock[28]
+ io_dataLastBlock[29] io_dataLastBlock[2] io_dataLastBlock[30] io_dataLastBlock[31]
+ io_dataLastBlock[32] io_dataLastBlock[33] io_dataLastBlock[34] io_dataLastBlock[35]
+ io_dataLastBlock[36] io_dataLastBlock[37] io_dataLastBlock[38] io_dataLastBlock[39]
+ io_dataLastBlock[3] io_dataLastBlock[40] io_dataLastBlock[41] io_dataLastBlock[42]
+ io_dataLastBlock[43] io_dataLastBlock[44] io_dataLastBlock[45] io_dataLastBlock[46]
+ io_dataLastBlock[47] io_dataLastBlock[48] io_dataLastBlock[49] io_dataLastBlock[4]
+ io_dataLastBlock[50] io_dataLastBlock[51] io_dataLastBlock[52] io_dataLastBlock[53]
+ io_dataLastBlock[54] io_dataLastBlock[55] io_dataLastBlock[56] io_dataLastBlock[57]
+ io_dataLastBlock[58] io_dataLastBlock[59] io_dataLastBlock[5] io_dataLastBlock[60]
+ io_dataLastBlock[61] io_dataLastBlock[62] io_dataLastBlock[63] io_dataLastBlock[6]
+ io_dataLastBlock[7] io_dataLastBlock[8] io_dataLastBlock[9] io_dsi_in[0] io_dsi_in[1]
+ io_dsi_in[2] io_dsi_in[3] io_dsi_in[4] io_dsi_in[5] io_dsi_in[6] io_dsi_in[7] io_dsi_o
+ io_irq io_vout[0] io_vout[10] io_vout[1] io_vout[2] io_vout[3] io_vout[4] io_vout[5]
+ io_vout[6] io_vout[7] io_vout[8] io_vout[9] io_we_i wb_clk_i wb_rst_i vccd1 vssd1
.ends

* Black-box entry subcircuit for wb_local abstract view
.subckt wb_local dsi[0] dsi[1] dsi[2] dsi[3] dsi[4] dsi[5] dsi[6] dsi[7] io_in[0]
+ io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] irq[0] irq[1] irq[2]
+ m_irqs[0] m_irqs[10] m_irqs[11] m_irqs[1] m_irqs[2] m_irqs[3] m_irqs[4] m_irqs[5]
+ m_irqs[6] m_irqs[7] m_irqs[8] m_irqs[9] m_wb_clk_i m_wb_rst_i m_wbs_ack_o[0] m_wbs_ack_o[10]
+ m_wbs_ack_o[11] m_wbs_ack_o[1] m_wbs_ack_o[2] m_wbs_ack_o[3] m_wbs_ack_o[4] m_wbs_ack_o[5]
+ m_wbs_ack_o[6] m_wbs_ack_o[7] m_wbs_ack_o[8] m_wbs_ack_o[9] m_wbs_adr_i[0] m_wbs_adr_i[10]
+ m_wbs_adr_i[11] m_wbs_adr_i[1] m_wbs_adr_i[2] m_wbs_adr_i[3] m_wbs_adr_i[4] m_wbs_adr_i[5]
+ m_wbs_adr_i[6] m_wbs_adr_i[7] m_wbs_adr_i[8] m_wbs_adr_i[9] m_wbs_cs_i[0] m_wbs_cs_i[10]
+ m_wbs_cs_i[11] m_wbs_cs_i[1] m_wbs_cs_i[2] m_wbs_cs_i[3] m_wbs_cs_i[4] m_wbs_cs_i[5]
+ m_wbs_cs_i[6] m_wbs_cs_i[7] m_wbs_cs_i[8] m_wbs_cs_i[9] m_wbs_dat_i[0] m_wbs_dat_i[10]
+ m_wbs_dat_i[11] m_wbs_dat_i[12] m_wbs_dat_i[13] m_wbs_dat_i[14] m_wbs_dat_i[15]
+ m_wbs_dat_i[16] m_wbs_dat_i[17] m_wbs_dat_i[18] m_wbs_dat_i[19] m_wbs_dat_i[1] m_wbs_dat_i[20]
+ m_wbs_dat_i[21] m_wbs_dat_i[22] m_wbs_dat_i[23] m_wbs_dat_i[24] m_wbs_dat_i[25]
+ m_wbs_dat_i[26] m_wbs_dat_i[27] m_wbs_dat_i[28] m_wbs_dat_i[29] m_wbs_dat_i[2] m_wbs_dat_i[30]
+ m_wbs_dat_i[31] m_wbs_dat_i[3] m_wbs_dat_i[4] m_wbs_dat_i[5] m_wbs_dat_i[6] m_wbs_dat_i[7]
+ m_wbs_dat_i[8] m_wbs_dat_i[9] m_wbs_dat_o_0[0] m_wbs_dat_o_0[10] m_wbs_dat_o_0[11]
+ m_wbs_dat_o_0[12] m_wbs_dat_o_0[13] m_wbs_dat_o_0[14] m_wbs_dat_o_0[15] m_wbs_dat_o_0[16]
+ m_wbs_dat_o_0[17] m_wbs_dat_o_0[18] m_wbs_dat_o_0[19] m_wbs_dat_o_0[1] m_wbs_dat_o_0[20]
+ m_wbs_dat_o_0[21] m_wbs_dat_o_0[22] m_wbs_dat_o_0[23] m_wbs_dat_o_0[24] m_wbs_dat_o_0[25]
+ m_wbs_dat_o_0[26] m_wbs_dat_o_0[27] m_wbs_dat_o_0[28] m_wbs_dat_o_0[29] m_wbs_dat_o_0[2]
+ m_wbs_dat_o_0[30] m_wbs_dat_o_0[31] m_wbs_dat_o_0[3] m_wbs_dat_o_0[4] m_wbs_dat_o_0[5]
+ m_wbs_dat_o_0[6] m_wbs_dat_o_0[7] m_wbs_dat_o_0[8] m_wbs_dat_o_0[9] m_wbs_dat_o_10[0]
+ m_wbs_dat_o_10[10] m_wbs_dat_o_10[11] m_wbs_dat_o_10[12] m_wbs_dat_o_10[13] m_wbs_dat_o_10[14]
+ m_wbs_dat_o_10[15] m_wbs_dat_o_10[16] m_wbs_dat_o_10[17] m_wbs_dat_o_10[18] m_wbs_dat_o_10[19]
+ m_wbs_dat_o_10[1] m_wbs_dat_o_10[20] m_wbs_dat_o_10[21] m_wbs_dat_o_10[22] m_wbs_dat_o_10[23]
+ m_wbs_dat_o_10[24] m_wbs_dat_o_10[25] m_wbs_dat_o_10[26] m_wbs_dat_o_10[27] m_wbs_dat_o_10[28]
+ m_wbs_dat_o_10[29] m_wbs_dat_o_10[2] m_wbs_dat_o_10[30] m_wbs_dat_o_10[31] m_wbs_dat_o_10[3]
+ m_wbs_dat_o_10[4] m_wbs_dat_o_10[5] m_wbs_dat_o_10[6] m_wbs_dat_o_10[7] m_wbs_dat_o_10[8]
+ m_wbs_dat_o_10[9] m_wbs_dat_o_11[0] m_wbs_dat_o_11[10] m_wbs_dat_o_11[11] m_wbs_dat_o_11[12]
+ m_wbs_dat_o_11[13] m_wbs_dat_o_11[14] m_wbs_dat_o_11[15] m_wbs_dat_o_11[16] m_wbs_dat_o_11[17]
+ m_wbs_dat_o_11[18] m_wbs_dat_o_11[19] m_wbs_dat_o_11[1] m_wbs_dat_o_11[20] m_wbs_dat_o_11[21]
+ m_wbs_dat_o_11[22] m_wbs_dat_o_11[23] m_wbs_dat_o_11[24] m_wbs_dat_o_11[25] m_wbs_dat_o_11[26]
+ m_wbs_dat_o_11[27] m_wbs_dat_o_11[28] m_wbs_dat_o_11[29] m_wbs_dat_o_11[2] m_wbs_dat_o_11[30]
+ m_wbs_dat_o_11[31] m_wbs_dat_o_11[3] m_wbs_dat_o_11[4] m_wbs_dat_o_11[5] m_wbs_dat_o_11[6]
+ m_wbs_dat_o_11[7] m_wbs_dat_o_11[8] m_wbs_dat_o_11[9] m_wbs_dat_o_1[0] m_wbs_dat_o_1[10]
+ m_wbs_dat_o_1[11] m_wbs_dat_o_1[12] m_wbs_dat_o_1[13] m_wbs_dat_o_1[14] m_wbs_dat_o_1[15]
+ m_wbs_dat_o_1[16] m_wbs_dat_o_1[17] m_wbs_dat_o_1[18] m_wbs_dat_o_1[19] m_wbs_dat_o_1[1]
+ m_wbs_dat_o_1[20] m_wbs_dat_o_1[21] m_wbs_dat_o_1[22] m_wbs_dat_o_1[23] m_wbs_dat_o_1[24]
+ m_wbs_dat_o_1[25] m_wbs_dat_o_1[26] m_wbs_dat_o_1[27] m_wbs_dat_o_1[28] m_wbs_dat_o_1[29]
+ m_wbs_dat_o_1[2] m_wbs_dat_o_1[30] m_wbs_dat_o_1[31] m_wbs_dat_o_1[3] m_wbs_dat_o_1[4]
+ m_wbs_dat_o_1[5] m_wbs_dat_o_1[6] m_wbs_dat_o_1[7] m_wbs_dat_o_1[8] m_wbs_dat_o_1[9]
+ m_wbs_dat_o_2[0] m_wbs_dat_o_2[10] m_wbs_dat_o_2[11] m_wbs_dat_o_2[12] m_wbs_dat_o_2[13]
+ m_wbs_dat_o_2[14] m_wbs_dat_o_2[15] m_wbs_dat_o_2[16] m_wbs_dat_o_2[17] m_wbs_dat_o_2[18]
+ m_wbs_dat_o_2[19] m_wbs_dat_o_2[1] m_wbs_dat_o_2[20] m_wbs_dat_o_2[21] m_wbs_dat_o_2[22]
+ m_wbs_dat_o_2[23] m_wbs_dat_o_2[24] m_wbs_dat_o_2[25] m_wbs_dat_o_2[26] m_wbs_dat_o_2[27]
+ m_wbs_dat_o_2[28] m_wbs_dat_o_2[29] m_wbs_dat_o_2[2] m_wbs_dat_o_2[30] m_wbs_dat_o_2[31]
+ m_wbs_dat_o_2[3] m_wbs_dat_o_2[4] m_wbs_dat_o_2[5] m_wbs_dat_o_2[6] m_wbs_dat_o_2[7]
+ m_wbs_dat_o_2[8] m_wbs_dat_o_2[9] m_wbs_dat_o_3[0] m_wbs_dat_o_3[10] m_wbs_dat_o_3[11]
+ m_wbs_dat_o_3[12] m_wbs_dat_o_3[13] m_wbs_dat_o_3[14] m_wbs_dat_o_3[15] m_wbs_dat_o_3[16]
+ m_wbs_dat_o_3[17] m_wbs_dat_o_3[18] m_wbs_dat_o_3[19] m_wbs_dat_o_3[1] m_wbs_dat_o_3[20]
+ m_wbs_dat_o_3[21] m_wbs_dat_o_3[22] m_wbs_dat_o_3[23] m_wbs_dat_o_3[24] m_wbs_dat_o_3[25]
+ m_wbs_dat_o_3[26] m_wbs_dat_o_3[27] m_wbs_dat_o_3[28] m_wbs_dat_o_3[29] m_wbs_dat_o_3[2]
+ m_wbs_dat_o_3[30] m_wbs_dat_o_3[31] m_wbs_dat_o_3[3] m_wbs_dat_o_3[4] m_wbs_dat_o_3[5]
+ m_wbs_dat_o_3[6] m_wbs_dat_o_3[7] m_wbs_dat_o_3[8] m_wbs_dat_o_3[9] m_wbs_dat_o_4[0]
+ m_wbs_dat_o_4[10] m_wbs_dat_o_4[11] m_wbs_dat_o_4[12] m_wbs_dat_o_4[13] m_wbs_dat_o_4[14]
+ m_wbs_dat_o_4[15] m_wbs_dat_o_4[16] m_wbs_dat_o_4[17] m_wbs_dat_o_4[18] m_wbs_dat_o_4[19]
+ m_wbs_dat_o_4[1] m_wbs_dat_o_4[20] m_wbs_dat_o_4[21] m_wbs_dat_o_4[22] m_wbs_dat_o_4[23]
+ m_wbs_dat_o_4[24] m_wbs_dat_o_4[25] m_wbs_dat_o_4[26] m_wbs_dat_o_4[27] m_wbs_dat_o_4[28]
+ m_wbs_dat_o_4[29] m_wbs_dat_o_4[2] m_wbs_dat_o_4[30] m_wbs_dat_o_4[31] m_wbs_dat_o_4[3]
+ m_wbs_dat_o_4[4] m_wbs_dat_o_4[5] m_wbs_dat_o_4[6] m_wbs_dat_o_4[7] m_wbs_dat_o_4[8]
+ m_wbs_dat_o_4[9] m_wbs_dat_o_5[0] m_wbs_dat_o_5[10] m_wbs_dat_o_5[11] m_wbs_dat_o_5[12]
+ m_wbs_dat_o_5[13] m_wbs_dat_o_5[14] m_wbs_dat_o_5[15] m_wbs_dat_o_5[16] m_wbs_dat_o_5[17]
+ m_wbs_dat_o_5[18] m_wbs_dat_o_5[19] m_wbs_dat_o_5[1] m_wbs_dat_o_5[20] m_wbs_dat_o_5[21]
+ m_wbs_dat_o_5[22] m_wbs_dat_o_5[23] m_wbs_dat_o_5[24] m_wbs_dat_o_5[25] m_wbs_dat_o_5[26]
+ m_wbs_dat_o_5[27] m_wbs_dat_o_5[28] m_wbs_dat_o_5[29] m_wbs_dat_o_5[2] m_wbs_dat_o_5[30]
+ m_wbs_dat_o_5[31] m_wbs_dat_o_5[3] m_wbs_dat_o_5[4] m_wbs_dat_o_5[5] m_wbs_dat_o_5[6]
+ m_wbs_dat_o_5[7] m_wbs_dat_o_5[8] m_wbs_dat_o_5[9] m_wbs_dat_o_6[0] m_wbs_dat_o_6[10]
+ m_wbs_dat_o_6[11] m_wbs_dat_o_6[12] m_wbs_dat_o_6[13] m_wbs_dat_o_6[14] m_wbs_dat_o_6[15]
+ m_wbs_dat_o_6[16] m_wbs_dat_o_6[17] m_wbs_dat_o_6[18] m_wbs_dat_o_6[19] m_wbs_dat_o_6[1]
+ m_wbs_dat_o_6[20] m_wbs_dat_o_6[21] m_wbs_dat_o_6[22] m_wbs_dat_o_6[23] m_wbs_dat_o_6[24]
+ m_wbs_dat_o_6[25] m_wbs_dat_o_6[26] m_wbs_dat_o_6[27] m_wbs_dat_o_6[28] m_wbs_dat_o_6[29]
+ m_wbs_dat_o_6[2] m_wbs_dat_o_6[30] m_wbs_dat_o_6[31] m_wbs_dat_o_6[3] m_wbs_dat_o_6[4]
+ m_wbs_dat_o_6[5] m_wbs_dat_o_6[6] m_wbs_dat_o_6[7] m_wbs_dat_o_6[8] m_wbs_dat_o_6[9]
+ m_wbs_dat_o_7[0] m_wbs_dat_o_7[10] m_wbs_dat_o_7[11] m_wbs_dat_o_7[12] m_wbs_dat_o_7[13]
+ m_wbs_dat_o_7[14] m_wbs_dat_o_7[15] m_wbs_dat_o_7[16] m_wbs_dat_o_7[17] m_wbs_dat_o_7[18]
+ m_wbs_dat_o_7[19] m_wbs_dat_o_7[1] m_wbs_dat_o_7[20] m_wbs_dat_o_7[21] m_wbs_dat_o_7[22]
+ m_wbs_dat_o_7[23] m_wbs_dat_o_7[24] m_wbs_dat_o_7[25] m_wbs_dat_o_7[26] m_wbs_dat_o_7[27]
+ m_wbs_dat_o_7[28] m_wbs_dat_o_7[29] m_wbs_dat_o_7[2] m_wbs_dat_o_7[30] m_wbs_dat_o_7[31]
+ m_wbs_dat_o_7[3] m_wbs_dat_o_7[4] m_wbs_dat_o_7[5] m_wbs_dat_o_7[6] m_wbs_dat_o_7[7]
+ m_wbs_dat_o_7[8] m_wbs_dat_o_7[9] m_wbs_dat_o_8[0] m_wbs_dat_o_8[10] m_wbs_dat_o_8[11]
+ m_wbs_dat_o_8[12] m_wbs_dat_o_8[13] m_wbs_dat_o_8[14] m_wbs_dat_o_8[15] m_wbs_dat_o_8[16]
+ m_wbs_dat_o_8[17] m_wbs_dat_o_8[18] m_wbs_dat_o_8[19] m_wbs_dat_o_8[1] m_wbs_dat_o_8[20]
+ m_wbs_dat_o_8[21] m_wbs_dat_o_8[22] m_wbs_dat_o_8[23] m_wbs_dat_o_8[24] m_wbs_dat_o_8[25]
+ m_wbs_dat_o_8[26] m_wbs_dat_o_8[27] m_wbs_dat_o_8[28] m_wbs_dat_o_8[29] m_wbs_dat_o_8[2]
+ m_wbs_dat_o_8[30] m_wbs_dat_o_8[31] m_wbs_dat_o_8[3] m_wbs_dat_o_8[4] m_wbs_dat_o_8[5]
+ m_wbs_dat_o_8[6] m_wbs_dat_o_8[7] m_wbs_dat_o_8[8] m_wbs_dat_o_8[9] m_wbs_dat_o_9[0]
+ m_wbs_dat_o_9[10] m_wbs_dat_o_9[11] m_wbs_dat_o_9[12] m_wbs_dat_o_9[13] m_wbs_dat_o_9[14]
+ m_wbs_dat_o_9[15] m_wbs_dat_o_9[16] m_wbs_dat_o_9[17] m_wbs_dat_o_9[18] m_wbs_dat_o_9[19]
+ m_wbs_dat_o_9[1] m_wbs_dat_o_9[20] m_wbs_dat_o_9[21] m_wbs_dat_o_9[22] m_wbs_dat_o_9[23]
+ m_wbs_dat_o_9[24] m_wbs_dat_o_9[25] m_wbs_dat_o_9[26] m_wbs_dat_o_9[27] m_wbs_dat_o_9[28]
+ m_wbs_dat_o_9[29] m_wbs_dat_o_9[2] m_wbs_dat_o_9[30] m_wbs_dat_o_9[31] m_wbs_dat_o_9[3]
+ m_wbs_dat_o_9[4] m_wbs_dat_o_9[5] m_wbs_dat_o_9[6] m_wbs_dat_o_9[7] m_wbs_dat_o_9[8]
+ m_wbs_dat_o_9[9] m_wbs_we_i mt_QEI_ChA_0 mt_QEI_ChA_1 mt_QEI_ChA_2 mt_QEI_ChA_3
+ mt_QEI_ChB_0 mt_QEI_ChB_1 mt_QEI_ChB_2 mt_QEI_ChB_3 mt_pwm_h_0 mt_pwm_h_1 mt_pwm_h_2
+ mt_pwm_h_3 mt_pwm_l_0 mt_pwm_l_1 mt_pwm_l_2 mt_pwm_l_3 wb_clk_i wb_rst_i wbs_ack_o
+ wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ vccd1 vssd1 vccd2 vssd2 vdda1 vssa1 vdda2 vssa2 vdda2_uq0 vdda2_uq1 vdda2_uq2 vdda2_uq3
+ vdda2_uq4 vdda2_uq5 vdda2_uq6 vdda2_uq7 vdda2_uq8 vdda2_uq9 vdda2_uq10 vdda2_uq11
+ vdda2_uq12 vdda2_uq13 vdda2_uq14 vdda2_uq15 vdda2_uq16 vdda2_uq17 vdda2_uq18 vdda2_uq19
+ vdda2_uq20 vdda2_uq21 vdda2_uq22 vdda2_uq23 vdda2_uq24 vdda2_uq25 vdda2_uq26 vdda2_uq27
+ vdda2_uq28 vdda2_uq29 vdda2_uq30 vdda2_uq31 vdda2_uq32 vdda2_uq33 vdda2_uq34 vdda2_uq35
+ vdda2_uq36 vdda2_uq37 vdda2_uq38 vdda2_uq39 vdda2_uq40 vdda2_uq41 vdda2_uq42 vdda2_uq43
+ vdda2_uq44 vdda2_uq45 vdda2_uq46 vdda2_uq47 vdda2_uq48 vdda2_uq49 vdda2_uq50 vdda2_uq51
+ vdda2_uq52 vdda2_uq53 vdda2_uq54 vdda2_uq55 vdda2_uq56 vdda2_uq57 vdda2_uq58 vdda2_uq59
+ vdda2_uq60 vdda2_uq61 vdda2_uq62 vdda2_uq63 vdda2_uq64 vdda2_uq65 vdda1_uq0 vdda1_uq1
+ vdda1_uq2 vdda1_uq3 vdda1_uq4 vdda1_uq5 vdda1_uq6 vdda1_uq7 vdda1_uq8 vdda1_uq9
+ vdda1_uq10 vdda1_uq11 vdda1_uq12 vdda1_uq13 vdda1_uq14 vdda1_uq15 vdda1_uq16 vdda1_uq17
+ vdda1_uq18 vdda1_uq19 vdda1_uq20 vdda1_uq21 vdda1_uq22 vdda1_uq23 vdda1_uq24 vdda1_uq25
+ vdda1_uq26 vdda1_uq27 vdda1_uq28 vdda1_uq29 vdda1_uq30 vdda1_uq31 vdda1_uq32 vdda1_uq33
+ vdda1_uq34 vdda1_uq35 vdda1_uq36 vdda1_uq37 vdda1_uq38 vdda1_uq39 vdda1_uq40 vdda1_uq41
+ vdda1_uq42 vdda1_uq43 vdda1_uq44 vdda1_uq45 vdda1_uq46 vdda1_uq47 vdda1_uq48 vdda1_uq49
+ vdda1_uq50 vdda1_uq51 vdda1_uq52 vdda1_uq53 vdda1_uq54 vdda1_uq55 vdda1_uq56 vdda1_uq57
+ vdda1_uq58 vdda1_uq59 vdda1_uq60 vdda1_uq61 vdda1_uq62 vdda1_uq63 vdda1_uq64 vdda1_uq65
+ vdda1_uq66 vdda1_uq67 vdda1_uq68 vdda1_uq69 vdda1_uq70 vdda1_uq71 vdda1_uq72 vdda1_uq73
+ vdda1_uq74 vdda1_uq75 vdda1_uq76 vdda1_uq77 vdda1_uq78 vdda1_uq79 vdda1_uq80 vdda1_uq81
+ vdda1_uq82 vdda1_uq83 vccd2_uq0 vccd2_uq1 vccd2_uq2 vccd2_uq3 vccd2_uq4 vccd2_uq5
+ vccd2_uq6 vccd2_uq7 vccd2_uq8 vccd2_uq9 vccd2_uq10 vccd2_uq11 vccd2_uq12 vccd2_uq13
+ vccd2_uq14 vccd2_uq15 vccd2_uq16 vccd2_uq17 vccd2_uq18 vccd2_uq19 vccd2_uq20 vccd2_uq21
+ vccd2_uq22 vccd2_uq23 vccd2_uq24 vccd2_uq25 vccd2_uq26 vccd2_uq27 vccd2_uq28 vccd2_uq29
+ vccd2_uq30 vccd2_uq31 vccd2_uq32 vccd2_uq33 vccd2_uq34 vccd2_uq35 vccd2_uq36 vccd2_uq37
+ vccd2_uq38 vccd2_uq39 vccd2_uq40 vccd2_uq41 vccd2_uq42 vccd2_uq43 vccd2_uq44 vccd2_uq45
+ vccd2_uq46 vccd2_uq47 vccd2_uq48 vccd2_uq49 vccd2_uq50 vccd2_uq51 vccd2_uq52 vccd2_uq53
+ vccd2_uq54 vccd2_uq55 vccd2_uq56 vccd2_uq57 vccd2_uq58 vccd2_uq59 vccd2_uq60 vccd2_uq61
+ vccd2_uq62 vccd2_uq63 vccd2_uq64 vccd2_uq65 vccd2_uq66 vccd2_uq67 vccd2_uq68 vccd2_uq69
+ vccd2_uq70 vccd2_uq71 vccd2_uq72 vccd2_uq73 vccd2_uq74 vccd2_uq75 vccd2_uq76 vccd2_uq77
+ vccd2_uq78 vccd2_uq79 vccd2_uq80 vccd2_uq81 vccd2_uq82 vccd2_uq83 vccd2_uq84 vccd2_uq85
+ vccd2_uq86 vccd2_uq87 vccd2_uq88 vccd2_uq89 vccd2_uq90 vccd2_uq91 vccd2_uq92 vccd2_uq93
+ vccd2_uq94 vccd2_uq95 vccd2_uq96 vccd2_uq97 vccd2_uq98 vccd2_uq99 vccd2_uq100 vccd2_uq101
+ vccd2_uq102 vccd2_uq103 vssa2_uq0 vssa2_uq1 vssa2_uq2 vssa2_uq3 vssa2_uq4 vssa2_uq5
+ vssa2_uq6 vssa2_uq7 vssa2_uq8 vssa2_uq9 vssa2_uq10 vssa2_uq11 vssa2_uq12 vssa2_uq13
+ vssa2_uq14 vssa2_uq15 vssa2_uq16 vssa2_uq17 vssa2_uq18 vssa2_uq19 vssa2_uq20 vssa2_uq21
+ vssa2_uq22 vssa2_uq23 vssa2_uq24 vssa2_uq25 vssa2_uq26 vssa2_uq27 vssa2_uq28 vssa2_uq29
+ vssa2_uq30 vssa2_uq31 vssa2_uq32 vssa2_uq33 vssa2_uq34 vssa2_uq35 vssa2_uq36 vssa2_uq37
+ vssa2_uq38 vssa2_uq39 vssa2_uq40 vssa2_uq41 vssa2_uq42 vssa2_uq43 vssa2_uq44 vssa2_uq45
+ vssa2_uq46 vssa2_uq47 vssa2_uq48 vssa2_uq49 vssa2_uq50 vssa2_uq51 vssa2_uq52 vssa2_uq53
+ vssa2_uq54 vssa2_uq55 vssa2_uq56 vssa2_uq57 vssa2_uq58 vssa2_uq59 vssa2_uq60 vssa2_uq61
+ vssa2_uq62 vssa2_uq63 vssa2_uq64 vssa2_uq65 vssa2_uq66 vssa2_uq67 vssa2_uq68 vssa2_uq69
+ vssa2_uq70 vssa2_uq71 vssa2_uq72 vssa2_uq73 vssa2_uq74 vssa2_uq75 vssa2_uq76 vssa2_uq77
+ vssa1_uq0 vssa1_uq1 vssa1_uq2 vssa1_uq3 vssa1_uq4 vssa1_uq5 vssa1_uq6 vssa1_uq7
+ vssa1_uq8 vssa1_uq9 vssa1_uq10 vssa1_uq11 vssa1_uq12 vssa1_uq13 vssa1_uq14 vssa1_uq15
+ vssa1_uq16 vssa1_uq17 vssa1_uq18 vssa1_uq19 vssa1_uq20 vssa1_uq21 vssa1_uq22 vssa1_uq23
+ vssa1_uq24 vssa1_uq25 vssa1_uq26 vssa1_uq27 vssa1_uq28 vssa1_uq29 vssa1_uq30 vssa1_uq31
+ vssa1_uq32 vssa1_uq33 vssa1_uq34 vssa1_uq35 vssa1_uq36 vssa1_uq37 vssa1_uq38 vssa1_uq39
+ vssa1_uq40 vssa1_uq41 vssa1_uq42 vssa1_uq43 vssa1_uq44 vssa1_uq45 vssa1_uq46 vssa1_uq47
+ vssa1_uq48 vssa1_uq49 vssa1_uq50 vssa1_uq51 vssd2_uq0 vssd2_uq1 vssd2_uq2 vssd2_uq3
+ vssd2_uq4 vssd2_uq5 vssd2_uq6 vssd2_uq7 vssd2_uq8 vssd2_uq9 vssd2_uq10 vssd2_uq11
+ vssd2_uq12 vssd2_uq13 vssd2_uq14 vssd2_uq15 vssd2_uq16 vssd2_uq17 vssd2_uq18 vssd2_uq19
+ vssd2_uq20 vssd2_uq21 vssd2_uq22 vssd2_uq23 vssd2_uq24 vssd2_uq25 vssd2_uq26 vssd2_uq27
+ vssd2_uq28 vssd2_uq29 vssd2_uq30 vssd2_uq31 vssd2_uq32 vssd2_uq33 vssd2_uq34 vssd2_uq35
+ vssd2_uq36 vssd2_uq37 vssd2_uq38 vssd2_uq39 vssd2_uq40 vssd2_uq41 vssd2_uq42 vssd2_uq43
+ vssd2_uq44 vssd2_uq45 vssd2_uq46 vssd2_uq47 vssd2_uq48 vssd2_uq49 vssd2_uq50 vssd2_uq51
Xcb_1_10 cb_1_9/io_adr_i[0] cb_1_9/io_adr_i[1] cb_1_10/io_cs_i cb_1_9/io_dat_i[0]
+ cb_1_9/io_dat_i[10] cb_1_9/io_dat_i[11] cb_1_9/io_dat_i[12] cb_1_9/io_dat_i[13]
+ cb_1_9/io_dat_i[14] cb_1_9/io_dat_i[15] cb_1_9/io_dat_i[1] cb_1_9/io_dat_i[2] cb_1_9/io_dat_i[3]
+ cb_1_9/io_dat_i[4] cb_1_9/io_dat_i[5] cb_1_9/io_dat_i[6] cb_1_9/io_dat_i[7] cb_1_9/io_dat_i[8]
+ cb_1_9/io_dat_i[9] cb_1_10/io_dat_o[0] cb_1_10/io_dat_o[10] cb_1_10/io_dat_o[11]
+ cb_1_10/io_dat_o[12] cb_1_10/io_dat_o[13] cb_1_10/io_dat_o[14] cb_1_10/io_dat_o[15]
+ cb_1_10/io_dat_o[1] cb_1_10/io_dat_o[2] cb_1_10/io_dat_o[3] cb_1_10/io_dat_o[4]
+ cb_1_10/io_dat_o[5] cb_1_10/io_dat_o[6] cb_1_10/io_dat_o[7] cb_1_10/io_dat_o[8]
+ cb_1_10/io_dat_o[9] cb_1_10/io_eo[0] cb_1_10/io_eo[10] cb_1_10/io_eo[11] cb_1_10/io_eo[12]
+ cb_1_10/io_eo[13] cb_1_10/io_eo[14] cb_1_10/io_eo[15] cb_1_10/io_eo[16] cb_1_10/io_eo[17]
+ cb_1_10/io_eo[18] cb_1_10/io_eo[19] cb_1_10/io_eo[1] cb_1_10/io_eo[20] cb_1_10/io_eo[21]
+ cb_1_10/io_eo[22] cb_1_10/io_eo[23] cb_1_10/io_eo[24] cb_1_10/io_eo[25] cb_1_10/io_eo[26]
+ cb_1_10/io_eo[27] cb_1_10/io_eo[28] cb_1_10/io_eo[29] cb_1_10/io_eo[2] cb_1_10/io_eo[30]
+ cb_1_10/io_eo[31] cb_1_10/io_eo[32] cb_1_10/io_eo[33] cb_1_10/io_eo[34] cb_1_10/io_eo[35]
+ cb_1_10/io_eo[36] cb_1_10/io_eo[37] cb_1_10/io_eo[38] cb_1_10/io_eo[39] cb_1_10/io_eo[3]
+ cb_1_10/io_eo[40] cb_1_10/io_eo[41] cb_1_10/io_eo[42] cb_1_10/io_eo[43] cb_1_10/io_eo[44]
+ cb_1_10/io_eo[45] cb_1_10/io_eo[46] cb_1_10/io_eo[47] cb_1_10/io_eo[48] cb_1_10/io_eo[49]
+ cb_1_10/io_eo[4] cb_1_10/io_eo[50] cb_1_10/io_eo[51] cb_1_10/io_eo[52] cb_1_10/io_eo[53]
+ cb_1_10/io_eo[54] cb_1_10/io_eo[55] cb_1_10/io_eo[56] cb_1_10/io_eo[57] cb_1_10/io_eo[58]
+ cb_1_10/io_eo[59] cb_1_10/io_eo[5] cb_1_10/io_eo[60] cb_1_10/io_eo[61] cb_1_10/io_eo[62]
+ cb_1_10/io_eo[63] cb_1_10/io_eo[6] cb_1_10/io_eo[7] cb_1_10/io_eo[8] cb_1_10/io_eo[9]
+ cb_1_9/io_o_0_co cb_1_9/io_o_0_out[0] cb_1_9/io_o_0_out[1] cb_1_9/io_o_0_out[2]
+ cb_1_9/io_o_0_out[3] cb_1_9/io_o_0_out[4] cb_1_9/io_o_0_out[5] cb_1_9/io_o_0_out[6]
+ cb_1_9/io_o_0_out[7] cb_1_9/io_o_1_co cb_1_9/io_o_1_out[0] cb_1_9/io_o_1_out[1]
+ cb_1_9/io_o_1_out[2] cb_1_9/io_o_1_out[3] cb_1_9/io_o_1_out[4] cb_1_9/io_o_1_out[5]
+ cb_1_9/io_o_1_out[6] cb_1_9/io_o_1_out[7] cb_1_9/io_o_2_co cb_1_9/io_o_2_out[0]
+ cb_1_9/io_o_2_out[1] cb_1_9/io_o_2_out[2] cb_1_9/io_o_2_out[3] cb_1_9/io_o_2_out[4]
+ cb_1_9/io_o_2_out[5] cb_1_9/io_o_2_out[6] cb_1_9/io_o_2_out[7] cb_1_9/io_o_3_co
+ cb_1_9/io_o_3_out[0] cb_1_9/io_o_3_out[1] cb_1_9/io_o_3_out[2] cb_1_9/io_o_3_out[3]
+ cb_1_9/io_o_3_out[4] cb_1_9/io_o_3_out[5] cb_1_9/io_o_3_out[6] cb_1_9/io_o_3_out[7]
+ cb_1_9/io_o_4_co cb_1_9/io_o_4_out[0] cb_1_9/io_o_4_out[1] cb_1_9/io_o_4_out[2]
+ cb_1_9/io_o_4_out[3] cb_1_9/io_o_4_out[4] cb_1_9/io_o_4_out[5] cb_1_9/io_o_4_out[6]
+ cb_1_9/io_o_4_out[7] cb_1_9/io_o_5_co cb_1_9/io_o_5_out[0] cb_1_9/io_o_5_out[1]
+ cb_1_9/io_o_5_out[2] cb_1_9/io_o_5_out[3] cb_1_9/io_o_5_out[4] cb_1_9/io_o_5_out[5]
+ cb_1_9/io_o_5_out[6] cb_1_9/io_o_5_out[7] cb_1_9/io_o_6_co cb_1_9/io_o_6_out[0]
+ cb_1_9/io_o_6_out[1] cb_1_9/io_o_6_out[2] cb_1_9/io_o_6_out[3] cb_1_9/io_o_6_out[4]
+ cb_1_9/io_o_6_out[5] cb_1_9/io_o_6_out[6] cb_1_9/io_o_6_out[7] cb_1_9/io_o_7_co
+ cb_1_9/io_o_7_out[0] cb_1_9/io_o_7_out[1] cb_1_9/io_o_7_out[2] cb_1_9/io_o_7_out[3]
+ cb_1_9/io_o_7_out[4] cb_1_9/io_o_7_out[5] cb_1_9/io_o_7_out[6] cb_1_9/io_o_7_out[7]
+ cb_1_10/io_o_0_co cb_1_10/io_eo[0] cb_1_10/io_eo[1] cb_1_10/io_eo[2] cb_1_10/io_eo[3]
+ cb_1_10/io_eo[4] cb_1_10/io_eo[5] cb_1_10/io_eo[6] cb_1_10/io_eo[7] cb_1_10/io_o_1_co
+ cb_1_10/io_eo[8] cb_1_10/io_eo[9] cb_1_10/io_eo[10] cb_1_10/io_eo[11] cb_1_10/io_eo[12]
+ cb_1_10/io_eo[13] cb_1_10/io_eo[14] cb_1_10/io_eo[15] cb_1_10/io_o_2_co cb_1_10/io_eo[16]
+ cb_1_10/io_eo[17] cb_1_10/io_eo[18] cb_1_10/io_eo[19] cb_1_10/io_eo[20] cb_1_10/io_eo[21]
+ cb_1_10/io_eo[22] cb_1_10/io_eo[23] cb_1_10/io_o_3_co cb_1_10/io_eo[24] cb_1_10/io_eo[25]
+ cb_1_10/io_eo[26] cb_1_10/io_eo[27] cb_1_10/io_eo[28] cb_1_10/io_eo[29] cb_1_10/io_eo[30]
+ cb_1_10/io_eo[31] cb_1_10/io_o_4_co cb_1_10/io_eo[32] cb_1_10/io_eo[33] cb_1_10/io_eo[34]
+ cb_1_10/io_eo[35] cb_1_10/io_eo[36] cb_1_10/io_eo[37] cb_1_10/io_eo[38] cb_1_10/io_eo[39]
+ cb_1_10/io_o_5_co cb_1_10/io_eo[40] cb_1_10/io_eo[41] cb_1_10/io_eo[42] cb_1_10/io_eo[43]
+ cb_1_10/io_eo[44] cb_1_10/io_eo[45] cb_1_10/io_eo[46] cb_1_10/io_eo[47] cb_1_10/io_o_6_co
+ cb_1_10/io_eo[48] cb_1_10/io_eo[49] cb_1_10/io_eo[50] cb_1_10/io_eo[51] cb_1_10/io_eo[52]
+ cb_1_10/io_eo[53] cb_1_10/io_eo[54] cb_1_10/io_eo[55] cb_1_10/io_o_7_co cb_1_10/io_eo[56]
+ cb_1_10/io_eo[57] cb_1_10/io_eo[58] cb_1_10/io_eo[59] cb_1_10/io_eo[60] cb_1_10/io_eo[61]
+ cb_1_10/io_eo[62] cb_1_10/io_eo[63] cb_1_9/io_vco cb_1_10/io_vco cb_1_10/io_vi cb_1_9/io_we_i
+ cb_1_9/io_eo[0] cb_1_9/io_eo[10] cb_1_9/io_eo[11] cb_1_9/io_eo[12] cb_1_9/io_eo[13]
+ cb_1_9/io_eo[14] cb_1_9/io_eo[15] cb_1_9/io_eo[16] cb_1_9/io_eo[17] cb_1_9/io_eo[18]
+ cb_1_9/io_eo[19] cb_1_9/io_eo[1] cb_1_9/io_eo[20] cb_1_9/io_eo[21] cb_1_9/io_eo[22]
+ cb_1_9/io_eo[23] cb_1_9/io_eo[24] cb_1_9/io_eo[25] cb_1_9/io_eo[26] cb_1_9/io_eo[27]
+ cb_1_9/io_eo[28] cb_1_9/io_eo[29] cb_1_9/io_eo[2] cb_1_9/io_eo[30] cb_1_9/io_eo[31]
+ cb_1_9/io_eo[32] cb_1_9/io_eo[33] cb_1_9/io_eo[34] cb_1_9/io_eo[35] cb_1_9/io_eo[36]
+ cb_1_9/io_eo[37] cb_1_9/io_eo[38] cb_1_9/io_eo[39] cb_1_9/io_eo[3] cb_1_9/io_eo[40]
+ cb_1_9/io_eo[41] cb_1_9/io_eo[42] cb_1_9/io_eo[43] cb_1_9/io_eo[44] cb_1_9/io_eo[45]
+ cb_1_9/io_eo[46] cb_1_9/io_eo[47] cb_1_9/io_eo[48] cb_1_9/io_eo[49] cb_1_9/io_eo[4]
+ cb_1_9/io_eo[50] cb_1_9/io_eo[51] cb_1_9/io_eo[52] cb_1_9/io_eo[53] cb_1_9/io_eo[54]
+ cb_1_9/io_eo[55] cb_1_9/io_eo[56] cb_1_9/io_eo[57] cb_1_9/io_eo[58] cb_1_9/io_eo[59]
+ cb_1_9/io_eo[5] cb_1_9/io_eo[60] cb_1_9/io_eo[61] cb_1_9/io_eo[62] cb_1_9/io_eo[63]
+ cb_1_9/io_eo[6] cb_1_9/io_eo[7] cb_1_9/io_eo[8] cb_1_9/io_eo[9] mcons_3/clock mcons_3/reset
+ vccd1 vssd1 cic_block
Xmcons_1 mcons_3/clock icon/mt_QEI_ChA_1 icon/mt_QEI_ChB_1 mcons_1/io_irq icon/mt_pwm_h_1
+ icon/mt_pwm_l_1 mcons_1/io_wb_ack_o ccon_7/io_adr_i[0] ccon_7/io_adr_i[10] ccon_7/io_adr_i[11]
+ ccon_7/io_adr_i[1] ccon_7/io_adr_i[2] ccon_7/io_adr_i[3] ccon_7/io_adr_i[4] ccon_7/io_adr_i[5]
+ ccon_7/io_adr_i[6] ccon_7/io_adr_i[7] ccon_7/io_adr_i[8] ccon_7/io_adr_i[9] mcons_1/io_wb_cs_i
+ ccon_7/io_dat_i[0] ccon_7/io_dat_i[10] ccon_7/io_dat_i[11] ccon_7/io_dat_i[12] ccon_7/io_dat_i[13]
+ ccon_7/io_dat_i[14] ccon_7/io_dat_i[15] ccon_7/io_dat_i[16] ccon_7/io_dat_i[17]
+ ccon_7/io_dat_i[18] ccon_7/io_dat_i[19] ccon_7/io_dat_i[1] ccon_7/io_dat_i[20] ccon_7/io_dat_i[21]
+ ccon_7/io_dat_i[22] ccon_7/io_dat_i[23] ccon_7/io_dat_i[24] ccon_7/io_dat_i[25]
+ ccon_7/io_dat_i[26] ccon_7/io_dat_i[27] ccon_7/io_dat_i[28] ccon_7/io_dat_i[29]
+ ccon_7/io_dat_i[2] ccon_7/io_dat_i[30] ccon_7/io_dat_i[31] ccon_7/io_dat_i[3] ccon_7/io_dat_i[4]
+ ccon_7/io_dat_i[5] ccon_7/io_dat_i[6] ccon_7/io_dat_i[7] ccon_7/io_dat_i[8] ccon_7/io_dat_i[9]
+ icon/m_wbs_dat_o_1[0] icon/m_wbs_dat_o_1[10] icon/m_wbs_dat_o_1[11] icon/m_wbs_dat_o_1[12]
+ icon/m_wbs_dat_o_1[13] icon/m_wbs_dat_o_1[14] icon/m_wbs_dat_o_1[15] icon/m_wbs_dat_o_1[16]
+ icon/m_wbs_dat_o_1[17] icon/m_wbs_dat_o_1[18] icon/m_wbs_dat_o_1[19] icon/m_wbs_dat_o_1[1]
+ icon/m_wbs_dat_o_1[20] icon/m_wbs_dat_o_1[21] icon/m_wbs_dat_o_1[22] icon/m_wbs_dat_o_1[23]
+ icon/m_wbs_dat_o_1[24] icon/m_wbs_dat_o_1[25] icon/m_wbs_dat_o_1[26] icon/m_wbs_dat_o_1[27]
+ icon/m_wbs_dat_o_1[28] icon/m_wbs_dat_o_1[29] icon/m_wbs_dat_o_1[2] icon/m_wbs_dat_o_1[30]
+ icon/m_wbs_dat_o_1[31] icon/m_wbs_dat_o_1[3] icon/m_wbs_dat_o_1[4] icon/m_wbs_dat_o_1[5]
+ icon/m_wbs_dat_o_1[6] icon/m_wbs_dat_o_1[7] icon/m_wbs_dat_o_1[8] icon/m_wbs_dat_o_1[9]
+ ccon_7/io_we_i mcons_3/reset vccd1 vssd1 motor_top
Xcb_6_2 cb_6_9/io_adr_i[0] cb_6_9/io_adr_i[1] cb_6_2/io_cs_i cb_6_9/io_dat_i[0] cb_6_9/io_dat_i[10]
+ cb_6_9/io_dat_i[11] cb_6_9/io_dat_i[12] cb_6_9/io_dat_i[13] cb_6_9/io_dat_i[14]
+ cb_6_9/io_dat_i[15] cb_6_9/io_dat_i[1] cb_6_9/io_dat_i[2] cb_6_9/io_dat_i[3] cb_6_9/io_dat_i[4]
+ cb_6_9/io_dat_i[5] cb_6_9/io_dat_i[6] cb_6_9/io_dat_i[7] cb_6_9/io_dat_i[8] cb_6_9/io_dat_i[9]
+ cb_6_2/io_dat_o[0] cb_6_2/io_dat_o[10] cb_6_2/io_dat_o[11] cb_6_2/io_dat_o[12] cb_6_2/io_dat_o[13]
+ cb_6_2/io_dat_o[14] cb_6_2/io_dat_o[15] cb_6_2/io_dat_o[1] cb_6_2/io_dat_o[2] cb_6_2/io_dat_o[3]
+ cb_6_2/io_dat_o[4] cb_6_2/io_dat_o[5] cb_6_2/io_dat_o[6] cb_6_2/io_dat_o[7] cb_6_2/io_dat_o[8]
+ cb_6_2/io_dat_o[9] cb_6_3/io_wo[0] cb_6_3/io_wo[10] cb_6_3/io_wo[11] cb_6_3/io_wo[12]
+ cb_6_3/io_wo[13] cb_6_3/io_wo[14] cb_6_3/io_wo[15] cb_6_3/io_wo[16] cb_6_3/io_wo[17]
+ cb_6_3/io_wo[18] cb_6_3/io_wo[19] cb_6_3/io_wo[1] cb_6_3/io_wo[20] cb_6_3/io_wo[21]
+ cb_6_3/io_wo[22] cb_6_3/io_wo[23] cb_6_3/io_wo[24] cb_6_3/io_wo[25] cb_6_3/io_wo[26]
+ cb_6_3/io_wo[27] cb_6_3/io_wo[28] cb_6_3/io_wo[29] cb_6_3/io_wo[2] cb_6_3/io_wo[30]
+ cb_6_3/io_wo[31] cb_6_3/io_wo[32] cb_6_3/io_wo[33] cb_6_3/io_wo[34] cb_6_3/io_wo[35]
+ cb_6_3/io_wo[36] cb_6_3/io_wo[37] cb_6_3/io_wo[38] cb_6_3/io_wo[39] cb_6_3/io_wo[3]
+ cb_6_3/io_wo[40] cb_6_3/io_wo[41] cb_6_3/io_wo[42] cb_6_3/io_wo[43] cb_6_3/io_wo[44]
+ cb_6_3/io_wo[45] cb_6_3/io_wo[46] cb_6_3/io_wo[47] cb_6_3/io_wo[48] cb_6_3/io_wo[49]
+ cb_6_3/io_wo[4] cb_6_3/io_wo[50] cb_6_3/io_wo[51] cb_6_3/io_wo[52] cb_6_3/io_wo[53]
+ cb_6_3/io_wo[54] cb_6_3/io_wo[55] cb_6_3/io_wo[56] cb_6_3/io_wo[57] cb_6_3/io_wo[58]
+ cb_6_3/io_wo[59] cb_6_3/io_wo[5] cb_6_3/io_wo[60] cb_6_3/io_wo[61] cb_6_3/io_wo[62]
+ cb_6_3/io_wo[63] cb_6_3/io_wo[6] cb_6_3/io_wo[7] cb_6_3/io_wo[8] cb_6_3/io_wo[9]
+ cb_6_2/io_i_0_ci cb_6_2/io_i_0_in1[0] cb_6_2/io_i_0_in1[1] cb_6_2/io_i_0_in1[2]
+ cb_6_2/io_i_0_in1[3] cb_6_2/io_i_0_in1[4] cb_6_2/io_i_0_in1[5] cb_6_2/io_i_0_in1[6]
+ cb_6_2/io_i_0_in1[7] cb_6_2/io_i_1_ci cb_6_2/io_i_1_in1[0] cb_6_2/io_i_1_in1[1]
+ cb_6_2/io_i_1_in1[2] cb_6_2/io_i_1_in1[3] cb_6_2/io_i_1_in1[4] cb_6_2/io_i_1_in1[5]
+ cb_6_2/io_i_1_in1[6] cb_6_2/io_i_1_in1[7] cb_6_2/io_i_2_ci cb_6_2/io_i_2_in1[0]
+ cb_6_2/io_i_2_in1[1] cb_6_2/io_i_2_in1[2] cb_6_2/io_i_2_in1[3] cb_6_2/io_i_2_in1[4]
+ cb_6_2/io_i_2_in1[5] cb_6_2/io_i_2_in1[6] cb_6_2/io_i_2_in1[7] cb_6_2/io_i_3_ci
+ cb_6_2/io_i_3_in1[0] cb_6_2/io_i_3_in1[1] cb_6_2/io_i_3_in1[2] cb_6_2/io_i_3_in1[3]
+ cb_6_2/io_i_3_in1[4] cb_6_2/io_i_3_in1[5] cb_6_2/io_i_3_in1[6] cb_6_2/io_i_3_in1[7]
+ cb_6_2/io_i_4_ci cb_6_2/io_i_4_in1[0] cb_6_2/io_i_4_in1[1] cb_6_2/io_i_4_in1[2]
+ cb_6_2/io_i_4_in1[3] cb_6_2/io_i_4_in1[4] cb_6_2/io_i_4_in1[5] cb_6_2/io_i_4_in1[6]
+ cb_6_2/io_i_4_in1[7] cb_6_2/io_i_5_ci cb_6_2/io_i_5_in1[0] cb_6_2/io_i_5_in1[1]
+ cb_6_2/io_i_5_in1[2] cb_6_2/io_i_5_in1[3] cb_6_2/io_i_5_in1[4] cb_6_2/io_i_5_in1[5]
+ cb_6_2/io_i_5_in1[6] cb_6_2/io_i_5_in1[7] cb_6_2/io_i_6_ci cb_6_2/io_i_6_in1[0]
+ cb_6_2/io_i_6_in1[1] cb_6_2/io_i_6_in1[2] cb_6_2/io_i_6_in1[3] cb_6_2/io_i_6_in1[4]
+ cb_6_2/io_i_6_in1[5] cb_6_2/io_i_6_in1[6] cb_6_2/io_i_6_in1[7] cb_6_2/io_i_7_ci
+ cb_6_2/io_i_7_in1[0] cb_6_2/io_i_7_in1[1] cb_6_2/io_i_7_in1[2] cb_6_2/io_i_7_in1[3]
+ cb_6_2/io_i_7_in1[4] cb_6_2/io_i_7_in1[5] cb_6_2/io_i_7_in1[6] cb_6_2/io_i_7_in1[7]
+ cb_6_3/io_i_0_ci cb_6_3/io_i_0_in1[0] cb_6_3/io_i_0_in1[1] cb_6_3/io_i_0_in1[2]
+ cb_6_3/io_i_0_in1[3] cb_6_3/io_i_0_in1[4] cb_6_3/io_i_0_in1[5] cb_6_3/io_i_0_in1[6]
+ cb_6_3/io_i_0_in1[7] cb_6_3/io_i_1_ci cb_6_3/io_i_1_in1[0] cb_6_3/io_i_1_in1[1]
+ cb_6_3/io_i_1_in1[2] cb_6_3/io_i_1_in1[3] cb_6_3/io_i_1_in1[4] cb_6_3/io_i_1_in1[5]
+ cb_6_3/io_i_1_in1[6] cb_6_3/io_i_1_in1[7] cb_6_3/io_i_2_ci cb_6_3/io_i_2_in1[0]
+ cb_6_3/io_i_2_in1[1] cb_6_3/io_i_2_in1[2] cb_6_3/io_i_2_in1[3] cb_6_3/io_i_2_in1[4]
+ cb_6_3/io_i_2_in1[5] cb_6_3/io_i_2_in1[6] cb_6_3/io_i_2_in1[7] cb_6_3/io_i_3_ci
+ cb_6_3/io_i_3_in1[0] cb_6_3/io_i_3_in1[1] cb_6_3/io_i_3_in1[2] cb_6_3/io_i_3_in1[3]
+ cb_6_3/io_i_3_in1[4] cb_6_3/io_i_3_in1[5] cb_6_3/io_i_3_in1[6] cb_6_3/io_i_3_in1[7]
+ cb_6_3/io_i_4_ci cb_6_3/io_i_4_in1[0] cb_6_3/io_i_4_in1[1] cb_6_3/io_i_4_in1[2]
+ cb_6_3/io_i_4_in1[3] cb_6_3/io_i_4_in1[4] cb_6_3/io_i_4_in1[5] cb_6_3/io_i_4_in1[6]
+ cb_6_3/io_i_4_in1[7] cb_6_3/io_i_5_ci cb_6_3/io_i_5_in1[0] cb_6_3/io_i_5_in1[1]
+ cb_6_3/io_i_5_in1[2] cb_6_3/io_i_5_in1[3] cb_6_3/io_i_5_in1[4] cb_6_3/io_i_5_in1[5]
+ cb_6_3/io_i_5_in1[6] cb_6_3/io_i_5_in1[7] cb_6_3/io_i_6_ci cb_6_3/io_i_6_in1[0]
+ cb_6_3/io_i_6_in1[1] cb_6_3/io_i_6_in1[2] cb_6_3/io_i_6_in1[3] cb_6_3/io_i_6_in1[4]
+ cb_6_3/io_i_6_in1[5] cb_6_3/io_i_6_in1[6] cb_6_3/io_i_6_in1[7] cb_6_3/io_i_7_ci
+ cb_6_3/io_i_7_in1[0] cb_6_3/io_i_7_in1[1] cb_6_3/io_i_7_in1[2] cb_6_3/io_i_7_in1[3]
+ cb_6_3/io_i_7_in1[4] cb_6_3/io_i_7_in1[5] cb_6_3/io_i_7_in1[6] cb_6_3/io_i_7_in1[7]
+ cb_6_2/io_vci cb_6_3/io_vci cb_6_2/io_vi cb_6_9/io_we_i cb_6_2/io_wo[0] cb_6_2/io_wo[10]
+ cb_6_2/io_wo[11] cb_6_2/io_wo[12] cb_6_2/io_wo[13] cb_6_2/io_wo[14] cb_6_2/io_wo[15]
+ cb_6_2/io_wo[16] cb_6_2/io_wo[17] cb_6_2/io_wo[18] cb_6_2/io_wo[19] cb_6_2/io_wo[1]
+ cb_6_2/io_wo[20] cb_6_2/io_wo[21] cb_6_2/io_wo[22] cb_6_2/io_wo[23] cb_6_2/io_wo[24]
+ cb_6_2/io_wo[25] cb_6_2/io_wo[26] cb_6_2/io_wo[27] cb_6_2/io_wo[28] cb_6_2/io_wo[29]
+ cb_6_2/io_wo[2] cb_6_2/io_wo[30] cb_6_2/io_wo[31] cb_6_2/io_wo[32] cb_6_2/io_wo[33]
+ cb_6_2/io_wo[34] cb_6_2/io_wo[35] cb_6_2/io_wo[36] cb_6_2/io_wo[37] cb_6_2/io_wo[38]
+ cb_6_2/io_wo[39] cb_6_2/io_wo[3] cb_6_2/io_wo[40] cb_6_2/io_wo[41] cb_6_2/io_wo[42]
+ cb_6_2/io_wo[43] cb_6_2/io_wo[44] cb_6_2/io_wo[45] cb_6_2/io_wo[46] cb_6_2/io_wo[47]
+ cb_6_2/io_wo[48] cb_6_2/io_wo[49] cb_6_2/io_wo[4] cb_6_2/io_wo[50] cb_6_2/io_wo[51]
+ cb_6_2/io_wo[52] cb_6_2/io_wo[53] cb_6_2/io_wo[54] cb_6_2/io_wo[55] cb_6_2/io_wo[56]
+ cb_6_2/io_wo[57] cb_6_2/io_wo[58] cb_6_2/io_wo[59] cb_6_2/io_wo[5] cb_6_2/io_wo[60]
+ cb_6_2/io_wo[61] cb_6_2/io_wo[62] cb_6_2/io_wo[63] cb_6_2/io_wo[6] cb_6_2/io_wo[7]
+ cb_6_2/io_wo[8] cb_6_2/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_4_10 cb_4_9/io_adr_i[0] cb_4_9/io_adr_i[1] cb_4_10/io_cs_i cb_4_9/io_dat_i[0]
+ cb_4_9/io_dat_i[10] cb_4_9/io_dat_i[11] cb_4_9/io_dat_i[12] cb_4_9/io_dat_i[13]
+ cb_4_9/io_dat_i[14] cb_4_9/io_dat_i[15] cb_4_9/io_dat_i[1] cb_4_9/io_dat_i[2] cb_4_9/io_dat_i[3]
+ cb_4_9/io_dat_i[4] cb_4_9/io_dat_i[5] cb_4_9/io_dat_i[6] cb_4_9/io_dat_i[7] cb_4_9/io_dat_i[8]
+ cb_4_9/io_dat_i[9] cb_4_10/io_dat_o[0] cb_4_10/io_dat_o[10] cb_4_10/io_dat_o[11]
+ cb_4_10/io_dat_o[12] cb_4_10/io_dat_o[13] cb_4_10/io_dat_o[14] cb_4_10/io_dat_o[15]
+ cb_4_10/io_dat_o[1] cb_4_10/io_dat_o[2] cb_4_10/io_dat_o[3] cb_4_10/io_dat_o[4]
+ cb_4_10/io_dat_o[5] cb_4_10/io_dat_o[6] cb_4_10/io_dat_o[7] cb_4_10/io_dat_o[8]
+ cb_4_10/io_dat_o[9] cb_4_10/io_eo[0] cb_4_10/io_eo[10] cb_4_10/io_eo[11] cb_4_10/io_eo[12]
+ cb_4_10/io_eo[13] cb_4_10/io_eo[14] cb_4_10/io_eo[15] cb_4_10/io_eo[16] cb_4_10/io_eo[17]
+ cb_4_10/io_eo[18] cb_4_10/io_eo[19] cb_4_10/io_eo[1] cb_4_10/io_eo[20] cb_4_10/io_eo[21]
+ cb_4_10/io_eo[22] cb_4_10/io_eo[23] cb_4_10/io_eo[24] cb_4_10/io_eo[25] cb_4_10/io_eo[26]
+ cb_4_10/io_eo[27] cb_4_10/io_eo[28] cb_4_10/io_eo[29] cb_4_10/io_eo[2] cb_4_10/io_eo[30]
+ cb_4_10/io_eo[31] cb_4_10/io_eo[32] cb_4_10/io_eo[33] cb_4_10/io_eo[34] cb_4_10/io_eo[35]
+ cb_4_10/io_eo[36] cb_4_10/io_eo[37] cb_4_10/io_eo[38] cb_4_10/io_eo[39] cb_4_10/io_eo[3]
+ cb_4_10/io_eo[40] cb_4_10/io_eo[41] cb_4_10/io_eo[42] cb_4_10/io_eo[43] cb_4_10/io_eo[44]
+ cb_4_10/io_eo[45] cb_4_10/io_eo[46] cb_4_10/io_eo[47] cb_4_10/io_eo[48] cb_4_10/io_eo[49]
+ cb_4_10/io_eo[4] cb_4_10/io_eo[50] cb_4_10/io_eo[51] cb_4_10/io_eo[52] cb_4_10/io_eo[53]
+ cb_4_10/io_eo[54] cb_4_10/io_eo[55] cb_4_10/io_eo[56] cb_4_10/io_eo[57] cb_4_10/io_eo[58]
+ cb_4_10/io_eo[59] cb_4_10/io_eo[5] cb_4_10/io_eo[60] cb_4_10/io_eo[61] cb_4_10/io_eo[62]
+ cb_4_10/io_eo[63] cb_4_10/io_eo[6] cb_4_10/io_eo[7] cb_4_10/io_eo[8] cb_4_10/io_eo[9]
+ cb_4_9/io_o_0_co cb_4_9/io_o_0_out[0] cb_4_9/io_o_0_out[1] cb_4_9/io_o_0_out[2]
+ cb_4_9/io_o_0_out[3] cb_4_9/io_o_0_out[4] cb_4_9/io_o_0_out[5] cb_4_9/io_o_0_out[6]
+ cb_4_9/io_o_0_out[7] cb_4_9/io_o_1_co cb_4_9/io_o_1_out[0] cb_4_9/io_o_1_out[1]
+ cb_4_9/io_o_1_out[2] cb_4_9/io_o_1_out[3] cb_4_9/io_o_1_out[4] cb_4_9/io_o_1_out[5]
+ cb_4_9/io_o_1_out[6] cb_4_9/io_o_1_out[7] cb_4_9/io_o_2_co cb_4_9/io_o_2_out[0]
+ cb_4_9/io_o_2_out[1] cb_4_9/io_o_2_out[2] cb_4_9/io_o_2_out[3] cb_4_9/io_o_2_out[4]
+ cb_4_9/io_o_2_out[5] cb_4_9/io_o_2_out[6] cb_4_9/io_o_2_out[7] cb_4_9/io_o_3_co
+ cb_4_9/io_o_3_out[0] cb_4_9/io_o_3_out[1] cb_4_9/io_o_3_out[2] cb_4_9/io_o_3_out[3]
+ cb_4_9/io_o_3_out[4] cb_4_9/io_o_3_out[5] cb_4_9/io_o_3_out[6] cb_4_9/io_o_3_out[7]
+ cb_4_9/io_o_4_co cb_4_9/io_o_4_out[0] cb_4_9/io_o_4_out[1] cb_4_9/io_o_4_out[2]
+ cb_4_9/io_o_4_out[3] cb_4_9/io_o_4_out[4] cb_4_9/io_o_4_out[5] cb_4_9/io_o_4_out[6]
+ cb_4_9/io_o_4_out[7] cb_4_9/io_o_5_co cb_4_9/io_o_5_out[0] cb_4_9/io_o_5_out[1]
+ cb_4_9/io_o_5_out[2] cb_4_9/io_o_5_out[3] cb_4_9/io_o_5_out[4] cb_4_9/io_o_5_out[5]
+ cb_4_9/io_o_5_out[6] cb_4_9/io_o_5_out[7] cb_4_9/io_o_6_co cb_4_9/io_o_6_out[0]
+ cb_4_9/io_o_6_out[1] cb_4_9/io_o_6_out[2] cb_4_9/io_o_6_out[3] cb_4_9/io_o_6_out[4]
+ cb_4_9/io_o_6_out[5] cb_4_9/io_o_6_out[6] cb_4_9/io_o_6_out[7] cb_4_9/io_o_7_co
+ cb_4_9/io_o_7_out[0] cb_4_9/io_o_7_out[1] cb_4_9/io_o_7_out[2] cb_4_9/io_o_7_out[3]
+ cb_4_9/io_o_7_out[4] cb_4_9/io_o_7_out[5] cb_4_9/io_o_7_out[6] cb_4_9/io_o_7_out[7]
+ cb_4_10/io_o_0_co cb_4_10/io_eo[0] cb_4_10/io_eo[1] cb_4_10/io_eo[2] cb_4_10/io_eo[3]
+ cb_4_10/io_eo[4] cb_4_10/io_eo[5] cb_4_10/io_eo[6] cb_4_10/io_eo[7] cb_4_10/io_o_1_co
+ cb_4_10/io_eo[8] cb_4_10/io_eo[9] cb_4_10/io_eo[10] cb_4_10/io_eo[11] cb_4_10/io_eo[12]
+ cb_4_10/io_eo[13] cb_4_10/io_eo[14] cb_4_10/io_eo[15] cb_4_10/io_o_2_co cb_4_10/io_eo[16]
+ cb_4_10/io_eo[17] cb_4_10/io_eo[18] cb_4_10/io_eo[19] cb_4_10/io_eo[20] cb_4_10/io_eo[21]
+ cb_4_10/io_eo[22] cb_4_10/io_eo[23] cb_4_10/io_o_3_co cb_4_10/io_eo[24] cb_4_10/io_eo[25]
+ cb_4_10/io_eo[26] cb_4_10/io_eo[27] cb_4_10/io_eo[28] cb_4_10/io_eo[29] cb_4_10/io_eo[30]
+ cb_4_10/io_eo[31] cb_4_10/io_o_4_co cb_4_10/io_eo[32] cb_4_10/io_eo[33] cb_4_10/io_eo[34]
+ cb_4_10/io_eo[35] cb_4_10/io_eo[36] cb_4_10/io_eo[37] cb_4_10/io_eo[38] cb_4_10/io_eo[39]
+ cb_4_10/io_o_5_co cb_4_10/io_eo[40] cb_4_10/io_eo[41] cb_4_10/io_eo[42] cb_4_10/io_eo[43]
+ cb_4_10/io_eo[44] cb_4_10/io_eo[45] cb_4_10/io_eo[46] cb_4_10/io_eo[47] cb_4_10/io_o_6_co
+ cb_4_10/io_eo[48] cb_4_10/io_eo[49] cb_4_10/io_eo[50] cb_4_10/io_eo[51] cb_4_10/io_eo[52]
+ cb_4_10/io_eo[53] cb_4_10/io_eo[54] cb_4_10/io_eo[55] cb_4_10/io_o_7_co cb_4_10/io_eo[56]
+ cb_4_10/io_eo[57] cb_4_10/io_eo[58] cb_4_10/io_eo[59] cb_4_10/io_eo[60] cb_4_10/io_eo[61]
+ cb_4_10/io_eo[62] cb_4_10/io_eo[63] cb_4_9/io_vco cb_4_10/io_vco cb_4_10/io_vi cb_4_9/io_we_i
+ cb_4_9/io_eo[0] cb_4_9/io_eo[10] cb_4_9/io_eo[11] cb_4_9/io_eo[12] cb_4_9/io_eo[13]
+ cb_4_9/io_eo[14] cb_4_9/io_eo[15] cb_4_9/io_eo[16] cb_4_9/io_eo[17] cb_4_9/io_eo[18]
+ cb_4_9/io_eo[19] cb_4_9/io_eo[1] cb_4_9/io_eo[20] cb_4_9/io_eo[21] cb_4_9/io_eo[22]
+ cb_4_9/io_eo[23] cb_4_9/io_eo[24] cb_4_9/io_eo[25] cb_4_9/io_eo[26] cb_4_9/io_eo[27]
+ cb_4_9/io_eo[28] cb_4_9/io_eo[29] cb_4_9/io_eo[2] cb_4_9/io_eo[30] cb_4_9/io_eo[31]
+ cb_4_9/io_eo[32] cb_4_9/io_eo[33] cb_4_9/io_eo[34] cb_4_9/io_eo[35] cb_4_9/io_eo[36]
+ cb_4_9/io_eo[37] cb_4_9/io_eo[38] cb_4_9/io_eo[39] cb_4_9/io_eo[3] cb_4_9/io_eo[40]
+ cb_4_9/io_eo[41] cb_4_9/io_eo[42] cb_4_9/io_eo[43] cb_4_9/io_eo[44] cb_4_9/io_eo[45]
+ cb_4_9/io_eo[46] cb_4_9/io_eo[47] cb_4_9/io_eo[48] cb_4_9/io_eo[49] cb_4_9/io_eo[4]
+ cb_4_9/io_eo[50] cb_4_9/io_eo[51] cb_4_9/io_eo[52] cb_4_9/io_eo[53] cb_4_9/io_eo[54]
+ cb_4_9/io_eo[55] cb_4_9/io_eo[56] cb_4_9/io_eo[57] cb_4_9/io_eo[58] cb_4_9/io_eo[59]
+ cb_4_9/io_eo[5] cb_4_9/io_eo[60] cb_4_9/io_eo[61] cb_4_9/io_eo[62] cb_4_9/io_eo[63]
+ cb_4_9/io_eo[6] cb_4_9/io_eo[7] cb_4_9/io_eo[8] cb_4_9/io_eo[9] mcons_3/clock mcons_3/reset
+ vccd1 vssd1 cic_block
Xmcons_2 mcons_3/clock icon/mt_QEI_ChA_2 icon/mt_QEI_ChB_2 mcons_2/io_irq icon/mt_pwm_h_2
+ icon/mt_pwm_l_2 mcons_2/io_wb_ack_o ccon_7/io_adr_i[0] ccon_7/io_adr_i[10] ccon_7/io_adr_i[11]
+ ccon_7/io_adr_i[1] ccon_7/io_adr_i[2] ccon_7/io_adr_i[3] ccon_7/io_adr_i[4] ccon_7/io_adr_i[5]
+ ccon_7/io_adr_i[6] ccon_7/io_adr_i[7] ccon_7/io_adr_i[8] ccon_7/io_adr_i[9] mcons_2/io_wb_cs_i
+ ccon_7/io_dat_i[0] ccon_7/io_dat_i[10] ccon_7/io_dat_i[11] ccon_7/io_dat_i[12] ccon_7/io_dat_i[13]
+ ccon_7/io_dat_i[14] ccon_7/io_dat_i[15] ccon_7/io_dat_i[16] ccon_7/io_dat_i[17]
+ ccon_7/io_dat_i[18] ccon_7/io_dat_i[19] ccon_7/io_dat_i[1] ccon_7/io_dat_i[20] ccon_7/io_dat_i[21]
+ ccon_7/io_dat_i[22] ccon_7/io_dat_i[23] ccon_7/io_dat_i[24] ccon_7/io_dat_i[25]
+ ccon_7/io_dat_i[26] ccon_7/io_dat_i[27] ccon_7/io_dat_i[28] ccon_7/io_dat_i[29]
+ ccon_7/io_dat_i[2] ccon_7/io_dat_i[30] ccon_7/io_dat_i[31] ccon_7/io_dat_i[3] ccon_7/io_dat_i[4]
+ ccon_7/io_dat_i[5] ccon_7/io_dat_i[6] ccon_7/io_dat_i[7] ccon_7/io_dat_i[8] ccon_7/io_dat_i[9]
+ icon/m_wbs_dat_o_2[0] icon/m_wbs_dat_o_2[10] icon/m_wbs_dat_o_2[11] icon/m_wbs_dat_o_2[12]
+ icon/m_wbs_dat_o_2[13] icon/m_wbs_dat_o_2[14] icon/m_wbs_dat_o_2[15] icon/m_wbs_dat_o_2[16]
+ icon/m_wbs_dat_o_2[17] icon/m_wbs_dat_o_2[18] icon/m_wbs_dat_o_2[19] icon/m_wbs_dat_o_2[1]
+ icon/m_wbs_dat_o_2[20] icon/m_wbs_dat_o_2[21] icon/m_wbs_dat_o_2[22] icon/m_wbs_dat_o_2[23]
+ icon/m_wbs_dat_o_2[24] icon/m_wbs_dat_o_2[25] icon/m_wbs_dat_o_2[26] icon/m_wbs_dat_o_2[27]
+ icon/m_wbs_dat_o_2[28] icon/m_wbs_dat_o_2[29] icon/m_wbs_dat_o_2[2] icon/m_wbs_dat_o_2[30]
+ icon/m_wbs_dat_o_2[31] icon/m_wbs_dat_o_2[3] icon/m_wbs_dat_o_2[4] icon/m_wbs_dat_o_2[5]
+ icon/m_wbs_dat_o_2[6] icon/m_wbs_dat_o_2[7] icon/m_wbs_dat_o_2[8] icon/m_wbs_dat_o_2[9]
+ ccon_7/io_we_i mcons_3/reset vccd1 vssd1 motor_top
Xcb_6_3 cb_6_9/io_adr_i[0] cb_6_9/io_adr_i[1] cb_6_3/io_cs_i cb_6_9/io_dat_i[0] cb_6_9/io_dat_i[10]
+ cb_6_9/io_dat_i[11] cb_6_9/io_dat_i[12] cb_6_9/io_dat_i[13] cb_6_9/io_dat_i[14]
+ cb_6_9/io_dat_i[15] cb_6_9/io_dat_i[1] cb_6_9/io_dat_i[2] cb_6_9/io_dat_i[3] cb_6_9/io_dat_i[4]
+ cb_6_9/io_dat_i[5] cb_6_9/io_dat_i[6] cb_6_9/io_dat_i[7] cb_6_9/io_dat_i[8] cb_6_9/io_dat_i[9]
+ cb_6_3/io_dat_o[0] cb_6_3/io_dat_o[10] cb_6_3/io_dat_o[11] cb_6_3/io_dat_o[12] cb_6_3/io_dat_o[13]
+ cb_6_3/io_dat_o[14] cb_6_3/io_dat_o[15] cb_6_3/io_dat_o[1] cb_6_3/io_dat_o[2] cb_6_3/io_dat_o[3]
+ cb_6_3/io_dat_o[4] cb_6_3/io_dat_o[5] cb_6_3/io_dat_o[6] cb_6_3/io_dat_o[7] cb_6_3/io_dat_o[8]
+ cb_6_3/io_dat_o[9] cb_6_4/io_wo[0] cb_6_4/io_wo[10] cb_6_4/io_wo[11] cb_6_4/io_wo[12]
+ cb_6_4/io_wo[13] cb_6_4/io_wo[14] cb_6_4/io_wo[15] cb_6_4/io_wo[16] cb_6_4/io_wo[17]
+ cb_6_4/io_wo[18] cb_6_4/io_wo[19] cb_6_4/io_wo[1] cb_6_4/io_wo[20] cb_6_4/io_wo[21]
+ cb_6_4/io_wo[22] cb_6_4/io_wo[23] cb_6_4/io_wo[24] cb_6_4/io_wo[25] cb_6_4/io_wo[26]
+ cb_6_4/io_wo[27] cb_6_4/io_wo[28] cb_6_4/io_wo[29] cb_6_4/io_wo[2] cb_6_4/io_wo[30]
+ cb_6_4/io_wo[31] cb_6_4/io_wo[32] cb_6_4/io_wo[33] cb_6_4/io_wo[34] cb_6_4/io_wo[35]
+ cb_6_4/io_wo[36] cb_6_4/io_wo[37] cb_6_4/io_wo[38] cb_6_4/io_wo[39] cb_6_4/io_wo[3]
+ cb_6_4/io_wo[40] cb_6_4/io_wo[41] cb_6_4/io_wo[42] cb_6_4/io_wo[43] cb_6_4/io_wo[44]
+ cb_6_4/io_wo[45] cb_6_4/io_wo[46] cb_6_4/io_wo[47] cb_6_4/io_wo[48] cb_6_4/io_wo[49]
+ cb_6_4/io_wo[4] cb_6_4/io_wo[50] cb_6_4/io_wo[51] cb_6_4/io_wo[52] cb_6_4/io_wo[53]
+ cb_6_4/io_wo[54] cb_6_4/io_wo[55] cb_6_4/io_wo[56] cb_6_4/io_wo[57] cb_6_4/io_wo[58]
+ cb_6_4/io_wo[59] cb_6_4/io_wo[5] cb_6_4/io_wo[60] cb_6_4/io_wo[61] cb_6_4/io_wo[62]
+ cb_6_4/io_wo[63] cb_6_4/io_wo[6] cb_6_4/io_wo[7] cb_6_4/io_wo[8] cb_6_4/io_wo[9]
+ cb_6_3/io_i_0_ci cb_6_3/io_i_0_in1[0] cb_6_3/io_i_0_in1[1] cb_6_3/io_i_0_in1[2]
+ cb_6_3/io_i_0_in1[3] cb_6_3/io_i_0_in1[4] cb_6_3/io_i_0_in1[5] cb_6_3/io_i_0_in1[6]
+ cb_6_3/io_i_0_in1[7] cb_6_3/io_i_1_ci cb_6_3/io_i_1_in1[0] cb_6_3/io_i_1_in1[1]
+ cb_6_3/io_i_1_in1[2] cb_6_3/io_i_1_in1[3] cb_6_3/io_i_1_in1[4] cb_6_3/io_i_1_in1[5]
+ cb_6_3/io_i_1_in1[6] cb_6_3/io_i_1_in1[7] cb_6_3/io_i_2_ci cb_6_3/io_i_2_in1[0]
+ cb_6_3/io_i_2_in1[1] cb_6_3/io_i_2_in1[2] cb_6_3/io_i_2_in1[3] cb_6_3/io_i_2_in1[4]
+ cb_6_3/io_i_2_in1[5] cb_6_3/io_i_2_in1[6] cb_6_3/io_i_2_in1[7] cb_6_3/io_i_3_ci
+ cb_6_3/io_i_3_in1[0] cb_6_3/io_i_3_in1[1] cb_6_3/io_i_3_in1[2] cb_6_3/io_i_3_in1[3]
+ cb_6_3/io_i_3_in1[4] cb_6_3/io_i_3_in1[5] cb_6_3/io_i_3_in1[6] cb_6_3/io_i_3_in1[7]
+ cb_6_3/io_i_4_ci cb_6_3/io_i_4_in1[0] cb_6_3/io_i_4_in1[1] cb_6_3/io_i_4_in1[2]
+ cb_6_3/io_i_4_in1[3] cb_6_3/io_i_4_in1[4] cb_6_3/io_i_4_in1[5] cb_6_3/io_i_4_in1[6]
+ cb_6_3/io_i_4_in1[7] cb_6_3/io_i_5_ci cb_6_3/io_i_5_in1[0] cb_6_3/io_i_5_in1[1]
+ cb_6_3/io_i_5_in1[2] cb_6_3/io_i_5_in1[3] cb_6_3/io_i_5_in1[4] cb_6_3/io_i_5_in1[5]
+ cb_6_3/io_i_5_in1[6] cb_6_3/io_i_5_in1[7] cb_6_3/io_i_6_ci cb_6_3/io_i_6_in1[0]
+ cb_6_3/io_i_6_in1[1] cb_6_3/io_i_6_in1[2] cb_6_3/io_i_6_in1[3] cb_6_3/io_i_6_in1[4]
+ cb_6_3/io_i_6_in1[5] cb_6_3/io_i_6_in1[6] cb_6_3/io_i_6_in1[7] cb_6_3/io_i_7_ci
+ cb_6_3/io_i_7_in1[0] cb_6_3/io_i_7_in1[1] cb_6_3/io_i_7_in1[2] cb_6_3/io_i_7_in1[3]
+ cb_6_3/io_i_7_in1[4] cb_6_3/io_i_7_in1[5] cb_6_3/io_i_7_in1[6] cb_6_3/io_i_7_in1[7]
+ cb_6_4/io_i_0_ci cb_6_4/io_i_0_in1[0] cb_6_4/io_i_0_in1[1] cb_6_4/io_i_0_in1[2]
+ cb_6_4/io_i_0_in1[3] cb_6_4/io_i_0_in1[4] cb_6_4/io_i_0_in1[5] cb_6_4/io_i_0_in1[6]
+ cb_6_4/io_i_0_in1[7] cb_6_4/io_i_1_ci cb_6_4/io_i_1_in1[0] cb_6_4/io_i_1_in1[1]
+ cb_6_4/io_i_1_in1[2] cb_6_4/io_i_1_in1[3] cb_6_4/io_i_1_in1[4] cb_6_4/io_i_1_in1[5]
+ cb_6_4/io_i_1_in1[6] cb_6_4/io_i_1_in1[7] cb_6_4/io_i_2_ci cb_6_4/io_i_2_in1[0]
+ cb_6_4/io_i_2_in1[1] cb_6_4/io_i_2_in1[2] cb_6_4/io_i_2_in1[3] cb_6_4/io_i_2_in1[4]
+ cb_6_4/io_i_2_in1[5] cb_6_4/io_i_2_in1[6] cb_6_4/io_i_2_in1[7] cb_6_4/io_i_3_ci
+ cb_6_4/io_i_3_in1[0] cb_6_4/io_i_3_in1[1] cb_6_4/io_i_3_in1[2] cb_6_4/io_i_3_in1[3]
+ cb_6_4/io_i_3_in1[4] cb_6_4/io_i_3_in1[5] cb_6_4/io_i_3_in1[6] cb_6_4/io_i_3_in1[7]
+ cb_6_4/io_i_4_ci cb_6_4/io_i_4_in1[0] cb_6_4/io_i_4_in1[1] cb_6_4/io_i_4_in1[2]
+ cb_6_4/io_i_4_in1[3] cb_6_4/io_i_4_in1[4] cb_6_4/io_i_4_in1[5] cb_6_4/io_i_4_in1[6]
+ cb_6_4/io_i_4_in1[7] cb_6_4/io_i_5_ci cb_6_4/io_i_5_in1[0] cb_6_4/io_i_5_in1[1]
+ cb_6_4/io_i_5_in1[2] cb_6_4/io_i_5_in1[3] cb_6_4/io_i_5_in1[4] cb_6_4/io_i_5_in1[5]
+ cb_6_4/io_i_5_in1[6] cb_6_4/io_i_5_in1[7] cb_6_4/io_i_6_ci cb_6_4/io_i_6_in1[0]
+ cb_6_4/io_i_6_in1[1] cb_6_4/io_i_6_in1[2] cb_6_4/io_i_6_in1[3] cb_6_4/io_i_6_in1[4]
+ cb_6_4/io_i_6_in1[5] cb_6_4/io_i_6_in1[6] cb_6_4/io_i_6_in1[7] cb_6_4/io_i_7_ci
+ cb_6_4/io_i_7_in1[0] cb_6_4/io_i_7_in1[1] cb_6_4/io_i_7_in1[2] cb_6_4/io_i_7_in1[3]
+ cb_6_4/io_i_7_in1[4] cb_6_4/io_i_7_in1[5] cb_6_4/io_i_7_in1[6] cb_6_4/io_i_7_in1[7]
+ cb_6_3/io_vci cb_6_4/io_vci cb_6_3/io_vi cb_6_9/io_we_i cb_6_3/io_wo[0] cb_6_3/io_wo[10]
+ cb_6_3/io_wo[11] cb_6_3/io_wo[12] cb_6_3/io_wo[13] cb_6_3/io_wo[14] cb_6_3/io_wo[15]
+ cb_6_3/io_wo[16] cb_6_3/io_wo[17] cb_6_3/io_wo[18] cb_6_3/io_wo[19] cb_6_3/io_wo[1]
+ cb_6_3/io_wo[20] cb_6_3/io_wo[21] cb_6_3/io_wo[22] cb_6_3/io_wo[23] cb_6_3/io_wo[24]
+ cb_6_3/io_wo[25] cb_6_3/io_wo[26] cb_6_3/io_wo[27] cb_6_3/io_wo[28] cb_6_3/io_wo[29]
+ cb_6_3/io_wo[2] cb_6_3/io_wo[30] cb_6_3/io_wo[31] cb_6_3/io_wo[32] cb_6_3/io_wo[33]
+ cb_6_3/io_wo[34] cb_6_3/io_wo[35] cb_6_3/io_wo[36] cb_6_3/io_wo[37] cb_6_3/io_wo[38]
+ cb_6_3/io_wo[39] cb_6_3/io_wo[3] cb_6_3/io_wo[40] cb_6_3/io_wo[41] cb_6_3/io_wo[42]
+ cb_6_3/io_wo[43] cb_6_3/io_wo[44] cb_6_3/io_wo[45] cb_6_3/io_wo[46] cb_6_3/io_wo[47]
+ cb_6_3/io_wo[48] cb_6_3/io_wo[49] cb_6_3/io_wo[4] cb_6_3/io_wo[50] cb_6_3/io_wo[51]
+ cb_6_3/io_wo[52] cb_6_3/io_wo[53] cb_6_3/io_wo[54] cb_6_3/io_wo[55] cb_6_3/io_wo[56]
+ cb_6_3/io_wo[57] cb_6_3/io_wo[58] cb_6_3/io_wo[59] cb_6_3/io_wo[5] cb_6_3/io_wo[60]
+ cb_6_3/io_wo[61] cb_6_3/io_wo[62] cb_6_3/io_wo[63] cb_6_3/io_wo[6] cb_6_3/io_wo[7]
+ cb_6_3/io_wo[8] cb_6_3/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_7_10 cb_7_9/io_adr_i[0] cb_7_9/io_adr_i[1] cb_7_10/io_cs_i cb_7_9/io_dat_i[0]
+ cb_7_9/io_dat_i[10] cb_7_9/io_dat_i[11] cb_7_9/io_dat_i[12] cb_7_9/io_dat_i[13]
+ cb_7_9/io_dat_i[14] cb_7_9/io_dat_i[15] cb_7_9/io_dat_i[1] cb_7_9/io_dat_i[2] cb_7_9/io_dat_i[3]
+ cb_7_9/io_dat_i[4] cb_7_9/io_dat_i[5] cb_7_9/io_dat_i[6] cb_7_9/io_dat_i[7] cb_7_9/io_dat_i[8]
+ cb_7_9/io_dat_i[9] cb_7_10/io_dat_o[0] cb_7_10/io_dat_o[10] cb_7_10/io_dat_o[11]
+ cb_7_10/io_dat_o[12] cb_7_10/io_dat_o[13] cb_7_10/io_dat_o[14] cb_7_10/io_dat_o[15]
+ cb_7_10/io_dat_o[1] cb_7_10/io_dat_o[2] cb_7_10/io_dat_o[3] cb_7_10/io_dat_o[4]
+ cb_7_10/io_dat_o[5] cb_7_10/io_dat_o[6] cb_7_10/io_dat_o[7] cb_7_10/io_dat_o[8]
+ cb_7_10/io_dat_o[9] cb_7_10/io_eo[0] cb_7_10/io_eo[10] cb_7_10/io_eo[11] cb_7_10/io_eo[12]
+ cb_7_10/io_eo[13] cb_7_10/io_eo[14] cb_7_10/io_eo[15] cb_7_10/io_eo[16] cb_7_10/io_eo[17]
+ cb_7_10/io_eo[18] cb_7_10/io_eo[19] cb_7_10/io_eo[1] cb_7_10/io_eo[20] cb_7_10/io_eo[21]
+ cb_7_10/io_eo[22] cb_7_10/io_eo[23] cb_7_10/io_eo[24] cb_7_10/io_eo[25] cb_7_10/io_eo[26]
+ cb_7_10/io_eo[27] cb_7_10/io_eo[28] cb_7_10/io_eo[29] cb_7_10/io_eo[2] cb_7_10/io_eo[30]
+ cb_7_10/io_eo[31] cb_7_10/io_eo[32] cb_7_10/io_eo[33] cb_7_10/io_eo[34] cb_7_10/io_eo[35]
+ cb_7_10/io_eo[36] cb_7_10/io_eo[37] cb_7_10/io_eo[38] cb_7_10/io_eo[39] cb_7_10/io_eo[3]
+ cb_7_10/io_eo[40] cb_7_10/io_eo[41] cb_7_10/io_eo[42] cb_7_10/io_eo[43] cb_7_10/io_eo[44]
+ cb_7_10/io_eo[45] cb_7_10/io_eo[46] cb_7_10/io_eo[47] cb_7_10/io_eo[48] cb_7_10/io_eo[49]
+ cb_7_10/io_eo[4] cb_7_10/io_eo[50] cb_7_10/io_eo[51] cb_7_10/io_eo[52] cb_7_10/io_eo[53]
+ cb_7_10/io_eo[54] cb_7_10/io_eo[55] cb_7_10/io_eo[56] cb_7_10/io_eo[57] cb_7_10/io_eo[58]
+ cb_7_10/io_eo[59] cb_7_10/io_eo[5] cb_7_10/io_eo[60] cb_7_10/io_eo[61] cb_7_10/io_eo[62]
+ cb_7_10/io_eo[63] cb_7_10/io_eo[6] cb_7_10/io_eo[7] cb_7_10/io_eo[8] cb_7_10/io_eo[9]
+ cb_7_9/io_o_0_co cb_7_9/io_o_0_out[0] cb_7_9/io_o_0_out[1] cb_7_9/io_o_0_out[2]
+ cb_7_9/io_o_0_out[3] cb_7_9/io_o_0_out[4] cb_7_9/io_o_0_out[5] cb_7_9/io_o_0_out[6]
+ cb_7_9/io_o_0_out[7] cb_7_9/io_o_1_co cb_7_9/io_o_1_out[0] cb_7_9/io_o_1_out[1]
+ cb_7_9/io_o_1_out[2] cb_7_9/io_o_1_out[3] cb_7_9/io_o_1_out[4] cb_7_9/io_o_1_out[5]
+ cb_7_9/io_o_1_out[6] cb_7_9/io_o_1_out[7] cb_7_9/io_o_2_co cb_7_9/io_o_2_out[0]
+ cb_7_9/io_o_2_out[1] cb_7_9/io_o_2_out[2] cb_7_9/io_o_2_out[3] cb_7_9/io_o_2_out[4]
+ cb_7_9/io_o_2_out[5] cb_7_9/io_o_2_out[6] cb_7_9/io_o_2_out[7] cb_7_9/io_o_3_co
+ cb_7_9/io_o_3_out[0] cb_7_9/io_o_3_out[1] cb_7_9/io_o_3_out[2] cb_7_9/io_o_3_out[3]
+ cb_7_9/io_o_3_out[4] cb_7_9/io_o_3_out[5] cb_7_9/io_o_3_out[6] cb_7_9/io_o_3_out[7]
+ cb_7_9/io_o_4_co cb_7_9/io_o_4_out[0] cb_7_9/io_o_4_out[1] cb_7_9/io_o_4_out[2]
+ cb_7_9/io_o_4_out[3] cb_7_9/io_o_4_out[4] cb_7_9/io_o_4_out[5] cb_7_9/io_o_4_out[6]
+ cb_7_9/io_o_4_out[7] cb_7_9/io_o_5_co cb_7_9/io_o_5_out[0] cb_7_9/io_o_5_out[1]
+ cb_7_9/io_o_5_out[2] cb_7_9/io_o_5_out[3] cb_7_9/io_o_5_out[4] cb_7_9/io_o_5_out[5]
+ cb_7_9/io_o_5_out[6] cb_7_9/io_o_5_out[7] cb_7_9/io_o_6_co cb_7_9/io_o_6_out[0]
+ cb_7_9/io_o_6_out[1] cb_7_9/io_o_6_out[2] cb_7_9/io_o_6_out[3] cb_7_9/io_o_6_out[4]
+ cb_7_9/io_o_6_out[5] cb_7_9/io_o_6_out[6] cb_7_9/io_o_6_out[7] cb_7_9/io_o_7_co
+ cb_7_9/io_o_7_out[0] cb_7_9/io_o_7_out[1] cb_7_9/io_o_7_out[2] cb_7_9/io_o_7_out[3]
+ cb_7_9/io_o_7_out[4] cb_7_9/io_o_7_out[5] cb_7_9/io_o_7_out[6] cb_7_9/io_o_7_out[7]
+ cb_7_10/io_o_0_co cb_7_10/io_eo[0] cb_7_10/io_eo[1] cb_7_10/io_eo[2] cb_7_10/io_eo[3]
+ cb_7_10/io_eo[4] cb_7_10/io_eo[5] cb_7_10/io_eo[6] cb_7_10/io_eo[7] cb_7_10/io_o_1_co
+ cb_7_10/io_eo[8] cb_7_10/io_eo[9] cb_7_10/io_eo[10] cb_7_10/io_eo[11] cb_7_10/io_eo[12]
+ cb_7_10/io_eo[13] cb_7_10/io_eo[14] cb_7_10/io_eo[15] cb_7_10/io_o_2_co cb_7_10/io_eo[16]
+ cb_7_10/io_eo[17] cb_7_10/io_eo[18] cb_7_10/io_eo[19] cb_7_10/io_eo[20] cb_7_10/io_eo[21]
+ cb_7_10/io_eo[22] cb_7_10/io_eo[23] cb_7_10/io_o_3_co cb_7_10/io_eo[24] cb_7_10/io_eo[25]
+ cb_7_10/io_eo[26] cb_7_10/io_eo[27] cb_7_10/io_eo[28] cb_7_10/io_eo[29] cb_7_10/io_eo[30]
+ cb_7_10/io_eo[31] cb_7_10/io_o_4_co cb_7_10/io_eo[32] cb_7_10/io_eo[33] cb_7_10/io_eo[34]
+ cb_7_10/io_eo[35] cb_7_10/io_eo[36] cb_7_10/io_eo[37] cb_7_10/io_eo[38] cb_7_10/io_eo[39]
+ cb_7_10/io_o_5_co cb_7_10/io_eo[40] cb_7_10/io_eo[41] cb_7_10/io_eo[42] cb_7_10/io_eo[43]
+ cb_7_10/io_eo[44] cb_7_10/io_eo[45] cb_7_10/io_eo[46] cb_7_10/io_eo[47] cb_7_10/io_o_6_co
+ cb_7_10/io_eo[48] cb_7_10/io_eo[49] cb_7_10/io_eo[50] cb_7_10/io_eo[51] cb_7_10/io_eo[52]
+ cb_7_10/io_eo[53] cb_7_10/io_eo[54] cb_7_10/io_eo[55] cb_7_10/io_o_7_co cb_7_10/io_eo[56]
+ cb_7_10/io_eo[57] cb_7_10/io_eo[58] cb_7_10/io_eo[59] cb_7_10/io_eo[60] cb_7_10/io_eo[61]
+ cb_7_10/io_eo[62] cb_7_10/io_eo[63] cb_7_9/io_vco cb_7_10/io_vco cb_7_10/io_vi cb_7_9/io_we_i
+ cb_7_9/io_eo[0] cb_7_9/io_eo[10] cb_7_9/io_eo[11] cb_7_9/io_eo[12] cb_7_9/io_eo[13]
+ cb_7_9/io_eo[14] cb_7_9/io_eo[15] cb_7_9/io_eo[16] cb_7_9/io_eo[17] cb_7_9/io_eo[18]
+ cb_7_9/io_eo[19] cb_7_9/io_eo[1] cb_7_9/io_eo[20] cb_7_9/io_eo[21] cb_7_9/io_eo[22]
+ cb_7_9/io_eo[23] cb_7_9/io_eo[24] cb_7_9/io_eo[25] cb_7_9/io_eo[26] cb_7_9/io_eo[27]
+ cb_7_9/io_eo[28] cb_7_9/io_eo[29] cb_7_9/io_eo[2] cb_7_9/io_eo[30] cb_7_9/io_eo[31]
+ cb_7_9/io_eo[32] cb_7_9/io_eo[33] cb_7_9/io_eo[34] cb_7_9/io_eo[35] cb_7_9/io_eo[36]
+ cb_7_9/io_eo[37] cb_7_9/io_eo[38] cb_7_9/io_eo[39] cb_7_9/io_eo[3] cb_7_9/io_eo[40]
+ cb_7_9/io_eo[41] cb_7_9/io_eo[42] cb_7_9/io_eo[43] cb_7_9/io_eo[44] cb_7_9/io_eo[45]
+ cb_7_9/io_eo[46] cb_7_9/io_eo[47] cb_7_9/io_eo[48] cb_7_9/io_eo[49] cb_7_9/io_eo[4]
+ cb_7_9/io_eo[50] cb_7_9/io_eo[51] cb_7_9/io_eo[52] cb_7_9/io_eo[53] cb_7_9/io_eo[54]
+ cb_7_9/io_eo[55] cb_7_9/io_eo[56] cb_7_9/io_eo[57] cb_7_9/io_eo[58] cb_7_9/io_eo[59]
+ cb_7_9/io_eo[5] cb_7_9/io_eo[60] cb_7_9/io_eo[61] cb_7_9/io_eo[62] cb_7_9/io_eo[63]
+ cb_7_9/io_eo[6] cb_7_9/io_eo[7] cb_7_9/io_eo[8] cb_7_9/io_eo[9] mcons_3/clock mcons_3/reset
+ vccd1 vssd1 cic_block
Xcb_4_0 cb_4_9/io_adr_i[0] cb_4_9/io_adr_i[1] cb_4_0/io_cs_i cb_4_9/io_dat_i[0] cb_4_9/io_dat_i[10]
+ cb_4_9/io_dat_i[11] cb_4_9/io_dat_i[12] cb_4_9/io_dat_i[13] cb_4_9/io_dat_i[14]
+ cb_4_9/io_dat_i[15] cb_4_9/io_dat_i[1] cb_4_9/io_dat_i[2] cb_4_9/io_dat_i[3] cb_4_9/io_dat_i[4]
+ cb_4_9/io_dat_i[5] cb_4_9/io_dat_i[6] cb_4_9/io_dat_i[7] cb_4_9/io_dat_i[8] cb_4_9/io_dat_i[9]
+ cb_4_0/io_dat_o[0] cb_4_0/io_dat_o[10] cb_4_0/io_dat_o[11] cb_4_0/io_dat_o[12] cb_4_0/io_dat_o[13]
+ cb_4_0/io_dat_o[14] cb_4_0/io_dat_o[15] cb_4_0/io_dat_o[1] cb_4_0/io_dat_o[2] cb_4_0/io_dat_o[3]
+ cb_4_0/io_dat_o[4] cb_4_0/io_dat_o[5] cb_4_0/io_dat_o[6] cb_4_0/io_dat_o[7] cb_4_0/io_dat_o[8]
+ cb_4_0/io_dat_o[9] cb_4_1/io_wo[0] cb_4_1/io_wo[10] cb_4_1/io_wo[11] cb_4_1/io_wo[12]
+ cb_4_1/io_wo[13] cb_4_1/io_wo[14] cb_4_1/io_wo[15] cb_4_1/io_wo[16] cb_4_1/io_wo[17]
+ cb_4_1/io_wo[18] cb_4_1/io_wo[19] cb_4_1/io_wo[1] cb_4_1/io_wo[20] cb_4_1/io_wo[21]
+ cb_4_1/io_wo[22] cb_4_1/io_wo[23] cb_4_1/io_wo[24] cb_4_1/io_wo[25] cb_4_1/io_wo[26]
+ cb_4_1/io_wo[27] cb_4_1/io_wo[28] cb_4_1/io_wo[29] cb_4_1/io_wo[2] cb_4_1/io_wo[30]
+ cb_4_1/io_wo[31] cb_4_1/io_wo[32] cb_4_1/io_wo[33] cb_4_1/io_wo[34] cb_4_1/io_wo[35]
+ cb_4_1/io_wo[36] cb_4_1/io_wo[37] cb_4_1/io_wo[38] cb_4_1/io_wo[39] cb_4_1/io_wo[3]
+ cb_4_1/io_wo[40] cb_4_1/io_wo[41] cb_4_1/io_wo[42] cb_4_1/io_wo[43] cb_4_1/io_wo[44]
+ cb_4_1/io_wo[45] cb_4_1/io_wo[46] cb_4_1/io_wo[47] cb_4_1/io_wo[48] cb_4_1/io_wo[49]
+ cb_4_1/io_wo[4] cb_4_1/io_wo[50] cb_4_1/io_wo[51] cb_4_1/io_wo[52] cb_4_1/io_wo[53]
+ cb_4_1/io_wo[54] cb_4_1/io_wo[55] cb_4_1/io_wo[56] cb_4_1/io_wo[57] cb_4_1/io_wo[58]
+ cb_4_1/io_wo[59] cb_4_1/io_wo[5] cb_4_1/io_wo[60] cb_4_1/io_wo[61] cb_4_1/io_wo[62]
+ cb_4_1/io_wo[63] cb_4_1/io_wo[6] cb_4_1/io_wo[7] cb_4_1/io_wo[8] cb_4_1/io_wo[9]
+ ccon_4/io_dsi_o cb_4_0/io_i_0_in1[0] cb_4_0/io_i_0_in1[1] cb_4_0/io_i_0_in1[2] cb_4_0/io_i_0_in1[3]
+ cb_4_0/io_i_0_in1[4] cb_4_0/io_i_0_in1[5] cb_4_0/io_i_0_in1[6] cb_4_0/io_i_0_in1[7]
+ cb_4_0/io_i_1_ci cb_4_0/io_i_1_in1[0] cb_4_0/io_i_1_in1[1] cb_4_0/io_i_1_in1[2]
+ cb_4_0/io_i_1_in1[3] cb_4_0/io_i_1_in1[4] cb_4_0/io_i_1_in1[5] cb_4_0/io_i_1_in1[6]
+ cb_4_0/io_i_1_in1[7] cb_4_0/io_i_2_ci cb_4_0/io_i_2_in1[0] cb_4_0/io_i_2_in1[1]
+ cb_4_0/io_i_2_in1[2] cb_4_0/io_i_2_in1[3] cb_4_0/io_i_2_in1[4] cb_4_0/io_i_2_in1[5]
+ cb_4_0/io_i_2_in1[6] cb_4_0/io_i_2_in1[7] cb_4_0/io_i_3_ci cb_4_0/io_i_3_in1[0]
+ cb_4_0/io_i_3_in1[1] cb_4_0/io_i_3_in1[2] cb_4_0/io_i_3_in1[3] cb_4_0/io_i_3_in1[4]
+ cb_4_0/io_i_3_in1[5] cb_4_0/io_i_3_in1[6] cb_4_0/io_i_3_in1[7] cb_4_0/io_i_4_ci
+ cb_4_0/io_i_4_in1[0] cb_4_0/io_i_4_in1[1] cb_4_0/io_i_4_in1[2] cb_4_0/io_i_4_in1[3]
+ cb_4_0/io_i_4_in1[4] cb_4_0/io_i_4_in1[5] cb_4_0/io_i_4_in1[6] cb_4_0/io_i_4_in1[7]
+ cb_4_0/io_i_5_ci cb_4_0/io_i_5_in1[0] cb_4_0/io_i_5_in1[1] cb_4_0/io_i_5_in1[2]
+ cb_4_0/io_i_5_in1[3] cb_4_0/io_i_5_in1[4] cb_4_0/io_i_5_in1[5] cb_4_0/io_i_5_in1[6]
+ cb_4_0/io_i_5_in1[7] cb_4_0/io_i_6_ci cb_4_0/io_i_6_in1[0] cb_4_0/io_i_6_in1[1]
+ cb_4_0/io_i_6_in1[2] cb_4_0/io_i_6_in1[3] cb_4_0/io_i_6_in1[4] cb_4_0/io_i_6_in1[5]
+ cb_4_0/io_i_6_in1[6] cb_4_0/io_i_6_in1[7] cb_4_0/io_i_7_ci cb_4_0/io_i_7_in1[0]
+ cb_4_0/io_i_7_in1[1] cb_4_0/io_i_7_in1[2] cb_4_0/io_i_7_in1[3] cb_4_0/io_i_7_in1[4]
+ cb_4_0/io_i_7_in1[5] cb_4_0/io_i_7_in1[6] cb_4_0/io_i_7_in1[7] cb_4_1/io_i_0_ci
+ cb_4_1/io_i_0_in1[0] cb_4_1/io_i_0_in1[1] cb_4_1/io_i_0_in1[2] cb_4_1/io_i_0_in1[3]
+ cb_4_1/io_i_0_in1[4] cb_4_1/io_i_0_in1[5] cb_4_1/io_i_0_in1[6] cb_4_1/io_i_0_in1[7]
+ cb_4_1/io_i_1_ci cb_4_1/io_i_1_in1[0] cb_4_1/io_i_1_in1[1] cb_4_1/io_i_1_in1[2]
+ cb_4_1/io_i_1_in1[3] cb_4_1/io_i_1_in1[4] cb_4_1/io_i_1_in1[5] cb_4_1/io_i_1_in1[6]
+ cb_4_1/io_i_1_in1[7] cb_4_1/io_i_2_ci cb_4_1/io_i_2_in1[0] cb_4_1/io_i_2_in1[1]
+ cb_4_1/io_i_2_in1[2] cb_4_1/io_i_2_in1[3] cb_4_1/io_i_2_in1[4] cb_4_1/io_i_2_in1[5]
+ cb_4_1/io_i_2_in1[6] cb_4_1/io_i_2_in1[7] cb_4_1/io_i_3_ci cb_4_1/io_i_3_in1[0]
+ cb_4_1/io_i_3_in1[1] cb_4_1/io_i_3_in1[2] cb_4_1/io_i_3_in1[3] cb_4_1/io_i_3_in1[4]
+ cb_4_1/io_i_3_in1[5] cb_4_1/io_i_3_in1[6] cb_4_1/io_i_3_in1[7] cb_4_1/io_i_4_ci
+ cb_4_1/io_i_4_in1[0] cb_4_1/io_i_4_in1[1] cb_4_1/io_i_4_in1[2] cb_4_1/io_i_4_in1[3]
+ cb_4_1/io_i_4_in1[4] cb_4_1/io_i_4_in1[5] cb_4_1/io_i_4_in1[6] cb_4_1/io_i_4_in1[7]
+ cb_4_1/io_i_5_ci cb_4_1/io_i_5_in1[0] cb_4_1/io_i_5_in1[1] cb_4_1/io_i_5_in1[2]
+ cb_4_1/io_i_5_in1[3] cb_4_1/io_i_5_in1[4] cb_4_1/io_i_5_in1[5] cb_4_1/io_i_5_in1[6]
+ cb_4_1/io_i_5_in1[7] cb_4_1/io_i_6_ci cb_4_1/io_i_6_in1[0] cb_4_1/io_i_6_in1[1]
+ cb_4_1/io_i_6_in1[2] cb_4_1/io_i_6_in1[3] cb_4_1/io_i_6_in1[4] cb_4_1/io_i_6_in1[5]
+ cb_4_1/io_i_6_in1[6] cb_4_1/io_i_6_in1[7] cb_4_1/io_i_7_ci cb_4_1/io_i_7_in1[0]
+ cb_4_1/io_i_7_in1[1] cb_4_1/io_i_7_in1[2] cb_4_1/io_i_7_in1[3] cb_4_1/io_i_7_in1[4]
+ cb_4_1/io_i_7_in1[5] cb_4_1/io_i_7_in1[6] cb_4_1/io_i_7_in1[7] cb_4_0/io_vci cb_4_1/io_vci
+ cb_4_0/io_vi cb_4_9/io_we_i cb_4_0/io_wo[0] cb_4_0/io_wo[10] cb_4_0/io_wo[11] cb_4_0/io_wo[12]
+ cb_4_0/io_wo[13] cb_4_0/io_wo[14] cb_4_0/io_wo[15] cb_4_0/io_wo[16] cb_4_0/io_wo[17]
+ cb_4_0/io_wo[18] cb_4_0/io_wo[19] cb_4_0/io_wo[1] cb_4_0/io_wo[20] cb_4_0/io_wo[21]
+ cb_4_0/io_wo[22] cb_4_0/io_wo[23] cb_4_0/io_wo[24] cb_4_0/io_wo[25] cb_4_0/io_wo[26]
+ cb_4_0/io_wo[27] cb_4_0/io_wo[28] cb_4_0/io_wo[29] cb_4_0/io_wo[2] cb_4_0/io_wo[30]
+ cb_4_0/io_wo[31] cb_4_0/io_wo[32] cb_4_0/io_wo[33] cb_4_0/io_wo[34] cb_4_0/io_wo[35]
+ cb_4_0/io_wo[36] cb_4_0/io_wo[37] cb_4_0/io_wo[38] cb_4_0/io_wo[39] cb_4_0/io_wo[3]
+ cb_4_0/io_wo[40] cb_4_0/io_wo[41] cb_4_0/io_wo[42] cb_4_0/io_wo[43] cb_4_0/io_wo[44]
+ cb_4_0/io_wo[45] cb_4_0/io_wo[46] cb_4_0/io_wo[47] cb_4_0/io_wo[48] cb_4_0/io_wo[49]
+ cb_4_0/io_wo[4] cb_4_0/io_wo[50] cb_4_0/io_wo[51] cb_4_0/io_wo[52] cb_4_0/io_wo[53]
+ cb_4_0/io_wo[54] cb_4_0/io_wo[55] cb_4_0/io_wo[56] cb_4_0/io_wo[57] cb_4_0/io_wo[58]
+ cb_4_0/io_wo[59] cb_4_0/io_wo[5] cb_4_0/io_wo[60] cb_4_0/io_wo[61] cb_4_0/io_wo[62]
+ cb_4_0/io_wo[63] cb_4_0/io_wo[6] cb_4_0/io_wo[7] cb_4_0/io_wo[8] cb_4_0/io_wo[9]
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xmcons_3 mcons_3/clock icon/mt_QEI_ChA_3 icon/mt_QEI_ChB_3 mcons_3/io_irq icon/mt_pwm_h_3
+ icon/mt_pwm_l_3 mcons_3/io_wb_ack_o ccon_7/io_adr_i[0] ccon_7/io_adr_i[10] ccon_7/io_adr_i[11]
+ ccon_7/io_adr_i[1] ccon_7/io_adr_i[2] ccon_7/io_adr_i[3] ccon_7/io_adr_i[4] ccon_7/io_adr_i[5]
+ ccon_7/io_adr_i[6] ccon_7/io_adr_i[7] ccon_7/io_adr_i[8] ccon_7/io_adr_i[9] mcons_3/io_wb_cs_i
+ ccon_7/io_dat_i[0] ccon_7/io_dat_i[10] ccon_7/io_dat_i[11] ccon_7/io_dat_i[12] ccon_7/io_dat_i[13]
+ ccon_7/io_dat_i[14] ccon_7/io_dat_i[15] ccon_7/io_dat_i[16] ccon_7/io_dat_i[17]
+ ccon_7/io_dat_i[18] ccon_7/io_dat_i[19] ccon_7/io_dat_i[1] ccon_7/io_dat_i[20] ccon_7/io_dat_i[21]
+ ccon_7/io_dat_i[22] ccon_7/io_dat_i[23] ccon_7/io_dat_i[24] ccon_7/io_dat_i[25]
+ ccon_7/io_dat_i[26] ccon_7/io_dat_i[27] ccon_7/io_dat_i[28] ccon_7/io_dat_i[29]
+ ccon_7/io_dat_i[2] ccon_7/io_dat_i[30] ccon_7/io_dat_i[31] ccon_7/io_dat_i[3] ccon_7/io_dat_i[4]
+ ccon_7/io_dat_i[5] ccon_7/io_dat_i[6] ccon_7/io_dat_i[7] ccon_7/io_dat_i[8] ccon_7/io_dat_i[9]
+ icon/m_wbs_dat_o_3[0] icon/m_wbs_dat_o_3[10] icon/m_wbs_dat_o_3[11] icon/m_wbs_dat_o_3[12]
+ icon/m_wbs_dat_o_3[13] icon/m_wbs_dat_o_3[14] icon/m_wbs_dat_o_3[15] icon/m_wbs_dat_o_3[16]
+ icon/m_wbs_dat_o_3[17] icon/m_wbs_dat_o_3[18] icon/m_wbs_dat_o_3[19] icon/m_wbs_dat_o_3[1]
+ icon/m_wbs_dat_o_3[20] icon/m_wbs_dat_o_3[21] icon/m_wbs_dat_o_3[22] icon/m_wbs_dat_o_3[23]
+ icon/m_wbs_dat_o_3[24] icon/m_wbs_dat_o_3[25] icon/m_wbs_dat_o_3[26] icon/m_wbs_dat_o_3[27]
+ icon/m_wbs_dat_o_3[28] icon/m_wbs_dat_o_3[29] icon/m_wbs_dat_o_3[2] icon/m_wbs_dat_o_3[30]
+ icon/m_wbs_dat_o_3[31] icon/m_wbs_dat_o_3[3] icon/m_wbs_dat_o_3[4] icon/m_wbs_dat_o_3[5]
+ icon/m_wbs_dat_o_3[6] icon/m_wbs_dat_o_3[7] icon/m_wbs_dat_o_3[8] icon/m_wbs_dat_o_3[9]
+ ccon_7/io_we_i mcons_3/reset vccd1 vssd1 motor_top
Xcb_6_4 cb_6_9/io_adr_i[0] cb_6_9/io_adr_i[1] cb_6_4/io_cs_i cb_6_9/io_dat_i[0] cb_6_9/io_dat_i[10]
+ cb_6_9/io_dat_i[11] cb_6_9/io_dat_i[12] cb_6_9/io_dat_i[13] cb_6_9/io_dat_i[14]
+ cb_6_9/io_dat_i[15] cb_6_9/io_dat_i[1] cb_6_9/io_dat_i[2] cb_6_9/io_dat_i[3] cb_6_9/io_dat_i[4]
+ cb_6_9/io_dat_i[5] cb_6_9/io_dat_i[6] cb_6_9/io_dat_i[7] cb_6_9/io_dat_i[8] cb_6_9/io_dat_i[9]
+ cb_6_4/io_dat_o[0] cb_6_4/io_dat_o[10] cb_6_4/io_dat_o[11] cb_6_4/io_dat_o[12] cb_6_4/io_dat_o[13]
+ cb_6_4/io_dat_o[14] cb_6_4/io_dat_o[15] cb_6_4/io_dat_o[1] cb_6_4/io_dat_o[2] cb_6_4/io_dat_o[3]
+ cb_6_4/io_dat_o[4] cb_6_4/io_dat_o[5] cb_6_4/io_dat_o[6] cb_6_4/io_dat_o[7] cb_6_4/io_dat_o[8]
+ cb_6_4/io_dat_o[9] cb_6_5/io_wo[0] cb_6_5/io_wo[10] cb_6_5/io_wo[11] cb_6_5/io_wo[12]
+ cb_6_5/io_wo[13] cb_6_5/io_wo[14] cb_6_5/io_wo[15] cb_6_5/io_wo[16] cb_6_5/io_wo[17]
+ cb_6_5/io_wo[18] cb_6_5/io_wo[19] cb_6_5/io_wo[1] cb_6_5/io_wo[20] cb_6_5/io_wo[21]
+ cb_6_5/io_wo[22] cb_6_5/io_wo[23] cb_6_5/io_wo[24] cb_6_5/io_wo[25] cb_6_5/io_wo[26]
+ cb_6_5/io_wo[27] cb_6_5/io_wo[28] cb_6_5/io_wo[29] cb_6_5/io_wo[2] cb_6_5/io_wo[30]
+ cb_6_5/io_wo[31] cb_6_5/io_wo[32] cb_6_5/io_wo[33] cb_6_5/io_wo[34] cb_6_5/io_wo[35]
+ cb_6_5/io_wo[36] cb_6_5/io_wo[37] cb_6_5/io_wo[38] cb_6_5/io_wo[39] cb_6_5/io_wo[3]
+ cb_6_5/io_wo[40] cb_6_5/io_wo[41] cb_6_5/io_wo[42] cb_6_5/io_wo[43] cb_6_5/io_wo[44]
+ cb_6_5/io_wo[45] cb_6_5/io_wo[46] cb_6_5/io_wo[47] cb_6_5/io_wo[48] cb_6_5/io_wo[49]
+ cb_6_5/io_wo[4] cb_6_5/io_wo[50] cb_6_5/io_wo[51] cb_6_5/io_wo[52] cb_6_5/io_wo[53]
+ cb_6_5/io_wo[54] cb_6_5/io_wo[55] cb_6_5/io_wo[56] cb_6_5/io_wo[57] cb_6_5/io_wo[58]
+ cb_6_5/io_wo[59] cb_6_5/io_wo[5] cb_6_5/io_wo[60] cb_6_5/io_wo[61] cb_6_5/io_wo[62]
+ cb_6_5/io_wo[63] cb_6_5/io_wo[6] cb_6_5/io_wo[7] cb_6_5/io_wo[8] cb_6_5/io_wo[9]
+ cb_6_4/io_i_0_ci cb_6_4/io_i_0_in1[0] cb_6_4/io_i_0_in1[1] cb_6_4/io_i_0_in1[2]
+ cb_6_4/io_i_0_in1[3] cb_6_4/io_i_0_in1[4] cb_6_4/io_i_0_in1[5] cb_6_4/io_i_0_in1[6]
+ cb_6_4/io_i_0_in1[7] cb_6_4/io_i_1_ci cb_6_4/io_i_1_in1[0] cb_6_4/io_i_1_in1[1]
+ cb_6_4/io_i_1_in1[2] cb_6_4/io_i_1_in1[3] cb_6_4/io_i_1_in1[4] cb_6_4/io_i_1_in1[5]
+ cb_6_4/io_i_1_in1[6] cb_6_4/io_i_1_in1[7] cb_6_4/io_i_2_ci cb_6_4/io_i_2_in1[0]
+ cb_6_4/io_i_2_in1[1] cb_6_4/io_i_2_in1[2] cb_6_4/io_i_2_in1[3] cb_6_4/io_i_2_in1[4]
+ cb_6_4/io_i_2_in1[5] cb_6_4/io_i_2_in1[6] cb_6_4/io_i_2_in1[7] cb_6_4/io_i_3_ci
+ cb_6_4/io_i_3_in1[0] cb_6_4/io_i_3_in1[1] cb_6_4/io_i_3_in1[2] cb_6_4/io_i_3_in1[3]
+ cb_6_4/io_i_3_in1[4] cb_6_4/io_i_3_in1[5] cb_6_4/io_i_3_in1[6] cb_6_4/io_i_3_in1[7]
+ cb_6_4/io_i_4_ci cb_6_4/io_i_4_in1[0] cb_6_4/io_i_4_in1[1] cb_6_4/io_i_4_in1[2]
+ cb_6_4/io_i_4_in1[3] cb_6_4/io_i_4_in1[4] cb_6_4/io_i_4_in1[5] cb_6_4/io_i_4_in1[6]
+ cb_6_4/io_i_4_in1[7] cb_6_4/io_i_5_ci cb_6_4/io_i_5_in1[0] cb_6_4/io_i_5_in1[1]
+ cb_6_4/io_i_5_in1[2] cb_6_4/io_i_5_in1[3] cb_6_4/io_i_5_in1[4] cb_6_4/io_i_5_in1[5]
+ cb_6_4/io_i_5_in1[6] cb_6_4/io_i_5_in1[7] cb_6_4/io_i_6_ci cb_6_4/io_i_6_in1[0]
+ cb_6_4/io_i_6_in1[1] cb_6_4/io_i_6_in1[2] cb_6_4/io_i_6_in1[3] cb_6_4/io_i_6_in1[4]
+ cb_6_4/io_i_6_in1[5] cb_6_4/io_i_6_in1[6] cb_6_4/io_i_6_in1[7] cb_6_4/io_i_7_ci
+ cb_6_4/io_i_7_in1[0] cb_6_4/io_i_7_in1[1] cb_6_4/io_i_7_in1[2] cb_6_4/io_i_7_in1[3]
+ cb_6_4/io_i_7_in1[4] cb_6_4/io_i_7_in1[5] cb_6_4/io_i_7_in1[6] cb_6_4/io_i_7_in1[7]
+ cb_6_5/io_i_0_ci cb_6_5/io_i_0_in1[0] cb_6_5/io_i_0_in1[1] cb_6_5/io_i_0_in1[2]
+ cb_6_5/io_i_0_in1[3] cb_6_5/io_i_0_in1[4] cb_6_5/io_i_0_in1[5] cb_6_5/io_i_0_in1[6]
+ cb_6_5/io_i_0_in1[7] cb_6_5/io_i_1_ci cb_6_5/io_i_1_in1[0] cb_6_5/io_i_1_in1[1]
+ cb_6_5/io_i_1_in1[2] cb_6_5/io_i_1_in1[3] cb_6_5/io_i_1_in1[4] cb_6_5/io_i_1_in1[5]
+ cb_6_5/io_i_1_in1[6] cb_6_5/io_i_1_in1[7] cb_6_5/io_i_2_ci cb_6_5/io_i_2_in1[0]
+ cb_6_5/io_i_2_in1[1] cb_6_5/io_i_2_in1[2] cb_6_5/io_i_2_in1[3] cb_6_5/io_i_2_in1[4]
+ cb_6_5/io_i_2_in1[5] cb_6_5/io_i_2_in1[6] cb_6_5/io_i_2_in1[7] cb_6_5/io_i_3_ci
+ cb_6_5/io_i_3_in1[0] cb_6_5/io_i_3_in1[1] cb_6_5/io_i_3_in1[2] cb_6_5/io_i_3_in1[3]
+ cb_6_5/io_i_3_in1[4] cb_6_5/io_i_3_in1[5] cb_6_5/io_i_3_in1[6] cb_6_5/io_i_3_in1[7]
+ cb_6_5/io_i_4_ci cb_6_5/io_i_4_in1[0] cb_6_5/io_i_4_in1[1] cb_6_5/io_i_4_in1[2]
+ cb_6_5/io_i_4_in1[3] cb_6_5/io_i_4_in1[4] cb_6_5/io_i_4_in1[5] cb_6_5/io_i_4_in1[6]
+ cb_6_5/io_i_4_in1[7] cb_6_5/io_i_5_ci cb_6_5/io_i_5_in1[0] cb_6_5/io_i_5_in1[1]
+ cb_6_5/io_i_5_in1[2] cb_6_5/io_i_5_in1[3] cb_6_5/io_i_5_in1[4] cb_6_5/io_i_5_in1[5]
+ cb_6_5/io_i_5_in1[6] cb_6_5/io_i_5_in1[7] cb_6_5/io_i_6_ci cb_6_5/io_i_6_in1[0]
+ cb_6_5/io_i_6_in1[1] cb_6_5/io_i_6_in1[2] cb_6_5/io_i_6_in1[3] cb_6_5/io_i_6_in1[4]
+ cb_6_5/io_i_6_in1[5] cb_6_5/io_i_6_in1[6] cb_6_5/io_i_6_in1[7] cb_6_5/io_i_7_ci
+ cb_6_5/io_i_7_in1[0] cb_6_5/io_i_7_in1[1] cb_6_5/io_i_7_in1[2] cb_6_5/io_i_7_in1[3]
+ cb_6_5/io_i_7_in1[4] cb_6_5/io_i_7_in1[5] cb_6_5/io_i_7_in1[6] cb_6_5/io_i_7_in1[7]
+ cb_6_4/io_vci cb_6_5/io_vci cb_6_4/io_vi cb_6_9/io_we_i cb_6_4/io_wo[0] cb_6_4/io_wo[10]
+ cb_6_4/io_wo[11] cb_6_4/io_wo[12] cb_6_4/io_wo[13] cb_6_4/io_wo[14] cb_6_4/io_wo[15]
+ cb_6_4/io_wo[16] cb_6_4/io_wo[17] cb_6_4/io_wo[18] cb_6_4/io_wo[19] cb_6_4/io_wo[1]
+ cb_6_4/io_wo[20] cb_6_4/io_wo[21] cb_6_4/io_wo[22] cb_6_4/io_wo[23] cb_6_4/io_wo[24]
+ cb_6_4/io_wo[25] cb_6_4/io_wo[26] cb_6_4/io_wo[27] cb_6_4/io_wo[28] cb_6_4/io_wo[29]
+ cb_6_4/io_wo[2] cb_6_4/io_wo[30] cb_6_4/io_wo[31] cb_6_4/io_wo[32] cb_6_4/io_wo[33]
+ cb_6_4/io_wo[34] cb_6_4/io_wo[35] cb_6_4/io_wo[36] cb_6_4/io_wo[37] cb_6_4/io_wo[38]
+ cb_6_4/io_wo[39] cb_6_4/io_wo[3] cb_6_4/io_wo[40] cb_6_4/io_wo[41] cb_6_4/io_wo[42]
+ cb_6_4/io_wo[43] cb_6_4/io_wo[44] cb_6_4/io_wo[45] cb_6_4/io_wo[46] cb_6_4/io_wo[47]
+ cb_6_4/io_wo[48] cb_6_4/io_wo[49] cb_6_4/io_wo[4] cb_6_4/io_wo[50] cb_6_4/io_wo[51]
+ cb_6_4/io_wo[52] cb_6_4/io_wo[53] cb_6_4/io_wo[54] cb_6_4/io_wo[55] cb_6_4/io_wo[56]
+ cb_6_4/io_wo[57] cb_6_4/io_wo[58] cb_6_4/io_wo[59] cb_6_4/io_wo[5] cb_6_4/io_wo[60]
+ cb_6_4/io_wo[61] cb_6_4/io_wo[62] cb_6_4/io_wo[63] cb_6_4/io_wo[6] cb_6_4/io_wo[7]
+ cb_6_4/io_wo[8] cb_6_4/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_4_1 cb_4_9/io_adr_i[0] cb_4_9/io_adr_i[1] cb_4_1/io_cs_i cb_4_9/io_dat_i[0] cb_4_9/io_dat_i[10]
+ cb_4_9/io_dat_i[11] cb_4_9/io_dat_i[12] cb_4_9/io_dat_i[13] cb_4_9/io_dat_i[14]
+ cb_4_9/io_dat_i[15] cb_4_9/io_dat_i[1] cb_4_9/io_dat_i[2] cb_4_9/io_dat_i[3] cb_4_9/io_dat_i[4]
+ cb_4_9/io_dat_i[5] cb_4_9/io_dat_i[6] cb_4_9/io_dat_i[7] cb_4_9/io_dat_i[8] cb_4_9/io_dat_i[9]
+ cb_4_1/io_dat_o[0] cb_4_1/io_dat_o[10] cb_4_1/io_dat_o[11] cb_4_1/io_dat_o[12] cb_4_1/io_dat_o[13]
+ cb_4_1/io_dat_o[14] cb_4_1/io_dat_o[15] cb_4_1/io_dat_o[1] cb_4_1/io_dat_o[2] cb_4_1/io_dat_o[3]
+ cb_4_1/io_dat_o[4] cb_4_1/io_dat_o[5] cb_4_1/io_dat_o[6] cb_4_1/io_dat_o[7] cb_4_1/io_dat_o[8]
+ cb_4_1/io_dat_o[9] cb_4_2/io_wo[0] cb_4_2/io_wo[10] cb_4_2/io_wo[11] cb_4_2/io_wo[12]
+ cb_4_2/io_wo[13] cb_4_2/io_wo[14] cb_4_2/io_wo[15] cb_4_2/io_wo[16] cb_4_2/io_wo[17]
+ cb_4_2/io_wo[18] cb_4_2/io_wo[19] cb_4_2/io_wo[1] cb_4_2/io_wo[20] cb_4_2/io_wo[21]
+ cb_4_2/io_wo[22] cb_4_2/io_wo[23] cb_4_2/io_wo[24] cb_4_2/io_wo[25] cb_4_2/io_wo[26]
+ cb_4_2/io_wo[27] cb_4_2/io_wo[28] cb_4_2/io_wo[29] cb_4_2/io_wo[2] cb_4_2/io_wo[30]
+ cb_4_2/io_wo[31] cb_4_2/io_wo[32] cb_4_2/io_wo[33] cb_4_2/io_wo[34] cb_4_2/io_wo[35]
+ cb_4_2/io_wo[36] cb_4_2/io_wo[37] cb_4_2/io_wo[38] cb_4_2/io_wo[39] cb_4_2/io_wo[3]
+ cb_4_2/io_wo[40] cb_4_2/io_wo[41] cb_4_2/io_wo[42] cb_4_2/io_wo[43] cb_4_2/io_wo[44]
+ cb_4_2/io_wo[45] cb_4_2/io_wo[46] cb_4_2/io_wo[47] cb_4_2/io_wo[48] cb_4_2/io_wo[49]
+ cb_4_2/io_wo[4] cb_4_2/io_wo[50] cb_4_2/io_wo[51] cb_4_2/io_wo[52] cb_4_2/io_wo[53]
+ cb_4_2/io_wo[54] cb_4_2/io_wo[55] cb_4_2/io_wo[56] cb_4_2/io_wo[57] cb_4_2/io_wo[58]
+ cb_4_2/io_wo[59] cb_4_2/io_wo[5] cb_4_2/io_wo[60] cb_4_2/io_wo[61] cb_4_2/io_wo[62]
+ cb_4_2/io_wo[63] cb_4_2/io_wo[6] cb_4_2/io_wo[7] cb_4_2/io_wo[8] cb_4_2/io_wo[9]
+ cb_4_1/io_i_0_ci cb_4_1/io_i_0_in1[0] cb_4_1/io_i_0_in1[1] cb_4_1/io_i_0_in1[2]
+ cb_4_1/io_i_0_in1[3] cb_4_1/io_i_0_in1[4] cb_4_1/io_i_0_in1[5] cb_4_1/io_i_0_in1[6]
+ cb_4_1/io_i_0_in1[7] cb_4_1/io_i_1_ci cb_4_1/io_i_1_in1[0] cb_4_1/io_i_1_in1[1]
+ cb_4_1/io_i_1_in1[2] cb_4_1/io_i_1_in1[3] cb_4_1/io_i_1_in1[4] cb_4_1/io_i_1_in1[5]
+ cb_4_1/io_i_1_in1[6] cb_4_1/io_i_1_in1[7] cb_4_1/io_i_2_ci cb_4_1/io_i_2_in1[0]
+ cb_4_1/io_i_2_in1[1] cb_4_1/io_i_2_in1[2] cb_4_1/io_i_2_in1[3] cb_4_1/io_i_2_in1[4]
+ cb_4_1/io_i_2_in1[5] cb_4_1/io_i_2_in1[6] cb_4_1/io_i_2_in1[7] cb_4_1/io_i_3_ci
+ cb_4_1/io_i_3_in1[0] cb_4_1/io_i_3_in1[1] cb_4_1/io_i_3_in1[2] cb_4_1/io_i_3_in1[3]
+ cb_4_1/io_i_3_in1[4] cb_4_1/io_i_3_in1[5] cb_4_1/io_i_3_in1[6] cb_4_1/io_i_3_in1[7]
+ cb_4_1/io_i_4_ci cb_4_1/io_i_4_in1[0] cb_4_1/io_i_4_in1[1] cb_4_1/io_i_4_in1[2]
+ cb_4_1/io_i_4_in1[3] cb_4_1/io_i_4_in1[4] cb_4_1/io_i_4_in1[5] cb_4_1/io_i_4_in1[6]
+ cb_4_1/io_i_4_in1[7] cb_4_1/io_i_5_ci cb_4_1/io_i_5_in1[0] cb_4_1/io_i_5_in1[1]
+ cb_4_1/io_i_5_in1[2] cb_4_1/io_i_5_in1[3] cb_4_1/io_i_5_in1[4] cb_4_1/io_i_5_in1[5]
+ cb_4_1/io_i_5_in1[6] cb_4_1/io_i_5_in1[7] cb_4_1/io_i_6_ci cb_4_1/io_i_6_in1[0]
+ cb_4_1/io_i_6_in1[1] cb_4_1/io_i_6_in1[2] cb_4_1/io_i_6_in1[3] cb_4_1/io_i_6_in1[4]
+ cb_4_1/io_i_6_in1[5] cb_4_1/io_i_6_in1[6] cb_4_1/io_i_6_in1[7] cb_4_1/io_i_7_ci
+ cb_4_1/io_i_7_in1[0] cb_4_1/io_i_7_in1[1] cb_4_1/io_i_7_in1[2] cb_4_1/io_i_7_in1[3]
+ cb_4_1/io_i_7_in1[4] cb_4_1/io_i_7_in1[5] cb_4_1/io_i_7_in1[6] cb_4_1/io_i_7_in1[7]
+ cb_4_2/io_i_0_ci cb_4_2/io_i_0_in1[0] cb_4_2/io_i_0_in1[1] cb_4_2/io_i_0_in1[2]
+ cb_4_2/io_i_0_in1[3] cb_4_2/io_i_0_in1[4] cb_4_2/io_i_0_in1[5] cb_4_2/io_i_0_in1[6]
+ cb_4_2/io_i_0_in1[7] cb_4_2/io_i_1_ci cb_4_2/io_i_1_in1[0] cb_4_2/io_i_1_in1[1]
+ cb_4_2/io_i_1_in1[2] cb_4_2/io_i_1_in1[3] cb_4_2/io_i_1_in1[4] cb_4_2/io_i_1_in1[5]
+ cb_4_2/io_i_1_in1[6] cb_4_2/io_i_1_in1[7] cb_4_2/io_i_2_ci cb_4_2/io_i_2_in1[0]
+ cb_4_2/io_i_2_in1[1] cb_4_2/io_i_2_in1[2] cb_4_2/io_i_2_in1[3] cb_4_2/io_i_2_in1[4]
+ cb_4_2/io_i_2_in1[5] cb_4_2/io_i_2_in1[6] cb_4_2/io_i_2_in1[7] cb_4_2/io_i_3_ci
+ cb_4_2/io_i_3_in1[0] cb_4_2/io_i_3_in1[1] cb_4_2/io_i_3_in1[2] cb_4_2/io_i_3_in1[3]
+ cb_4_2/io_i_3_in1[4] cb_4_2/io_i_3_in1[5] cb_4_2/io_i_3_in1[6] cb_4_2/io_i_3_in1[7]
+ cb_4_2/io_i_4_ci cb_4_2/io_i_4_in1[0] cb_4_2/io_i_4_in1[1] cb_4_2/io_i_4_in1[2]
+ cb_4_2/io_i_4_in1[3] cb_4_2/io_i_4_in1[4] cb_4_2/io_i_4_in1[5] cb_4_2/io_i_4_in1[6]
+ cb_4_2/io_i_4_in1[7] cb_4_2/io_i_5_ci cb_4_2/io_i_5_in1[0] cb_4_2/io_i_5_in1[1]
+ cb_4_2/io_i_5_in1[2] cb_4_2/io_i_5_in1[3] cb_4_2/io_i_5_in1[4] cb_4_2/io_i_5_in1[5]
+ cb_4_2/io_i_5_in1[6] cb_4_2/io_i_5_in1[7] cb_4_2/io_i_6_ci cb_4_2/io_i_6_in1[0]
+ cb_4_2/io_i_6_in1[1] cb_4_2/io_i_6_in1[2] cb_4_2/io_i_6_in1[3] cb_4_2/io_i_6_in1[4]
+ cb_4_2/io_i_6_in1[5] cb_4_2/io_i_6_in1[6] cb_4_2/io_i_6_in1[7] cb_4_2/io_i_7_ci
+ cb_4_2/io_i_7_in1[0] cb_4_2/io_i_7_in1[1] cb_4_2/io_i_7_in1[2] cb_4_2/io_i_7_in1[3]
+ cb_4_2/io_i_7_in1[4] cb_4_2/io_i_7_in1[5] cb_4_2/io_i_7_in1[6] cb_4_2/io_i_7_in1[7]
+ cb_4_1/io_vci cb_4_2/io_vci cb_4_1/io_vi cb_4_9/io_we_i cb_4_1/io_wo[0] cb_4_1/io_wo[10]
+ cb_4_1/io_wo[11] cb_4_1/io_wo[12] cb_4_1/io_wo[13] cb_4_1/io_wo[14] cb_4_1/io_wo[15]
+ cb_4_1/io_wo[16] cb_4_1/io_wo[17] cb_4_1/io_wo[18] cb_4_1/io_wo[19] cb_4_1/io_wo[1]
+ cb_4_1/io_wo[20] cb_4_1/io_wo[21] cb_4_1/io_wo[22] cb_4_1/io_wo[23] cb_4_1/io_wo[24]
+ cb_4_1/io_wo[25] cb_4_1/io_wo[26] cb_4_1/io_wo[27] cb_4_1/io_wo[28] cb_4_1/io_wo[29]
+ cb_4_1/io_wo[2] cb_4_1/io_wo[30] cb_4_1/io_wo[31] cb_4_1/io_wo[32] cb_4_1/io_wo[33]
+ cb_4_1/io_wo[34] cb_4_1/io_wo[35] cb_4_1/io_wo[36] cb_4_1/io_wo[37] cb_4_1/io_wo[38]
+ cb_4_1/io_wo[39] cb_4_1/io_wo[3] cb_4_1/io_wo[40] cb_4_1/io_wo[41] cb_4_1/io_wo[42]
+ cb_4_1/io_wo[43] cb_4_1/io_wo[44] cb_4_1/io_wo[45] cb_4_1/io_wo[46] cb_4_1/io_wo[47]
+ cb_4_1/io_wo[48] cb_4_1/io_wo[49] cb_4_1/io_wo[4] cb_4_1/io_wo[50] cb_4_1/io_wo[51]
+ cb_4_1/io_wo[52] cb_4_1/io_wo[53] cb_4_1/io_wo[54] cb_4_1/io_wo[55] cb_4_1/io_wo[56]
+ cb_4_1/io_wo[57] cb_4_1/io_wo[58] cb_4_1/io_wo[59] cb_4_1/io_wo[5] cb_4_1/io_wo[60]
+ cb_4_1/io_wo[61] cb_4_1/io_wo[62] cb_4_1/io_wo[63] cb_4_1/io_wo[6] cb_4_1/io_wo[7]
+ cb_4_1/io_wo[8] cb_4_1/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_6_5 cb_6_9/io_adr_i[0] cb_6_9/io_adr_i[1] cb_6_5/io_cs_i cb_6_9/io_dat_i[0] cb_6_9/io_dat_i[10]
+ cb_6_9/io_dat_i[11] cb_6_9/io_dat_i[12] cb_6_9/io_dat_i[13] cb_6_9/io_dat_i[14]
+ cb_6_9/io_dat_i[15] cb_6_9/io_dat_i[1] cb_6_9/io_dat_i[2] cb_6_9/io_dat_i[3] cb_6_9/io_dat_i[4]
+ cb_6_9/io_dat_i[5] cb_6_9/io_dat_i[6] cb_6_9/io_dat_i[7] cb_6_9/io_dat_i[8] cb_6_9/io_dat_i[9]
+ cb_6_5/io_dat_o[0] cb_6_5/io_dat_o[10] cb_6_5/io_dat_o[11] cb_6_5/io_dat_o[12] cb_6_5/io_dat_o[13]
+ cb_6_5/io_dat_o[14] cb_6_5/io_dat_o[15] cb_6_5/io_dat_o[1] cb_6_5/io_dat_o[2] cb_6_5/io_dat_o[3]
+ cb_6_5/io_dat_o[4] cb_6_5/io_dat_o[5] cb_6_5/io_dat_o[6] cb_6_5/io_dat_o[7] cb_6_5/io_dat_o[8]
+ cb_6_5/io_dat_o[9] cb_6_6/io_wo[0] cb_6_6/io_wo[10] cb_6_6/io_wo[11] cb_6_6/io_wo[12]
+ cb_6_6/io_wo[13] cb_6_6/io_wo[14] cb_6_6/io_wo[15] cb_6_6/io_wo[16] cb_6_6/io_wo[17]
+ cb_6_6/io_wo[18] cb_6_6/io_wo[19] cb_6_6/io_wo[1] cb_6_6/io_wo[20] cb_6_6/io_wo[21]
+ cb_6_6/io_wo[22] cb_6_6/io_wo[23] cb_6_6/io_wo[24] cb_6_6/io_wo[25] cb_6_6/io_wo[26]
+ cb_6_6/io_wo[27] cb_6_6/io_wo[28] cb_6_6/io_wo[29] cb_6_6/io_wo[2] cb_6_6/io_wo[30]
+ cb_6_6/io_wo[31] cb_6_6/io_wo[32] cb_6_6/io_wo[33] cb_6_6/io_wo[34] cb_6_6/io_wo[35]
+ cb_6_6/io_wo[36] cb_6_6/io_wo[37] cb_6_6/io_wo[38] cb_6_6/io_wo[39] cb_6_6/io_wo[3]
+ cb_6_6/io_wo[40] cb_6_6/io_wo[41] cb_6_6/io_wo[42] cb_6_6/io_wo[43] cb_6_6/io_wo[44]
+ cb_6_6/io_wo[45] cb_6_6/io_wo[46] cb_6_6/io_wo[47] cb_6_6/io_wo[48] cb_6_6/io_wo[49]
+ cb_6_6/io_wo[4] cb_6_6/io_wo[50] cb_6_6/io_wo[51] cb_6_6/io_wo[52] cb_6_6/io_wo[53]
+ cb_6_6/io_wo[54] cb_6_6/io_wo[55] cb_6_6/io_wo[56] cb_6_6/io_wo[57] cb_6_6/io_wo[58]
+ cb_6_6/io_wo[59] cb_6_6/io_wo[5] cb_6_6/io_wo[60] cb_6_6/io_wo[61] cb_6_6/io_wo[62]
+ cb_6_6/io_wo[63] cb_6_6/io_wo[6] cb_6_6/io_wo[7] cb_6_6/io_wo[8] cb_6_6/io_wo[9]
+ cb_6_5/io_i_0_ci cb_6_5/io_i_0_in1[0] cb_6_5/io_i_0_in1[1] cb_6_5/io_i_0_in1[2]
+ cb_6_5/io_i_0_in1[3] cb_6_5/io_i_0_in1[4] cb_6_5/io_i_0_in1[5] cb_6_5/io_i_0_in1[6]
+ cb_6_5/io_i_0_in1[7] cb_6_5/io_i_1_ci cb_6_5/io_i_1_in1[0] cb_6_5/io_i_1_in1[1]
+ cb_6_5/io_i_1_in1[2] cb_6_5/io_i_1_in1[3] cb_6_5/io_i_1_in1[4] cb_6_5/io_i_1_in1[5]
+ cb_6_5/io_i_1_in1[6] cb_6_5/io_i_1_in1[7] cb_6_5/io_i_2_ci cb_6_5/io_i_2_in1[0]
+ cb_6_5/io_i_2_in1[1] cb_6_5/io_i_2_in1[2] cb_6_5/io_i_2_in1[3] cb_6_5/io_i_2_in1[4]
+ cb_6_5/io_i_2_in1[5] cb_6_5/io_i_2_in1[6] cb_6_5/io_i_2_in1[7] cb_6_5/io_i_3_ci
+ cb_6_5/io_i_3_in1[0] cb_6_5/io_i_3_in1[1] cb_6_5/io_i_3_in1[2] cb_6_5/io_i_3_in1[3]
+ cb_6_5/io_i_3_in1[4] cb_6_5/io_i_3_in1[5] cb_6_5/io_i_3_in1[6] cb_6_5/io_i_3_in1[7]
+ cb_6_5/io_i_4_ci cb_6_5/io_i_4_in1[0] cb_6_5/io_i_4_in1[1] cb_6_5/io_i_4_in1[2]
+ cb_6_5/io_i_4_in1[3] cb_6_5/io_i_4_in1[4] cb_6_5/io_i_4_in1[5] cb_6_5/io_i_4_in1[6]
+ cb_6_5/io_i_4_in1[7] cb_6_5/io_i_5_ci cb_6_5/io_i_5_in1[0] cb_6_5/io_i_5_in1[1]
+ cb_6_5/io_i_5_in1[2] cb_6_5/io_i_5_in1[3] cb_6_5/io_i_5_in1[4] cb_6_5/io_i_5_in1[5]
+ cb_6_5/io_i_5_in1[6] cb_6_5/io_i_5_in1[7] cb_6_5/io_i_6_ci cb_6_5/io_i_6_in1[0]
+ cb_6_5/io_i_6_in1[1] cb_6_5/io_i_6_in1[2] cb_6_5/io_i_6_in1[3] cb_6_5/io_i_6_in1[4]
+ cb_6_5/io_i_6_in1[5] cb_6_5/io_i_6_in1[6] cb_6_5/io_i_6_in1[7] cb_6_5/io_i_7_ci
+ cb_6_5/io_i_7_in1[0] cb_6_5/io_i_7_in1[1] cb_6_5/io_i_7_in1[2] cb_6_5/io_i_7_in1[3]
+ cb_6_5/io_i_7_in1[4] cb_6_5/io_i_7_in1[5] cb_6_5/io_i_7_in1[6] cb_6_5/io_i_7_in1[7]
+ cb_6_6/io_i_0_ci cb_6_6/io_i_0_in1[0] cb_6_6/io_i_0_in1[1] cb_6_6/io_i_0_in1[2]
+ cb_6_6/io_i_0_in1[3] cb_6_6/io_i_0_in1[4] cb_6_6/io_i_0_in1[5] cb_6_6/io_i_0_in1[6]
+ cb_6_6/io_i_0_in1[7] cb_6_6/io_i_1_ci cb_6_6/io_i_1_in1[0] cb_6_6/io_i_1_in1[1]
+ cb_6_6/io_i_1_in1[2] cb_6_6/io_i_1_in1[3] cb_6_6/io_i_1_in1[4] cb_6_6/io_i_1_in1[5]
+ cb_6_6/io_i_1_in1[6] cb_6_6/io_i_1_in1[7] cb_6_6/io_i_2_ci cb_6_6/io_i_2_in1[0]
+ cb_6_6/io_i_2_in1[1] cb_6_6/io_i_2_in1[2] cb_6_6/io_i_2_in1[3] cb_6_6/io_i_2_in1[4]
+ cb_6_6/io_i_2_in1[5] cb_6_6/io_i_2_in1[6] cb_6_6/io_i_2_in1[7] cb_6_6/io_i_3_ci
+ cb_6_6/io_i_3_in1[0] cb_6_6/io_i_3_in1[1] cb_6_6/io_i_3_in1[2] cb_6_6/io_i_3_in1[3]
+ cb_6_6/io_i_3_in1[4] cb_6_6/io_i_3_in1[5] cb_6_6/io_i_3_in1[6] cb_6_6/io_i_3_in1[7]
+ cb_6_6/io_i_4_ci cb_6_6/io_i_4_in1[0] cb_6_6/io_i_4_in1[1] cb_6_6/io_i_4_in1[2]
+ cb_6_6/io_i_4_in1[3] cb_6_6/io_i_4_in1[4] cb_6_6/io_i_4_in1[5] cb_6_6/io_i_4_in1[6]
+ cb_6_6/io_i_4_in1[7] cb_6_6/io_i_5_ci cb_6_6/io_i_5_in1[0] cb_6_6/io_i_5_in1[1]
+ cb_6_6/io_i_5_in1[2] cb_6_6/io_i_5_in1[3] cb_6_6/io_i_5_in1[4] cb_6_6/io_i_5_in1[5]
+ cb_6_6/io_i_5_in1[6] cb_6_6/io_i_5_in1[7] cb_6_6/io_i_6_ci cb_6_6/io_i_6_in1[0]
+ cb_6_6/io_i_6_in1[1] cb_6_6/io_i_6_in1[2] cb_6_6/io_i_6_in1[3] cb_6_6/io_i_6_in1[4]
+ cb_6_6/io_i_6_in1[5] cb_6_6/io_i_6_in1[6] cb_6_6/io_i_6_in1[7] cb_6_6/io_i_7_ci
+ cb_6_6/io_i_7_in1[0] cb_6_6/io_i_7_in1[1] cb_6_6/io_i_7_in1[2] cb_6_6/io_i_7_in1[3]
+ cb_6_6/io_i_7_in1[4] cb_6_6/io_i_7_in1[5] cb_6_6/io_i_7_in1[6] cb_6_6/io_i_7_in1[7]
+ cb_6_5/io_vci cb_6_6/io_vci cb_6_5/io_vi cb_6_9/io_we_i cb_6_5/io_wo[0] cb_6_5/io_wo[10]
+ cb_6_5/io_wo[11] cb_6_5/io_wo[12] cb_6_5/io_wo[13] cb_6_5/io_wo[14] cb_6_5/io_wo[15]
+ cb_6_5/io_wo[16] cb_6_5/io_wo[17] cb_6_5/io_wo[18] cb_6_5/io_wo[19] cb_6_5/io_wo[1]
+ cb_6_5/io_wo[20] cb_6_5/io_wo[21] cb_6_5/io_wo[22] cb_6_5/io_wo[23] cb_6_5/io_wo[24]
+ cb_6_5/io_wo[25] cb_6_5/io_wo[26] cb_6_5/io_wo[27] cb_6_5/io_wo[28] cb_6_5/io_wo[29]
+ cb_6_5/io_wo[2] cb_6_5/io_wo[30] cb_6_5/io_wo[31] cb_6_5/io_wo[32] cb_6_5/io_wo[33]
+ cb_6_5/io_wo[34] cb_6_5/io_wo[35] cb_6_5/io_wo[36] cb_6_5/io_wo[37] cb_6_5/io_wo[38]
+ cb_6_5/io_wo[39] cb_6_5/io_wo[3] cb_6_5/io_wo[40] cb_6_5/io_wo[41] cb_6_5/io_wo[42]
+ cb_6_5/io_wo[43] cb_6_5/io_wo[44] cb_6_5/io_wo[45] cb_6_5/io_wo[46] cb_6_5/io_wo[47]
+ cb_6_5/io_wo[48] cb_6_5/io_wo[49] cb_6_5/io_wo[4] cb_6_5/io_wo[50] cb_6_5/io_wo[51]
+ cb_6_5/io_wo[52] cb_6_5/io_wo[53] cb_6_5/io_wo[54] cb_6_5/io_wo[55] cb_6_5/io_wo[56]
+ cb_6_5/io_wo[57] cb_6_5/io_wo[58] cb_6_5/io_wo[59] cb_6_5/io_wo[5] cb_6_5/io_wo[60]
+ cb_6_5/io_wo[61] cb_6_5/io_wo[62] cb_6_5/io_wo[63] cb_6_5/io_wo[6] cb_6_5/io_wo[7]
+ cb_6_5/io_wo[8] cb_6_5/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_4_2 cb_4_9/io_adr_i[0] cb_4_9/io_adr_i[1] cb_4_2/io_cs_i cb_4_9/io_dat_i[0] cb_4_9/io_dat_i[10]
+ cb_4_9/io_dat_i[11] cb_4_9/io_dat_i[12] cb_4_9/io_dat_i[13] cb_4_9/io_dat_i[14]
+ cb_4_9/io_dat_i[15] cb_4_9/io_dat_i[1] cb_4_9/io_dat_i[2] cb_4_9/io_dat_i[3] cb_4_9/io_dat_i[4]
+ cb_4_9/io_dat_i[5] cb_4_9/io_dat_i[6] cb_4_9/io_dat_i[7] cb_4_9/io_dat_i[8] cb_4_9/io_dat_i[9]
+ cb_4_2/io_dat_o[0] cb_4_2/io_dat_o[10] cb_4_2/io_dat_o[11] cb_4_2/io_dat_o[12] cb_4_2/io_dat_o[13]
+ cb_4_2/io_dat_o[14] cb_4_2/io_dat_o[15] cb_4_2/io_dat_o[1] cb_4_2/io_dat_o[2] cb_4_2/io_dat_o[3]
+ cb_4_2/io_dat_o[4] cb_4_2/io_dat_o[5] cb_4_2/io_dat_o[6] cb_4_2/io_dat_o[7] cb_4_2/io_dat_o[8]
+ cb_4_2/io_dat_o[9] cb_4_3/io_wo[0] cb_4_3/io_wo[10] cb_4_3/io_wo[11] cb_4_3/io_wo[12]
+ cb_4_3/io_wo[13] cb_4_3/io_wo[14] cb_4_3/io_wo[15] cb_4_3/io_wo[16] cb_4_3/io_wo[17]
+ cb_4_3/io_wo[18] cb_4_3/io_wo[19] cb_4_3/io_wo[1] cb_4_3/io_wo[20] cb_4_3/io_wo[21]
+ cb_4_3/io_wo[22] cb_4_3/io_wo[23] cb_4_3/io_wo[24] cb_4_3/io_wo[25] cb_4_3/io_wo[26]
+ cb_4_3/io_wo[27] cb_4_3/io_wo[28] cb_4_3/io_wo[29] cb_4_3/io_wo[2] cb_4_3/io_wo[30]
+ cb_4_3/io_wo[31] cb_4_3/io_wo[32] cb_4_3/io_wo[33] cb_4_3/io_wo[34] cb_4_3/io_wo[35]
+ cb_4_3/io_wo[36] cb_4_3/io_wo[37] cb_4_3/io_wo[38] cb_4_3/io_wo[39] cb_4_3/io_wo[3]
+ cb_4_3/io_wo[40] cb_4_3/io_wo[41] cb_4_3/io_wo[42] cb_4_3/io_wo[43] cb_4_3/io_wo[44]
+ cb_4_3/io_wo[45] cb_4_3/io_wo[46] cb_4_3/io_wo[47] cb_4_3/io_wo[48] cb_4_3/io_wo[49]
+ cb_4_3/io_wo[4] cb_4_3/io_wo[50] cb_4_3/io_wo[51] cb_4_3/io_wo[52] cb_4_3/io_wo[53]
+ cb_4_3/io_wo[54] cb_4_3/io_wo[55] cb_4_3/io_wo[56] cb_4_3/io_wo[57] cb_4_3/io_wo[58]
+ cb_4_3/io_wo[59] cb_4_3/io_wo[5] cb_4_3/io_wo[60] cb_4_3/io_wo[61] cb_4_3/io_wo[62]
+ cb_4_3/io_wo[63] cb_4_3/io_wo[6] cb_4_3/io_wo[7] cb_4_3/io_wo[8] cb_4_3/io_wo[9]
+ cb_4_2/io_i_0_ci cb_4_2/io_i_0_in1[0] cb_4_2/io_i_0_in1[1] cb_4_2/io_i_0_in1[2]
+ cb_4_2/io_i_0_in1[3] cb_4_2/io_i_0_in1[4] cb_4_2/io_i_0_in1[5] cb_4_2/io_i_0_in1[6]
+ cb_4_2/io_i_0_in1[7] cb_4_2/io_i_1_ci cb_4_2/io_i_1_in1[0] cb_4_2/io_i_1_in1[1]
+ cb_4_2/io_i_1_in1[2] cb_4_2/io_i_1_in1[3] cb_4_2/io_i_1_in1[4] cb_4_2/io_i_1_in1[5]
+ cb_4_2/io_i_1_in1[6] cb_4_2/io_i_1_in1[7] cb_4_2/io_i_2_ci cb_4_2/io_i_2_in1[0]
+ cb_4_2/io_i_2_in1[1] cb_4_2/io_i_2_in1[2] cb_4_2/io_i_2_in1[3] cb_4_2/io_i_2_in1[4]
+ cb_4_2/io_i_2_in1[5] cb_4_2/io_i_2_in1[6] cb_4_2/io_i_2_in1[7] cb_4_2/io_i_3_ci
+ cb_4_2/io_i_3_in1[0] cb_4_2/io_i_3_in1[1] cb_4_2/io_i_3_in1[2] cb_4_2/io_i_3_in1[3]
+ cb_4_2/io_i_3_in1[4] cb_4_2/io_i_3_in1[5] cb_4_2/io_i_3_in1[6] cb_4_2/io_i_3_in1[7]
+ cb_4_2/io_i_4_ci cb_4_2/io_i_4_in1[0] cb_4_2/io_i_4_in1[1] cb_4_2/io_i_4_in1[2]
+ cb_4_2/io_i_4_in1[3] cb_4_2/io_i_4_in1[4] cb_4_2/io_i_4_in1[5] cb_4_2/io_i_4_in1[6]
+ cb_4_2/io_i_4_in1[7] cb_4_2/io_i_5_ci cb_4_2/io_i_5_in1[0] cb_4_2/io_i_5_in1[1]
+ cb_4_2/io_i_5_in1[2] cb_4_2/io_i_5_in1[3] cb_4_2/io_i_5_in1[4] cb_4_2/io_i_5_in1[5]
+ cb_4_2/io_i_5_in1[6] cb_4_2/io_i_5_in1[7] cb_4_2/io_i_6_ci cb_4_2/io_i_6_in1[0]
+ cb_4_2/io_i_6_in1[1] cb_4_2/io_i_6_in1[2] cb_4_2/io_i_6_in1[3] cb_4_2/io_i_6_in1[4]
+ cb_4_2/io_i_6_in1[5] cb_4_2/io_i_6_in1[6] cb_4_2/io_i_6_in1[7] cb_4_2/io_i_7_ci
+ cb_4_2/io_i_7_in1[0] cb_4_2/io_i_7_in1[1] cb_4_2/io_i_7_in1[2] cb_4_2/io_i_7_in1[3]
+ cb_4_2/io_i_7_in1[4] cb_4_2/io_i_7_in1[5] cb_4_2/io_i_7_in1[6] cb_4_2/io_i_7_in1[7]
+ cb_4_3/io_i_0_ci cb_4_3/io_i_0_in1[0] cb_4_3/io_i_0_in1[1] cb_4_3/io_i_0_in1[2]
+ cb_4_3/io_i_0_in1[3] cb_4_3/io_i_0_in1[4] cb_4_3/io_i_0_in1[5] cb_4_3/io_i_0_in1[6]
+ cb_4_3/io_i_0_in1[7] cb_4_3/io_i_1_ci cb_4_3/io_i_1_in1[0] cb_4_3/io_i_1_in1[1]
+ cb_4_3/io_i_1_in1[2] cb_4_3/io_i_1_in1[3] cb_4_3/io_i_1_in1[4] cb_4_3/io_i_1_in1[5]
+ cb_4_3/io_i_1_in1[6] cb_4_3/io_i_1_in1[7] cb_4_3/io_i_2_ci cb_4_3/io_i_2_in1[0]
+ cb_4_3/io_i_2_in1[1] cb_4_3/io_i_2_in1[2] cb_4_3/io_i_2_in1[3] cb_4_3/io_i_2_in1[4]
+ cb_4_3/io_i_2_in1[5] cb_4_3/io_i_2_in1[6] cb_4_3/io_i_2_in1[7] cb_4_3/io_i_3_ci
+ cb_4_3/io_i_3_in1[0] cb_4_3/io_i_3_in1[1] cb_4_3/io_i_3_in1[2] cb_4_3/io_i_3_in1[3]
+ cb_4_3/io_i_3_in1[4] cb_4_3/io_i_3_in1[5] cb_4_3/io_i_3_in1[6] cb_4_3/io_i_3_in1[7]
+ cb_4_3/io_i_4_ci cb_4_3/io_i_4_in1[0] cb_4_3/io_i_4_in1[1] cb_4_3/io_i_4_in1[2]
+ cb_4_3/io_i_4_in1[3] cb_4_3/io_i_4_in1[4] cb_4_3/io_i_4_in1[5] cb_4_3/io_i_4_in1[6]
+ cb_4_3/io_i_4_in1[7] cb_4_3/io_i_5_ci cb_4_3/io_i_5_in1[0] cb_4_3/io_i_5_in1[1]
+ cb_4_3/io_i_5_in1[2] cb_4_3/io_i_5_in1[3] cb_4_3/io_i_5_in1[4] cb_4_3/io_i_5_in1[5]
+ cb_4_3/io_i_5_in1[6] cb_4_3/io_i_5_in1[7] cb_4_3/io_i_6_ci cb_4_3/io_i_6_in1[0]
+ cb_4_3/io_i_6_in1[1] cb_4_3/io_i_6_in1[2] cb_4_3/io_i_6_in1[3] cb_4_3/io_i_6_in1[4]
+ cb_4_3/io_i_6_in1[5] cb_4_3/io_i_6_in1[6] cb_4_3/io_i_6_in1[7] cb_4_3/io_i_7_ci
+ cb_4_3/io_i_7_in1[0] cb_4_3/io_i_7_in1[1] cb_4_3/io_i_7_in1[2] cb_4_3/io_i_7_in1[3]
+ cb_4_3/io_i_7_in1[4] cb_4_3/io_i_7_in1[5] cb_4_3/io_i_7_in1[6] cb_4_3/io_i_7_in1[7]
+ cb_4_2/io_vci cb_4_3/io_vci cb_4_2/io_vi cb_4_9/io_we_i cb_4_2/io_wo[0] cb_4_2/io_wo[10]
+ cb_4_2/io_wo[11] cb_4_2/io_wo[12] cb_4_2/io_wo[13] cb_4_2/io_wo[14] cb_4_2/io_wo[15]
+ cb_4_2/io_wo[16] cb_4_2/io_wo[17] cb_4_2/io_wo[18] cb_4_2/io_wo[19] cb_4_2/io_wo[1]
+ cb_4_2/io_wo[20] cb_4_2/io_wo[21] cb_4_2/io_wo[22] cb_4_2/io_wo[23] cb_4_2/io_wo[24]
+ cb_4_2/io_wo[25] cb_4_2/io_wo[26] cb_4_2/io_wo[27] cb_4_2/io_wo[28] cb_4_2/io_wo[29]
+ cb_4_2/io_wo[2] cb_4_2/io_wo[30] cb_4_2/io_wo[31] cb_4_2/io_wo[32] cb_4_2/io_wo[33]
+ cb_4_2/io_wo[34] cb_4_2/io_wo[35] cb_4_2/io_wo[36] cb_4_2/io_wo[37] cb_4_2/io_wo[38]
+ cb_4_2/io_wo[39] cb_4_2/io_wo[3] cb_4_2/io_wo[40] cb_4_2/io_wo[41] cb_4_2/io_wo[42]
+ cb_4_2/io_wo[43] cb_4_2/io_wo[44] cb_4_2/io_wo[45] cb_4_2/io_wo[46] cb_4_2/io_wo[47]
+ cb_4_2/io_wo[48] cb_4_2/io_wo[49] cb_4_2/io_wo[4] cb_4_2/io_wo[50] cb_4_2/io_wo[51]
+ cb_4_2/io_wo[52] cb_4_2/io_wo[53] cb_4_2/io_wo[54] cb_4_2/io_wo[55] cb_4_2/io_wo[56]
+ cb_4_2/io_wo[57] cb_4_2/io_wo[58] cb_4_2/io_wo[59] cb_4_2/io_wo[5] cb_4_2/io_wo[60]
+ cb_4_2/io_wo[61] cb_4_2/io_wo[62] cb_4_2/io_wo[63] cb_4_2/io_wo[6] cb_4_2/io_wo[7]
+ cb_4_2/io_wo[8] cb_4_2/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_6_6 cb_6_9/io_adr_i[0] cb_6_9/io_adr_i[1] cb_6_6/io_cs_i cb_6_9/io_dat_i[0] cb_6_9/io_dat_i[10]
+ cb_6_9/io_dat_i[11] cb_6_9/io_dat_i[12] cb_6_9/io_dat_i[13] cb_6_9/io_dat_i[14]
+ cb_6_9/io_dat_i[15] cb_6_9/io_dat_i[1] cb_6_9/io_dat_i[2] cb_6_9/io_dat_i[3] cb_6_9/io_dat_i[4]
+ cb_6_9/io_dat_i[5] cb_6_9/io_dat_i[6] cb_6_9/io_dat_i[7] cb_6_9/io_dat_i[8] cb_6_9/io_dat_i[9]
+ cb_6_6/io_dat_o[0] cb_6_6/io_dat_o[10] cb_6_6/io_dat_o[11] cb_6_6/io_dat_o[12] cb_6_6/io_dat_o[13]
+ cb_6_6/io_dat_o[14] cb_6_6/io_dat_o[15] cb_6_6/io_dat_o[1] cb_6_6/io_dat_o[2] cb_6_6/io_dat_o[3]
+ cb_6_6/io_dat_o[4] cb_6_6/io_dat_o[5] cb_6_6/io_dat_o[6] cb_6_6/io_dat_o[7] cb_6_6/io_dat_o[8]
+ cb_6_6/io_dat_o[9] cb_6_7/io_wo[0] cb_6_7/io_wo[10] cb_6_7/io_wo[11] cb_6_7/io_wo[12]
+ cb_6_7/io_wo[13] cb_6_7/io_wo[14] cb_6_7/io_wo[15] cb_6_7/io_wo[16] cb_6_7/io_wo[17]
+ cb_6_7/io_wo[18] cb_6_7/io_wo[19] cb_6_7/io_wo[1] cb_6_7/io_wo[20] cb_6_7/io_wo[21]
+ cb_6_7/io_wo[22] cb_6_7/io_wo[23] cb_6_7/io_wo[24] cb_6_7/io_wo[25] cb_6_7/io_wo[26]
+ cb_6_7/io_wo[27] cb_6_7/io_wo[28] cb_6_7/io_wo[29] cb_6_7/io_wo[2] cb_6_7/io_wo[30]
+ cb_6_7/io_wo[31] cb_6_7/io_wo[32] cb_6_7/io_wo[33] cb_6_7/io_wo[34] cb_6_7/io_wo[35]
+ cb_6_7/io_wo[36] cb_6_7/io_wo[37] cb_6_7/io_wo[38] cb_6_7/io_wo[39] cb_6_7/io_wo[3]
+ cb_6_7/io_wo[40] cb_6_7/io_wo[41] cb_6_7/io_wo[42] cb_6_7/io_wo[43] cb_6_7/io_wo[44]
+ cb_6_7/io_wo[45] cb_6_7/io_wo[46] cb_6_7/io_wo[47] cb_6_7/io_wo[48] cb_6_7/io_wo[49]
+ cb_6_7/io_wo[4] cb_6_7/io_wo[50] cb_6_7/io_wo[51] cb_6_7/io_wo[52] cb_6_7/io_wo[53]
+ cb_6_7/io_wo[54] cb_6_7/io_wo[55] cb_6_7/io_wo[56] cb_6_7/io_wo[57] cb_6_7/io_wo[58]
+ cb_6_7/io_wo[59] cb_6_7/io_wo[5] cb_6_7/io_wo[60] cb_6_7/io_wo[61] cb_6_7/io_wo[62]
+ cb_6_7/io_wo[63] cb_6_7/io_wo[6] cb_6_7/io_wo[7] cb_6_7/io_wo[8] cb_6_7/io_wo[9]
+ cb_6_6/io_i_0_ci cb_6_6/io_i_0_in1[0] cb_6_6/io_i_0_in1[1] cb_6_6/io_i_0_in1[2]
+ cb_6_6/io_i_0_in1[3] cb_6_6/io_i_0_in1[4] cb_6_6/io_i_0_in1[5] cb_6_6/io_i_0_in1[6]
+ cb_6_6/io_i_0_in1[7] cb_6_6/io_i_1_ci cb_6_6/io_i_1_in1[0] cb_6_6/io_i_1_in1[1]
+ cb_6_6/io_i_1_in1[2] cb_6_6/io_i_1_in1[3] cb_6_6/io_i_1_in1[4] cb_6_6/io_i_1_in1[5]
+ cb_6_6/io_i_1_in1[6] cb_6_6/io_i_1_in1[7] cb_6_6/io_i_2_ci cb_6_6/io_i_2_in1[0]
+ cb_6_6/io_i_2_in1[1] cb_6_6/io_i_2_in1[2] cb_6_6/io_i_2_in1[3] cb_6_6/io_i_2_in1[4]
+ cb_6_6/io_i_2_in1[5] cb_6_6/io_i_2_in1[6] cb_6_6/io_i_2_in1[7] cb_6_6/io_i_3_ci
+ cb_6_6/io_i_3_in1[0] cb_6_6/io_i_3_in1[1] cb_6_6/io_i_3_in1[2] cb_6_6/io_i_3_in1[3]
+ cb_6_6/io_i_3_in1[4] cb_6_6/io_i_3_in1[5] cb_6_6/io_i_3_in1[6] cb_6_6/io_i_3_in1[7]
+ cb_6_6/io_i_4_ci cb_6_6/io_i_4_in1[0] cb_6_6/io_i_4_in1[1] cb_6_6/io_i_4_in1[2]
+ cb_6_6/io_i_4_in1[3] cb_6_6/io_i_4_in1[4] cb_6_6/io_i_4_in1[5] cb_6_6/io_i_4_in1[6]
+ cb_6_6/io_i_4_in1[7] cb_6_6/io_i_5_ci cb_6_6/io_i_5_in1[0] cb_6_6/io_i_5_in1[1]
+ cb_6_6/io_i_5_in1[2] cb_6_6/io_i_5_in1[3] cb_6_6/io_i_5_in1[4] cb_6_6/io_i_5_in1[5]
+ cb_6_6/io_i_5_in1[6] cb_6_6/io_i_5_in1[7] cb_6_6/io_i_6_ci cb_6_6/io_i_6_in1[0]
+ cb_6_6/io_i_6_in1[1] cb_6_6/io_i_6_in1[2] cb_6_6/io_i_6_in1[3] cb_6_6/io_i_6_in1[4]
+ cb_6_6/io_i_6_in1[5] cb_6_6/io_i_6_in1[6] cb_6_6/io_i_6_in1[7] cb_6_6/io_i_7_ci
+ cb_6_6/io_i_7_in1[0] cb_6_6/io_i_7_in1[1] cb_6_6/io_i_7_in1[2] cb_6_6/io_i_7_in1[3]
+ cb_6_6/io_i_7_in1[4] cb_6_6/io_i_7_in1[5] cb_6_6/io_i_7_in1[6] cb_6_6/io_i_7_in1[7]
+ cb_6_7/io_i_0_ci cb_6_7/io_i_0_in1[0] cb_6_7/io_i_0_in1[1] cb_6_7/io_i_0_in1[2]
+ cb_6_7/io_i_0_in1[3] cb_6_7/io_i_0_in1[4] cb_6_7/io_i_0_in1[5] cb_6_7/io_i_0_in1[6]
+ cb_6_7/io_i_0_in1[7] cb_6_7/io_i_1_ci cb_6_7/io_i_1_in1[0] cb_6_7/io_i_1_in1[1]
+ cb_6_7/io_i_1_in1[2] cb_6_7/io_i_1_in1[3] cb_6_7/io_i_1_in1[4] cb_6_7/io_i_1_in1[5]
+ cb_6_7/io_i_1_in1[6] cb_6_7/io_i_1_in1[7] cb_6_7/io_i_2_ci cb_6_7/io_i_2_in1[0]
+ cb_6_7/io_i_2_in1[1] cb_6_7/io_i_2_in1[2] cb_6_7/io_i_2_in1[3] cb_6_7/io_i_2_in1[4]
+ cb_6_7/io_i_2_in1[5] cb_6_7/io_i_2_in1[6] cb_6_7/io_i_2_in1[7] cb_6_7/io_i_3_ci
+ cb_6_7/io_i_3_in1[0] cb_6_7/io_i_3_in1[1] cb_6_7/io_i_3_in1[2] cb_6_7/io_i_3_in1[3]
+ cb_6_7/io_i_3_in1[4] cb_6_7/io_i_3_in1[5] cb_6_7/io_i_3_in1[6] cb_6_7/io_i_3_in1[7]
+ cb_6_7/io_i_4_ci cb_6_7/io_i_4_in1[0] cb_6_7/io_i_4_in1[1] cb_6_7/io_i_4_in1[2]
+ cb_6_7/io_i_4_in1[3] cb_6_7/io_i_4_in1[4] cb_6_7/io_i_4_in1[5] cb_6_7/io_i_4_in1[6]
+ cb_6_7/io_i_4_in1[7] cb_6_7/io_i_5_ci cb_6_7/io_i_5_in1[0] cb_6_7/io_i_5_in1[1]
+ cb_6_7/io_i_5_in1[2] cb_6_7/io_i_5_in1[3] cb_6_7/io_i_5_in1[4] cb_6_7/io_i_5_in1[5]
+ cb_6_7/io_i_5_in1[6] cb_6_7/io_i_5_in1[7] cb_6_7/io_i_6_ci cb_6_7/io_i_6_in1[0]
+ cb_6_7/io_i_6_in1[1] cb_6_7/io_i_6_in1[2] cb_6_7/io_i_6_in1[3] cb_6_7/io_i_6_in1[4]
+ cb_6_7/io_i_6_in1[5] cb_6_7/io_i_6_in1[6] cb_6_7/io_i_6_in1[7] cb_6_7/io_i_7_ci
+ cb_6_7/io_i_7_in1[0] cb_6_7/io_i_7_in1[1] cb_6_7/io_i_7_in1[2] cb_6_7/io_i_7_in1[3]
+ cb_6_7/io_i_7_in1[4] cb_6_7/io_i_7_in1[5] cb_6_7/io_i_7_in1[6] cb_6_7/io_i_7_in1[7]
+ cb_6_6/io_vci cb_6_7/io_vci cb_6_6/io_vi cb_6_9/io_we_i cb_6_6/io_wo[0] cb_6_6/io_wo[10]
+ cb_6_6/io_wo[11] cb_6_6/io_wo[12] cb_6_6/io_wo[13] cb_6_6/io_wo[14] cb_6_6/io_wo[15]
+ cb_6_6/io_wo[16] cb_6_6/io_wo[17] cb_6_6/io_wo[18] cb_6_6/io_wo[19] cb_6_6/io_wo[1]
+ cb_6_6/io_wo[20] cb_6_6/io_wo[21] cb_6_6/io_wo[22] cb_6_6/io_wo[23] cb_6_6/io_wo[24]
+ cb_6_6/io_wo[25] cb_6_6/io_wo[26] cb_6_6/io_wo[27] cb_6_6/io_wo[28] cb_6_6/io_wo[29]
+ cb_6_6/io_wo[2] cb_6_6/io_wo[30] cb_6_6/io_wo[31] cb_6_6/io_wo[32] cb_6_6/io_wo[33]
+ cb_6_6/io_wo[34] cb_6_6/io_wo[35] cb_6_6/io_wo[36] cb_6_6/io_wo[37] cb_6_6/io_wo[38]
+ cb_6_6/io_wo[39] cb_6_6/io_wo[3] cb_6_6/io_wo[40] cb_6_6/io_wo[41] cb_6_6/io_wo[42]
+ cb_6_6/io_wo[43] cb_6_6/io_wo[44] cb_6_6/io_wo[45] cb_6_6/io_wo[46] cb_6_6/io_wo[47]
+ cb_6_6/io_wo[48] cb_6_6/io_wo[49] cb_6_6/io_wo[4] cb_6_6/io_wo[50] cb_6_6/io_wo[51]
+ cb_6_6/io_wo[52] cb_6_6/io_wo[53] cb_6_6/io_wo[54] cb_6_6/io_wo[55] cb_6_6/io_wo[56]
+ cb_6_6/io_wo[57] cb_6_6/io_wo[58] cb_6_6/io_wo[59] cb_6_6/io_wo[5] cb_6_6/io_wo[60]
+ cb_6_6/io_wo[61] cb_6_6/io_wo[62] cb_6_6/io_wo[63] cb_6_6/io_wo[6] cb_6_6/io_wo[7]
+ cb_6_6/io_wo[8] cb_6_6/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_4_3 cb_4_9/io_adr_i[0] cb_4_9/io_adr_i[1] cb_4_3/io_cs_i cb_4_9/io_dat_i[0] cb_4_9/io_dat_i[10]
+ cb_4_9/io_dat_i[11] cb_4_9/io_dat_i[12] cb_4_9/io_dat_i[13] cb_4_9/io_dat_i[14]
+ cb_4_9/io_dat_i[15] cb_4_9/io_dat_i[1] cb_4_9/io_dat_i[2] cb_4_9/io_dat_i[3] cb_4_9/io_dat_i[4]
+ cb_4_9/io_dat_i[5] cb_4_9/io_dat_i[6] cb_4_9/io_dat_i[7] cb_4_9/io_dat_i[8] cb_4_9/io_dat_i[9]
+ cb_4_3/io_dat_o[0] cb_4_3/io_dat_o[10] cb_4_3/io_dat_o[11] cb_4_3/io_dat_o[12] cb_4_3/io_dat_o[13]
+ cb_4_3/io_dat_o[14] cb_4_3/io_dat_o[15] cb_4_3/io_dat_o[1] cb_4_3/io_dat_o[2] cb_4_3/io_dat_o[3]
+ cb_4_3/io_dat_o[4] cb_4_3/io_dat_o[5] cb_4_3/io_dat_o[6] cb_4_3/io_dat_o[7] cb_4_3/io_dat_o[8]
+ cb_4_3/io_dat_o[9] cb_4_4/io_wo[0] cb_4_4/io_wo[10] cb_4_4/io_wo[11] cb_4_4/io_wo[12]
+ cb_4_4/io_wo[13] cb_4_4/io_wo[14] cb_4_4/io_wo[15] cb_4_4/io_wo[16] cb_4_4/io_wo[17]
+ cb_4_4/io_wo[18] cb_4_4/io_wo[19] cb_4_4/io_wo[1] cb_4_4/io_wo[20] cb_4_4/io_wo[21]
+ cb_4_4/io_wo[22] cb_4_4/io_wo[23] cb_4_4/io_wo[24] cb_4_4/io_wo[25] cb_4_4/io_wo[26]
+ cb_4_4/io_wo[27] cb_4_4/io_wo[28] cb_4_4/io_wo[29] cb_4_4/io_wo[2] cb_4_4/io_wo[30]
+ cb_4_4/io_wo[31] cb_4_4/io_wo[32] cb_4_4/io_wo[33] cb_4_4/io_wo[34] cb_4_4/io_wo[35]
+ cb_4_4/io_wo[36] cb_4_4/io_wo[37] cb_4_4/io_wo[38] cb_4_4/io_wo[39] cb_4_4/io_wo[3]
+ cb_4_4/io_wo[40] cb_4_4/io_wo[41] cb_4_4/io_wo[42] cb_4_4/io_wo[43] cb_4_4/io_wo[44]
+ cb_4_4/io_wo[45] cb_4_4/io_wo[46] cb_4_4/io_wo[47] cb_4_4/io_wo[48] cb_4_4/io_wo[49]
+ cb_4_4/io_wo[4] cb_4_4/io_wo[50] cb_4_4/io_wo[51] cb_4_4/io_wo[52] cb_4_4/io_wo[53]
+ cb_4_4/io_wo[54] cb_4_4/io_wo[55] cb_4_4/io_wo[56] cb_4_4/io_wo[57] cb_4_4/io_wo[58]
+ cb_4_4/io_wo[59] cb_4_4/io_wo[5] cb_4_4/io_wo[60] cb_4_4/io_wo[61] cb_4_4/io_wo[62]
+ cb_4_4/io_wo[63] cb_4_4/io_wo[6] cb_4_4/io_wo[7] cb_4_4/io_wo[8] cb_4_4/io_wo[9]
+ cb_4_3/io_i_0_ci cb_4_3/io_i_0_in1[0] cb_4_3/io_i_0_in1[1] cb_4_3/io_i_0_in1[2]
+ cb_4_3/io_i_0_in1[3] cb_4_3/io_i_0_in1[4] cb_4_3/io_i_0_in1[5] cb_4_3/io_i_0_in1[6]
+ cb_4_3/io_i_0_in1[7] cb_4_3/io_i_1_ci cb_4_3/io_i_1_in1[0] cb_4_3/io_i_1_in1[1]
+ cb_4_3/io_i_1_in1[2] cb_4_3/io_i_1_in1[3] cb_4_3/io_i_1_in1[4] cb_4_3/io_i_1_in1[5]
+ cb_4_3/io_i_1_in1[6] cb_4_3/io_i_1_in1[7] cb_4_3/io_i_2_ci cb_4_3/io_i_2_in1[0]
+ cb_4_3/io_i_2_in1[1] cb_4_3/io_i_2_in1[2] cb_4_3/io_i_2_in1[3] cb_4_3/io_i_2_in1[4]
+ cb_4_3/io_i_2_in1[5] cb_4_3/io_i_2_in1[6] cb_4_3/io_i_2_in1[7] cb_4_3/io_i_3_ci
+ cb_4_3/io_i_3_in1[0] cb_4_3/io_i_3_in1[1] cb_4_3/io_i_3_in1[2] cb_4_3/io_i_3_in1[3]
+ cb_4_3/io_i_3_in1[4] cb_4_3/io_i_3_in1[5] cb_4_3/io_i_3_in1[6] cb_4_3/io_i_3_in1[7]
+ cb_4_3/io_i_4_ci cb_4_3/io_i_4_in1[0] cb_4_3/io_i_4_in1[1] cb_4_3/io_i_4_in1[2]
+ cb_4_3/io_i_4_in1[3] cb_4_3/io_i_4_in1[4] cb_4_3/io_i_4_in1[5] cb_4_3/io_i_4_in1[6]
+ cb_4_3/io_i_4_in1[7] cb_4_3/io_i_5_ci cb_4_3/io_i_5_in1[0] cb_4_3/io_i_5_in1[1]
+ cb_4_3/io_i_5_in1[2] cb_4_3/io_i_5_in1[3] cb_4_3/io_i_5_in1[4] cb_4_3/io_i_5_in1[5]
+ cb_4_3/io_i_5_in1[6] cb_4_3/io_i_5_in1[7] cb_4_3/io_i_6_ci cb_4_3/io_i_6_in1[0]
+ cb_4_3/io_i_6_in1[1] cb_4_3/io_i_6_in1[2] cb_4_3/io_i_6_in1[3] cb_4_3/io_i_6_in1[4]
+ cb_4_3/io_i_6_in1[5] cb_4_3/io_i_6_in1[6] cb_4_3/io_i_6_in1[7] cb_4_3/io_i_7_ci
+ cb_4_3/io_i_7_in1[0] cb_4_3/io_i_7_in1[1] cb_4_3/io_i_7_in1[2] cb_4_3/io_i_7_in1[3]
+ cb_4_3/io_i_7_in1[4] cb_4_3/io_i_7_in1[5] cb_4_3/io_i_7_in1[6] cb_4_3/io_i_7_in1[7]
+ cb_4_4/io_i_0_ci cb_4_4/io_i_0_in1[0] cb_4_4/io_i_0_in1[1] cb_4_4/io_i_0_in1[2]
+ cb_4_4/io_i_0_in1[3] cb_4_4/io_i_0_in1[4] cb_4_4/io_i_0_in1[5] cb_4_4/io_i_0_in1[6]
+ cb_4_4/io_i_0_in1[7] cb_4_4/io_i_1_ci cb_4_4/io_i_1_in1[0] cb_4_4/io_i_1_in1[1]
+ cb_4_4/io_i_1_in1[2] cb_4_4/io_i_1_in1[3] cb_4_4/io_i_1_in1[4] cb_4_4/io_i_1_in1[5]
+ cb_4_4/io_i_1_in1[6] cb_4_4/io_i_1_in1[7] cb_4_4/io_i_2_ci cb_4_4/io_i_2_in1[0]
+ cb_4_4/io_i_2_in1[1] cb_4_4/io_i_2_in1[2] cb_4_4/io_i_2_in1[3] cb_4_4/io_i_2_in1[4]
+ cb_4_4/io_i_2_in1[5] cb_4_4/io_i_2_in1[6] cb_4_4/io_i_2_in1[7] cb_4_4/io_i_3_ci
+ cb_4_4/io_i_3_in1[0] cb_4_4/io_i_3_in1[1] cb_4_4/io_i_3_in1[2] cb_4_4/io_i_3_in1[3]
+ cb_4_4/io_i_3_in1[4] cb_4_4/io_i_3_in1[5] cb_4_4/io_i_3_in1[6] cb_4_4/io_i_3_in1[7]
+ cb_4_4/io_i_4_ci cb_4_4/io_i_4_in1[0] cb_4_4/io_i_4_in1[1] cb_4_4/io_i_4_in1[2]
+ cb_4_4/io_i_4_in1[3] cb_4_4/io_i_4_in1[4] cb_4_4/io_i_4_in1[5] cb_4_4/io_i_4_in1[6]
+ cb_4_4/io_i_4_in1[7] cb_4_4/io_i_5_ci cb_4_4/io_i_5_in1[0] cb_4_4/io_i_5_in1[1]
+ cb_4_4/io_i_5_in1[2] cb_4_4/io_i_5_in1[3] cb_4_4/io_i_5_in1[4] cb_4_4/io_i_5_in1[5]
+ cb_4_4/io_i_5_in1[6] cb_4_4/io_i_5_in1[7] cb_4_4/io_i_6_ci cb_4_4/io_i_6_in1[0]
+ cb_4_4/io_i_6_in1[1] cb_4_4/io_i_6_in1[2] cb_4_4/io_i_6_in1[3] cb_4_4/io_i_6_in1[4]
+ cb_4_4/io_i_6_in1[5] cb_4_4/io_i_6_in1[6] cb_4_4/io_i_6_in1[7] cb_4_4/io_i_7_ci
+ cb_4_4/io_i_7_in1[0] cb_4_4/io_i_7_in1[1] cb_4_4/io_i_7_in1[2] cb_4_4/io_i_7_in1[3]
+ cb_4_4/io_i_7_in1[4] cb_4_4/io_i_7_in1[5] cb_4_4/io_i_7_in1[6] cb_4_4/io_i_7_in1[7]
+ cb_4_3/io_vci cb_4_4/io_vci cb_4_3/io_vi cb_4_9/io_we_i cb_4_3/io_wo[0] cb_4_3/io_wo[10]
+ cb_4_3/io_wo[11] cb_4_3/io_wo[12] cb_4_3/io_wo[13] cb_4_3/io_wo[14] cb_4_3/io_wo[15]
+ cb_4_3/io_wo[16] cb_4_3/io_wo[17] cb_4_3/io_wo[18] cb_4_3/io_wo[19] cb_4_3/io_wo[1]
+ cb_4_3/io_wo[20] cb_4_3/io_wo[21] cb_4_3/io_wo[22] cb_4_3/io_wo[23] cb_4_3/io_wo[24]
+ cb_4_3/io_wo[25] cb_4_3/io_wo[26] cb_4_3/io_wo[27] cb_4_3/io_wo[28] cb_4_3/io_wo[29]
+ cb_4_3/io_wo[2] cb_4_3/io_wo[30] cb_4_3/io_wo[31] cb_4_3/io_wo[32] cb_4_3/io_wo[33]
+ cb_4_3/io_wo[34] cb_4_3/io_wo[35] cb_4_3/io_wo[36] cb_4_3/io_wo[37] cb_4_3/io_wo[38]
+ cb_4_3/io_wo[39] cb_4_3/io_wo[3] cb_4_3/io_wo[40] cb_4_3/io_wo[41] cb_4_3/io_wo[42]
+ cb_4_3/io_wo[43] cb_4_3/io_wo[44] cb_4_3/io_wo[45] cb_4_3/io_wo[46] cb_4_3/io_wo[47]
+ cb_4_3/io_wo[48] cb_4_3/io_wo[49] cb_4_3/io_wo[4] cb_4_3/io_wo[50] cb_4_3/io_wo[51]
+ cb_4_3/io_wo[52] cb_4_3/io_wo[53] cb_4_3/io_wo[54] cb_4_3/io_wo[55] cb_4_3/io_wo[56]
+ cb_4_3/io_wo[57] cb_4_3/io_wo[58] cb_4_3/io_wo[59] cb_4_3/io_wo[5] cb_4_3/io_wo[60]
+ cb_4_3/io_wo[61] cb_4_3/io_wo[62] cb_4_3/io_wo[63] cb_4_3/io_wo[6] cb_4_3/io_wo[7]
+ cb_4_3/io_wo[8] cb_4_3/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_2_0 cb_2_9/io_adr_i[0] cb_2_9/io_adr_i[1] cb_2_0/io_cs_i cb_2_9/io_dat_i[0] cb_2_9/io_dat_i[10]
+ cb_2_9/io_dat_i[11] cb_2_9/io_dat_i[12] cb_2_9/io_dat_i[13] cb_2_9/io_dat_i[14]
+ cb_2_9/io_dat_i[15] cb_2_9/io_dat_i[1] cb_2_9/io_dat_i[2] cb_2_9/io_dat_i[3] cb_2_9/io_dat_i[4]
+ cb_2_9/io_dat_i[5] cb_2_9/io_dat_i[6] cb_2_9/io_dat_i[7] cb_2_9/io_dat_i[8] cb_2_9/io_dat_i[9]
+ cb_2_0/io_dat_o[0] cb_2_0/io_dat_o[10] cb_2_0/io_dat_o[11] cb_2_0/io_dat_o[12] cb_2_0/io_dat_o[13]
+ cb_2_0/io_dat_o[14] cb_2_0/io_dat_o[15] cb_2_0/io_dat_o[1] cb_2_0/io_dat_o[2] cb_2_0/io_dat_o[3]
+ cb_2_0/io_dat_o[4] cb_2_0/io_dat_o[5] cb_2_0/io_dat_o[6] cb_2_0/io_dat_o[7] cb_2_0/io_dat_o[8]
+ cb_2_0/io_dat_o[9] cb_2_1/io_wo[0] cb_2_1/io_wo[10] cb_2_1/io_wo[11] cb_2_1/io_wo[12]
+ cb_2_1/io_wo[13] cb_2_1/io_wo[14] cb_2_1/io_wo[15] cb_2_1/io_wo[16] cb_2_1/io_wo[17]
+ cb_2_1/io_wo[18] cb_2_1/io_wo[19] cb_2_1/io_wo[1] cb_2_1/io_wo[20] cb_2_1/io_wo[21]
+ cb_2_1/io_wo[22] cb_2_1/io_wo[23] cb_2_1/io_wo[24] cb_2_1/io_wo[25] cb_2_1/io_wo[26]
+ cb_2_1/io_wo[27] cb_2_1/io_wo[28] cb_2_1/io_wo[29] cb_2_1/io_wo[2] cb_2_1/io_wo[30]
+ cb_2_1/io_wo[31] cb_2_1/io_wo[32] cb_2_1/io_wo[33] cb_2_1/io_wo[34] cb_2_1/io_wo[35]
+ cb_2_1/io_wo[36] cb_2_1/io_wo[37] cb_2_1/io_wo[38] cb_2_1/io_wo[39] cb_2_1/io_wo[3]
+ cb_2_1/io_wo[40] cb_2_1/io_wo[41] cb_2_1/io_wo[42] cb_2_1/io_wo[43] cb_2_1/io_wo[44]
+ cb_2_1/io_wo[45] cb_2_1/io_wo[46] cb_2_1/io_wo[47] cb_2_1/io_wo[48] cb_2_1/io_wo[49]
+ cb_2_1/io_wo[4] cb_2_1/io_wo[50] cb_2_1/io_wo[51] cb_2_1/io_wo[52] cb_2_1/io_wo[53]
+ cb_2_1/io_wo[54] cb_2_1/io_wo[55] cb_2_1/io_wo[56] cb_2_1/io_wo[57] cb_2_1/io_wo[58]
+ cb_2_1/io_wo[59] cb_2_1/io_wo[5] cb_2_1/io_wo[60] cb_2_1/io_wo[61] cb_2_1/io_wo[62]
+ cb_2_1/io_wo[63] cb_2_1/io_wo[6] cb_2_1/io_wo[7] cb_2_1/io_wo[8] cb_2_1/io_wo[9]
+ ccon_2/io_dsi_o cb_2_0/io_i_0_in1[0] cb_2_0/io_i_0_in1[1] cb_2_0/io_i_0_in1[2] cb_2_0/io_i_0_in1[3]
+ cb_2_0/io_i_0_in1[4] cb_2_0/io_i_0_in1[5] cb_2_0/io_i_0_in1[6] cb_2_0/io_i_0_in1[7]
+ cb_2_0/io_i_1_ci cb_2_0/io_i_1_in1[0] cb_2_0/io_i_1_in1[1] cb_2_0/io_i_1_in1[2]
+ cb_2_0/io_i_1_in1[3] cb_2_0/io_i_1_in1[4] cb_2_0/io_i_1_in1[5] cb_2_0/io_i_1_in1[6]
+ cb_2_0/io_i_1_in1[7] cb_2_0/io_i_2_ci cb_2_0/io_i_2_in1[0] cb_2_0/io_i_2_in1[1]
+ cb_2_0/io_i_2_in1[2] cb_2_0/io_i_2_in1[3] cb_2_0/io_i_2_in1[4] cb_2_0/io_i_2_in1[5]
+ cb_2_0/io_i_2_in1[6] cb_2_0/io_i_2_in1[7] cb_2_0/io_i_3_ci cb_2_0/io_i_3_in1[0]
+ cb_2_0/io_i_3_in1[1] cb_2_0/io_i_3_in1[2] cb_2_0/io_i_3_in1[3] cb_2_0/io_i_3_in1[4]
+ cb_2_0/io_i_3_in1[5] cb_2_0/io_i_3_in1[6] cb_2_0/io_i_3_in1[7] cb_2_0/io_i_4_ci
+ cb_2_0/io_i_4_in1[0] cb_2_0/io_i_4_in1[1] cb_2_0/io_i_4_in1[2] cb_2_0/io_i_4_in1[3]
+ cb_2_0/io_i_4_in1[4] cb_2_0/io_i_4_in1[5] cb_2_0/io_i_4_in1[6] cb_2_0/io_i_4_in1[7]
+ cb_2_0/io_i_5_ci cb_2_0/io_i_5_in1[0] cb_2_0/io_i_5_in1[1] cb_2_0/io_i_5_in1[2]
+ cb_2_0/io_i_5_in1[3] cb_2_0/io_i_5_in1[4] cb_2_0/io_i_5_in1[5] cb_2_0/io_i_5_in1[6]
+ cb_2_0/io_i_5_in1[7] cb_2_0/io_i_6_ci cb_2_0/io_i_6_in1[0] cb_2_0/io_i_6_in1[1]
+ cb_2_0/io_i_6_in1[2] cb_2_0/io_i_6_in1[3] cb_2_0/io_i_6_in1[4] cb_2_0/io_i_6_in1[5]
+ cb_2_0/io_i_6_in1[6] cb_2_0/io_i_6_in1[7] cb_2_0/io_i_7_ci cb_2_0/io_i_7_in1[0]
+ cb_2_0/io_i_7_in1[1] cb_2_0/io_i_7_in1[2] cb_2_0/io_i_7_in1[3] cb_2_0/io_i_7_in1[4]
+ cb_2_0/io_i_7_in1[5] cb_2_0/io_i_7_in1[6] cb_2_0/io_i_7_in1[7] cb_2_1/io_i_0_ci
+ cb_2_1/io_i_0_in1[0] cb_2_1/io_i_0_in1[1] cb_2_1/io_i_0_in1[2] cb_2_1/io_i_0_in1[3]
+ cb_2_1/io_i_0_in1[4] cb_2_1/io_i_0_in1[5] cb_2_1/io_i_0_in1[6] cb_2_1/io_i_0_in1[7]
+ cb_2_1/io_i_1_ci cb_2_1/io_i_1_in1[0] cb_2_1/io_i_1_in1[1] cb_2_1/io_i_1_in1[2]
+ cb_2_1/io_i_1_in1[3] cb_2_1/io_i_1_in1[4] cb_2_1/io_i_1_in1[5] cb_2_1/io_i_1_in1[6]
+ cb_2_1/io_i_1_in1[7] cb_2_1/io_i_2_ci cb_2_1/io_i_2_in1[0] cb_2_1/io_i_2_in1[1]
+ cb_2_1/io_i_2_in1[2] cb_2_1/io_i_2_in1[3] cb_2_1/io_i_2_in1[4] cb_2_1/io_i_2_in1[5]
+ cb_2_1/io_i_2_in1[6] cb_2_1/io_i_2_in1[7] cb_2_1/io_i_3_ci cb_2_1/io_i_3_in1[0]
+ cb_2_1/io_i_3_in1[1] cb_2_1/io_i_3_in1[2] cb_2_1/io_i_3_in1[3] cb_2_1/io_i_3_in1[4]
+ cb_2_1/io_i_3_in1[5] cb_2_1/io_i_3_in1[6] cb_2_1/io_i_3_in1[7] cb_2_1/io_i_4_ci
+ cb_2_1/io_i_4_in1[0] cb_2_1/io_i_4_in1[1] cb_2_1/io_i_4_in1[2] cb_2_1/io_i_4_in1[3]
+ cb_2_1/io_i_4_in1[4] cb_2_1/io_i_4_in1[5] cb_2_1/io_i_4_in1[6] cb_2_1/io_i_4_in1[7]
+ cb_2_1/io_i_5_ci cb_2_1/io_i_5_in1[0] cb_2_1/io_i_5_in1[1] cb_2_1/io_i_5_in1[2]
+ cb_2_1/io_i_5_in1[3] cb_2_1/io_i_5_in1[4] cb_2_1/io_i_5_in1[5] cb_2_1/io_i_5_in1[6]
+ cb_2_1/io_i_5_in1[7] cb_2_1/io_i_6_ci cb_2_1/io_i_6_in1[0] cb_2_1/io_i_6_in1[1]
+ cb_2_1/io_i_6_in1[2] cb_2_1/io_i_6_in1[3] cb_2_1/io_i_6_in1[4] cb_2_1/io_i_6_in1[5]
+ cb_2_1/io_i_6_in1[6] cb_2_1/io_i_6_in1[7] cb_2_1/io_i_7_ci cb_2_1/io_i_7_in1[0]
+ cb_2_1/io_i_7_in1[1] cb_2_1/io_i_7_in1[2] cb_2_1/io_i_7_in1[3] cb_2_1/io_i_7_in1[4]
+ cb_2_1/io_i_7_in1[5] cb_2_1/io_i_7_in1[6] cb_2_1/io_i_7_in1[7] cb_2_0/io_vci cb_2_1/io_vci
+ cb_2_0/io_vi cb_2_9/io_we_i cb_2_0/io_wo[0] cb_2_0/io_wo[10] cb_2_0/io_wo[11] cb_2_0/io_wo[12]
+ cb_2_0/io_wo[13] cb_2_0/io_wo[14] cb_2_0/io_wo[15] cb_2_0/io_wo[16] cb_2_0/io_wo[17]
+ cb_2_0/io_wo[18] cb_2_0/io_wo[19] cb_2_0/io_wo[1] cb_2_0/io_wo[20] cb_2_0/io_wo[21]
+ cb_2_0/io_wo[22] cb_2_0/io_wo[23] cb_2_0/io_wo[24] cb_2_0/io_wo[25] cb_2_0/io_wo[26]
+ cb_2_0/io_wo[27] cb_2_0/io_wo[28] cb_2_0/io_wo[29] cb_2_0/io_wo[2] cb_2_0/io_wo[30]
+ cb_2_0/io_wo[31] cb_2_0/io_wo[32] cb_2_0/io_wo[33] cb_2_0/io_wo[34] cb_2_0/io_wo[35]
+ cb_2_0/io_wo[36] cb_2_0/io_wo[37] cb_2_0/io_wo[38] cb_2_0/io_wo[39] cb_2_0/io_wo[3]
+ cb_2_0/io_wo[40] cb_2_0/io_wo[41] cb_2_0/io_wo[42] cb_2_0/io_wo[43] cb_2_0/io_wo[44]
+ cb_2_0/io_wo[45] cb_2_0/io_wo[46] cb_2_0/io_wo[47] cb_2_0/io_wo[48] cb_2_0/io_wo[49]
+ cb_2_0/io_wo[4] cb_2_0/io_wo[50] cb_2_0/io_wo[51] cb_2_0/io_wo[52] cb_2_0/io_wo[53]
+ cb_2_0/io_wo[54] cb_2_0/io_wo[55] cb_2_0/io_wo[56] cb_2_0/io_wo[57] cb_2_0/io_wo[58]
+ cb_2_0/io_wo[59] cb_2_0/io_wo[5] cb_2_0/io_wo[60] cb_2_0/io_wo[61] cb_2_0/io_wo[62]
+ cb_2_0/io_wo[63] cb_2_0/io_wo[6] cb_2_0/io_wo[7] cb_2_0/io_wo[8] cb_2_0/io_wo[9]
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_6_7 cb_6_9/io_adr_i[0] cb_6_9/io_adr_i[1] cb_6_7/io_cs_i cb_6_9/io_dat_i[0] cb_6_9/io_dat_i[10]
+ cb_6_9/io_dat_i[11] cb_6_9/io_dat_i[12] cb_6_9/io_dat_i[13] cb_6_9/io_dat_i[14]
+ cb_6_9/io_dat_i[15] cb_6_9/io_dat_i[1] cb_6_9/io_dat_i[2] cb_6_9/io_dat_i[3] cb_6_9/io_dat_i[4]
+ cb_6_9/io_dat_i[5] cb_6_9/io_dat_i[6] cb_6_9/io_dat_i[7] cb_6_9/io_dat_i[8] cb_6_9/io_dat_i[9]
+ cb_6_7/io_dat_o[0] cb_6_7/io_dat_o[10] cb_6_7/io_dat_o[11] cb_6_7/io_dat_o[12] cb_6_7/io_dat_o[13]
+ cb_6_7/io_dat_o[14] cb_6_7/io_dat_o[15] cb_6_7/io_dat_o[1] cb_6_7/io_dat_o[2] cb_6_7/io_dat_o[3]
+ cb_6_7/io_dat_o[4] cb_6_7/io_dat_o[5] cb_6_7/io_dat_o[6] cb_6_7/io_dat_o[7] cb_6_7/io_dat_o[8]
+ cb_6_7/io_dat_o[9] cb_6_8/io_wo[0] cb_6_8/io_wo[10] cb_6_8/io_wo[11] cb_6_8/io_wo[12]
+ cb_6_8/io_wo[13] cb_6_8/io_wo[14] cb_6_8/io_wo[15] cb_6_8/io_wo[16] cb_6_8/io_wo[17]
+ cb_6_8/io_wo[18] cb_6_8/io_wo[19] cb_6_8/io_wo[1] cb_6_8/io_wo[20] cb_6_8/io_wo[21]
+ cb_6_8/io_wo[22] cb_6_8/io_wo[23] cb_6_8/io_wo[24] cb_6_8/io_wo[25] cb_6_8/io_wo[26]
+ cb_6_8/io_wo[27] cb_6_8/io_wo[28] cb_6_8/io_wo[29] cb_6_8/io_wo[2] cb_6_8/io_wo[30]
+ cb_6_8/io_wo[31] cb_6_8/io_wo[32] cb_6_8/io_wo[33] cb_6_8/io_wo[34] cb_6_8/io_wo[35]
+ cb_6_8/io_wo[36] cb_6_8/io_wo[37] cb_6_8/io_wo[38] cb_6_8/io_wo[39] cb_6_8/io_wo[3]
+ cb_6_8/io_wo[40] cb_6_8/io_wo[41] cb_6_8/io_wo[42] cb_6_8/io_wo[43] cb_6_8/io_wo[44]
+ cb_6_8/io_wo[45] cb_6_8/io_wo[46] cb_6_8/io_wo[47] cb_6_8/io_wo[48] cb_6_8/io_wo[49]
+ cb_6_8/io_wo[4] cb_6_8/io_wo[50] cb_6_8/io_wo[51] cb_6_8/io_wo[52] cb_6_8/io_wo[53]
+ cb_6_8/io_wo[54] cb_6_8/io_wo[55] cb_6_8/io_wo[56] cb_6_8/io_wo[57] cb_6_8/io_wo[58]
+ cb_6_8/io_wo[59] cb_6_8/io_wo[5] cb_6_8/io_wo[60] cb_6_8/io_wo[61] cb_6_8/io_wo[62]
+ cb_6_8/io_wo[63] cb_6_8/io_wo[6] cb_6_8/io_wo[7] cb_6_8/io_wo[8] cb_6_8/io_wo[9]
+ cb_6_7/io_i_0_ci cb_6_7/io_i_0_in1[0] cb_6_7/io_i_0_in1[1] cb_6_7/io_i_0_in1[2]
+ cb_6_7/io_i_0_in1[3] cb_6_7/io_i_0_in1[4] cb_6_7/io_i_0_in1[5] cb_6_7/io_i_0_in1[6]
+ cb_6_7/io_i_0_in1[7] cb_6_7/io_i_1_ci cb_6_7/io_i_1_in1[0] cb_6_7/io_i_1_in1[1]
+ cb_6_7/io_i_1_in1[2] cb_6_7/io_i_1_in1[3] cb_6_7/io_i_1_in1[4] cb_6_7/io_i_1_in1[5]
+ cb_6_7/io_i_1_in1[6] cb_6_7/io_i_1_in1[7] cb_6_7/io_i_2_ci cb_6_7/io_i_2_in1[0]
+ cb_6_7/io_i_2_in1[1] cb_6_7/io_i_2_in1[2] cb_6_7/io_i_2_in1[3] cb_6_7/io_i_2_in1[4]
+ cb_6_7/io_i_2_in1[5] cb_6_7/io_i_2_in1[6] cb_6_7/io_i_2_in1[7] cb_6_7/io_i_3_ci
+ cb_6_7/io_i_3_in1[0] cb_6_7/io_i_3_in1[1] cb_6_7/io_i_3_in1[2] cb_6_7/io_i_3_in1[3]
+ cb_6_7/io_i_3_in1[4] cb_6_7/io_i_3_in1[5] cb_6_7/io_i_3_in1[6] cb_6_7/io_i_3_in1[7]
+ cb_6_7/io_i_4_ci cb_6_7/io_i_4_in1[0] cb_6_7/io_i_4_in1[1] cb_6_7/io_i_4_in1[2]
+ cb_6_7/io_i_4_in1[3] cb_6_7/io_i_4_in1[4] cb_6_7/io_i_4_in1[5] cb_6_7/io_i_4_in1[6]
+ cb_6_7/io_i_4_in1[7] cb_6_7/io_i_5_ci cb_6_7/io_i_5_in1[0] cb_6_7/io_i_5_in1[1]
+ cb_6_7/io_i_5_in1[2] cb_6_7/io_i_5_in1[3] cb_6_7/io_i_5_in1[4] cb_6_7/io_i_5_in1[5]
+ cb_6_7/io_i_5_in1[6] cb_6_7/io_i_5_in1[7] cb_6_7/io_i_6_ci cb_6_7/io_i_6_in1[0]
+ cb_6_7/io_i_6_in1[1] cb_6_7/io_i_6_in1[2] cb_6_7/io_i_6_in1[3] cb_6_7/io_i_6_in1[4]
+ cb_6_7/io_i_6_in1[5] cb_6_7/io_i_6_in1[6] cb_6_7/io_i_6_in1[7] cb_6_7/io_i_7_ci
+ cb_6_7/io_i_7_in1[0] cb_6_7/io_i_7_in1[1] cb_6_7/io_i_7_in1[2] cb_6_7/io_i_7_in1[3]
+ cb_6_7/io_i_7_in1[4] cb_6_7/io_i_7_in1[5] cb_6_7/io_i_7_in1[6] cb_6_7/io_i_7_in1[7]
+ cb_6_8/io_i_0_ci cb_6_8/io_i_0_in1[0] cb_6_8/io_i_0_in1[1] cb_6_8/io_i_0_in1[2]
+ cb_6_8/io_i_0_in1[3] cb_6_8/io_i_0_in1[4] cb_6_8/io_i_0_in1[5] cb_6_8/io_i_0_in1[6]
+ cb_6_8/io_i_0_in1[7] cb_6_8/io_i_1_ci cb_6_8/io_i_1_in1[0] cb_6_8/io_i_1_in1[1]
+ cb_6_8/io_i_1_in1[2] cb_6_8/io_i_1_in1[3] cb_6_8/io_i_1_in1[4] cb_6_8/io_i_1_in1[5]
+ cb_6_8/io_i_1_in1[6] cb_6_8/io_i_1_in1[7] cb_6_8/io_i_2_ci cb_6_8/io_i_2_in1[0]
+ cb_6_8/io_i_2_in1[1] cb_6_8/io_i_2_in1[2] cb_6_8/io_i_2_in1[3] cb_6_8/io_i_2_in1[4]
+ cb_6_8/io_i_2_in1[5] cb_6_8/io_i_2_in1[6] cb_6_8/io_i_2_in1[7] cb_6_8/io_i_3_ci
+ cb_6_8/io_i_3_in1[0] cb_6_8/io_i_3_in1[1] cb_6_8/io_i_3_in1[2] cb_6_8/io_i_3_in1[3]
+ cb_6_8/io_i_3_in1[4] cb_6_8/io_i_3_in1[5] cb_6_8/io_i_3_in1[6] cb_6_8/io_i_3_in1[7]
+ cb_6_8/io_i_4_ci cb_6_8/io_i_4_in1[0] cb_6_8/io_i_4_in1[1] cb_6_8/io_i_4_in1[2]
+ cb_6_8/io_i_4_in1[3] cb_6_8/io_i_4_in1[4] cb_6_8/io_i_4_in1[5] cb_6_8/io_i_4_in1[6]
+ cb_6_8/io_i_4_in1[7] cb_6_8/io_i_5_ci cb_6_8/io_i_5_in1[0] cb_6_8/io_i_5_in1[1]
+ cb_6_8/io_i_5_in1[2] cb_6_8/io_i_5_in1[3] cb_6_8/io_i_5_in1[4] cb_6_8/io_i_5_in1[5]
+ cb_6_8/io_i_5_in1[6] cb_6_8/io_i_5_in1[7] cb_6_8/io_i_6_ci cb_6_8/io_i_6_in1[0]
+ cb_6_8/io_i_6_in1[1] cb_6_8/io_i_6_in1[2] cb_6_8/io_i_6_in1[3] cb_6_8/io_i_6_in1[4]
+ cb_6_8/io_i_6_in1[5] cb_6_8/io_i_6_in1[6] cb_6_8/io_i_6_in1[7] cb_6_8/io_i_7_ci
+ cb_6_8/io_i_7_in1[0] cb_6_8/io_i_7_in1[1] cb_6_8/io_i_7_in1[2] cb_6_8/io_i_7_in1[3]
+ cb_6_8/io_i_7_in1[4] cb_6_8/io_i_7_in1[5] cb_6_8/io_i_7_in1[6] cb_6_8/io_i_7_in1[7]
+ cb_6_7/io_vci cb_6_8/io_vci cb_6_7/io_vi cb_6_9/io_we_i cb_6_7/io_wo[0] cb_6_7/io_wo[10]
+ cb_6_7/io_wo[11] cb_6_7/io_wo[12] cb_6_7/io_wo[13] cb_6_7/io_wo[14] cb_6_7/io_wo[15]
+ cb_6_7/io_wo[16] cb_6_7/io_wo[17] cb_6_7/io_wo[18] cb_6_7/io_wo[19] cb_6_7/io_wo[1]
+ cb_6_7/io_wo[20] cb_6_7/io_wo[21] cb_6_7/io_wo[22] cb_6_7/io_wo[23] cb_6_7/io_wo[24]
+ cb_6_7/io_wo[25] cb_6_7/io_wo[26] cb_6_7/io_wo[27] cb_6_7/io_wo[28] cb_6_7/io_wo[29]
+ cb_6_7/io_wo[2] cb_6_7/io_wo[30] cb_6_7/io_wo[31] cb_6_7/io_wo[32] cb_6_7/io_wo[33]
+ cb_6_7/io_wo[34] cb_6_7/io_wo[35] cb_6_7/io_wo[36] cb_6_7/io_wo[37] cb_6_7/io_wo[38]
+ cb_6_7/io_wo[39] cb_6_7/io_wo[3] cb_6_7/io_wo[40] cb_6_7/io_wo[41] cb_6_7/io_wo[42]
+ cb_6_7/io_wo[43] cb_6_7/io_wo[44] cb_6_7/io_wo[45] cb_6_7/io_wo[46] cb_6_7/io_wo[47]
+ cb_6_7/io_wo[48] cb_6_7/io_wo[49] cb_6_7/io_wo[4] cb_6_7/io_wo[50] cb_6_7/io_wo[51]
+ cb_6_7/io_wo[52] cb_6_7/io_wo[53] cb_6_7/io_wo[54] cb_6_7/io_wo[55] cb_6_7/io_wo[56]
+ cb_6_7/io_wo[57] cb_6_7/io_wo[58] cb_6_7/io_wo[59] cb_6_7/io_wo[5] cb_6_7/io_wo[60]
+ cb_6_7/io_wo[61] cb_6_7/io_wo[62] cb_6_7/io_wo[63] cb_6_7/io_wo[6] cb_6_7/io_wo[7]
+ cb_6_7/io_wo[8] cb_6_7/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_4_4 cb_4_9/io_adr_i[0] cb_4_9/io_adr_i[1] cb_4_4/io_cs_i cb_4_9/io_dat_i[0] cb_4_9/io_dat_i[10]
+ cb_4_9/io_dat_i[11] cb_4_9/io_dat_i[12] cb_4_9/io_dat_i[13] cb_4_9/io_dat_i[14]
+ cb_4_9/io_dat_i[15] cb_4_9/io_dat_i[1] cb_4_9/io_dat_i[2] cb_4_9/io_dat_i[3] cb_4_9/io_dat_i[4]
+ cb_4_9/io_dat_i[5] cb_4_9/io_dat_i[6] cb_4_9/io_dat_i[7] cb_4_9/io_dat_i[8] cb_4_9/io_dat_i[9]
+ cb_4_4/io_dat_o[0] cb_4_4/io_dat_o[10] cb_4_4/io_dat_o[11] cb_4_4/io_dat_o[12] cb_4_4/io_dat_o[13]
+ cb_4_4/io_dat_o[14] cb_4_4/io_dat_o[15] cb_4_4/io_dat_o[1] cb_4_4/io_dat_o[2] cb_4_4/io_dat_o[3]
+ cb_4_4/io_dat_o[4] cb_4_4/io_dat_o[5] cb_4_4/io_dat_o[6] cb_4_4/io_dat_o[7] cb_4_4/io_dat_o[8]
+ cb_4_4/io_dat_o[9] cb_4_5/io_wo[0] cb_4_5/io_wo[10] cb_4_5/io_wo[11] cb_4_5/io_wo[12]
+ cb_4_5/io_wo[13] cb_4_5/io_wo[14] cb_4_5/io_wo[15] cb_4_5/io_wo[16] cb_4_5/io_wo[17]
+ cb_4_5/io_wo[18] cb_4_5/io_wo[19] cb_4_5/io_wo[1] cb_4_5/io_wo[20] cb_4_5/io_wo[21]
+ cb_4_5/io_wo[22] cb_4_5/io_wo[23] cb_4_5/io_wo[24] cb_4_5/io_wo[25] cb_4_5/io_wo[26]
+ cb_4_5/io_wo[27] cb_4_5/io_wo[28] cb_4_5/io_wo[29] cb_4_5/io_wo[2] cb_4_5/io_wo[30]
+ cb_4_5/io_wo[31] cb_4_5/io_wo[32] cb_4_5/io_wo[33] cb_4_5/io_wo[34] cb_4_5/io_wo[35]
+ cb_4_5/io_wo[36] cb_4_5/io_wo[37] cb_4_5/io_wo[38] cb_4_5/io_wo[39] cb_4_5/io_wo[3]
+ cb_4_5/io_wo[40] cb_4_5/io_wo[41] cb_4_5/io_wo[42] cb_4_5/io_wo[43] cb_4_5/io_wo[44]
+ cb_4_5/io_wo[45] cb_4_5/io_wo[46] cb_4_5/io_wo[47] cb_4_5/io_wo[48] cb_4_5/io_wo[49]
+ cb_4_5/io_wo[4] cb_4_5/io_wo[50] cb_4_5/io_wo[51] cb_4_5/io_wo[52] cb_4_5/io_wo[53]
+ cb_4_5/io_wo[54] cb_4_5/io_wo[55] cb_4_5/io_wo[56] cb_4_5/io_wo[57] cb_4_5/io_wo[58]
+ cb_4_5/io_wo[59] cb_4_5/io_wo[5] cb_4_5/io_wo[60] cb_4_5/io_wo[61] cb_4_5/io_wo[62]
+ cb_4_5/io_wo[63] cb_4_5/io_wo[6] cb_4_5/io_wo[7] cb_4_5/io_wo[8] cb_4_5/io_wo[9]
+ cb_4_4/io_i_0_ci cb_4_4/io_i_0_in1[0] cb_4_4/io_i_0_in1[1] cb_4_4/io_i_0_in1[2]
+ cb_4_4/io_i_0_in1[3] cb_4_4/io_i_0_in1[4] cb_4_4/io_i_0_in1[5] cb_4_4/io_i_0_in1[6]
+ cb_4_4/io_i_0_in1[7] cb_4_4/io_i_1_ci cb_4_4/io_i_1_in1[0] cb_4_4/io_i_1_in1[1]
+ cb_4_4/io_i_1_in1[2] cb_4_4/io_i_1_in1[3] cb_4_4/io_i_1_in1[4] cb_4_4/io_i_1_in1[5]
+ cb_4_4/io_i_1_in1[6] cb_4_4/io_i_1_in1[7] cb_4_4/io_i_2_ci cb_4_4/io_i_2_in1[0]
+ cb_4_4/io_i_2_in1[1] cb_4_4/io_i_2_in1[2] cb_4_4/io_i_2_in1[3] cb_4_4/io_i_2_in1[4]
+ cb_4_4/io_i_2_in1[5] cb_4_4/io_i_2_in1[6] cb_4_4/io_i_2_in1[7] cb_4_4/io_i_3_ci
+ cb_4_4/io_i_3_in1[0] cb_4_4/io_i_3_in1[1] cb_4_4/io_i_3_in1[2] cb_4_4/io_i_3_in1[3]
+ cb_4_4/io_i_3_in1[4] cb_4_4/io_i_3_in1[5] cb_4_4/io_i_3_in1[6] cb_4_4/io_i_3_in1[7]
+ cb_4_4/io_i_4_ci cb_4_4/io_i_4_in1[0] cb_4_4/io_i_4_in1[1] cb_4_4/io_i_4_in1[2]
+ cb_4_4/io_i_4_in1[3] cb_4_4/io_i_4_in1[4] cb_4_4/io_i_4_in1[5] cb_4_4/io_i_4_in1[6]
+ cb_4_4/io_i_4_in1[7] cb_4_4/io_i_5_ci cb_4_4/io_i_5_in1[0] cb_4_4/io_i_5_in1[1]
+ cb_4_4/io_i_5_in1[2] cb_4_4/io_i_5_in1[3] cb_4_4/io_i_5_in1[4] cb_4_4/io_i_5_in1[5]
+ cb_4_4/io_i_5_in1[6] cb_4_4/io_i_5_in1[7] cb_4_4/io_i_6_ci cb_4_4/io_i_6_in1[0]
+ cb_4_4/io_i_6_in1[1] cb_4_4/io_i_6_in1[2] cb_4_4/io_i_6_in1[3] cb_4_4/io_i_6_in1[4]
+ cb_4_4/io_i_6_in1[5] cb_4_4/io_i_6_in1[6] cb_4_4/io_i_6_in1[7] cb_4_4/io_i_7_ci
+ cb_4_4/io_i_7_in1[0] cb_4_4/io_i_7_in1[1] cb_4_4/io_i_7_in1[2] cb_4_4/io_i_7_in1[3]
+ cb_4_4/io_i_7_in1[4] cb_4_4/io_i_7_in1[5] cb_4_4/io_i_7_in1[6] cb_4_4/io_i_7_in1[7]
+ cb_4_5/io_i_0_ci cb_4_5/io_i_0_in1[0] cb_4_5/io_i_0_in1[1] cb_4_5/io_i_0_in1[2]
+ cb_4_5/io_i_0_in1[3] cb_4_5/io_i_0_in1[4] cb_4_5/io_i_0_in1[5] cb_4_5/io_i_0_in1[6]
+ cb_4_5/io_i_0_in1[7] cb_4_5/io_i_1_ci cb_4_5/io_i_1_in1[0] cb_4_5/io_i_1_in1[1]
+ cb_4_5/io_i_1_in1[2] cb_4_5/io_i_1_in1[3] cb_4_5/io_i_1_in1[4] cb_4_5/io_i_1_in1[5]
+ cb_4_5/io_i_1_in1[6] cb_4_5/io_i_1_in1[7] cb_4_5/io_i_2_ci cb_4_5/io_i_2_in1[0]
+ cb_4_5/io_i_2_in1[1] cb_4_5/io_i_2_in1[2] cb_4_5/io_i_2_in1[3] cb_4_5/io_i_2_in1[4]
+ cb_4_5/io_i_2_in1[5] cb_4_5/io_i_2_in1[6] cb_4_5/io_i_2_in1[7] cb_4_5/io_i_3_ci
+ cb_4_5/io_i_3_in1[0] cb_4_5/io_i_3_in1[1] cb_4_5/io_i_3_in1[2] cb_4_5/io_i_3_in1[3]
+ cb_4_5/io_i_3_in1[4] cb_4_5/io_i_3_in1[5] cb_4_5/io_i_3_in1[6] cb_4_5/io_i_3_in1[7]
+ cb_4_5/io_i_4_ci cb_4_5/io_i_4_in1[0] cb_4_5/io_i_4_in1[1] cb_4_5/io_i_4_in1[2]
+ cb_4_5/io_i_4_in1[3] cb_4_5/io_i_4_in1[4] cb_4_5/io_i_4_in1[5] cb_4_5/io_i_4_in1[6]
+ cb_4_5/io_i_4_in1[7] cb_4_5/io_i_5_ci cb_4_5/io_i_5_in1[0] cb_4_5/io_i_5_in1[1]
+ cb_4_5/io_i_5_in1[2] cb_4_5/io_i_5_in1[3] cb_4_5/io_i_5_in1[4] cb_4_5/io_i_5_in1[5]
+ cb_4_5/io_i_5_in1[6] cb_4_5/io_i_5_in1[7] cb_4_5/io_i_6_ci cb_4_5/io_i_6_in1[0]
+ cb_4_5/io_i_6_in1[1] cb_4_5/io_i_6_in1[2] cb_4_5/io_i_6_in1[3] cb_4_5/io_i_6_in1[4]
+ cb_4_5/io_i_6_in1[5] cb_4_5/io_i_6_in1[6] cb_4_5/io_i_6_in1[7] cb_4_5/io_i_7_ci
+ cb_4_5/io_i_7_in1[0] cb_4_5/io_i_7_in1[1] cb_4_5/io_i_7_in1[2] cb_4_5/io_i_7_in1[3]
+ cb_4_5/io_i_7_in1[4] cb_4_5/io_i_7_in1[5] cb_4_5/io_i_7_in1[6] cb_4_5/io_i_7_in1[7]
+ cb_4_4/io_vci cb_4_5/io_vci cb_4_4/io_vi cb_4_9/io_we_i cb_4_4/io_wo[0] cb_4_4/io_wo[10]
+ cb_4_4/io_wo[11] cb_4_4/io_wo[12] cb_4_4/io_wo[13] cb_4_4/io_wo[14] cb_4_4/io_wo[15]
+ cb_4_4/io_wo[16] cb_4_4/io_wo[17] cb_4_4/io_wo[18] cb_4_4/io_wo[19] cb_4_4/io_wo[1]
+ cb_4_4/io_wo[20] cb_4_4/io_wo[21] cb_4_4/io_wo[22] cb_4_4/io_wo[23] cb_4_4/io_wo[24]
+ cb_4_4/io_wo[25] cb_4_4/io_wo[26] cb_4_4/io_wo[27] cb_4_4/io_wo[28] cb_4_4/io_wo[29]
+ cb_4_4/io_wo[2] cb_4_4/io_wo[30] cb_4_4/io_wo[31] cb_4_4/io_wo[32] cb_4_4/io_wo[33]
+ cb_4_4/io_wo[34] cb_4_4/io_wo[35] cb_4_4/io_wo[36] cb_4_4/io_wo[37] cb_4_4/io_wo[38]
+ cb_4_4/io_wo[39] cb_4_4/io_wo[3] cb_4_4/io_wo[40] cb_4_4/io_wo[41] cb_4_4/io_wo[42]
+ cb_4_4/io_wo[43] cb_4_4/io_wo[44] cb_4_4/io_wo[45] cb_4_4/io_wo[46] cb_4_4/io_wo[47]
+ cb_4_4/io_wo[48] cb_4_4/io_wo[49] cb_4_4/io_wo[4] cb_4_4/io_wo[50] cb_4_4/io_wo[51]
+ cb_4_4/io_wo[52] cb_4_4/io_wo[53] cb_4_4/io_wo[54] cb_4_4/io_wo[55] cb_4_4/io_wo[56]
+ cb_4_4/io_wo[57] cb_4_4/io_wo[58] cb_4_4/io_wo[59] cb_4_4/io_wo[5] cb_4_4/io_wo[60]
+ cb_4_4/io_wo[61] cb_4_4/io_wo[62] cb_4_4/io_wo[63] cb_4_4/io_wo[6] cb_4_4/io_wo[7]
+ cb_4_4/io_wo[8] cb_4_4/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_2_1 cb_2_9/io_adr_i[0] cb_2_9/io_adr_i[1] cb_2_1/io_cs_i cb_2_9/io_dat_i[0] cb_2_9/io_dat_i[10]
+ cb_2_9/io_dat_i[11] cb_2_9/io_dat_i[12] cb_2_9/io_dat_i[13] cb_2_9/io_dat_i[14]
+ cb_2_9/io_dat_i[15] cb_2_9/io_dat_i[1] cb_2_9/io_dat_i[2] cb_2_9/io_dat_i[3] cb_2_9/io_dat_i[4]
+ cb_2_9/io_dat_i[5] cb_2_9/io_dat_i[6] cb_2_9/io_dat_i[7] cb_2_9/io_dat_i[8] cb_2_9/io_dat_i[9]
+ cb_2_1/io_dat_o[0] cb_2_1/io_dat_o[10] cb_2_1/io_dat_o[11] cb_2_1/io_dat_o[12] cb_2_1/io_dat_o[13]
+ cb_2_1/io_dat_o[14] cb_2_1/io_dat_o[15] cb_2_1/io_dat_o[1] cb_2_1/io_dat_o[2] cb_2_1/io_dat_o[3]
+ cb_2_1/io_dat_o[4] cb_2_1/io_dat_o[5] cb_2_1/io_dat_o[6] cb_2_1/io_dat_o[7] cb_2_1/io_dat_o[8]
+ cb_2_1/io_dat_o[9] cb_2_2/io_wo[0] cb_2_2/io_wo[10] cb_2_2/io_wo[11] cb_2_2/io_wo[12]
+ cb_2_2/io_wo[13] cb_2_2/io_wo[14] cb_2_2/io_wo[15] cb_2_2/io_wo[16] cb_2_2/io_wo[17]
+ cb_2_2/io_wo[18] cb_2_2/io_wo[19] cb_2_2/io_wo[1] cb_2_2/io_wo[20] cb_2_2/io_wo[21]
+ cb_2_2/io_wo[22] cb_2_2/io_wo[23] cb_2_2/io_wo[24] cb_2_2/io_wo[25] cb_2_2/io_wo[26]
+ cb_2_2/io_wo[27] cb_2_2/io_wo[28] cb_2_2/io_wo[29] cb_2_2/io_wo[2] cb_2_2/io_wo[30]
+ cb_2_2/io_wo[31] cb_2_2/io_wo[32] cb_2_2/io_wo[33] cb_2_2/io_wo[34] cb_2_2/io_wo[35]
+ cb_2_2/io_wo[36] cb_2_2/io_wo[37] cb_2_2/io_wo[38] cb_2_2/io_wo[39] cb_2_2/io_wo[3]
+ cb_2_2/io_wo[40] cb_2_2/io_wo[41] cb_2_2/io_wo[42] cb_2_2/io_wo[43] cb_2_2/io_wo[44]
+ cb_2_2/io_wo[45] cb_2_2/io_wo[46] cb_2_2/io_wo[47] cb_2_2/io_wo[48] cb_2_2/io_wo[49]
+ cb_2_2/io_wo[4] cb_2_2/io_wo[50] cb_2_2/io_wo[51] cb_2_2/io_wo[52] cb_2_2/io_wo[53]
+ cb_2_2/io_wo[54] cb_2_2/io_wo[55] cb_2_2/io_wo[56] cb_2_2/io_wo[57] cb_2_2/io_wo[58]
+ cb_2_2/io_wo[59] cb_2_2/io_wo[5] cb_2_2/io_wo[60] cb_2_2/io_wo[61] cb_2_2/io_wo[62]
+ cb_2_2/io_wo[63] cb_2_2/io_wo[6] cb_2_2/io_wo[7] cb_2_2/io_wo[8] cb_2_2/io_wo[9]
+ cb_2_1/io_i_0_ci cb_2_1/io_i_0_in1[0] cb_2_1/io_i_0_in1[1] cb_2_1/io_i_0_in1[2]
+ cb_2_1/io_i_0_in1[3] cb_2_1/io_i_0_in1[4] cb_2_1/io_i_0_in1[5] cb_2_1/io_i_0_in1[6]
+ cb_2_1/io_i_0_in1[7] cb_2_1/io_i_1_ci cb_2_1/io_i_1_in1[0] cb_2_1/io_i_1_in1[1]
+ cb_2_1/io_i_1_in1[2] cb_2_1/io_i_1_in1[3] cb_2_1/io_i_1_in1[4] cb_2_1/io_i_1_in1[5]
+ cb_2_1/io_i_1_in1[6] cb_2_1/io_i_1_in1[7] cb_2_1/io_i_2_ci cb_2_1/io_i_2_in1[0]
+ cb_2_1/io_i_2_in1[1] cb_2_1/io_i_2_in1[2] cb_2_1/io_i_2_in1[3] cb_2_1/io_i_2_in1[4]
+ cb_2_1/io_i_2_in1[5] cb_2_1/io_i_2_in1[6] cb_2_1/io_i_2_in1[7] cb_2_1/io_i_3_ci
+ cb_2_1/io_i_3_in1[0] cb_2_1/io_i_3_in1[1] cb_2_1/io_i_3_in1[2] cb_2_1/io_i_3_in1[3]
+ cb_2_1/io_i_3_in1[4] cb_2_1/io_i_3_in1[5] cb_2_1/io_i_3_in1[6] cb_2_1/io_i_3_in1[7]
+ cb_2_1/io_i_4_ci cb_2_1/io_i_4_in1[0] cb_2_1/io_i_4_in1[1] cb_2_1/io_i_4_in1[2]
+ cb_2_1/io_i_4_in1[3] cb_2_1/io_i_4_in1[4] cb_2_1/io_i_4_in1[5] cb_2_1/io_i_4_in1[6]
+ cb_2_1/io_i_4_in1[7] cb_2_1/io_i_5_ci cb_2_1/io_i_5_in1[0] cb_2_1/io_i_5_in1[1]
+ cb_2_1/io_i_5_in1[2] cb_2_1/io_i_5_in1[3] cb_2_1/io_i_5_in1[4] cb_2_1/io_i_5_in1[5]
+ cb_2_1/io_i_5_in1[6] cb_2_1/io_i_5_in1[7] cb_2_1/io_i_6_ci cb_2_1/io_i_6_in1[0]
+ cb_2_1/io_i_6_in1[1] cb_2_1/io_i_6_in1[2] cb_2_1/io_i_6_in1[3] cb_2_1/io_i_6_in1[4]
+ cb_2_1/io_i_6_in1[5] cb_2_1/io_i_6_in1[6] cb_2_1/io_i_6_in1[7] cb_2_1/io_i_7_ci
+ cb_2_1/io_i_7_in1[0] cb_2_1/io_i_7_in1[1] cb_2_1/io_i_7_in1[2] cb_2_1/io_i_7_in1[3]
+ cb_2_1/io_i_7_in1[4] cb_2_1/io_i_7_in1[5] cb_2_1/io_i_7_in1[6] cb_2_1/io_i_7_in1[7]
+ cb_2_2/io_i_0_ci cb_2_2/io_i_0_in1[0] cb_2_2/io_i_0_in1[1] cb_2_2/io_i_0_in1[2]
+ cb_2_2/io_i_0_in1[3] cb_2_2/io_i_0_in1[4] cb_2_2/io_i_0_in1[5] cb_2_2/io_i_0_in1[6]
+ cb_2_2/io_i_0_in1[7] cb_2_2/io_i_1_ci cb_2_2/io_i_1_in1[0] cb_2_2/io_i_1_in1[1]
+ cb_2_2/io_i_1_in1[2] cb_2_2/io_i_1_in1[3] cb_2_2/io_i_1_in1[4] cb_2_2/io_i_1_in1[5]
+ cb_2_2/io_i_1_in1[6] cb_2_2/io_i_1_in1[7] cb_2_2/io_i_2_ci cb_2_2/io_i_2_in1[0]
+ cb_2_2/io_i_2_in1[1] cb_2_2/io_i_2_in1[2] cb_2_2/io_i_2_in1[3] cb_2_2/io_i_2_in1[4]
+ cb_2_2/io_i_2_in1[5] cb_2_2/io_i_2_in1[6] cb_2_2/io_i_2_in1[7] cb_2_2/io_i_3_ci
+ cb_2_2/io_i_3_in1[0] cb_2_2/io_i_3_in1[1] cb_2_2/io_i_3_in1[2] cb_2_2/io_i_3_in1[3]
+ cb_2_2/io_i_3_in1[4] cb_2_2/io_i_3_in1[5] cb_2_2/io_i_3_in1[6] cb_2_2/io_i_3_in1[7]
+ cb_2_2/io_i_4_ci cb_2_2/io_i_4_in1[0] cb_2_2/io_i_4_in1[1] cb_2_2/io_i_4_in1[2]
+ cb_2_2/io_i_4_in1[3] cb_2_2/io_i_4_in1[4] cb_2_2/io_i_4_in1[5] cb_2_2/io_i_4_in1[6]
+ cb_2_2/io_i_4_in1[7] cb_2_2/io_i_5_ci cb_2_2/io_i_5_in1[0] cb_2_2/io_i_5_in1[1]
+ cb_2_2/io_i_5_in1[2] cb_2_2/io_i_5_in1[3] cb_2_2/io_i_5_in1[4] cb_2_2/io_i_5_in1[5]
+ cb_2_2/io_i_5_in1[6] cb_2_2/io_i_5_in1[7] cb_2_2/io_i_6_ci cb_2_2/io_i_6_in1[0]
+ cb_2_2/io_i_6_in1[1] cb_2_2/io_i_6_in1[2] cb_2_2/io_i_6_in1[3] cb_2_2/io_i_6_in1[4]
+ cb_2_2/io_i_6_in1[5] cb_2_2/io_i_6_in1[6] cb_2_2/io_i_6_in1[7] cb_2_2/io_i_7_ci
+ cb_2_2/io_i_7_in1[0] cb_2_2/io_i_7_in1[1] cb_2_2/io_i_7_in1[2] cb_2_2/io_i_7_in1[3]
+ cb_2_2/io_i_7_in1[4] cb_2_2/io_i_7_in1[5] cb_2_2/io_i_7_in1[6] cb_2_2/io_i_7_in1[7]
+ cb_2_1/io_vci cb_2_2/io_vci cb_2_1/io_vi cb_2_9/io_we_i cb_2_1/io_wo[0] cb_2_1/io_wo[10]
+ cb_2_1/io_wo[11] cb_2_1/io_wo[12] cb_2_1/io_wo[13] cb_2_1/io_wo[14] cb_2_1/io_wo[15]
+ cb_2_1/io_wo[16] cb_2_1/io_wo[17] cb_2_1/io_wo[18] cb_2_1/io_wo[19] cb_2_1/io_wo[1]
+ cb_2_1/io_wo[20] cb_2_1/io_wo[21] cb_2_1/io_wo[22] cb_2_1/io_wo[23] cb_2_1/io_wo[24]
+ cb_2_1/io_wo[25] cb_2_1/io_wo[26] cb_2_1/io_wo[27] cb_2_1/io_wo[28] cb_2_1/io_wo[29]
+ cb_2_1/io_wo[2] cb_2_1/io_wo[30] cb_2_1/io_wo[31] cb_2_1/io_wo[32] cb_2_1/io_wo[33]
+ cb_2_1/io_wo[34] cb_2_1/io_wo[35] cb_2_1/io_wo[36] cb_2_1/io_wo[37] cb_2_1/io_wo[38]
+ cb_2_1/io_wo[39] cb_2_1/io_wo[3] cb_2_1/io_wo[40] cb_2_1/io_wo[41] cb_2_1/io_wo[42]
+ cb_2_1/io_wo[43] cb_2_1/io_wo[44] cb_2_1/io_wo[45] cb_2_1/io_wo[46] cb_2_1/io_wo[47]
+ cb_2_1/io_wo[48] cb_2_1/io_wo[49] cb_2_1/io_wo[4] cb_2_1/io_wo[50] cb_2_1/io_wo[51]
+ cb_2_1/io_wo[52] cb_2_1/io_wo[53] cb_2_1/io_wo[54] cb_2_1/io_wo[55] cb_2_1/io_wo[56]
+ cb_2_1/io_wo[57] cb_2_1/io_wo[58] cb_2_1/io_wo[59] cb_2_1/io_wo[5] cb_2_1/io_wo[60]
+ cb_2_1/io_wo[61] cb_2_1/io_wo[62] cb_2_1/io_wo[63] cb_2_1/io_wo[6] cb_2_1/io_wo[7]
+ cb_2_1/io_wo[8] cb_2_1/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_6_8 cb_6_9/io_adr_i[0] cb_6_9/io_adr_i[1] cb_6_8/io_cs_i cb_6_9/io_dat_i[0] cb_6_9/io_dat_i[10]
+ cb_6_9/io_dat_i[11] cb_6_9/io_dat_i[12] cb_6_9/io_dat_i[13] cb_6_9/io_dat_i[14]
+ cb_6_9/io_dat_i[15] cb_6_9/io_dat_i[1] cb_6_9/io_dat_i[2] cb_6_9/io_dat_i[3] cb_6_9/io_dat_i[4]
+ cb_6_9/io_dat_i[5] cb_6_9/io_dat_i[6] cb_6_9/io_dat_i[7] cb_6_9/io_dat_i[8] cb_6_9/io_dat_i[9]
+ cb_6_8/io_dat_o[0] cb_6_8/io_dat_o[10] cb_6_8/io_dat_o[11] cb_6_8/io_dat_o[12] cb_6_8/io_dat_o[13]
+ cb_6_8/io_dat_o[14] cb_6_8/io_dat_o[15] cb_6_8/io_dat_o[1] cb_6_8/io_dat_o[2] cb_6_8/io_dat_o[3]
+ cb_6_8/io_dat_o[4] cb_6_8/io_dat_o[5] cb_6_8/io_dat_o[6] cb_6_8/io_dat_o[7] cb_6_8/io_dat_o[8]
+ cb_6_8/io_dat_o[9] cb_6_9/io_wo[0] cb_6_9/io_wo[10] cb_6_9/io_wo[11] cb_6_9/io_wo[12]
+ cb_6_9/io_wo[13] cb_6_9/io_wo[14] cb_6_9/io_wo[15] cb_6_9/io_wo[16] cb_6_9/io_wo[17]
+ cb_6_9/io_wo[18] cb_6_9/io_wo[19] cb_6_9/io_wo[1] cb_6_9/io_wo[20] cb_6_9/io_wo[21]
+ cb_6_9/io_wo[22] cb_6_9/io_wo[23] cb_6_9/io_wo[24] cb_6_9/io_wo[25] cb_6_9/io_wo[26]
+ cb_6_9/io_wo[27] cb_6_9/io_wo[28] cb_6_9/io_wo[29] cb_6_9/io_wo[2] cb_6_9/io_wo[30]
+ cb_6_9/io_wo[31] cb_6_9/io_wo[32] cb_6_9/io_wo[33] cb_6_9/io_wo[34] cb_6_9/io_wo[35]
+ cb_6_9/io_wo[36] cb_6_9/io_wo[37] cb_6_9/io_wo[38] cb_6_9/io_wo[39] cb_6_9/io_wo[3]
+ cb_6_9/io_wo[40] cb_6_9/io_wo[41] cb_6_9/io_wo[42] cb_6_9/io_wo[43] cb_6_9/io_wo[44]
+ cb_6_9/io_wo[45] cb_6_9/io_wo[46] cb_6_9/io_wo[47] cb_6_9/io_wo[48] cb_6_9/io_wo[49]
+ cb_6_9/io_wo[4] cb_6_9/io_wo[50] cb_6_9/io_wo[51] cb_6_9/io_wo[52] cb_6_9/io_wo[53]
+ cb_6_9/io_wo[54] cb_6_9/io_wo[55] cb_6_9/io_wo[56] cb_6_9/io_wo[57] cb_6_9/io_wo[58]
+ cb_6_9/io_wo[59] cb_6_9/io_wo[5] cb_6_9/io_wo[60] cb_6_9/io_wo[61] cb_6_9/io_wo[62]
+ cb_6_9/io_wo[63] cb_6_9/io_wo[6] cb_6_9/io_wo[7] cb_6_9/io_wo[8] cb_6_9/io_wo[9]
+ cb_6_8/io_i_0_ci cb_6_8/io_i_0_in1[0] cb_6_8/io_i_0_in1[1] cb_6_8/io_i_0_in1[2]
+ cb_6_8/io_i_0_in1[3] cb_6_8/io_i_0_in1[4] cb_6_8/io_i_0_in1[5] cb_6_8/io_i_0_in1[6]
+ cb_6_8/io_i_0_in1[7] cb_6_8/io_i_1_ci cb_6_8/io_i_1_in1[0] cb_6_8/io_i_1_in1[1]
+ cb_6_8/io_i_1_in1[2] cb_6_8/io_i_1_in1[3] cb_6_8/io_i_1_in1[4] cb_6_8/io_i_1_in1[5]
+ cb_6_8/io_i_1_in1[6] cb_6_8/io_i_1_in1[7] cb_6_8/io_i_2_ci cb_6_8/io_i_2_in1[0]
+ cb_6_8/io_i_2_in1[1] cb_6_8/io_i_2_in1[2] cb_6_8/io_i_2_in1[3] cb_6_8/io_i_2_in1[4]
+ cb_6_8/io_i_2_in1[5] cb_6_8/io_i_2_in1[6] cb_6_8/io_i_2_in1[7] cb_6_8/io_i_3_ci
+ cb_6_8/io_i_3_in1[0] cb_6_8/io_i_3_in1[1] cb_6_8/io_i_3_in1[2] cb_6_8/io_i_3_in1[3]
+ cb_6_8/io_i_3_in1[4] cb_6_8/io_i_3_in1[5] cb_6_8/io_i_3_in1[6] cb_6_8/io_i_3_in1[7]
+ cb_6_8/io_i_4_ci cb_6_8/io_i_4_in1[0] cb_6_8/io_i_4_in1[1] cb_6_8/io_i_4_in1[2]
+ cb_6_8/io_i_4_in1[3] cb_6_8/io_i_4_in1[4] cb_6_8/io_i_4_in1[5] cb_6_8/io_i_4_in1[6]
+ cb_6_8/io_i_4_in1[7] cb_6_8/io_i_5_ci cb_6_8/io_i_5_in1[0] cb_6_8/io_i_5_in1[1]
+ cb_6_8/io_i_5_in1[2] cb_6_8/io_i_5_in1[3] cb_6_8/io_i_5_in1[4] cb_6_8/io_i_5_in1[5]
+ cb_6_8/io_i_5_in1[6] cb_6_8/io_i_5_in1[7] cb_6_8/io_i_6_ci cb_6_8/io_i_6_in1[0]
+ cb_6_8/io_i_6_in1[1] cb_6_8/io_i_6_in1[2] cb_6_8/io_i_6_in1[3] cb_6_8/io_i_6_in1[4]
+ cb_6_8/io_i_6_in1[5] cb_6_8/io_i_6_in1[6] cb_6_8/io_i_6_in1[7] cb_6_8/io_i_7_ci
+ cb_6_8/io_i_7_in1[0] cb_6_8/io_i_7_in1[1] cb_6_8/io_i_7_in1[2] cb_6_8/io_i_7_in1[3]
+ cb_6_8/io_i_7_in1[4] cb_6_8/io_i_7_in1[5] cb_6_8/io_i_7_in1[6] cb_6_8/io_i_7_in1[7]
+ cb_6_9/io_i_0_ci cb_6_9/io_i_0_in1[0] cb_6_9/io_i_0_in1[1] cb_6_9/io_i_0_in1[2]
+ cb_6_9/io_i_0_in1[3] cb_6_9/io_i_0_in1[4] cb_6_9/io_i_0_in1[5] cb_6_9/io_i_0_in1[6]
+ cb_6_9/io_i_0_in1[7] cb_6_9/io_i_1_ci cb_6_9/io_i_1_in1[0] cb_6_9/io_i_1_in1[1]
+ cb_6_9/io_i_1_in1[2] cb_6_9/io_i_1_in1[3] cb_6_9/io_i_1_in1[4] cb_6_9/io_i_1_in1[5]
+ cb_6_9/io_i_1_in1[6] cb_6_9/io_i_1_in1[7] cb_6_9/io_i_2_ci cb_6_9/io_i_2_in1[0]
+ cb_6_9/io_i_2_in1[1] cb_6_9/io_i_2_in1[2] cb_6_9/io_i_2_in1[3] cb_6_9/io_i_2_in1[4]
+ cb_6_9/io_i_2_in1[5] cb_6_9/io_i_2_in1[6] cb_6_9/io_i_2_in1[7] cb_6_9/io_i_3_ci
+ cb_6_9/io_i_3_in1[0] cb_6_9/io_i_3_in1[1] cb_6_9/io_i_3_in1[2] cb_6_9/io_i_3_in1[3]
+ cb_6_9/io_i_3_in1[4] cb_6_9/io_i_3_in1[5] cb_6_9/io_i_3_in1[6] cb_6_9/io_i_3_in1[7]
+ cb_6_9/io_i_4_ci cb_6_9/io_i_4_in1[0] cb_6_9/io_i_4_in1[1] cb_6_9/io_i_4_in1[2]
+ cb_6_9/io_i_4_in1[3] cb_6_9/io_i_4_in1[4] cb_6_9/io_i_4_in1[5] cb_6_9/io_i_4_in1[6]
+ cb_6_9/io_i_4_in1[7] cb_6_9/io_i_5_ci cb_6_9/io_i_5_in1[0] cb_6_9/io_i_5_in1[1]
+ cb_6_9/io_i_5_in1[2] cb_6_9/io_i_5_in1[3] cb_6_9/io_i_5_in1[4] cb_6_9/io_i_5_in1[5]
+ cb_6_9/io_i_5_in1[6] cb_6_9/io_i_5_in1[7] cb_6_9/io_i_6_ci cb_6_9/io_i_6_in1[0]
+ cb_6_9/io_i_6_in1[1] cb_6_9/io_i_6_in1[2] cb_6_9/io_i_6_in1[3] cb_6_9/io_i_6_in1[4]
+ cb_6_9/io_i_6_in1[5] cb_6_9/io_i_6_in1[6] cb_6_9/io_i_6_in1[7] cb_6_9/io_i_7_ci
+ cb_6_9/io_i_7_in1[0] cb_6_9/io_i_7_in1[1] cb_6_9/io_i_7_in1[2] cb_6_9/io_i_7_in1[3]
+ cb_6_9/io_i_7_in1[4] cb_6_9/io_i_7_in1[5] cb_6_9/io_i_7_in1[6] cb_6_9/io_i_7_in1[7]
+ cb_6_8/io_vci cb_6_9/io_vci cb_6_8/io_vi cb_6_9/io_we_i cb_6_8/io_wo[0] cb_6_8/io_wo[10]
+ cb_6_8/io_wo[11] cb_6_8/io_wo[12] cb_6_8/io_wo[13] cb_6_8/io_wo[14] cb_6_8/io_wo[15]
+ cb_6_8/io_wo[16] cb_6_8/io_wo[17] cb_6_8/io_wo[18] cb_6_8/io_wo[19] cb_6_8/io_wo[1]
+ cb_6_8/io_wo[20] cb_6_8/io_wo[21] cb_6_8/io_wo[22] cb_6_8/io_wo[23] cb_6_8/io_wo[24]
+ cb_6_8/io_wo[25] cb_6_8/io_wo[26] cb_6_8/io_wo[27] cb_6_8/io_wo[28] cb_6_8/io_wo[29]
+ cb_6_8/io_wo[2] cb_6_8/io_wo[30] cb_6_8/io_wo[31] cb_6_8/io_wo[32] cb_6_8/io_wo[33]
+ cb_6_8/io_wo[34] cb_6_8/io_wo[35] cb_6_8/io_wo[36] cb_6_8/io_wo[37] cb_6_8/io_wo[38]
+ cb_6_8/io_wo[39] cb_6_8/io_wo[3] cb_6_8/io_wo[40] cb_6_8/io_wo[41] cb_6_8/io_wo[42]
+ cb_6_8/io_wo[43] cb_6_8/io_wo[44] cb_6_8/io_wo[45] cb_6_8/io_wo[46] cb_6_8/io_wo[47]
+ cb_6_8/io_wo[48] cb_6_8/io_wo[49] cb_6_8/io_wo[4] cb_6_8/io_wo[50] cb_6_8/io_wo[51]
+ cb_6_8/io_wo[52] cb_6_8/io_wo[53] cb_6_8/io_wo[54] cb_6_8/io_wo[55] cb_6_8/io_wo[56]
+ cb_6_8/io_wo[57] cb_6_8/io_wo[58] cb_6_8/io_wo[59] cb_6_8/io_wo[5] cb_6_8/io_wo[60]
+ cb_6_8/io_wo[61] cb_6_8/io_wo[62] cb_6_8/io_wo[63] cb_6_8/io_wo[6] cb_6_8/io_wo[7]
+ cb_6_8/io_wo[8] cb_6_8/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_4_5 cb_4_9/io_adr_i[0] cb_4_9/io_adr_i[1] cb_4_5/io_cs_i cb_4_9/io_dat_i[0] cb_4_9/io_dat_i[10]
+ cb_4_9/io_dat_i[11] cb_4_9/io_dat_i[12] cb_4_9/io_dat_i[13] cb_4_9/io_dat_i[14]
+ cb_4_9/io_dat_i[15] cb_4_9/io_dat_i[1] cb_4_9/io_dat_i[2] cb_4_9/io_dat_i[3] cb_4_9/io_dat_i[4]
+ cb_4_9/io_dat_i[5] cb_4_9/io_dat_i[6] cb_4_9/io_dat_i[7] cb_4_9/io_dat_i[8] cb_4_9/io_dat_i[9]
+ cb_4_5/io_dat_o[0] cb_4_5/io_dat_o[10] cb_4_5/io_dat_o[11] cb_4_5/io_dat_o[12] cb_4_5/io_dat_o[13]
+ cb_4_5/io_dat_o[14] cb_4_5/io_dat_o[15] cb_4_5/io_dat_o[1] cb_4_5/io_dat_o[2] cb_4_5/io_dat_o[3]
+ cb_4_5/io_dat_o[4] cb_4_5/io_dat_o[5] cb_4_5/io_dat_o[6] cb_4_5/io_dat_o[7] cb_4_5/io_dat_o[8]
+ cb_4_5/io_dat_o[9] cb_4_6/io_wo[0] cb_4_6/io_wo[10] cb_4_6/io_wo[11] cb_4_6/io_wo[12]
+ cb_4_6/io_wo[13] cb_4_6/io_wo[14] cb_4_6/io_wo[15] cb_4_6/io_wo[16] cb_4_6/io_wo[17]
+ cb_4_6/io_wo[18] cb_4_6/io_wo[19] cb_4_6/io_wo[1] cb_4_6/io_wo[20] cb_4_6/io_wo[21]
+ cb_4_6/io_wo[22] cb_4_6/io_wo[23] cb_4_6/io_wo[24] cb_4_6/io_wo[25] cb_4_6/io_wo[26]
+ cb_4_6/io_wo[27] cb_4_6/io_wo[28] cb_4_6/io_wo[29] cb_4_6/io_wo[2] cb_4_6/io_wo[30]
+ cb_4_6/io_wo[31] cb_4_6/io_wo[32] cb_4_6/io_wo[33] cb_4_6/io_wo[34] cb_4_6/io_wo[35]
+ cb_4_6/io_wo[36] cb_4_6/io_wo[37] cb_4_6/io_wo[38] cb_4_6/io_wo[39] cb_4_6/io_wo[3]
+ cb_4_6/io_wo[40] cb_4_6/io_wo[41] cb_4_6/io_wo[42] cb_4_6/io_wo[43] cb_4_6/io_wo[44]
+ cb_4_6/io_wo[45] cb_4_6/io_wo[46] cb_4_6/io_wo[47] cb_4_6/io_wo[48] cb_4_6/io_wo[49]
+ cb_4_6/io_wo[4] cb_4_6/io_wo[50] cb_4_6/io_wo[51] cb_4_6/io_wo[52] cb_4_6/io_wo[53]
+ cb_4_6/io_wo[54] cb_4_6/io_wo[55] cb_4_6/io_wo[56] cb_4_6/io_wo[57] cb_4_6/io_wo[58]
+ cb_4_6/io_wo[59] cb_4_6/io_wo[5] cb_4_6/io_wo[60] cb_4_6/io_wo[61] cb_4_6/io_wo[62]
+ cb_4_6/io_wo[63] cb_4_6/io_wo[6] cb_4_6/io_wo[7] cb_4_6/io_wo[8] cb_4_6/io_wo[9]
+ cb_4_5/io_i_0_ci cb_4_5/io_i_0_in1[0] cb_4_5/io_i_0_in1[1] cb_4_5/io_i_0_in1[2]
+ cb_4_5/io_i_0_in1[3] cb_4_5/io_i_0_in1[4] cb_4_5/io_i_0_in1[5] cb_4_5/io_i_0_in1[6]
+ cb_4_5/io_i_0_in1[7] cb_4_5/io_i_1_ci cb_4_5/io_i_1_in1[0] cb_4_5/io_i_1_in1[1]
+ cb_4_5/io_i_1_in1[2] cb_4_5/io_i_1_in1[3] cb_4_5/io_i_1_in1[4] cb_4_5/io_i_1_in1[5]
+ cb_4_5/io_i_1_in1[6] cb_4_5/io_i_1_in1[7] cb_4_5/io_i_2_ci cb_4_5/io_i_2_in1[0]
+ cb_4_5/io_i_2_in1[1] cb_4_5/io_i_2_in1[2] cb_4_5/io_i_2_in1[3] cb_4_5/io_i_2_in1[4]
+ cb_4_5/io_i_2_in1[5] cb_4_5/io_i_2_in1[6] cb_4_5/io_i_2_in1[7] cb_4_5/io_i_3_ci
+ cb_4_5/io_i_3_in1[0] cb_4_5/io_i_3_in1[1] cb_4_5/io_i_3_in1[2] cb_4_5/io_i_3_in1[3]
+ cb_4_5/io_i_3_in1[4] cb_4_5/io_i_3_in1[5] cb_4_5/io_i_3_in1[6] cb_4_5/io_i_3_in1[7]
+ cb_4_5/io_i_4_ci cb_4_5/io_i_4_in1[0] cb_4_5/io_i_4_in1[1] cb_4_5/io_i_4_in1[2]
+ cb_4_5/io_i_4_in1[3] cb_4_5/io_i_4_in1[4] cb_4_5/io_i_4_in1[5] cb_4_5/io_i_4_in1[6]
+ cb_4_5/io_i_4_in1[7] cb_4_5/io_i_5_ci cb_4_5/io_i_5_in1[0] cb_4_5/io_i_5_in1[1]
+ cb_4_5/io_i_5_in1[2] cb_4_5/io_i_5_in1[3] cb_4_5/io_i_5_in1[4] cb_4_5/io_i_5_in1[5]
+ cb_4_5/io_i_5_in1[6] cb_4_5/io_i_5_in1[7] cb_4_5/io_i_6_ci cb_4_5/io_i_6_in1[0]
+ cb_4_5/io_i_6_in1[1] cb_4_5/io_i_6_in1[2] cb_4_5/io_i_6_in1[3] cb_4_5/io_i_6_in1[4]
+ cb_4_5/io_i_6_in1[5] cb_4_5/io_i_6_in1[6] cb_4_5/io_i_6_in1[7] cb_4_5/io_i_7_ci
+ cb_4_5/io_i_7_in1[0] cb_4_5/io_i_7_in1[1] cb_4_5/io_i_7_in1[2] cb_4_5/io_i_7_in1[3]
+ cb_4_5/io_i_7_in1[4] cb_4_5/io_i_7_in1[5] cb_4_5/io_i_7_in1[6] cb_4_5/io_i_7_in1[7]
+ cb_4_6/io_i_0_ci cb_4_6/io_i_0_in1[0] cb_4_6/io_i_0_in1[1] cb_4_6/io_i_0_in1[2]
+ cb_4_6/io_i_0_in1[3] cb_4_6/io_i_0_in1[4] cb_4_6/io_i_0_in1[5] cb_4_6/io_i_0_in1[6]
+ cb_4_6/io_i_0_in1[7] cb_4_6/io_i_1_ci cb_4_6/io_i_1_in1[0] cb_4_6/io_i_1_in1[1]
+ cb_4_6/io_i_1_in1[2] cb_4_6/io_i_1_in1[3] cb_4_6/io_i_1_in1[4] cb_4_6/io_i_1_in1[5]
+ cb_4_6/io_i_1_in1[6] cb_4_6/io_i_1_in1[7] cb_4_6/io_i_2_ci cb_4_6/io_i_2_in1[0]
+ cb_4_6/io_i_2_in1[1] cb_4_6/io_i_2_in1[2] cb_4_6/io_i_2_in1[3] cb_4_6/io_i_2_in1[4]
+ cb_4_6/io_i_2_in1[5] cb_4_6/io_i_2_in1[6] cb_4_6/io_i_2_in1[7] cb_4_6/io_i_3_ci
+ cb_4_6/io_i_3_in1[0] cb_4_6/io_i_3_in1[1] cb_4_6/io_i_3_in1[2] cb_4_6/io_i_3_in1[3]
+ cb_4_6/io_i_3_in1[4] cb_4_6/io_i_3_in1[5] cb_4_6/io_i_3_in1[6] cb_4_6/io_i_3_in1[7]
+ cb_4_6/io_i_4_ci cb_4_6/io_i_4_in1[0] cb_4_6/io_i_4_in1[1] cb_4_6/io_i_4_in1[2]
+ cb_4_6/io_i_4_in1[3] cb_4_6/io_i_4_in1[4] cb_4_6/io_i_4_in1[5] cb_4_6/io_i_4_in1[6]
+ cb_4_6/io_i_4_in1[7] cb_4_6/io_i_5_ci cb_4_6/io_i_5_in1[0] cb_4_6/io_i_5_in1[1]
+ cb_4_6/io_i_5_in1[2] cb_4_6/io_i_5_in1[3] cb_4_6/io_i_5_in1[4] cb_4_6/io_i_5_in1[5]
+ cb_4_6/io_i_5_in1[6] cb_4_6/io_i_5_in1[7] cb_4_6/io_i_6_ci cb_4_6/io_i_6_in1[0]
+ cb_4_6/io_i_6_in1[1] cb_4_6/io_i_6_in1[2] cb_4_6/io_i_6_in1[3] cb_4_6/io_i_6_in1[4]
+ cb_4_6/io_i_6_in1[5] cb_4_6/io_i_6_in1[6] cb_4_6/io_i_6_in1[7] cb_4_6/io_i_7_ci
+ cb_4_6/io_i_7_in1[0] cb_4_6/io_i_7_in1[1] cb_4_6/io_i_7_in1[2] cb_4_6/io_i_7_in1[3]
+ cb_4_6/io_i_7_in1[4] cb_4_6/io_i_7_in1[5] cb_4_6/io_i_7_in1[6] cb_4_6/io_i_7_in1[7]
+ cb_4_5/io_vci cb_4_6/io_vci cb_4_5/io_vi cb_4_9/io_we_i cb_4_5/io_wo[0] cb_4_5/io_wo[10]
+ cb_4_5/io_wo[11] cb_4_5/io_wo[12] cb_4_5/io_wo[13] cb_4_5/io_wo[14] cb_4_5/io_wo[15]
+ cb_4_5/io_wo[16] cb_4_5/io_wo[17] cb_4_5/io_wo[18] cb_4_5/io_wo[19] cb_4_5/io_wo[1]
+ cb_4_5/io_wo[20] cb_4_5/io_wo[21] cb_4_5/io_wo[22] cb_4_5/io_wo[23] cb_4_5/io_wo[24]
+ cb_4_5/io_wo[25] cb_4_5/io_wo[26] cb_4_5/io_wo[27] cb_4_5/io_wo[28] cb_4_5/io_wo[29]
+ cb_4_5/io_wo[2] cb_4_5/io_wo[30] cb_4_5/io_wo[31] cb_4_5/io_wo[32] cb_4_5/io_wo[33]
+ cb_4_5/io_wo[34] cb_4_5/io_wo[35] cb_4_5/io_wo[36] cb_4_5/io_wo[37] cb_4_5/io_wo[38]
+ cb_4_5/io_wo[39] cb_4_5/io_wo[3] cb_4_5/io_wo[40] cb_4_5/io_wo[41] cb_4_5/io_wo[42]
+ cb_4_5/io_wo[43] cb_4_5/io_wo[44] cb_4_5/io_wo[45] cb_4_5/io_wo[46] cb_4_5/io_wo[47]
+ cb_4_5/io_wo[48] cb_4_5/io_wo[49] cb_4_5/io_wo[4] cb_4_5/io_wo[50] cb_4_5/io_wo[51]
+ cb_4_5/io_wo[52] cb_4_5/io_wo[53] cb_4_5/io_wo[54] cb_4_5/io_wo[55] cb_4_5/io_wo[56]
+ cb_4_5/io_wo[57] cb_4_5/io_wo[58] cb_4_5/io_wo[59] cb_4_5/io_wo[5] cb_4_5/io_wo[60]
+ cb_4_5/io_wo[61] cb_4_5/io_wo[62] cb_4_5/io_wo[63] cb_4_5/io_wo[6] cb_4_5/io_wo[7]
+ cb_4_5/io_wo[8] cb_4_5/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_2_2 cb_2_9/io_adr_i[0] cb_2_9/io_adr_i[1] cb_2_2/io_cs_i cb_2_9/io_dat_i[0] cb_2_9/io_dat_i[10]
+ cb_2_9/io_dat_i[11] cb_2_9/io_dat_i[12] cb_2_9/io_dat_i[13] cb_2_9/io_dat_i[14]
+ cb_2_9/io_dat_i[15] cb_2_9/io_dat_i[1] cb_2_9/io_dat_i[2] cb_2_9/io_dat_i[3] cb_2_9/io_dat_i[4]
+ cb_2_9/io_dat_i[5] cb_2_9/io_dat_i[6] cb_2_9/io_dat_i[7] cb_2_9/io_dat_i[8] cb_2_9/io_dat_i[9]
+ cb_2_2/io_dat_o[0] cb_2_2/io_dat_o[10] cb_2_2/io_dat_o[11] cb_2_2/io_dat_o[12] cb_2_2/io_dat_o[13]
+ cb_2_2/io_dat_o[14] cb_2_2/io_dat_o[15] cb_2_2/io_dat_o[1] cb_2_2/io_dat_o[2] cb_2_2/io_dat_o[3]
+ cb_2_2/io_dat_o[4] cb_2_2/io_dat_o[5] cb_2_2/io_dat_o[6] cb_2_2/io_dat_o[7] cb_2_2/io_dat_o[8]
+ cb_2_2/io_dat_o[9] cb_2_3/io_wo[0] cb_2_3/io_wo[10] cb_2_3/io_wo[11] cb_2_3/io_wo[12]
+ cb_2_3/io_wo[13] cb_2_3/io_wo[14] cb_2_3/io_wo[15] cb_2_3/io_wo[16] cb_2_3/io_wo[17]
+ cb_2_3/io_wo[18] cb_2_3/io_wo[19] cb_2_3/io_wo[1] cb_2_3/io_wo[20] cb_2_3/io_wo[21]
+ cb_2_3/io_wo[22] cb_2_3/io_wo[23] cb_2_3/io_wo[24] cb_2_3/io_wo[25] cb_2_3/io_wo[26]
+ cb_2_3/io_wo[27] cb_2_3/io_wo[28] cb_2_3/io_wo[29] cb_2_3/io_wo[2] cb_2_3/io_wo[30]
+ cb_2_3/io_wo[31] cb_2_3/io_wo[32] cb_2_3/io_wo[33] cb_2_3/io_wo[34] cb_2_3/io_wo[35]
+ cb_2_3/io_wo[36] cb_2_3/io_wo[37] cb_2_3/io_wo[38] cb_2_3/io_wo[39] cb_2_3/io_wo[3]
+ cb_2_3/io_wo[40] cb_2_3/io_wo[41] cb_2_3/io_wo[42] cb_2_3/io_wo[43] cb_2_3/io_wo[44]
+ cb_2_3/io_wo[45] cb_2_3/io_wo[46] cb_2_3/io_wo[47] cb_2_3/io_wo[48] cb_2_3/io_wo[49]
+ cb_2_3/io_wo[4] cb_2_3/io_wo[50] cb_2_3/io_wo[51] cb_2_3/io_wo[52] cb_2_3/io_wo[53]
+ cb_2_3/io_wo[54] cb_2_3/io_wo[55] cb_2_3/io_wo[56] cb_2_3/io_wo[57] cb_2_3/io_wo[58]
+ cb_2_3/io_wo[59] cb_2_3/io_wo[5] cb_2_3/io_wo[60] cb_2_3/io_wo[61] cb_2_3/io_wo[62]
+ cb_2_3/io_wo[63] cb_2_3/io_wo[6] cb_2_3/io_wo[7] cb_2_3/io_wo[8] cb_2_3/io_wo[9]
+ cb_2_2/io_i_0_ci cb_2_2/io_i_0_in1[0] cb_2_2/io_i_0_in1[1] cb_2_2/io_i_0_in1[2]
+ cb_2_2/io_i_0_in1[3] cb_2_2/io_i_0_in1[4] cb_2_2/io_i_0_in1[5] cb_2_2/io_i_0_in1[6]
+ cb_2_2/io_i_0_in1[7] cb_2_2/io_i_1_ci cb_2_2/io_i_1_in1[0] cb_2_2/io_i_1_in1[1]
+ cb_2_2/io_i_1_in1[2] cb_2_2/io_i_1_in1[3] cb_2_2/io_i_1_in1[4] cb_2_2/io_i_1_in1[5]
+ cb_2_2/io_i_1_in1[6] cb_2_2/io_i_1_in1[7] cb_2_2/io_i_2_ci cb_2_2/io_i_2_in1[0]
+ cb_2_2/io_i_2_in1[1] cb_2_2/io_i_2_in1[2] cb_2_2/io_i_2_in1[3] cb_2_2/io_i_2_in1[4]
+ cb_2_2/io_i_2_in1[5] cb_2_2/io_i_2_in1[6] cb_2_2/io_i_2_in1[7] cb_2_2/io_i_3_ci
+ cb_2_2/io_i_3_in1[0] cb_2_2/io_i_3_in1[1] cb_2_2/io_i_3_in1[2] cb_2_2/io_i_3_in1[3]
+ cb_2_2/io_i_3_in1[4] cb_2_2/io_i_3_in1[5] cb_2_2/io_i_3_in1[6] cb_2_2/io_i_3_in1[7]
+ cb_2_2/io_i_4_ci cb_2_2/io_i_4_in1[0] cb_2_2/io_i_4_in1[1] cb_2_2/io_i_4_in1[2]
+ cb_2_2/io_i_4_in1[3] cb_2_2/io_i_4_in1[4] cb_2_2/io_i_4_in1[5] cb_2_2/io_i_4_in1[6]
+ cb_2_2/io_i_4_in1[7] cb_2_2/io_i_5_ci cb_2_2/io_i_5_in1[0] cb_2_2/io_i_5_in1[1]
+ cb_2_2/io_i_5_in1[2] cb_2_2/io_i_5_in1[3] cb_2_2/io_i_5_in1[4] cb_2_2/io_i_5_in1[5]
+ cb_2_2/io_i_5_in1[6] cb_2_2/io_i_5_in1[7] cb_2_2/io_i_6_ci cb_2_2/io_i_6_in1[0]
+ cb_2_2/io_i_6_in1[1] cb_2_2/io_i_6_in1[2] cb_2_2/io_i_6_in1[3] cb_2_2/io_i_6_in1[4]
+ cb_2_2/io_i_6_in1[5] cb_2_2/io_i_6_in1[6] cb_2_2/io_i_6_in1[7] cb_2_2/io_i_7_ci
+ cb_2_2/io_i_7_in1[0] cb_2_2/io_i_7_in1[1] cb_2_2/io_i_7_in1[2] cb_2_2/io_i_7_in1[3]
+ cb_2_2/io_i_7_in1[4] cb_2_2/io_i_7_in1[5] cb_2_2/io_i_7_in1[6] cb_2_2/io_i_7_in1[7]
+ cb_2_3/io_i_0_ci cb_2_3/io_i_0_in1[0] cb_2_3/io_i_0_in1[1] cb_2_3/io_i_0_in1[2]
+ cb_2_3/io_i_0_in1[3] cb_2_3/io_i_0_in1[4] cb_2_3/io_i_0_in1[5] cb_2_3/io_i_0_in1[6]
+ cb_2_3/io_i_0_in1[7] cb_2_3/io_i_1_ci cb_2_3/io_i_1_in1[0] cb_2_3/io_i_1_in1[1]
+ cb_2_3/io_i_1_in1[2] cb_2_3/io_i_1_in1[3] cb_2_3/io_i_1_in1[4] cb_2_3/io_i_1_in1[5]
+ cb_2_3/io_i_1_in1[6] cb_2_3/io_i_1_in1[7] cb_2_3/io_i_2_ci cb_2_3/io_i_2_in1[0]
+ cb_2_3/io_i_2_in1[1] cb_2_3/io_i_2_in1[2] cb_2_3/io_i_2_in1[3] cb_2_3/io_i_2_in1[4]
+ cb_2_3/io_i_2_in1[5] cb_2_3/io_i_2_in1[6] cb_2_3/io_i_2_in1[7] cb_2_3/io_i_3_ci
+ cb_2_3/io_i_3_in1[0] cb_2_3/io_i_3_in1[1] cb_2_3/io_i_3_in1[2] cb_2_3/io_i_3_in1[3]
+ cb_2_3/io_i_3_in1[4] cb_2_3/io_i_3_in1[5] cb_2_3/io_i_3_in1[6] cb_2_3/io_i_3_in1[7]
+ cb_2_3/io_i_4_ci cb_2_3/io_i_4_in1[0] cb_2_3/io_i_4_in1[1] cb_2_3/io_i_4_in1[2]
+ cb_2_3/io_i_4_in1[3] cb_2_3/io_i_4_in1[4] cb_2_3/io_i_4_in1[5] cb_2_3/io_i_4_in1[6]
+ cb_2_3/io_i_4_in1[7] cb_2_3/io_i_5_ci cb_2_3/io_i_5_in1[0] cb_2_3/io_i_5_in1[1]
+ cb_2_3/io_i_5_in1[2] cb_2_3/io_i_5_in1[3] cb_2_3/io_i_5_in1[4] cb_2_3/io_i_5_in1[5]
+ cb_2_3/io_i_5_in1[6] cb_2_3/io_i_5_in1[7] cb_2_3/io_i_6_ci cb_2_3/io_i_6_in1[0]
+ cb_2_3/io_i_6_in1[1] cb_2_3/io_i_6_in1[2] cb_2_3/io_i_6_in1[3] cb_2_3/io_i_6_in1[4]
+ cb_2_3/io_i_6_in1[5] cb_2_3/io_i_6_in1[6] cb_2_3/io_i_6_in1[7] cb_2_3/io_i_7_ci
+ cb_2_3/io_i_7_in1[0] cb_2_3/io_i_7_in1[1] cb_2_3/io_i_7_in1[2] cb_2_3/io_i_7_in1[3]
+ cb_2_3/io_i_7_in1[4] cb_2_3/io_i_7_in1[5] cb_2_3/io_i_7_in1[6] cb_2_3/io_i_7_in1[7]
+ cb_2_2/io_vci cb_2_3/io_vci cb_2_2/io_vi cb_2_9/io_we_i cb_2_2/io_wo[0] cb_2_2/io_wo[10]
+ cb_2_2/io_wo[11] cb_2_2/io_wo[12] cb_2_2/io_wo[13] cb_2_2/io_wo[14] cb_2_2/io_wo[15]
+ cb_2_2/io_wo[16] cb_2_2/io_wo[17] cb_2_2/io_wo[18] cb_2_2/io_wo[19] cb_2_2/io_wo[1]
+ cb_2_2/io_wo[20] cb_2_2/io_wo[21] cb_2_2/io_wo[22] cb_2_2/io_wo[23] cb_2_2/io_wo[24]
+ cb_2_2/io_wo[25] cb_2_2/io_wo[26] cb_2_2/io_wo[27] cb_2_2/io_wo[28] cb_2_2/io_wo[29]
+ cb_2_2/io_wo[2] cb_2_2/io_wo[30] cb_2_2/io_wo[31] cb_2_2/io_wo[32] cb_2_2/io_wo[33]
+ cb_2_2/io_wo[34] cb_2_2/io_wo[35] cb_2_2/io_wo[36] cb_2_2/io_wo[37] cb_2_2/io_wo[38]
+ cb_2_2/io_wo[39] cb_2_2/io_wo[3] cb_2_2/io_wo[40] cb_2_2/io_wo[41] cb_2_2/io_wo[42]
+ cb_2_2/io_wo[43] cb_2_2/io_wo[44] cb_2_2/io_wo[45] cb_2_2/io_wo[46] cb_2_2/io_wo[47]
+ cb_2_2/io_wo[48] cb_2_2/io_wo[49] cb_2_2/io_wo[4] cb_2_2/io_wo[50] cb_2_2/io_wo[51]
+ cb_2_2/io_wo[52] cb_2_2/io_wo[53] cb_2_2/io_wo[54] cb_2_2/io_wo[55] cb_2_2/io_wo[56]
+ cb_2_2/io_wo[57] cb_2_2/io_wo[58] cb_2_2/io_wo[59] cb_2_2/io_wo[5] cb_2_2/io_wo[60]
+ cb_2_2/io_wo[61] cb_2_2/io_wo[62] cb_2_2/io_wo[63] cb_2_2/io_wo[6] cb_2_2/io_wo[7]
+ cb_2_2/io_wo[8] cb_2_2/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_6_9 cb_6_9/io_adr_i[0] cb_6_9/io_adr_i[1] cb_6_9/io_cs_i cb_6_9/io_dat_i[0] cb_6_9/io_dat_i[10]
+ cb_6_9/io_dat_i[11] cb_6_9/io_dat_i[12] cb_6_9/io_dat_i[13] cb_6_9/io_dat_i[14]
+ cb_6_9/io_dat_i[15] cb_6_9/io_dat_i[1] cb_6_9/io_dat_i[2] cb_6_9/io_dat_i[3] cb_6_9/io_dat_i[4]
+ cb_6_9/io_dat_i[5] cb_6_9/io_dat_i[6] cb_6_9/io_dat_i[7] cb_6_9/io_dat_i[8] cb_6_9/io_dat_i[9]
+ cb_6_9/io_dat_o[0] cb_6_9/io_dat_o[10] cb_6_9/io_dat_o[11] cb_6_9/io_dat_o[12] cb_6_9/io_dat_o[13]
+ cb_6_9/io_dat_o[14] cb_6_9/io_dat_o[15] cb_6_9/io_dat_o[1] cb_6_9/io_dat_o[2] cb_6_9/io_dat_o[3]
+ cb_6_9/io_dat_o[4] cb_6_9/io_dat_o[5] cb_6_9/io_dat_o[6] cb_6_9/io_dat_o[7] cb_6_9/io_dat_o[8]
+ cb_6_9/io_dat_o[9] cb_6_9/io_eo[0] cb_6_9/io_eo[10] cb_6_9/io_eo[11] cb_6_9/io_eo[12]
+ cb_6_9/io_eo[13] cb_6_9/io_eo[14] cb_6_9/io_eo[15] cb_6_9/io_eo[16] cb_6_9/io_eo[17]
+ cb_6_9/io_eo[18] cb_6_9/io_eo[19] cb_6_9/io_eo[1] cb_6_9/io_eo[20] cb_6_9/io_eo[21]
+ cb_6_9/io_eo[22] cb_6_9/io_eo[23] cb_6_9/io_eo[24] cb_6_9/io_eo[25] cb_6_9/io_eo[26]
+ cb_6_9/io_eo[27] cb_6_9/io_eo[28] cb_6_9/io_eo[29] cb_6_9/io_eo[2] cb_6_9/io_eo[30]
+ cb_6_9/io_eo[31] cb_6_9/io_eo[32] cb_6_9/io_eo[33] cb_6_9/io_eo[34] cb_6_9/io_eo[35]
+ cb_6_9/io_eo[36] cb_6_9/io_eo[37] cb_6_9/io_eo[38] cb_6_9/io_eo[39] cb_6_9/io_eo[3]
+ cb_6_9/io_eo[40] cb_6_9/io_eo[41] cb_6_9/io_eo[42] cb_6_9/io_eo[43] cb_6_9/io_eo[44]
+ cb_6_9/io_eo[45] cb_6_9/io_eo[46] cb_6_9/io_eo[47] cb_6_9/io_eo[48] cb_6_9/io_eo[49]
+ cb_6_9/io_eo[4] cb_6_9/io_eo[50] cb_6_9/io_eo[51] cb_6_9/io_eo[52] cb_6_9/io_eo[53]
+ cb_6_9/io_eo[54] cb_6_9/io_eo[55] cb_6_9/io_eo[56] cb_6_9/io_eo[57] cb_6_9/io_eo[58]
+ cb_6_9/io_eo[59] cb_6_9/io_eo[5] cb_6_9/io_eo[60] cb_6_9/io_eo[61] cb_6_9/io_eo[62]
+ cb_6_9/io_eo[63] cb_6_9/io_eo[6] cb_6_9/io_eo[7] cb_6_9/io_eo[8] cb_6_9/io_eo[9]
+ cb_6_9/io_i_0_ci cb_6_9/io_i_0_in1[0] cb_6_9/io_i_0_in1[1] cb_6_9/io_i_0_in1[2]
+ cb_6_9/io_i_0_in1[3] cb_6_9/io_i_0_in1[4] cb_6_9/io_i_0_in1[5] cb_6_9/io_i_0_in1[6]
+ cb_6_9/io_i_0_in1[7] cb_6_9/io_i_1_ci cb_6_9/io_i_1_in1[0] cb_6_9/io_i_1_in1[1]
+ cb_6_9/io_i_1_in1[2] cb_6_9/io_i_1_in1[3] cb_6_9/io_i_1_in1[4] cb_6_9/io_i_1_in1[5]
+ cb_6_9/io_i_1_in1[6] cb_6_9/io_i_1_in1[7] cb_6_9/io_i_2_ci cb_6_9/io_i_2_in1[0]
+ cb_6_9/io_i_2_in1[1] cb_6_9/io_i_2_in1[2] cb_6_9/io_i_2_in1[3] cb_6_9/io_i_2_in1[4]
+ cb_6_9/io_i_2_in1[5] cb_6_9/io_i_2_in1[6] cb_6_9/io_i_2_in1[7] cb_6_9/io_i_3_ci
+ cb_6_9/io_i_3_in1[0] cb_6_9/io_i_3_in1[1] cb_6_9/io_i_3_in1[2] cb_6_9/io_i_3_in1[3]
+ cb_6_9/io_i_3_in1[4] cb_6_9/io_i_3_in1[5] cb_6_9/io_i_3_in1[6] cb_6_9/io_i_3_in1[7]
+ cb_6_9/io_i_4_ci cb_6_9/io_i_4_in1[0] cb_6_9/io_i_4_in1[1] cb_6_9/io_i_4_in1[2]
+ cb_6_9/io_i_4_in1[3] cb_6_9/io_i_4_in1[4] cb_6_9/io_i_4_in1[5] cb_6_9/io_i_4_in1[6]
+ cb_6_9/io_i_4_in1[7] cb_6_9/io_i_5_ci cb_6_9/io_i_5_in1[0] cb_6_9/io_i_5_in1[1]
+ cb_6_9/io_i_5_in1[2] cb_6_9/io_i_5_in1[3] cb_6_9/io_i_5_in1[4] cb_6_9/io_i_5_in1[5]
+ cb_6_9/io_i_5_in1[6] cb_6_9/io_i_5_in1[7] cb_6_9/io_i_6_ci cb_6_9/io_i_6_in1[0]
+ cb_6_9/io_i_6_in1[1] cb_6_9/io_i_6_in1[2] cb_6_9/io_i_6_in1[3] cb_6_9/io_i_6_in1[4]
+ cb_6_9/io_i_6_in1[5] cb_6_9/io_i_6_in1[6] cb_6_9/io_i_6_in1[7] cb_6_9/io_i_7_ci
+ cb_6_9/io_i_7_in1[0] cb_6_9/io_i_7_in1[1] cb_6_9/io_i_7_in1[2] cb_6_9/io_i_7_in1[3]
+ cb_6_9/io_i_7_in1[4] cb_6_9/io_i_7_in1[5] cb_6_9/io_i_7_in1[6] cb_6_9/io_i_7_in1[7]
+ cb_6_9/io_o_0_co cb_6_9/io_o_0_out[0] cb_6_9/io_o_0_out[1] cb_6_9/io_o_0_out[2]
+ cb_6_9/io_o_0_out[3] cb_6_9/io_o_0_out[4] cb_6_9/io_o_0_out[5] cb_6_9/io_o_0_out[6]
+ cb_6_9/io_o_0_out[7] cb_6_9/io_o_1_co cb_6_9/io_o_1_out[0] cb_6_9/io_o_1_out[1]
+ cb_6_9/io_o_1_out[2] cb_6_9/io_o_1_out[3] cb_6_9/io_o_1_out[4] cb_6_9/io_o_1_out[5]
+ cb_6_9/io_o_1_out[6] cb_6_9/io_o_1_out[7] cb_6_9/io_o_2_co cb_6_9/io_o_2_out[0]
+ cb_6_9/io_o_2_out[1] cb_6_9/io_o_2_out[2] cb_6_9/io_o_2_out[3] cb_6_9/io_o_2_out[4]
+ cb_6_9/io_o_2_out[5] cb_6_9/io_o_2_out[6] cb_6_9/io_o_2_out[7] cb_6_9/io_o_3_co
+ cb_6_9/io_o_3_out[0] cb_6_9/io_o_3_out[1] cb_6_9/io_o_3_out[2] cb_6_9/io_o_3_out[3]
+ cb_6_9/io_o_3_out[4] cb_6_9/io_o_3_out[5] cb_6_9/io_o_3_out[6] cb_6_9/io_o_3_out[7]
+ cb_6_9/io_o_4_co cb_6_9/io_o_4_out[0] cb_6_9/io_o_4_out[1] cb_6_9/io_o_4_out[2]
+ cb_6_9/io_o_4_out[3] cb_6_9/io_o_4_out[4] cb_6_9/io_o_4_out[5] cb_6_9/io_o_4_out[6]
+ cb_6_9/io_o_4_out[7] cb_6_9/io_o_5_co cb_6_9/io_o_5_out[0] cb_6_9/io_o_5_out[1]
+ cb_6_9/io_o_5_out[2] cb_6_9/io_o_5_out[3] cb_6_9/io_o_5_out[4] cb_6_9/io_o_5_out[5]
+ cb_6_9/io_o_5_out[6] cb_6_9/io_o_5_out[7] cb_6_9/io_o_6_co cb_6_9/io_o_6_out[0]
+ cb_6_9/io_o_6_out[1] cb_6_9/io_o_6_out[2] cb_6_9/io_o_6_out[3] cb_6_9/io_o_6_out[4]
+ cb_6_9/io_o_6_out[5] cb_6_9/io_o_6_out[6] cb_6_9/io_o_6_out[7] cb_6_9/io_o_7_co
+ cb_6_9/io_o_7_out[0] cb_6_9/io_o_7_out[1] cb_6_9/io_o_7_out[2] cb_6_9/io_o_7_out[3]
+ cb_6_9/io_o_7_out[4] cb_6_9/io_o_7_out[5] cb_6_9/io_o_7_out[6] cb_6_9/io_o_7_out[7]
+ cb_6_9/io_vci cb_6_9/io_vco cb_6_9/io_vi cb_6_9/io_we_i cb_6_9/io_wo[0] cb_6_9/io_wo[10]
+ cb_6_9/io_wo[11] cb_6_9/io_wo[12] cb_6_9/io_wo[13] cb_6_9/io_wo[14] cb_6_9/io_wo[15]
+ cb_6_9/io_wo[16] cb_6_9/io_wo[17] cb_6_9/io_wo[18] cb_6_9/io_wo[19] cb_6_9/io_wo[1]
+ cb_6_9/io_wo[20] cb_6_9/io_wo[21] cb_6_9/io_wo[22] cb_6_9/io_wo[23] cb_6_9/io_wo[24]
+ cb_6_9/io_wo[25] cb_6_9/io_wo[26] cb_6_9/io_wo[27] cb_6_9/io_wo[28] cb_6_9/io_wo[29]
+ cb_6_9/io_wo[2] cb_6_9/io_wo[30] cb_6_9/io_wo[31] cb_6_9/io_wo[32] cb_6_9/io_wo[33]
+ cb_6_9/io_wo[34] cb_6_9/io_wo[35] cb_6_9/io_wo[36] cb_6_9/io_wo[37] cb_6_9/io_wo[38]
+ cb_6_9/io_wo[39] cb_6_9/io_wo[3] cb_6_9/io_wo[40] cb_6_9/io_wo[41] cb_6_9/io_wo[42]
+ cb_6_9/io_wo[43] cb_6_9/io_wo[44] cb_6_9/io_wo[45] cb_6_9/io_wo[46] cb_6_9/io_wo[47]
+ cb_6_9/io_wo[48] cb_6_9/io_wo[49] cb_6_9/io_wo[4] cb_6_9/io_wo[50] cb_6_9/io_wo[51]
+ cb_6_9/io_wo[52] cb_6_9/io_wo[53] cb_6_9/io_wo[54] cb_6_9/io_wo[55] cb_6_9/io_wo[56]
+ cb_6_9/io_wo[57] cb_6_9/io_wo[58] cb_6_9/io_wo[59] cb_6_9/io_wo[5] cb_6_9/io_wo[60]
+ cb_6_9/io_wo[61] cb_6_9/io_wo[62] cb_6_9/io_wo[63] cb_6_9/io_wo[6] cb_6_9/io_wo[7]
+ cb_6_9/io_wo[8] cb_6_9/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_4_6 cb_4_9/io_adr_i[0] cb_4_9/io_adr_i[1] cb_4_6/io_cs_i cb_4_9/io_dat_i[0] cb_4_9/io_dat_i[10]
+ cb_4_9/io_dat_i[11] cb_4_9/io_dat_i[12] cb_4_9/io_dat_i[13] cb_4_9/io_dat_i[14]
+ cb_4_9/io_dat_i[15] cb_4_9/io_dat_i[1] cb_4_9/io_dat_i[2] cb_4_9/io_dat_i[3] cb_4_9/io_dat_i[4]
+ cb_4_9/io_dat_i[5] cb_4_9/io_dat_i[6] cb_4_9/io_dat_i[7] cb_4_9/io_dat_i[8] cb_4_9/io_dat_i[9]
+ cb_4_6/io_dat_o[0] cb_4_6/io_dat_o[10] cb_4_6/io_dat_o[11] cb_4_6/io_dat_o[12] cb_4_6/io_dat_o[13]
+ cb_4_6/io_dat_o[14] cb_4_6/io_dat_o[15] cb_4_6/io_dat_o[1] cb_4_6/io_dat_o[2] cb_4_6/io_dat_o[3]
+ cb_4_6/io_dat_o[4] cb_4_6/io_dat_o[5] cb_4_6/io_dat_o[6] cb_4_6/io_dat_o[7] cb_4_6/io_dat_o[8]
+ cb_4_6/io_dat_o[9] cb_4_7/io_wo[0] cb_4_7/io_wo[10] cb_4_7/io_wo[11] cb_4_7/io_wo[12]
+ cb_4_7/io_wo[13] cb_4_7/io_wo[14] cb_4_7/io_wo[15] cb_4_7/io_wo[16] cb_4_7/io_wo[17]
+ cb_4_7/io_wo[18] cb_4_7/io_wo[19] cb_4_7/io_wo[1] cb_4_7/io_wo[20] cb_4_7/io_wo[21]
+ cb_4_7/io_wo[22] cb_4_7/io_wo[23] cb_4_7/io_wo[24] cb_4_7/io_wo[25] cb_4_7/io_wo[26]
+ cb_4_7/io_wo[27] cb_4_7/io_wo[28] cb_4_7/io_wo[29] cb_4_7/io_wo[2] cb_4_7/io_wo[30]
+ cb_4_7/io_wo[31] cb_4_7/io_wo[32] cb_4_7/io_wo[33] cb_4_7/io_wo[34] cb_4_7/io_wo[35]
+ cb_4_7/io_wo[36] cb_4_7/io_wo[37] cb_4_7/io_wo[38] cb_4_7/io_wo[39] cb_4_7/io_wo[3]
+ cb_4_7/io_wo[40] cb_4_7/io_wo[41] cb_4_7/io_wo[42] cb_4_7/io_wo[43] cb_4_7/io_wo[44]
+ cb_4_7/io_wo[45] cb_4_7/io_wo[46] cb_4_7/io_wo[47] cb_4_7/io_wo[48] cb_4_7/io_wo[49]
+ cb_4_7/io_wo[4] cb_4_7/io_wo[50] cb_4_7/io_wo[51] cb_4_7/io_wo[52] cb_4_7/io_wo[53]
+ cb_4_7/io_wo[54] cb_4_7/io_wo[55] cb_4_7/io_wo[56] cb_4_7/io_wo[57] cb_4_7/io_wo[58]
+ cb_4_7/io_wo[59] cb_4_7/io_wo[5] cb_4_7/io_wo[60] cb_4_7/io_wo[61] cb_4_7/io_wo[62]
+ cb_4_7/io_wo[63] cb_4_7/io_wo[6] cb_4_7/io_wo[7] cb_4_7/io_wo[8] cb_4_7/io_wo[9]
+ cb_4_6/io_i_0_ci cb_4_6/io_i_0_in1[0] cb_4_6/io_i_0_in1[1] cb_4_6/io_i_0_in1[2]
+ cb_4_6/io_i_0_in1[3] cb_4_6/io_i_0_in1[4] cb_4_6/io_i_0_in1[5] cb_4_6/io_i_0_in1[6]
+ cb_4_6/io_i_0_in1[7] cb_4_6/io_i_1_ci cb_4_6/io_i_1_in1[0] cb_4_6/io_i_1_in1[1]
+ cb_4_6/io_i_1_in1[2] cb_4_6/io_i_1_in1[3] cb_4_6/io_i_1_in1[4] cb_4_6/io_i_1_in1[5]
+ cb_4_6/io_i_1_in1[6] cb_4_6/io_i_1_in1[7] cb_4_6/io_i_2_ci cb_4_6/io_i_2_in1[0]
+ cb_4_6/io_i_2_in1[1] cb_4_6/io_i_2_in1[2] cb_4_6/io_i_2_in1[3] cb_4_6/io_i_2_in1[4]
+ cb_4_6/io_i_2_in1[5] cb_4_6/io_i_2_in1[6] cb_4_6/io_i_2_in1[7] cb_4_6/io_i_3_ci
+ cb_4_6/io_i_3_in1[0] cb_4_6/io_i_3_in1[1] cb_4_6/io_i_3_in1[2] cb_4_6/io_i_3_in1[3]
+ cb_4_6/io_i_3_in1[4] cb_4_6/io_i_3_in1[5] cb_4_6/io_i_3_in1[6] cb_4_6/io_i_3_in1[7]
+ cb_4_6/io_i_4_ci cb_4_6/io_i_4_in1[0] cb_4_6/io_i_4_in1[1] cb_4_6/io_i_4_in1[2]
+ cb_4_6/io_i_4_in1[3] cb_4_6/io_i_4_in1[4] cb_4_6/io_i_4_in1[5] cb_4_6/io_i_4_in1[6]
+ cb_4_6/io_i_4_in1[7] cb_4_6/io_i_5_ci cb_4_6/io_i_5_in1[0] cb_4_6/io_i_5_in1[1]
+ cb_4_6/io_i_5_in1[2] cb_4_6/io_i_5_in1[3] cb_4_6/io_i_5_in1[4] cb_4_6/io_i_5_in1[5]
+ cb_4_6/io_i_5_in1[6] cb_4_6/io_i_5_in1[7] cb_4_6/io_i_6_ci cb_4_6/io_i_6_in1[0]
+ cb_4_6/io_i_6_in1[1] cb_4_6/io_i_6_in1[2] cb_4_6/io_i_6_in1[3] cb_4_6/io_i_6_in1[4]
+ cb_4_6/io_i_6_in1[5] cb_4_6/io_i_6_in1[6] cb_4_6/io_i_6_in1[7] cb_4_6/io_i_7_ci
+ cb_4_6/io_i_7_in1[0] cb_4_6/io_i_7_in1[1] cb_4_6/io_i_7_in1[2] cb_4_6/io_i_7_in1[3]
+ cb_4_6/io_i_7_in1[4] cb_4_6/io_i_7_in1[5] cb_4_6/io_i_7_in1[6] cb_4_6/io_i_7_in1[7]
+ cb_4_7/io_i_0_ci cb_4_7/io_i_0_in1[0] cb_4_7/io_i_0_in1[1] cb_4_7/io_i_0_in1[2]
+ cb_4_7/io_i_0_in1[3] cb_4_7/io_i_0_in1[4] cb_4_7/io_i_0_in1[5] cb_4_7/io_i_0_in1[6]
+ cb_4_7/io_i_0_in1[7] cb_4_7/io_i_1_ci cb_4_7/io_i_1_in1[0] cb_4_7/io_i_1_in1[1]
+ cb_4_7/io_i_1_in1[2] cb_4_7/io_i_1_in1[3] cb_4_7/io_i_1_in1[4] cb_4_7/io_i_1_in1[5]
+ cb_4_7/io_i_1_in1[6] cb_4_7/io_i_1_in1[7] cb_4_7/io_i_2_ci cb_4_7/io_i_2_in1[0]
+ cb_4_7/io_i_2_in1[1] cb_4_7/io_i_2_in1[2] cb_4_7/io_i_2_in1[3] cb_4_7/io_i_2_in1[4]
+ cb_4_7/io_i_2_in1[5] cb_4_7/io_i_2_in1[6] cb_4_7/io_i_2_in1[7] cb_4_7/io_i_3_ci
+ cb_4_7/io_i_3_in1[0] cb_4_7/io_i_3_in1[1] cb_4_7/io_i_3_in1[2] cb_4_7/io_i_3_in1[3]
+ cb_4_7/io_i_3_in1[4] cb_4_7/io_i_3_in1[5] cb_4_7/io_i_3_in1[6] cb_4_7/io_i_3_in1[7]
+ cb_4_7/io_i_4_ci cb_4_7/io_i_4_in1[0] cb_4_7/io_i_4_in1[1] cb_4_7/io_i_4_in1[2]
+ cb_4_7/io_i_4_in1[3] cb_4_7/io_i_4_in1[4] cb_4_7/io_i_4_in1[5] cb_4_7/io_i_4_in1[6]
+ cb_4_7/io_i_4_in1[7] cb_4_7/io_i_5_ci cb_4_7/io_i_5_in1[0] cb_4_7/io_i_5_in1[1]
+ cb_4_7/io_i_5_in1[2] cb_4_7/io_i_5_in1[3] cb_4_7/io_i_5_in1[4] cb_4_7/io_i_5_in1[5]
+ cb_4_7/io_i_5_in1[6] cb_4_7/io_i_5_in1[7] cb_4_7/io_i_6_ci cb_4_7/io_i_6_in1[0]
+ cb_4_7/io_i_6_in1[1] cb_4_7/io_i_6_in1[2] cb_4_7/io_i_6_in1[3] cb_4_7/io_i_6_in1[4]
+ cb_4_7/io_i_6_in1[5] cb_4_7/io_i_6_in1[6] cb_4_7/io_i_6_in1[7] cb_4_7/io_i_7_ci
+ cb_4_7/io_i_7_in1[0] cb_4_7/io_i_7_in1[1] cb_4_7/io_i_7_in1[2] cb_4_7/io_i_7_in1[3]
+ cb_4_7/io_i_7_in1[4] cb_4_7/io_i_7_in1[5] cb_4_7/io_i_7_in1[6] cb_4_7/io_i_7_in1[7]
+ cb_4_6/io_vci cb_4_7/io_vci cb_4_6/io_vi cb_4_9/io_we_i cb_4_6/io_wo[0] cb_4_6/io_wo[10]
+ cb_4_6/io_wo[11] cb_4_6/io_wo[12] cb_4_6/io_wo[13] cb_4_6/io_wo[14] cb_4_6/io_wo[15]
+ cb_4_6/io_wo[16] cb_4_6/io_wo[17] cb_4_6/io_wo[18] cb_4_6/io_wo[19] cb_4_6/io_wo[1]
+ cb_4_6/io_wo[20] cb_4_6/io_wo[21] cb_4_6/io_wo[22] cb_4_6/io_wo[23] cb_4_6/io_wo[24]
+ cb_4_6/io_wo[25] cb_4_6/io_wo[26] cb_4_6/io_wo[27] cb_4_6/io_wo[28] cb_4_6/io_wo[29]
+ cb_4_6/io_wo[2] cb_4_6/io_wo[30] cb_4_6/io_wo[31] cb_4_6/io_wo[32] cb_4_6/io_wo[33]
+ cb_4_6/io_wo[34] cb_4_6/io_wo[35] cb_4_6/io_wo[36] cb_4_6/io_wo[37] cb_4_6/io_wo[38]
+ cb_4_6/io_wo[39] cb_4_6/io_wo[3] cb_4_6/io_wo[40] cb_4_6/io_wo[41] cb_4_6/io_wo[42]
+ cb_4_6/io_wo[43] cb_4_6/io_wo[44] cb_4_6/io_wo[45] cb_4_6/io_wo[46] cb_4_6/io_wo[47]
+ cb_4_6/io_wo[48] cb_4_6/io_wo[49] cb_4_6/io_wo[4] cb_4_6/io_wo[50] cb_4_6/io_wo[51]
+ cb_4_6/io_wo[52] cb_4_6/io_wo[53] cb_4_6/io_wo[54] cb_4_6/io_wo[55] cb_4_6/io_wo[56]
+ cb_4_6/io_wo[57] cb_4_6/io_wo[58] cb_4_6/io_wo[59] cb_4_6/io_wo[5] cb_4_6/io_wo[60]
+ cb_4_6/io_wo[61] cb_4_6/io_wo[62] cb_4_6/io_wo[63] cb_4_6/io_wo[6] cb_4_6/io_wo[7]
+ cb_4_6/io_wo[8] cb_4_6/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_2_3 cb_2_9/io_adr_i[0] cb_2_9/io_adr_i[1] cb_2_3/io_cs_i cb_2_9/io_dat_i[0] cb_2_9/io_dat_i[10]
+ cb_2_9/io_dat_i[11] cb_2_9/io_dat_i[12] cb_2_9/io_dat_i[13] cb_2_9/io_dat_i[14]
+ cb_2_9/io_dat_i[15] cb_2_9/io_dat_i[1] cb_2_9/io_dat_i[2] cb_2_9/io_dat_i[3] cb_2_9/io_dat_i[4]
+ cb_2_9/io_dat_i[5] cb_2_9/io_dat_i[6] cb_2_9/io_dat_i[7] cb_2_9/io_dat_i[8] cb_2_9/io_dat_i[9]
+ cb_2_3/io_dat_o[0] cb_2_3/io_dat_o[10] cb_2_3/io_dat_o[11] cb_2_3/io_dat_o[12] cb_2_3/io_dat_o[13]
+ cb_2_3/io_dat_o[14] cb_2_3/io_dat_o[15] cb_2_3/io_dat_o[1] cb_2_3/io_dat_o[2] cb_2_3/io_dat_o[3]
+ cb_2_3/io_dat_o[4] cb_2_3/io_dat_o[5] cb_2_3/io_dat_o[6] cb_2_3/io_dat_o[7] cb_2_3/io_dat_o[8]
+ cb_2_3/io_dat_o[9] cb_2_4/io_wo[0] cb_2_4/io_wo[10] cb_2_4/io_wo[11] cb_2_4/io_wo[12]
+ cb_2_4/io_wo[13] cb_2_4/io_wo[14] cb_2_4/io_wo[15] cb_2_4/io_wo[16] cb_2_4/io_wo[17]
+ cb_2_4/io_wo[18] cb_2_4/io_wo[19] cb_2_4/io_wo[1] cb_2_4/io_wo[20] cb_2_4/io_wo[21]
+ cb_2_4/io_wo[22] cb_2_4/io_wo[23] cb_2_4/io_wo[24] cb_2_4/io_wo[25] cb_2_4/io_wo[26]
+ cb_2_4/io_wo[27] cb_2_4/io_wo[28] cb_2_4/io_wo[29] cb_2_4/io_wo[2] cb_2_4/io_wo[30]
+ cb_2_4/io_wo[31] cb_2_4/io_wo[32] cb_2_4/io_wo[33] cb_2_4/io_wo[34] cb_2_4/io_wo[35]
+ cb_2_4/io_wo[36] cb_2_4/io_wo[37] cb_2_4/io_wo[38] cb_2_4/io_wo[39] cb_2_4/io_wo[3]
+ cb_2_4/io_wo[40] cb_2_4/io_wo[41] cb_2_4/io_wo[42] cb_2_4/io_wo[43] cb_2_4/io_wo[44]
+ cb_2_4/io_wo[45] cb_2_4/io_wo[46] cb_2_4/io_wo[47] cb_2_4/io_wo[48] cb_2_4/io_wo[49]
+ cb_2_4/io_wo[4] cb_2_4/io_wo[50] cb_2_4/io_wo[51] cb_2_4/io_wo[52] cb_2_4/io_wo[53]
+ cb_2_4/io_wo[54] cb_2_4/io_wo[55] cb_2_4/io_wo[56] cb_2_4/io_wo[57] cb_2_4/io_wo[58]
+ cb_2_4/io_wo[59] cb_2_4/io_wo[5] cb_2_4/io_wo[60] cb_2_4/io_wo[61] cb_2_4/io_wo[62]
+ cb_2_4/io_wo[63] cb_2_4/io_wo[6] cb_2_4/io_wo[7] cb_2_4/io_wo[8] cb_2_4/io_wo[9]
+ cb_2_3/io_i_0_ci cb_2_3/io_i_0_in1[0] cb_2_3/io_i_0_in1[1] cb_2_3/io_i_0_in1[2]
+ cb_2_3/io_i_0_in1[3] cb_2_3/io_i_0_in1[4] cb_2_3/io_i_0_in1[5] cb_2_3/io_i_0_in1[6]
+ cb_2_3/io_i_0_in1[7] cb_2_3/io_i_1_ci cb_2_3/io_i_1_in1[0] cb_2_3/io_i_1_in1[1]
+ cb_2_3/io_i_1_in1[2] cb_2_3/io_i_1_in1[3] cb_2_3/io_i_1_in1[4] cb_2_3/io_i_1_in1[5]
+ cb_2_3/io_i_1_in1[6] cb_2_3/io_i_1_in1[7] cb_2_3/io_i_2_ci cb_2_3/io_i_2_in1[0]
+ cb_2_3/io_i_2_in1[1] cb_2_3/io_i_2_in1[2] cb_2_3/io_i_2_in1[3] cb_2_3/io_i_2_in1[4]
+ cb_2_3/io_i_2_in1[5] cb_2_3/io_i_2_in1[6] cb_2_3/io_i_2_in1[7] cb_2_3/io_i_3_ci
+ cb_2_3/io_i_3_in1[0] cb_2_3/io_i_3_in1[1] cb_2_3/io_i_3_in1[2] cb_2_3/io_i_3_in1[3]
+ cb_2_3/io_i_3_in1[4] cb_2_3/io_i_3_in1[5] cb_2_3/io_i_3_in1[6] cb_2_3/io_i_3_in1[7]
+ cb_2_3/io_i_4_ci cb_2_3/io_i_4_in1[0] cb_2_3/io_i_4_in1[1] cb_2_3/io_i_4_in1[2]
+ cb_2_3/io_i_4_in1[3] cb_2_3/io_i_4_in1[4] cb_2_3/io_i_4_in1[5] cb_2_3/io_i_4_in1[6]
+ cb_2_3/io_i_4_in1[7] cb_2_3/io_i_5_ci cb_2_3/io_i_5_in1[0] cb_2_3/io_i_5_in1[1]
+ cb_2_3/io_i_5_in1[2] cb_2_3/io_i_5_in1[3] cb_2_3/io_i_5_in1[4] cb_2_3/io_i_5_in1[5]
+ cb_2_3/io_i_5_in1[6] cb_2_3/io_i_5_in1[7] cb_2_3/io_i_6_ci cb_2_3/io_i_6_in1[0]
+ cb_2_3/io_i_6_in1[1] cb_2_3/io_i_6_in1[2] cb_2_3/io_i_6_in1[3] cb_2_3/io_i_6_in1[4]
+ cb_2_3/io_i_6_in1[5] cb_2_3/io_i_6_in1[6] cb_2_3/io_i_6_in1[7] cb_2_3/io_i_7_ci
+ cb_2_3/io_i_7_in1[0] cb_2_3/io_i_7_in1[1] cb_2_3/io_i_7_in1[2] cb_2_3/io_i_7_in1[3]
+ cb_2_3/io_i_7_in1[4] cb_2_3/io_i_7_in1[5] cb_2_3/io_i_7_in1[6] cb_2_3/io_i_7_in1[7]
+ cb_2_4/io_i_0_ci cb_2_4/io_i_0_in1[0] cb_2_4/io_i_0_in1[1] cb_2_4/io_i_0_in1[2]
+ cb_2_4/io_i_0_in1[3] cb_2_4/io_i_0_in1[4] cb_2_4/io_i_0_in1[5] cb_2_4/io_i_0_in1[6]
+ cb_2_4/io_i_0_in1[7] cb_2_4/io_i_1_ci cb_2_4/io_i_1_in1[0] cb_2_4/io_i_1_in1[1]
+ cb_2_4/io_i_1_in1[2] cb_2_4/io_i_1_in1[3] cb_2_4/io_i_1_in1[4] cb_2_4/io_i_1_in1[5]
+ cb_2_4/io_i_1_in1[6] cb_2_4/io_i_1_in1[7] cb_2_4/io_i_2_ci cb_2_4/io_i_2_in1[0]
+ cb_2_4/io_i_2_in1[1] cb_2_4/io_i_2_in1[2] cb_2_4/io_i_2_in1[3] cb_2_4/io_i_2_in1[4]
+ cb_2_4/io_i_2_in1[5] cb_2_4/io_i_2_in1[6] cb_2_4/io_i_2_in1[7] cb_2_4/io_i_3_ci
+ cb_2_4/io_i_3_in1[0] cb_2_4/io_i_3_in1[1] cb_2_4/io_i_3_in1[2] cb_2_4/io_i_3_in1[3]
+ cb_2_4/io_i_3_in1[4] cb_2_4/io_i_3_in1[5] cb_2_4/io_i_3_in1[6] cb_2_4/io_i_3_in1[7]
+ cb_2_4/io_i_4_ci cb_2_4/io_i_4_in1[0] cb_2_4/io_i_4_in1[1] cb_2_4/io_i_4_in1[2]
+ cb_2_4/io_i_4_in1[3] cb_2_4/io_i_4_in1[4] cb_2_4/io_i_4_in1[5] cb_2_4/io_i_4_in1[6]
+ cb_2_4/io_i_4_in1[7] cb_2_4/io_i_5_ci cb_2_4/io_i_5_in1[0] cb_2_4/io_i_5_in1[1]
+ cb_2_4/io_i_5_in1[2] cb_2_4/io_i_5_in1[3] cb_2_4/io_i_5_in1[4] cb_2_4/io_i_5_in1[5]
+ cb_2_4/io_i_5_in1[6] cb_2_4/io_i_5_in1[7] cb_2_4/io_i_6_ci cb_2_4/io_i_6_in1[0]
+ cb_2_4/io_i_6_in1[1] cb_2_4/io_i_6_in1[2] cb_2_4/io_i_6_in1[3] cb_2_4/io_i_6_in1[4]
+ cb_2_4/io_i_6_in1[5] cb_2_4/io_i_6_in1[6] cb_2_4/io_i_6_in1[7] cb_2_4/io_i_7_ci
+ cb_2_4/io_i_7_in1[0] cb_2_4/io_i_7_in1[1] cb_2_4/io_i_7_in1[2] cb_2_4/io_i_7_in1[3]
+ cb_2_4/io_i_7_in1[4] cb_2_4/io_i_7_in1[5] cb_2_4/io_i_7_in1[6] cb_2_4/io_i_7_in1[7]
+ cb_2_3/io_vci cb_2_4/io_vci cb_2_3/io_vi cb_2_9/io_we_i cb_2_3/io_wo[0] cb_2_3/io_wo[10]
+ cb_2_3/io_wo[11] cb_2_3/io_wo[12] cb_2_3/io_wo[13] cb_2_3/io_wo[14] cb_2_3/io_wo[15]
+ cb_2_3/io_wo[16] cb_2_3/io_wo[17] cb_2_3/io_wo[18] cb_2_3/io_wo[19] cb_2_3/io_wo[1]
+ cb_2_3/io_wo[20] cb_2_3/io_wo[21] cb_2_3/io_wo[22] cb_2_3/io_wo[23] cb_2_3/io_wo[24]
+ cb_2_3/io_wo[25] cb_2_3/io_wo[26] cb_2_3/io_wo[27] cb_2_3/io_wo[28] cb_2_3/io_wo[29]
+ cb_2_3/io_wo[2] cb_2_3/io_wo[30] cb_2_3/io_wo[31] cb_2_3/io_wo[32] cb_2_3/io_wo[33]
+ cb_2_3/io_wo[34] cb_2_3/io_wo[35] cb_2_3/io_wo[36] cb_2_3/io_wo[37] cb_2_3/io_wo[38]
+ cb_2_3/io_wo[39] cb_2_3/io_wo[3] cb_2_3/io_wo[40] cb_2_3/io_wo[41] cb_2_3/io_wo[42]
+ cb_2_3/io_wo[43] cb_2_3/io_wo[44] cb_2_3/io_wo[45] cb_2_3/io_wo[46] cb_2_3/io_wo[47]
+ cb_2_3/io_wo[48] cb_2_3/io_wo[49] cb_2_3/io_wo[4] cb_2_3/io_wo[50] cb_2_3/io_wo[51]
+ cb_2_3/io_wo[52] cb_2_3/io_wo[53] cb_2_3/io_wo[54] cb_2_3/io_wo[55] cb_2_3/io_wo[56]
+ cb_2_3/io_wo[57] cb_2_3/io_wo[58] cb_2_3/io_wo[59] cb_2_3/io_wo[5] cb_2_3/io_wo[60]
+ cb_2_3/io_wo[61] cb_2_3/io_wo[62] cb_2_3/io_wo[63] cb_2_3/io_wo[6] cb_2_3/io_wo[7]
+ cb_2_3/io_wo[8] cb_2_3/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_0_0 cb_0_9/io_adr_i[0] cb_0_9/io_adr_i[1] cb_0_0/io_cs_i cb_0_9/io_dat_i[0] cb_0_9/io_dat_i[10]
+ cb_0_9/io_dat_i[11] cb_0_9/io_dat_i[12] cb_0_9/io_dat_i[13] cb_0_9/io_dat_i[14]
+ cb_0_9/io_dat_i[15] cb_0_9/io_dat_i[1] cb_0_9/io_dat_i[2] cb_0_9/io_dat_i[3] cb_0_9/io_dat_i[4]
+ cb_0_9/io_dat_i[5] cb_0_9/io_dat_i[6] cb_0_9/io_dat_i[7] cb_0_9/io_dat_i[8] cb_0_9/io_dat_i[9]
+ cb_0_0/io_dat_o[0] cb_0_0/io_dat_o[10] cb_0_0/io_dat_o[11] cb_0_0/io_dat_o[12] cb_0_0/io_dat_o[13]
+ cb_0_0/io_dat_o[14] cb_0_0/io_dat_o[15] cb_0_0/io_dat_o[1] cb_0_0/io_dat_o[2] cb_0_0/io_dat_o[3]
+ cb_0_0/io_dat_o[4] cb_0_0/io_dat_o[5] cb_0_0/io_dat_o[6] cb_0_0/io_dat_o[7] cb_0_0/io_dat_o[8]
+ cb_0_0/io_dat_o[9] cb_0_1/io_wo[0] cb_0_1/io_wo[10] cb_0_1/io_wo[11] cb_0_1/io_wo[12]
+ cb_0_1/io_wo[13] cb_0_1/io_wo[14] cb_0_1/io_wo[15] cb_0_1/io_wo[16] cb_0_1/io_wo[17]
+ cb_0_1/io_wo[18] cb_0_1/io_wo[19] cb_0_1/io_wo[1] cb_0_1/io_wo[20] cb_0_1/io_wo[21]
+ cb_0_1/io_wo[22] cb_0_1/io_wo[23] cb_0_1/io_wo[24] cb_0_1/io_wo[25] cb_0_1/io_wo[26]
+ cb_0_1/io_wo[27] cb_0_1/io_wo[28] cb_0_1/io_wo[29] cb_0_1/io_wo[2] cb_0_1/io_wo[30]
+ cb_0_1/io_wo[31] cb_0_1/io_wo[32] cb_0_1/io_wo[33] cb_0_1/io_wo[34] cb_0_1/io_wo[35]
+ cb_0_1/io_wo[36] cb_0_1/io_wo[37] cb_0_1/io_wo[38] cb_0_1/io_wo[39] cb_0_1/io_wo[3]
+ cb_0_1/io_wo[40] cb_0_1/io_wo[41] cb_0_1/io_wo[42] cb_0_1/io_wo[43] cb_0_1/io_wo[44]
+ cb_0_1/io_wo[45] cb_0_1/io_wo[46] cb_0_1/io_wo[47] cb_0_1/io_wo[48] cb_0_1/io_wo[49]
+ cb_0_1/io_wo[4] cb_0_1/io_wo[50] cb_0_1/io_wo[51] cb_0_1/io_wo[52] cb_0_1/io_wo[53]
+ cb_0_1/io_wo[54] cb_0_1/io_wo[55] cb_0_1/io_wo[56] cb_0_1/io_wo[57] cb_0_1/io_wo[58]
+ cb_0_1/io_wo[59] cb_0_1/io_wo[5] cb_0_1/io_wo[60] cb_0_1/io_wo[61] cb_0_1/io_wo[62]
+ cb_0_1/io_wo[63] cb_0_1/io_wo[6] cb_0_1/io_wo[7] cb_0_1/io_wo[8] cb_0_1/io_wo[9]
+ ccon_0/io_dsi_o cb_0_0/io_i_0_in1[0] cb_0_0/io_i_0_in1[1] cb_0_0/io_i_0_in1[2] cb_0_0/io_i_0_in1[3]
+ cb_0_0/io_i_0_in1[4] cb_0_0/io_i_0_in1[5] cb_0_0/io_i_0_in1[6] cb_0_0/io_i_0_in1[7]
+ cb_0_0/io_i_1_ci cb_0_0/io_i_1_in1[0] cb_0_0/io_i_1_in1[1] cb_0_0/io_i_1_in1[2]
+ cb_0_0/io_i_1_in1[3] cb_0_0/io_i_1_in1[4] cb_0_0/io_i_1_in1[5] cb_0_0/io_i_1_in1[6]
+ cb_0_0/io_i_1_in1[7] cb_0_0/io_i_2_ci cb_0_0/io_i_2_in1[0] cb_0_0/io_i_2_in1[1]
+ cb_0_0/io_i_2_in1[2] cb_0_0/io_i_2_in1[3] cb_0_0/io_i_2_in1[4] cb_0_0/io_i_2_in1[5]
+ cb_0_0/io_i_2_in1[6] cb_0_0/io_i_2_in1[7] cb_0_0/io_i_3_ci cb_0_0/io_i_3_in1[0]
+ cb_0_0/io_i_3_in1[1] cb_0_0/io_i_3_in1[2] cb_0_0/io_i_3_in1[3] cb_0_0/io_i_3_in1[4]
+ cb_0_0/io_i_3_in1[5] cb_0_0/io_i_3_in1[6] cb_0_0/io_i_3_in1[7] cb_0_0/io_i_4_ci
+ cb_0_0/io_i_4_in1[0] cb_0_0/io_i_4_in1[1] cb_0_0/io_i_4_in1[2] cb_0_0/io_i_4_in1[3]
+ cb_0_0/io_i_4_in1[4] cb_0_0/io_i_4_in1[5] cb_0_0/io_i_4_in1[6] cb_0_0/io_i_4_in1[7]
+ cb_0_0/io_i_5_ci cb_0_0/io_i_5_in1[0] cb_0_0/io_i_5_in1[1] cb_0_0/io_i_5_in1[2]
+ cb_0_0/io_i_5_in1[3] cb_0_0/io_i_5_in1[4] cb_0_0/io_i_5_in1[5] cb_0_0/io_i_5_in1[6]
+ cb_0_0/io_i_5_in1[7] cb_0_0/io_i_6_ci cb_0_0/io_i_6_in1[0] cb_0_0/io_i_6_in1[1]
+ cb_0_0/io_i_6_in1[2] cb_0_0/io_i_6_in1[3] cb_0_0/io_i_6_in1[4] cb_0_0/io_i_6_in1[5]
+ cb_0_0/io_i_6_in1[6] cb_0_0/io_i_6_in1[7] cb_0_0/io_i_7_ci cb_0_0/io_i_7_in1[0]
+ cb_0_0/io_i_7_in1[1] cb_0_0/io_i_7_in1[2] cb_0_0/io_i_7_in1[3] cb_0_0/io_i_7_in1[4]
+ cb_0_0/io_i_7_in1[5] cb_0_0/io_i_7_in1[6] cb_0_0/io_i_7_in1[7] cb_0_1/io_i_0_ci
+ cb_0_1/io_i_0_in1[0] cb_0_1/io_i_0_in1[1] cb_0_1/io_i_0_in1[2] cb_0_1/io_i_0_in1[3]
+ cb_0_1/io_i_0_in1[4] cb_0_1/io_i_0_in1[5] cb_0_1/io_i_0_in1[6] cb_0_1/io_i_0_in1[7]
+ cb_0_1/io_i_1_ci cb_0_1/io_i_1_in1[0] cb_0_1/io_i_1_in1[1] cb_0_1/io_i_1_in1[2]
+ cb_0_1/io_i_1_in1[3] cb_0_1/io_i_1_in1[4] cb_0_1/io_i_1_in1[5] cb_0_1/io_i_1_in1[6]
+ cb_0_1/io_i_1_in1[7] cb_0_1/io_i_2_ci cb_0_1/io_i_2_in1[0] cb_0_1/io_i_2_in1[1]
+ cb_0_1/io_i_2_in1[2] cb_0_1/io_i_2_in1[3] cb_0_1/io_i_2_in1[4] cb_0_1/io_i_2_in1[5]
+ cb_0_1/io_i_2_in1[6] cb_0_1/io_i_2_in1[7] cb_0_1/io_i_3_ci cb_0_1/io_i_3_in1[0]
+ cb_0_1/io_i_3_in1[1] cb_0_1/io_i_3_in1[2] cb_0_1/io_i_3_in1[3] cb_0_1/io_i_3_in1[4]
+ cb_0_1/io_i_3_in1[5] cb_0_1/io_i_3_in1[6] cb_0_1/io_i_3_in1[7] cb_0_1/io_i_4_ci
+ cb_0_1/io_i_4_in1[0] cb_0_1/io_i_4_in1[1] cb_0_1/io_i_4_in1[2] cb_0_1/io_i_4_in1[3]
+ cb_0_1/io_i_4_in1[4] cb_0_1/io_i_4_in1[5] cb_0_1/io_i_4_in1[6] cb_0_1/io_i_4_in1[7]
+ cb_0_1/io_i_5_ci cb_0_1/io_i_5_in1[0] cb_0_1/io_i_5_in1[1] cb_0_1/io_i_5_in1[2]
+ cb_0_1/io_i_5_in1[3] cb_0_1/io_i_5_in1[4] cb_0_1/io_i_5_in1[5] cb_0_1/io_i_5_in1[6]
+ cb_0_1/io_i_5_in1[7] cb_0_1/io_i_6_ci cb_0_1/io_i_6_in1[0] cb_0_1/io_i_6_in1[1]
+ cb_0_1/io_i_6_in1[2] cb_0_1/io_i_6_in1[3] cb_0_1/io_i_6_in1[4] cb_0_1/io_i_6_in1[5]
+ cb_0_1/io_i_6_in1[6] cb_0_1/io_i_6_in1[7] cb_0_1/io_i_7_ci cb_0_1/io_i_7_in1[0]
+ cb_0_1/io_i_7_in1[1] cb_0_1/io_i_7_in1[2] cb_0_1/io_i_7_in1[3] cb_0_1/io_i_7_in1[4]
+ cb_0_1/io_i_7_in1[5] cb_0_1/io_i_7_in1[6] cb_0_1/io_i_7_in1[7] cb_0_0/io_vci cb_0_1/io_vci
+ cb_0_0/io_vi cb_0_9/io_we_i cb_0_0/io_wo[0] cb_0_0/io_wo[10] cb_0_0/io_wo[11] cb_0_0/io_wo[12]
+ cb_0_0/io_wo[13] cb_0_0/io_wo[14] cb_0_0/io_wo[15] cb_0_0/io_wo[16] cb_0_0/io_wo[17]
+ cb_0_0/io_wo[18] cb_0_0/io_wo[19] cb_0_0/io_wo[1] cb_0_0/io_wo[20] cb_0_0/io_wo[21]
+ cb_0_0/io_wo[22] cb_0_0/io_wo[23] cb_0_0/io_wo[24] cb_0_0/io_wo[25] cb_0_0/io_wo[26]
+ cb_0_0/io_wo[27] cb_0_0/io_wo[28] cb_0_0/io_wo[29] cb_0_0/io_wo[2] cb_0_0/io_wo[30]
+ cb_0_0/io_wo[31] cb_0_0/io_wo[32] cb_0_0/io_wo[33] cb_0_0/io_wo[34] cb_0_0/io_wo[35]
+ cb_0_0/io_wo[36] cb_0_0/io_wo[37] cb_0_0/io_wo[38] cb_0_0/io_wo[39] cb_0_0/io_wo[3]
+ cb_0_0/io_wo[40] cb_0_0/io_wo[41] cb_0_0/io_wo[42] cb_0_0/io_wo[43] cb_0_0/io_wo[44]
+ cb_0_0/io_wo[45] cb_0_0/io_wo[46] cb_0_0/io_wo[47] cb_0_0/io_wo[48] cb_0_0/io_wo[49]
+ cb_0_0/io_wo[4] cb_0_0/io_wo[50] cb_0_0/io_wo[51] cb_0_0/io_wo[52] cb_0_0/io_wo[53]
+ cb_0_0/io_wo[54] cb_0_0/io_wo[55] cb_0_0/io_wo[56] cb_0_0/io_wo[57] cb_0_0/io_wo[58]
+ cb_0_0/io_wo[59] cb_0_0/io_wo[5] cb_0_0/io_wo[60] cb_0_0/io_wo[61] cb_0_0/io_wo[62]
+ cb_0_0/io_wo[63] cb_0_0/io_wo[6] cb_0_0/io_wo[7] cb_0_0/io_wo[8] cb_0_0/io_wo[9]
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_4_7 cb_4_9/io_adr_i[0] cb_4_9/io_adr_i[1] cb_4_7/io_cs_i cb_4_9/io_dat_i[0] cb_4_9/io_dat_i[10]
+ cb_4_9/io_dat_i[11] cb_4_9/io_dat_i[12] cb_4_9/io_dat_i[13] cb_4_9/io_dat_i[14]
+ cb_4_9/io_dat_i[15] cb_4_9/io_dat_i[1] cb_4_9/io_dat_i[2] cb_4_9/io_dat_i[3] cb_4_9/io_dat_i[4]
+ cb_4_9/io_dat_i[5] cb_4_9/io_dat_i[6] cb_4_9/io_dat_i[7] cb_4_9/io_dat_i[8] cb_4_9/io_dat_i[9]
+ cb_4_7/io_dat_o[0] cb_4_7/io_dat_o[10] cb_4_7/io_dat_o[11] cb_4_7/io_dat_o[12] cb_4_7/io_dat_o[13]
+ cb_4_7/io_dat_o[14] cb_4_7/io_dat_o[15] cb_4_7/io_dat_o[1] cb_4_7/io_dat_o[2] cb_4_7/io_dat_o[3]
+ cb_4_7/io_dat_o[4] cb_4_7/io_dat_o[5] cb_4_7/io_dat_o[6] cb_4_7/io_dat_o[7] cb_4_7/io_dat_o[8]
+ cb_4_7/io_dat_o[9] cb_4_8/io_wo[0] cb_4_8/io_wo[10] cb_4_8/io_wo[11] cb_4_8/io_wo[12]
+ cb_4_8/io_wo[13] cb_4_8/io_wo[14] cb_4_8/io_wo[15] cb_4_8/io_wo[16] cb_4_8/io_wo[17]
+ cb_4_8/io_wo[18] cb_4_8/io_wo[19] cb_4_8/io_wo[1] cb_4_8/io_wo[20] cb_4_8/io_wo[21]
+ cb_4_8/io_wo[22] cb_4_8/io_wo[23] cb_4_8/io_wo[24] cb_4_8/io_wo[25] cb_4_8/io_wo[26]
+ cb_4_8/io_wo[27] cb_4_8/io_wo[28] cb_4_8/io_wo[29] cb_4_8/io_wo[2] cb_4_8/io_wo[30]
+ cb_4_8/io_wo[31] cb_4_8/io_wo[32] cb_4_8/io_wo[33] cb_4_8/io_wo[34] cb_4_8/io_wo[35]
+ cb_4_8/io_wo[36] cb_4_8/io_wo[37] cb_4_8/io_wo[38] cb_4_8/io_wo[39] cb_4_8/io_wo[3]
+ cb_4_8/io_wo[40] cb_4_8/io_wo[41] cb_4_8/io_wo[42] cb_4_8/io_wo[43] cb_4_8/io_wo[44]
+ cb_4_8/io_wo[45] cb_4_8/io_wo[46] cb_4_8/io_wo[47] cb_4_8/io_wo[48] cb_4_8/io_wo[49]
+ cb_4_8/io_wo[4] cb_4_8/io_wo[50] cb_4_8/io_wo[51] cb_4_8/io_wo[52] cb_4_8/io_wo[53]
+ cb_4_8/io_wo[54] cb_4_8/io_wo[55] cb_4_8/io_wo[56] cb_4_8/io_wo[57] cb_4_8/io_wo[58]
+ cb_4_8/io_wo[59] cb_4_8/io_wo[5] cb_4_8/io_wo[60] cb_4_8/io_wo[61] cb_4_8/io_wo[62]
+ cb_4_8/io_wo[63] cb_4_8/io_wo[6] cb_4_8/io_wo[7] cb_4_8/io_wo[8] cb_4_8/io_wo[9]
+ cb_4_7/io_i_0_ci cb_4_7/io_i_0_in1[0] cb_4_7/io_i_0_in1[1] cb_4_7/io_i_0_in1[2]
+ cb_4_7/io_i_0_in1[3] cb_4_7/io_i_0_in1[4] cb_4_7/io_i_0_in1[5] cb_4_7/io_i_0_in1[6]
+ cb_4_7/io_i_0_in1[7] cb_4_7/io_i_1_ci cb_4_7/io_i_1_in1[0] cb_4_7/io_i_1_in1[1]
+ cb_4_7/io_i_1_in1[2] cb_4_7/io_i_1_in1[3] cb_4_7/io_i_1_in1[4] cb_4_7/io_i_1_in1[5]
+ cb_4_7/io_i_1_in1[6] cb_4_7/io_i_1_in1[7] cb_4_7/io_i_2_ci cb_4_7/io_i_2_in1[0]
+ cb_4_7/io_i_2_in1[1] cb_4_7/io_i_2_in1[2] cb_4_7/io_i_2_in1[3] cb_4_7/io_i_2_in1[4]
+ cb_4_7/io_i_2_in1[5] cb_4_7/io_i_2_in1[6] cb_4_7/io_i_2_in1[7] cb_4_7/io_i_3_ci
+ cb_4_7/io_i_3_in1[0] cb_4_7/io_i_3_in1[1] cb_4_7/io_i_3_in1[2] cb_4_7/io_i_3_in1[3]
+ cb_4_7/io_i_3_in1[4] cb_4_7/io_i_3_in1[5] cb_4_7/io_i_3_in1[6] cb_4_7/io_i_3_in1[7]
+ cb_4_7/io_i_4_ci cb_4_7/io_i_4_in1[0] cb_4_7/io_i_4_in1[1] cb_4_7/io_i_4_in1[2]
+ cb_4_7/io_i_4_in1[3] cb_4_7/io_i_4_in1[4] cb_4_7/io_i_4_in1[5] cb_4_7/io_i_4_in1[6]
+ cb_4_7/io_i_4_in1[7] cb_4_7/io_i_5_ci cb_4_7/io_i_5_in1[0] cb_4_7/io_i_5_in1[1]
+ cb_4_7/io_i_5_in1[2] cb_4_7/io_i_5_in1[3] cb_4_7/io_i_5_in1[4] cb_4_7/io_i_5_in1[5]
+ cb_4_7/io_i_5_in1[6] cb_4_7/io_i_5_in1[7] cb_4_7/io_i_6_ci cb_4_7/io_i_6_in1[0]
+ cb_4_7/io_i_6_in1[1] cb_4_7/io_i_6_in1[2] cb_4_7/io_i_6_in1[3] cb_4_7/io_i_6_in1[4]
+ cb_4_7/io_i_6_in1[5] cb_4_7/io_i_6_in1[6] cb_4_7/io_i_6_in1[7] cb_4_7/io_i_7_ci
+ cb_4_7/io_i_7_in1[0] cb_4_7/io_i_7_in1[1] cb_4_7/io_i_7_in1[2] cb_4_7/io_i_7_in1[3]
+ cb_4_7/io_i_7_in1[4] cb_4_7/io_i_7_in1[5] cb_4_7/io_i_7_in1[6] cb_4_7/io_i_7_in1[7]
+ cb_4_8/io_i_0_ci cb_4_8/io_i_0_in1[0] cb_4_8/io_i_0_in1[1] cb_4_8/io_i_0_in1[2]
+ cb_4_8/io_i_0_in1[3] cb_4_8/io_i_0_in1[4] cb_4_8/io_i_0_in1[5] cb_4_8/io_i_0_in1[6]
+ cb_4_8/io_i_0_in1[7] cb_4_8/io_i_1_ci cb_4_8/io_i_1_in1[0] cb_4_8/io_i_1_in1[1]
+ cb_4_8/io_i_1_in1[2] cb_4_8/io_i_1_in1[3] cb_4_8/io_i_1_in1[4] cb_4_8/io_i_1_in1[5]
+ cb_4_8/io_i_1_in1[6] cb_4_8/io_i_1_in1[7] cb_4_8/io_i_2_ci cb_4_8/io_i_2_in1[0]
+ cb_4_8/io_i_2_in1[1] cb_4_8/io_i_2_in1[2] cb_4_8/io_i_2_in1[3] cb_4_8/io_i_2_in1[4]
+ cb_4_8/io_i_2_in1[5] cb_4_8/io_i_2_in1[6] cb_4_8/io_i_2_in1[7] cb_4_8/io_i_3_ci
+ cb_4_8/io_i_3_in1[0] cb_4_8/io_i_3_in1[1] cb_4_8/io_i_3_in1[2] cb_4_8/io_i_3_in1[3]
+ cb_4_8/io_i_3_in1[4] cb_4_8/io_i_3_in1[5] cb_4_8/io_i_3_in1[6] cb_4_8/io_i_3_in1[7]
+ cb_4_8/io_i_4_ci cb_4_8/io_i_4_in1[0] cb_4_8/io_i_4_in1[1] cb_4_8/io_i_4_in1[2]
+ cb_4_8/io_i_4_in1[3] cb_4_8/io_i_4_in1[4] cb_4_8/io_i_4_in1[5] cb_4_8/io_i_4_in1[6]
+ cb_4_8/io_i_4_in1[7] cb_4_8/io_i_5_ci cb_4_8/io_i_5_in1[0] cb_4_8/io_i_5_in1[1]
+ cb_4_8/io_i_5_in1[2] cb_4_8/io_i_5_in1[3] cb_4_8/io_i_5_in1[4] cb_4_8/io_i_5_in1[5]
+ cb_4_8/io_i_5_in1[6] cb_4_8/io_i_5_in1[7] cb_4_8/io_i_6_ci cb_4_8/io_i_6_in1[0]
+ cb_4_8/io_i_6_in1[1] cb_4_8/io_i_6_in1[2] cb_4_8/io_i_6_in1[3] cb_4_8/io_i_6_in1[4]
+ cb_4_8/io_i_6_in1[5] cb_4_8/io_i_6_in1[6] cb_4_8/io_i_6_in1[7] cb_4_8/io_i_7_ci
+ cb_4_8/io_i_7_in1[0] cb_4_8/io_i_7_in1[1] cb_4_8/io_i_7_in1[2] cb_4_8/io_i_7_in1[3]
+ cb_4_8/io_i_7_in1[4] cb_4_8/io_i_7_in1[5] cb_4_8/io_i_7_in1[6] cb_4_8/io_i_7_in1[7]
+ cb_4_7/io_vci cb_4_8/io_vci cb_4_7/io_vi cb_4_9/io_we_i cb_4_7/io_wo[0] cb_4_7/io_wo[10]
+ cb_4_7/io_wo[11] cb_4_7/io_wo[12] cb_4_7/io_wo[13] cb_4_7/io_wo[14] cb_4_7/io_wo[15]
+ cb_4_7/io_wo[16] cb_4_7/io_wo[17] cb_4_7/io_wo[18] cb_4_7/io_wo[19] cb_4_7/io_wo[1]
+ cb_4_7/io_wo[20] cb_4_7/io_wo[21] cb_4_7/io_wo[22] cb_4_7/io_wo[23] cb_4_7/io_wo[24]
+ cb_4_7/io_wo[25] cb_4_7/io_wo[26] cb_4_7/io_wo[27] cb_4_7/io_wo[28] cb_4_7/io_wo[29]
+ cb_4_7/io_wo[2] cb_4_7/io_wo[30] cb_4_7/io_wo[31] cb_4_7/io_wo[32] cb_4_7/io_wo[33]
+ cb_4_7/io_wo[34] cb_4_7/io_wo[35] cb_4_7/io_wo[36] cb_4_7/io_wo[37] cb_4_7/io_wo[38]
+ cb_4_7/io_wo[39] cb_4_7/io_wo[3] cb_4_7/io_wo[40] cb_4_7/io_wo[41] cb_4_7/io_wo[42]
+ cb_4_7/io_wo[43] cb_4_7/io_wo[44] cb_4_7/io_wo[45] cb_4_7/io_wo[46] cb_4_7/io_wo[47]
+ cb_4_7/io_wo[48] cb_4_7/io_wo[49] cb_4_7/io_wo[4] cb_4_7/io_wo[50] cb_4_7/io_wo[51]
+ cb_4_7/io_wo[52] cb_4_7/io_wo[53] cb_4_7/io_wo[54] cb_4_7/io_wo[55] cb_4_7/io_wo[56]
+ cb_4_7/io_wo[57] cb_4_7/io_wo[58] cb_4_7/io_wo[59] cb_4_7/io_wo[5] cb_4_7/io_wo[60]
+ cb_4_7/io_wo[61] cb_4_7/io_wo[62] cb_4_7/io_wo[63] cb_4_7/io_wo[6] cb_4_7/io_wo[7]
+ cb_4_7/io_wo[8] cb_4_7/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_2_4 cb_2_9/io_adr_i[0] cb_2_9/io_adr_i[1] cb_2_4/io_cs_i cb_2_9/io_dat_i[0] cb_2_9/io_dat_i[10]
+ cb_2_9/io_dat_i[11] cb_2_9/io_dat_i[12] cb_2_9/io_dat_i[13] cb_2_9/io_dat_i[14]
+ cb_2_9/io_dat_i[15] cb_2_9/io_dat_i[1] cb_2_9/io_dat_i[2] cb_2_9/io_dat_i[3] cb_2_9/io_dat_i[4]
+ cb_2_9/io_dat_i[5] cb_2_9/io_dat_i[6] cb_2_9/io_dat_i[7] cb_2_9/io_dat_i[8] cb_2_9/io_dat_i[9]
+ cb_2_4/io_dat_o[0] cb_2_4/io_dat_o[10] cb_2_4/io_dat_o[11] cb_2_4/io_dat_o[12] cb_2_4/io_dat_o[13]
+ cb_2_4/io_dat_o[14] cb_2_4/io_dat_o[15] cb_2_4/io_dat_o[1] cb_2_4/io_dat_o[2] cb_2_4/io_dat_o[3]
+ cb_2_4/io_dat_o[4] cb_2_4/io_dat_o[5] cb_2_4/io_dat_o[6] cb_2_4/io_dat_o[7] cb_2_4/io_dat_o[8]
+ cb_2_4/io_dat_o[9] cb_2_5/io_wo[0] cb_2_5/io_wo[10] cb_2_5/io_wo[11] cb_2_5/io_wo[12]
+ cb_2_5/io_wo[13] cb_2_5/io_wo[14] cb_2_5/io_wo[15] cb_2_5/io_wo[16] cb_2_5/io_wo[17]
+ cb_2_5/io_wo[18] cb_2_5/io_wo[19] cb_2_5/io_wo[1] cb_2_5/io_wo[20] cb_2_5/io_wo[21]
+ cb_2_5/io_wo[22] cb_2_5/io_wo[23] cb_2_5/io_wo[24] cb_2_5/io_wo[25] cb_2_5/io_wo[26]
+ cb_2_5/io_wo[27] cb_2_5/io_wo[28] cb_2_5/io_wo[29] cb_2_5/io_wo[2] cb_2_5/io_wo[30]
+ cb_2_5/io_wo[31] cb_2_5/io_wo[32] cb_2_5/io_wo[33] cb_2_5/io_wo[34] cb_2_5/io_wo[35]
+ cb_2_5/io_wo[36] cb_2_5/io_wo[37] cb_2_5/io_wo[38] cb_2_5/io_wo[39] cb_2_5/io_wo[3]
+ cb_2_5/io_wo[40] cb_2_5/io_wo[41] cb_2_5/io_wo[42] cb_2_5/io_wo[43] cb_2_5/io_wo[44]
+ cb_2_5/io_wo[45] cb_2_5/io_wo[46] cb_2_5/io_wo[47] cb_2_5/io_wo[48] cb_2_5/io_wo[49]
+ cb_2_5/io_wo[4] cb_2_5/io_wo[50] cb_2_5/io_wo[51] cb_2_5/io_wo[52] cb_2_5/io_wo[53]
+ cb_2_5/io_wo[54] cb_2_5/io_wo[55] cb_2_5/io_wo[56] cb_2_5/io_wo[57] cb_2_5/io_wo[58]
+ cb_2_5/io_wo[59] cb_2_5/io_wo[5] cb_2_5/io_wo[60] cb_2_5/io_wo[61] cb_2_5/io_wo[62]
+ cb_2_5/io_wo[63] cb_2_5/io_wo[6] cb_2_5/io_wo[7] cb_2_5/io_wo[8] cb_2_5/io_wo[9]
+ cb_2_4/io_i_0_ci cb_2_4/io_i_0_in1[0] cb_2_4/io_i_0_in1[1] cb_2_4/io_i_0_in1[2]
+ cb_2_4/io_i_0_in1[3] cb_2_4/io_i_0_in1[4] cb_2_4/io_i_0_in1[5] cb_2_4/io_i_0_in1[6]
+ cb_2_4/io_i_0_in1[7] cb_2_4/io_i_1_ci cb_2_4/io_i_1_in1[0] cb_2_4/io_i_1_in1[1]
+ cb_2_4/io_i_1_in1[2] cb_2_4/io_i_1_in1[3] cb_2_4/io_i_1_in1[4] cb_2_4/io_i_1_in1[5]
+ cb_2_4/io_i_1_in1[6] cb_2_4/io_i_1_in1[7] cb_2_4/io_i_2_ci cb_2_4/io_i_2_in1[0]
+ cb_2_4/io_i_2_in1[1] cb_2_4/io_i_2_in1[2] cb_2_4/io_i_2_in1[3] cb_2_4/io_i_2_in1[4]
+ cb_2_4/io_i_2_in1[5] cb_2_4/io_i_2_in1[6] cb_2_4/io_i_2_in1[7] cb_2_4/io_i_3_ci
+ cb_2_4/io_i_3_in1[0] cb_2_4/io_i_3_in1[1] cb_2_4/io_i_3_in1[2] cb_2_4/io_i_3_in1[3]
+ cb_2_4/io_i_3_in1[4] cb_2_4/io_i_3_in1[5] cb_2_4/io_i_3_in1[6] cb_2_4/io_i_3_in1[7]
+ cb_2_4/io_i_4_ci cb_2_4/io_i_4_in1[0] cb_2_4/io_i_4_in1[1] cb_2_4/io_i_4_in1[2]
+ cb_2_4/io_i_4_in1[3] cb_2_4/io_i_4_in1[4] cb_2_4/io_i_4_in1[5] cb_2_4/io_i_4_in1[6]
+ cb_2_4/io_i_4_in1[7] cb_2_4/io_i_5_ci cb_2_4/io_i_5_in1[0] cb_2_4/io_i_5_in1[1]
+ cb_2_4/io_i_5_in1[2] cb_2_4/io_i_5_in1[3] cb_2_4/io_i_5_in1[4] cb_2_4/io_i_5_in1[5]
+ cb_2_4/io_i_5_in1[6] cb_2_4/io_i_5_in1[7] cb_2_4/io_i_6_ci cb_2_4/io_i_6_in1[0]
+ cb_2_4/io_i_6_in1[1] cb_2_4/io_i_6_in1[2] cb_2_4/io_i_6_in1[3] cb_2_4/io_i_6_in1[4]
+ cb_2_4/io_i_6_in1[5] cb_2_4/io_i_6_in1[6] cb_2_4/io_i_6_in1[7] cb_2_4/io_i_7_ci
+ cb_2_4/io_i_7_in1[0] cb_2_4/io_i_7_in1[1] cb_2_4/io_i_7_in1[2] cb_2_4/io_i_7_in1[3]
+ cb_2_4/io_i_7_in1[4] cb_2_4/io_i_7_in1[5] cb_2_4/io_i_7_in1[6] cb_2_4/io_i_7_in1[7]
+ cb_2_5/io_i_0_ci cb_2_5/io_i_0_in1[0] cb_2_5/io_i_0_in1[1] cb_2_5/io_i_0_in1[2]
+ cb_2_5/io_i_0_in1[3] cb_2_5/io_i_0_in1[4] cb_2_5/io_i_0_in1[5] cb_2_5/io_i_0_in1[6]
+ cb_2_5/io_i_0_in1[7] cb_2_5/io_i_1_ci cb_2_5/io_i_1_in1[0] cb_2_5/io_i_1_in1[1]
+ cb_2_5/io_i_1_in1[2] cb_2_5/io_i_1_in1[3] cb_2_5/io_i_1_in1[4] cb_2_5/io_i_1_in1[5]
+ cb_2_5/io_i_1_in1[6] cb_2_5/io_i_1_in1[7] cb_2_5/io_i_2_ci cb_2_5/io_i_2_in1[0]
+ cb_2_5/io_i_2_in1[1] cb_2_5/io_i_2_in1[2] cb_2_5/io_i_2_in1[3] cb_2_5/io_i_2_in1[4]
+ cb_2_5/io_i_2_in1[5] cb_2_5/io_i_2_in1[6] cb_2_5/io_i_2_in1[7] cb_2_5/io_i_3_ci
+ cb_2_5/io_i_3_in1[0] cb_2_5/io_i_3_in1[1] cb_2_5/io_i_3_in1[2] cb_2_5/io_i_3_in1[3]
+ cb_2_5/io_i_3_in1[4] cb_2_5/io_i_3_in1[5] cb_2_5/io_i_3_in1[6] cb_2_5/io_i_3_in1[7]
+ cb_2_5/io_i_4_ci cb_2_5/io_i_4_in1[0] cb_2_5/io_i_4_in1[1] cb_2_5/io_i_4_in1[2]
+ cb_2_5/io_i_4_in1[3] cb_2_5/io_i_4_in1[4] cb_2_5/io_i_4_in1[5] cb_2_5/io_i_4_in1[6]
+ cb_2_5/io_i_4_in1[7] cb_2_5/io_i_5_ci cb_2_5/io_i_5_in1[0] cb_2_5/io_i_5_in1[1]
+ cb_2_5/io_i_5_in1[2] cb_2_5/io_i_5_in1[3] cb_2_5/io_i_5_in1[4] cb_2_5/io_i_5_in1[5]
+ cb_2_5/io_i_5_in1[6] cb_2_5/io_i_5_in1[7] cb_2_5/io_i_6_ci cb_2_5/io_i_6_in1[0]
+ cb_2_5/io_i_6_in1[1] cb_2_5/io_i_6_in1[2] cb_2_5/io_i_6_in1[3] cb_2_5/io_i_6_in1[4]
+ cb_2_5/io_i_6_in1[5] cb_2_5/io_i_6_in1[6] cb_2_5/io_i_6_in1[7] cb_2_5/io_i_7_ci
+ cb_2_5/io_i_7_in1[0] cb_2_5/io_i_7_in1[1] cb_2_5/io_i_7_in1[2] cb_2_5/io_i_7_in1[3]
+ cb_2_5/io_i_7_in1[4] cb_2_5/io_i_7_in1[5] cb_2_5/io_i_7_in1[6] cb_2_5/io_i_7_in1[7]
+ cb_2_4/io_vci cb_2_5/io_vci cb_2_4/io_vi cb_2_9/io_we_i cb_2_4/io_wo[0] cb_2_4/io_wo[10]
+ cb_2_4/io_wo[11] cb_2_4/io_wo[12] cb_2_4/io_wo[13] cb_2_4/io_wo[14] cb_2_4/io_wo[15]
+ cb_2_4/io_wo[16] cb_2_4/io_wo[17] cb_2_4/io_wo[18] cb_2_4/io_wo[19] cb_2_4/io_wo[1]
+ cb_2_4/io_wo[20] cb_2_4/io_wo[21] cb_2_4/io_wo[22] cb_2_4/io_wo[23] cb_2_4/io_wo[24]
+ cb_2_4/io_wo[25] cb_2_4/io_wo[26] cb_2_4/io_wo[27] cb_2_4/io_wo[28] cb_2_4/io_wo[29]
+ cb_2_4/io_wo[2] cb_2_4/io_wo[30] cb_2_4/io_wo[31] cb_2_4/io_wo[32] cb_2_4/io_wo[33]
+ cb_2_4/io_wo[34] cb_2_4/io_wo[35] cb_2_4/io_wo[36] cb_2_4/io_wo[37] cb_2_4/io_wo[38]
+ cb_2_4/io_wo[39] cb_2_4/io_wo[3] cb_2_4/io_wo[40] cb_2_4/io_wo[41] cb_2_4/io_wo[42]
+ cb_2_4/io_wo[43] cb_2_4/io_wo[44] cb_2_4/io_wo[45] cb_2_4/io_wo[46] cb_2_4/io_wo[47]
+ cb_2_4/io_wo[48] cb_2_4/io_wo[49] cb_2_4/io_wo[4] cb_2_4/io_wo[50] cb_2_4/io_wo[51]
+ cb_2_4/io_wo[52] cb_2_4/io_wo[53] cb_2_4/io_wo[54] cb_2_4/io_wo[55] cb_2_4/io_wo[56]
+ cb_2_4/io_wo[57] cb_2_4/io_wo[58] cb_2_4/io_wo[59] cb_2_4/io_wo[5] cb_2_4/io_wo[60]
+ cb_2_4/io_wo[61] cb_2_4/io_wo[62] cb_2_4/io_wo[63] cb_2_4/io_wo[6] cb_2_4/io_wo[7]
+ cb_2_4/io_wo[8] cb_2_4/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_0_1 cb_0_9/io_adr_i[0] cb_0_9/io_adr_i[1] cb_0_1/io_cs_i cb_0_9/io_dat_i[0] cb_0_9/io_dat_i[10]
+ cb_0_9/io_dat_i[11] cb_0_9/io_dat_i[12] cb_0_9/io_dat_i[13] cb_0_9/io_dat_i[14]
+ cb_0_9/io_dat_i[15] cb_0_9/io_dat_i[1] cb_0_9/io_dat_i[2] cb_0_9/io_dat_i[3] cb_0_9/io_dat_i[4]
+ cb_0_9/io_dat_i[5] cb_0_9/io_dat_i[6] cb_0_9/io_dat_i[7] cb_0_9/io_dat_i[8] cb_0_9/io_dat_i[9]
+ cb_0_1/io_dat_o[0] cb_0_1/io_dat_o[10] cb_0_1/io_dat_o[11] cb_0_1/io_dat_o[12] cb_0_1/io_dat_o[13]
+ cb_0_1/io_dat_o[14] cb_0_1/io_dat_o[15] cb_0_1/io_dat_o[1] cb_0_1/io_dat_o[2] cb_0_1/io_dat_o[3]
+ cb_0_1/io_dat_o[4] cb_0_1/io_dat_o[5] cb_0_1/io_dat_o[6] cb_0_1/io_dat_o[7] cb_0_1/io_dat_o[8]
+ cb_0_1/io_dat_o[9] cb_0_2/io_wo[0] cb_0_2/io_wo[10] cb_0_2/io_wo[11] cb_0_2/io_wo[12]
+ cb_0_2/io_wo[13] cb_0_2/io_wo[14] cb_0_2/io_wo[15] cb_0_2/io_wo[16] cb_0_2/io_wo[17]
+ cb_0_2/io_wo[18] cb_0_2/io_wo[19] cb_0_2/io_wo[1] cb_0_2/io_wo[20] cb_0_2/io_wo[21]
+ cb_0_2/io_wo[22] cb_0_2/io_wo[23] cb_0_2/io_wo[24] cb_0_2/io_wo[25] cb_0_2/io_wo[26]
+ cb_0_2/io_wo[27] cb_0_2/io_wo[28] cb_0_2/io_wo[29] cb_0_2/io_wo[2] cb_0_2/io_wo[30]
+ cb_0_2/io_wo[31] cb_0_2/io_wo[32] cb_0_2/io_wo[33] cb_0_2/io_wo[34] cb_0_2/io_wo[35]
+ cb_0_2/io_wo[36] cb_0_2/io_wo[37] cb_0_2/io_wo[38] cb_0_2/io_wo[39] cb_0_2/io_wo[3]
+ cb_0_2/io_wo[40] cb_0_2/io_wo[41] cb_0_2/io_wo[42] cb_0_2/io_wo[43] cb_0_2/io_wo[44]
+ cb_0_2/io_wo[45] cb_0_2/io_wo[46] cb_0_2/io_wo[47] cb_0_2/io_wo[48] cb_0_2/io_wo[49]
+ cb_0_2/io_wo[4] cb_0_2/io_wo[50] cb_0_2/io_wo[51] cb_0_2/io_wo[52] cb_0_2/io_wo[53]
+ cb_0_2/io_wo[54] cb_0_2/io_wo[55] cb_0_2/io_wo[56] cb_0_2/io_wo[57] cb_0_2/io_wo[58]
+ cb_0_2/io_wo[59] cb_0_2/io_wo[5] cb_0_2/io_wo[60] cb_0_2/io_wo[61] cb_0_2/io_wo[62]
+ cb_0_2/io_wo[63] cb_0_2/io_wo[6] cb_0_2/io_wo[7] cb_0_2/io_wo[8] cb_0_2/io_wo[9]
+ cb_0_1/io_i_0_ci cb_0_1/io_i_0_in1[0] cb_0_1/io_i_0_in1[1] cb_0_1/io_i_0_in1[2]
+ cb_0_1/io_i_0_in1[3] cb_0_1/io_i_0_in1[4] cb_0_1/io_i_0_in1[5] cb_0_1/io_i_0_in1[6]
+ cb_0_1/io_i_0_in1[7] cb_0_1/io_i_1_ci cb_0_1/io_i_1_in1[0] cb_0_1/io_i_1_in1[1]
+ cb_0_1/io_i_1_in1[2] cb_0_1/io_i_1_in1[3] cb_0_1/io_i_1_in1[4] cb_0_1/io_i_1_in1[5]
+ cb_0_1/io_i_1_in1[6] cb_0_1/io_i_1_in1[7] cb_0_1/io_i_2_ci cb_0_1/io_i_2_in1[0]
+ cb_0_1/io_i_2_in1[1] cb_0_1/io_i_2_in1[2] cb_0_1/io_i_2_in1[3] cb_0_1/io_i_2_in1[4]
+ cb_0_1/io_i_2_in1[5] cb_0_1/io_i_2_in1[6] cb_0_1/io_i_2_in1[7] cb_0_1/io_i_3_ci
+ cb_0_1/io_i_3_in1[0] cb_0_1/io_i_3_in1[1] cb_0_1/io_i_3_in1[2] cb_0_1/io_i_3_in1[3]
+ cb_0_1/io_i_3_in1[4] cb_0_1/io_i_3_in1[5] cb_0_1/io_i_3_in1[6] cb_0_1/io_i_3_in1[7]
+ cb_0_1/io_i_4_ci cb_0_1/io_i_4_in1[0] cb_0_1/io_i_4_in1[1] cb_0_1/io_i_4_in1[2]
+ cb_0_1/io_i_4_in1[3] cb_0_1/io_i_4_in1[4] cb_0_1/io_i_4_in1[5] cb_0_1/io_i_4_in1[6]
+ cb_0_1/io_i_4_in1[7] cb_0_1/io_i_5_ci cb_0_1/io_i_5_in1[0] cb_0_1/io_i_5_in1[1]
+ cb_0_1/io_i_5_in1[2] cb_0_1/io_i_5_in1[3] cb_0_1/io_i_5_in1[4] cb_0_1/io_i_5_in1[5]
+ cb_0_1/io_i_5_in1[6] cb_0_1/io_i_5_in1[7] cb_0_1/io_i_6_ci cb_0_1/io_i_6_in1[0]
+ cb_0_1/io_i_6_in1[1] cb_0_1/io_i_6_in1[2] cb_0_1/io_i_6_in1[3] cb_0_1/io_i_6_in1[4]
+ cb_0_1/io_i_6_in1[5] cb_0_1/io_i_6_in1[6] cb_0_1/io_i_6_in1[7] cb_0_1/io_i_7_ci
+ cb_0_1/io_i_7_in1[0] cb_0_1/io_i_7_in1[1] cb_0_1/io_i_7_in1[2] cb_0_1/io_i_7_in1[3]
+ cb_0_1/io_i_7_in1[4] cb_0_1/io_i_7_in1[5] cb_0_1/io_i_7_in1[6] cb_0_1/io_i_7_in1[7]
+ cb_0_2/io_i_0_ci cb_0_2/io_i_0_in1[0] cb_0_2/io_i_0_in1[1] cb_0_2/io_i_0_in1[2]
+ cb_0_2/io_i_0_in1[3] cb_0_2/io_i_0_in1[4] cb_0_2/io_i_0_in1[5] cb_0_2/io_i_0_in1[6]
+ cb_0_2/io_i_0_in1[7] cb_0_2/io_i_1_ci cb_0_2/io_i_1_in1[0] cb_0_2/io_i_1_in1[1]
+ cb_0_2/io_i_1_in1[2] cb_0_2/io_i_1_in1[3] cb_0_2/io_i_1_in1[4] cb_0_2/io_i_1_in1[5]
+ cb_0_2/io_i_1_in1[6] cb_0_2/io_i_1_in1[7] cb_0_2/io_i_2_ci cb_0_2/io_i_2_in1[0]
+ cb_0_2/io_i_2_in1[1] cb_0_2/io_i_2_in1[2] cb_0_2/io_i_2_in1[3] cb_0_2/io_i_2_in1[4]
+ cb_0_2/io_i_2_in1[5] cb_0_2/io_i_2_in1[6] cb_0_2/io_i_2_in1[7] cb_0_2/io_i_3_ci
+ cb_0_2/io_i_3_in1[0] cb_0_2/io_i_3_in1[1] cb_0_2/io_i_3_in1[2] cb_0_2/io_i_3_in1[3]
+ cb_0_2/io_i_3_in1[4] cb_0_2/io_i_3_in1[5] cb_0_2/io_i_3_in1[6] cb_0_2/io_i_3_in1[7]
+ cb_0_2/io_i_4_ci cb_0_2/io_i_4_in1[0] cb_0_2/io_i_4_in1[1] cb_0_2/io_i_4_in1[2]
+ cb_0_2/io_i_4_in1[3] cb_0_2/io_i_4_in1[4] cb_0_2/io_i_4_in1[5] cb_0_2/io_i_4_in1[6]
+ cb_0_2/io_i_4_in1[7] cb_0_2/io_i_5_ci cb_0_2/io_i_5_in1[0] cb_0_2/io_i_5_in1[1]
+ cb_0_2/io_i_5_in1[2] cb_0_2/io_i_5_in1[3] cb_0_2/io_i_5_in1[4] cb_0_2/io_i_5_in1[5]
+ cb_0_2/io_i_5_in1[6] cb_0_2/io_i_5_in1[7] cb_0_2/io_i_6_ci cb_0_2/io_i_6_in1[0]
+ cb_0_2/io_i_6_in1[1] cb_0_2/io_i_6_in1[2] cb_0_2/io_i_6_in1[3] cb_0_2/io_i_6_in1[4]
+ cb_0_2/io_i_6_in1[5] cb_0_2/io_i_6_in1[6] cb_0_2/io_i_6_in1[7] cb_0_2/io_i_7_ci
+ cb_0_2/io_i_7_in1[0] cb_0_2/io_i_7_in1[1] cb_0_2/io_i_7_in1[2] cb_0_2/io_i_7_in1[3]
+ cb_0_2/io_i_7_in1[4] cb_0_2/io_i_7_in1[5] cb_0_2/io_i_7_in1[6] cb_0_2/io_i_7_in1[7]
+ cb_0_1/io_vci cb_0_2/io_vci cb_0_1/io_vi cb_0_9/io_we_i cb_0_1/io_wo[0] cb_0_1/io_wo[10]
+ cb_0_1/io_wo[11] cb_0_1/io_wo[12] cb_0_1/io_wo[13] cb_0_1/io_wo[14] cb_0_1/io_wo[15]
+ cb_0_1/io_wo[16] cb_0_1/io_wo[17] cb_0_1/io_wo[18] cb_0_1/io_wo[19] cb_0_1/io_wo[1]
+ cb_0_1/io_wo[20] cb_0_1/io_wo[21] cb_0_1/io_wo[22] cb_0_1/io_wo[23] cb_0_1/io_wo[24]
+ cb_0_1/io_wo[25] cb_0_1/io_wo[26] cb_0_1/io_wo[27] cb_0_1/io_wo[28] cb_0_1/io_wo[29]
+ cb_0_1/io_wo[2] cb_0_1/io_wo[30] cb_0_1/io_wo[31] cb_0_1/io_wo[32] cb_0_1/io_wo[33]
+ cb_0_1/io_wo[34] cb_0_1/io_wo[35] cb_0_1/io_wo[36] cb_0_1/io_wo[37] cb_0_1/io_wo[38]
+ cb_0_1/io_wo[39] cb_0_1/io_wo[3] cb_0_1/io_wo[40] cb_0_1/io_wo[41] cb_0_1/io_wo[42]
+ cb_0_1/io_wo[43] cb_0_1/io_wo[44] cb_0_1/io_wo[45] cb_0_1/io_wo[46] cb_0_1/io_wo[47]
+ cb_0_1/io_wo[48] cb_0_1/io_wo[49] cb_0_1/io_wo[4] cb_0_1/io_wo[50] cb_0_1/io_wo[51]
+ cb_0_1/io_wo[52] cb_0_1/io_wo[53] cb_0_1/io_wo[54] cb_0_1/io_wo[55] cb_0_1/io_wo[56]
+ cb_0_1/io_wo[57] cb_0_1/io_wo[58] cb_0_1/io_wo[59] cb_0_1/io_wo[5] cb_0_1/io_wo[60]
+ cb_0_1/io_wo[61] cb_0_1/io_wo[62] cb_0_1/io_wo[63] cb_0_1/io_wo[6] cb_0_1/io_wo[7]
+ cb_0_1/io_wo[8] cb_0_1/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_4_8 cb_4_9/io_adr_i[0] cb_4_9/io_adr_i[1] cb_4_8/io_cs_i cb_4_9/io_dat_i[0] cb_4_9/io_dat_i[10]
+ cb_4_9/io_dat_i[11] cb_4_9/io_dat_i[12] cb_4_9/io_dat_i[13] cb_4_9/io_dat_i[14]
+ cb_4_9/io_dat_i[15] cb_4_9/io_dat_i[1] cb_4_9/io_dat_i[2] cb_4_9/io_dat_i[3] cb_4_9/io_dat_i[4]
+ cb_4_9/io_dat_i[5] cb_4_9/io_dat_i[6] cb_4_9/io_dat_i[7] cb_4_9/io_dat_i[8] cb_4_9/io_dat_i[9]
+ cb_4_8/io_dat_o[0] cb_4_8/io_dat_o[10] cb_4_8/io_dat_o[11] cb_4_8/io_dat_o[12] cb_4_8/io_dat_o[13]
+ cb_4_8/io_dat_o[14] cb_4_8/io_dat_o[15] cb_4_8/io_dat_o[1] cb_4_8/io_dat_o[2] cb_4_8/io_dat_o[3]
+ cb_4_8/io_dat_o[4] cb_4_8/io_dat_o[5] cb_4_8/io_dat_o[6] cb_4_8/io_dat_o[7] cb_4_8/io_dat_o[8]
+ cb_4_8/io_dat_o[9] cb_4_9/io_wo[0] cb_4_9/io_wo[10] cb_4_9/io_wo[11] cb_4_9/io_wo[12]
+ cb_4_9/io_wo[13] cb_4_9/io_wo[14] cb_4_9/io_wo[15] cb_4_9/io_wo[16] cb_4_9/io_wo[17]
+ cb_4_9/io_wo[18] cb_4_9/io_wo[19] cb_4_9/io_wo[1] cb_4_9/io_wo[20] cb_4_9/io_wo[21]
+ cb_4_9/io_wo[22] cb_4_9/io_wo[23] cb_4_9/io_wo[24] cb_4_9/io_wo[25] cb_4_9/io_wo[26]
+ cb_4_9/io_wo[27] cb_4_9/io_wo[28] cb_4_9/io_wo[29] cb_4_9/io_wo[2] cb_4_9/io_wo[30]
+ cb_4_9/io_wo[31] cb_4_9/io_wo[32] cb_4_9/io_wo[33] cb_4_9/io_wo[34] cb_4_9/io_wo[35]
+ cb_4_9/io_wo[36] cb_4_9/io_wo[37] cb_4_9/io_wo[38] cb_4_9/io_wo[39] cb_4_9/io_wo[3]
+ cb_4_9/io_wo[40] cb_4_9/io_wo[41] cb_4_9/io_wo[42] cb_4_9/io_wo[43] cb_4_9/io_wo[44]
+ cb_4_9/io_wo[45] cb_4_9/io_wo[46] cb_4_9/io_wo[47] cb_4_9/io_wo[48] cb_4_9/io_wo[49]
+ cb_4_9/io_wo[4] cb_4_9/io_wo[50] cb_4_9/io_wo[51] cb_4_9/io_wo[52] cb_4_9/io_wo[53]
+ cb_4_9/io_wo[54] cb_4_9/io_wo[55] cb_4_9/io_wo[56] cb_4_9/io_wo[57] cb_4_9/io_wo[58]
+ cb_4_9/io_wo[59] cb_4_9/io_wo[5] cb_4_9/io_wo[60] cb_4_9/io_wo[61] cb_4_9/io_wo[62]
+ cb_4_9/io_wo[63] cb_4_9/io_wo[6] cb_4_9/io_wo[7] cb_4_9/io_wo[8] cb_4_9/io_wo[9]
+ cb_4_8/io_i_0_ci cb_4_8/io_i_0_in1[0] cb_4_8/io_i_0_in1[1] cb_4_8/io_i_0_in1[2]
+ cb_4_8/io_i_0_in1[3] cb_4_8/io_i_0_in1[4] cb_4_8/io_i_0_in1[5] cb_4_8/io_i_0_in1[6]
+ cb_4_8/io_i_0_in1[7] cb_4_8/io_i_1_ci cb_4_8/io_i_1_in1[0] cb_4_8/io_i_1_in1[1]
+ cb_4_8/io_i_1_in1[2] cb_4_8/io_i_1_in1[3] cb_4_8/io_i_1_in1[4] cb_4_8/io_i_1_in1[5]
+ cb_4_8/io_i_1_in1[6] cb_4_8/io_i_1_in1[7] cb_4_8/io_i_2_ci cb_4_8/io_i_2_in1[0]
+ cb_4_8/io_i_2_in1[1] cb_4_8/io_i_2_in1[2] cb_4_8/io_i_2_in1[3] cb_4_8/io_i_2_in1[4]
+ cb_4_8/io_i_2_in1[5] cb_4_8/io_i_2_in1[6] cb_4_8/io_i_2_in1[7] cb_4_8/io_i_3_ci
+ cb_4_8/io_i_3_in1[0] cb_4_8/io_i_3_in1[1] cb_4_8/io_i_3_in1[2] cb_4_8/io_i_3_in1[3]
+ cb_4_8/io_i_3_in1[4] cb_4_8/io_i_3_in1[5] cb_4_8/io_i_3_in1[6] cb_4_8/io_i_3_in1[7]
+ cb_4_8/io_i_4_ci cb_4_8/io_i_4_in1[0] cb_4_8/io_i_4_in1[1] cb_4_8/io_i_4_in1[2]
+ cb_4_8/io_i_4_in1[3] cb_4_8/io_i_4_in1[4] cb_4_8/io_i_4_in1[5] cb_4_8/io_i_4_in1[6]
+ cb_4_8/io_i_4_in1[7] cb_4_8/io_i_5_ci cb_4_8/io_i_5_in1[0] cb_4_8/io_i_5_in1[1]
+ cb_4_8/io_i_5_in1[2] cb_4_8/io_i_5_in1[3] cb_4_8/io_i_5_in1[4] cb_4_8/io_i_5_in1[5]
+ cb_4_8/io_i_5_in1[6] cb_4_8/io_i_5_in1[7] cb_4_8/io_i_6_ci cb_4_8/io_i_6_in1[0]
+ cb_4_8/io_i_6_in1[1] cb_4_8/io_i_6_in1[2] cb_4_8/io_i_6_in1[3] cb_4_8/io_i_6_in1[4]
+ cb_4_8/io_i_6_in1[5] cb_4_8/io_i_6_in1[6] cb_4_8/io_i_6_in1[7] cb_4_8/io_i_7_ci
+ cb_4_8/io_i_7_in1[0] cb_4_8/io_i_7_in1[1] cb_4_8/io_i_7_in1[2] cb_4_8/io_i_7_in1[3]
+ cb_4_8/io_i_7_in1[4] cb_4_8/io_i_7_in1[5] cb_4_8/io_i_7_in1[6] cb_4_8/io_i_7_in1[7]
+ cb_4_9/io_i_0_ci cb_4_9/io_i_0_in1[0] cb_4_9/io_i_0_in1[1] cb_4_9/io_i_0_in1[2]
+ cb_4_9/io_i_0_in1[3] cb_4_9/io_i_0_in1[4] cb_4_9/io_i_0_in1[5] cb_4_9/io_i_0_in1[6]
+ cb_4_9/io_i_0_in1[7] cb_4_9/io_i_1_ci cb_4_9/io_i_1_in1[0] cb_4_9/io_i_1_in1[1]
+ cb_4_9/io_i_1_in1[2] cb_4_9/io_i_1_in1[3] cb_4_9/io_i_1_in1[4] cb_4_9/io_i_1_in1[5]
+ cb_4_9/io_i_1_in1[6] cb_4_9/io_i_1_in1[7] cb_4_9/io_i_2_ci cb_4_9/io_i_2_in1[0]
+ cb_4_9/io_i_2_in1[1] cb_4_9/io_i_2_in1[2] cb_4_9/io_i_2_in1[3] cb_4_9/io_i_2_in1[4]
+ cb_4_9/io_i_2_in1[5] cb_4_9/io_i_2_in1[6] cb_4_9/io_i_2_in1[7] cb_4_9/io_i_3_ci
+ cb_4_9/io_i_3_in1[0] cb_4_9/io_i_3_in1[1] cb_4_9/io_i_3_in1[2] cb_4_9/io_i_3_in1[3]
+ cb_4_9/io_i_3_in1[4] cb_4_9/io_i_3_in1[5] cb_4_9/io_i_3_in1[6] cb_4_9/io_i_3_in1[7]
+ cb_4_9/io_i_4_ci cb_4_9/io_i_4_in1[0] cb_4_9/io_i_4_in1[1] cb_4_9/io_i_4_in1[2]
+ cb_4_9/io_i_4_in1[3] cb_4_9/io_i_4_in1[4] cb_4_9/io_i_4_in1[5] cb_4_9/io_i_4_in1[6]
+ cb_4_9/io_i_4_in1[7] cb_4_9/io_i_5_ci cb_4_9/io_i_5_in1[0] cb_4_9/io_i_5_in1[1]
+ cb_4_9/io_i_5_in1[2] cb_4_9/io_i_5_in1[3] cb_4_9/io_i_5_in1[4] cb_4_9/io_i_5_in1[5]
+ cb_4_9/io_i_5_in1[6] cb_4_9/io_i_5_in1[7] cb_4_9/io_i_6_ci cb_4_9/io_i_6_in1[0]
+ cb_4_9/io_i_6_in1[1] cb_4_9/io_i_6_in1[2] cb_4_9/io_i_6_in1[3] cb_4_9/io_i_6_in1[4]
+ cb_4_9/io_i_6_in1[5] cb_4_9/io_i_6_in1[6] cb_4_9/io_i_6_in1[7] cb_4_9/io_i_7_ci
+ cb_4_9/io_i_7_in1[0] cb_4_9/io_i_7_in1[1] cb_4_9/io_i_7_in1[2] cb_4_9/io_i_7_in1[3]
+ cb_4_9/io_i_7_in1[4] cb_4_9/io_i_7_in1[5] cb_4_9/io_i_7_in1[6] cb_4_9/io_i_7_in1[7]
+ cb_4_8/io_vci cb_4_9/io_vci cb_4_8/io_vi cb_4_9/io_we_i cb_4_8/io_wo[0] cb_4_8/io_wo[10]
+ cb_4_8/io_wo[11] cb_4_8/io_wo[12] cb_4_8/io_wo[13] cb_4_8/io_wo[14] cb_4_8/io_wo[15]
+ cb_4_8/io_wo[16] cb_4_8/io_wo[17] cb_4_8/io_wo[18] cb_4_8/io_wo[19] cb_4_8/io_wo[1]
+ cb_4_8/io_wo[20] cb_4_8/io_wo[21] cb_4_8/io_wo[22] cb_4_8/io_wo[23] cb_4_8/io_wo[24]
+ cb_4_8/io_wo[25] cb_4_8/io_wo[26] cb_4_8/io_wo[27] cb_4_8/io_wo[28] cb_4_8/io_wo[29]
+ cb_4_8/io_wo[2] cb_4_8/io_wo[30] cb_4_8/io_wo[31] cb_4_8/io_wo[32] cb_4_8/io_wo[33]
+ cb_4_8/io_wo[34] cb_4_8/io_wo[35] cb_4_8/io_wo[36] cb_4_8/io_wo[37] cb_4_8/io_wo[38]
+ cb_4_8/io_wo[39] cb_4_8/io_wo[3] cb_4_8/io_wo[40] cb_4_8/io_wo[41] cb_4_8/io_wo[42]
+ cb_4_8/io_wo[43] cb_4_8/io_wo[44] cb_4_8/io_wo[45] cb_4_8/io_wo[46] cb_4_8/io_wo[47]
+ cb_4_8/io_wo[48] cb_4_8/io_wo[49] cb_4_8/io_wo[4] cb_4_8/io_wo[50] cb_4_8/io_wo[51]
+ cb_4_8/io_wo[52] cb_4_8/io_wo[53] cb_4_8/io_wo[54] cb_4_8/io_wo[55] cb_4_8/io_wo[56]
+ cb_4_8/io_wo[57] cb_4_8/io_wo[58] cb_4_8/io_wo[59] cb_4_8/io_wo[5] cb_4_8/io_wo[60]
+ cb_4_8/io_wo[61] cb_4_8/io_wo[62] cb_4_8/io_wo[63] cb_4_8/io_wo[6] cb_4_8/io_wo[7]
+ cb_4_8/io_wo[8] cb_4_8/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_2_5 cb_2_9/io_adr_i[0] cb_2_9/io_adr_i[1] cb_2_5/io_cs_i cb_2_9/io_dat_i[0] cb_2_9/io_dat_i[10]
+ cb_2_9/io_dat_i[11] cb_2_9/io_dat_i[12] cb_2_9/io_dat_i[13] cb_2_9/io_dat_i[14]
+ cb_2_9/io_dat_i[15] cb_2_9/io_dat_i[1] cb_2_9/io_dat_i[2] cb_2_9/io_dat_i[3] cb_2_9/io_dat_i[4]
+ cb_2_9/io_dat_i[5] cb_2_9/io_dat_i[6] cb_2_9/io_dat_i[7] cb_2_9/io_dat_i[8] cb_2_9/io_dat_i[9]
+ cb_2_5/io_dat_o[0] cb_2_5/io_dat_o[10] cb_2_5/io_dat_o[11] cb_2_5/io_dat_o[12] cb_2_5/io_dat_o[13]
+ cb_2_5/io_dat_o[14] cb_2_5/io_dat_o[15] cb_2_5/io_dat_o[1] cb_2_5/io_dat_o[2] cb_2_5/io_dat_o[3]
+ cb_2_5/io_dat_o[4] cb_2_5/io_dat_o[5] cb_2_5/io_dat_o[6] cb_2_5/io_dat_o[7] cb_2_5/io_dat_o[8]
+ cb_2_5/io_dat_o[9] cb_2_6/io_wo[0] cb_2_6/io_wo[10] cb_2_6/io_wo[11] cb_2_6/io_wo[12]
+ cb_2_6/io_wo[13] cb_2_6/io_wo[14] cb_2_6/io_wo[15] cb_2_6/io_wo[16] cb_2_6/io_wo[17]
+ cb_2_6/io_wo[18] cb_2_6/io_wo[19] cb_2_6/io_wo[1] cb_2_6/io_wo[20] cb_2_6/io_wo[21]
+ cb_2_6/io_wo[22] cb_2_6/io_wo[23] cb_2_6/io_wo[24] cb_2_6/io_wo[25] cb_2_6/io_wo[26]
+ cb_2_6/io_wo[27] cb_2_6/io_wo[28] cb_2_6/io_wo[29] cb_2_6/io_wo[2] cb_2_6/io_wo[30]
+ cb_2_6/io_wo[31] cb_2_6/io_wo[32] cb_2_6/io_wo[33] cb_2_6/io_wo[34] cb_2_6/io_wo[35]
+ cb_2_6/io_wo[36] cb_2_6/io_wo[37] cb_2_6/io_wo[38] cb_2_6/io_wo[39] cb_2_6/io_wo[3]
+ cb_2_6/io_wo[40] cb_2_6/io_wo[41] cb_2_6/io_wo[42] cb_2_6/io_wo[43] cb_2_6/io_wo[44]
+ cb_2_6/io_wo[45] cb_2_6/io_wo[46] cb_2_6/io_wo[47] cb_2_6/io_wo[48] cb_2_6/io_wo[49]
+ cb_2_6/io_wo[4] cb_2_6/io_wo[50] cb_2_6/io_wo[51] cb_2_6/io_wo[52] cb_2_6/io_wo[53]
+ cb_2_6/io_wo[54] cb_2_6/io_wo[55] cb_2_6/io_wo[56] cb_2_6/io_wo[57] cb_2_6/io_wo[58]
+ cb_2_6/io_wo[59] cb_2_6/io_wo[5] cb_2_6/io_wo[60] cb_2_6/io_wo[61] cb_2_6/io_wo[62]
+ cb_2_6/io_wo[63] cb_2_6/io_wo[6] cb_2_6/io_wo[7] cb_2_6/io_wo[8] cb_2_6/io_wo[9]
+ cb_2_5/io_i_0_ci cb_2_5/io_i_0_in1[0] cb_2_5/io_i_0_in1[1] cb_2_5/io_i_0_in1[2]
+ cb_2_5/io_i_0_in1[3] cb_2_5/io_i_0_in1[4] cb_2_5/io_i_0_in1[5] cb_2_5/io_i_0_in1[6]
+ cb_2_5/io_i_0_in1[7] cb_2_5/io_i_1_ci cb_2_5/io_i_1_in1[0] cb_2_5/io_i_1_in1[1]
+ cb_2_5/io_i_1_in1[2] cb_2_5/io_i_1_in1[3] cb_2_5/io_i_1_in1[4] cb_2_5/io_i_1_in1[5]
+ cb_2_5/io_i_1_in1[6] cb_2_5/io_i_1_in1[7] cb_2_5/io_i_2_ci cb_2_5/io_i_2_in1[0]
+ cb_2_5/io_i_2_in1[1] cb_2_5/io_i_2_in1[2] cb_2_5/io_i_2_in1[3] cb_2_5/io_i_2_in1[4]
+ cb_2_5/io_i_2_in1[5] cb_2_5/io_i_2_in1[6] cb_2_5/io_i_2_in1[7] cb_2_5/io_i_3_ci
+ cb_2_5/io_i_3_in1[0] cb_2_5/io_i_3_in1[1] cb_2_5/io_i_3_in1[2] cb_2_5/io_i_3_in1[3]
+ cb_2_5/io_i_3_in1[4] cb_2_5/io_i_3_in1[5] cb_2_5/io_i_3_in1[6] cb_2_5/io_i_3_in1[7]
+ cb_2_5/io_i_4_ci cb_2_5/io_i_4_in1[0] cb_2_5/io_i_4_in1[1] cb_2_5/io_i_4_in1[2]
+ cb_2_5/io_i_4_in1[3] cb_2_5/io_i_4_in1[4] cb_2_5/io_i_4_in1[5] cb_2_5/io_i_4_in1[6]
+ cb_2_5/io_i_4_in1[7] cb_2_5/io_i_5_ci cb_2_5/io_i_5_in1[0] cb_2_5/io_i_5_in1[1]
+ cb_2_5/io_i_5_in1[2] cb_2_5/io_i_5_in1[3] cb_2_5/io_i_5_in1[4] cb_2_5/io_i_5_in1[5]
+ cb_2_5/io_i_5_in1[6] cb_2_5/io_i_5_in1[7] cb_2_5/io_i_6_ci cb_2_5/io_i_6_in1[0]
+ cb_2_5/io_i_6_in1[1] cb_2_5/io_i_6_in1[2] cb_2_5/io_i_6_in1[3] cb_2_5/io_i_6_in1[4]
+ cb_2_5/io_i_6_in1[5] cb_2_5/io_i_6_in1[6] cb_2_5/io_i_6_in1[7] cb_2_5/io_i_7_ci
+ cb_2_5/io_i_7_in1[0] cb_2_5/io_i_7_in1[1] cb_2_5/io_i_7_in1[2] cb_2_5/io_i_7_in1[3]
+ cb_2_5/io_i_7_in1[4] cb_2_5/io_i_7_in1[5] cb_2_5/io_i_7_in1[6] cb_2_5/io_i_7_in1[7]
+ cb_2_6/io_i_0_ci cb_2_6/io_i_0_in1[0] cb_2_6/io_i_0_in1[1] cb_2_6/io_i_0_in1[2]
+ cb_2_6/io_i_0_in1[3] cb_2_6/io_i_0_in1[4] cb_2_6/io_i_0_in1[5] cb_2_6/io_i_0_in1[6]
+ cb_2_6/io_i_0_in1[7] cb_2_6/io_i_1_ci cb_2_6/io_i_1_in1[0] cb_2_6/io_i_1_in1[1]
+ cb_2_6/io_i_1_in1[2] cb_2_6/io_i_1_in1[3] cb_2_6/io_i_1_in1[4] cb_2_6/io_i_1_in1[5]
+ cb_2_6/io_i_1_in1[6] cb_2_6/io_i_1_in1[7] cb_2_6/io_i_2_ci cb_2_6/io_i_2_in1[0]
+ cb_2_6/io_i_2_in1[1] cb_2_6/io_i_2_in1[2] cb_2_6/io_i_2_in1[3] cb_2_6/io_i_2_in1[4]
+ cb_2_6/io_i_2_in1[5] cb_2_6/io_i_2_in1[6] cb_2_6/io_i_2_in1[7] cb_2_6/io_i_3_ci
+ cb_2_6/io_i_3_in1[0] cb_2_6/io_i_3_in1[1] cb_2_6/io_i_3_in1[2] cb_2_6/io_i_3_in1[3]
+ cb_2_6/io_i_3_in1[4] cb_2_6/io_i_3_in1[5] cb_2_6/io_i_3_in1[6] cb_2_6/io_i_3_in1[7]
+ cb_2_6/io_i_4_ci cb_2_6/io_i_4_in1[0] cb_2_6/io_i_4_in1[1] cb_2_6/io_i_4_in1[2]
+ cb_2_6/io_i_4_in1[3] cb_2_6/io_i_4_in1[4] cb_2_6/io_i_4_in1[5] cb_2_6/io_i_4_in1[6]
+ cb_2_6/io_i_4_in1[7] cb_2_6/io_i_5_ci cb_2_6/io_i_5_in1[0] cb_2_6/io_i_5_in1[1]
+ cb_2_6/io_i_5_in1[2] cb_2_6/io_i_5_in1[3] cb_2_6/io_i_5_in1[4] cb_2_6/io_i_5_in1[5]
+ cb_2_6/io_i_5_in1[6] cb_2_6/io_i_5_in1[7] cb_2_6/io_i_6_ci cb_2_6/io_i_6_in1[0]
+ cb_2_6/io_i_6_in1[1] cb_2_6/io_i_6_in1[2] cb_2_6/io_i_6_in1[3] cb_2_6/io_i_6_in1[4]
+ cb_2_6/io_i_6_in1[5] cb_2_6/io_i_6_in1[6] cb_2_6/io_i_6_in1[7] cb_2_6/io_i_7_ci
+ cb_2_6/io_i_7_in1[0] cb_2_6/io_i_7_in1[1] cb_2_6/io_i_7_in1[2] cb_2_6/io_i_7_in1[3]
+ cb_2_6/io_i_7_in1[4] cb_2_6/io_i_7_in1[5] cb_2_6/io_i_7_in1[6] cb_2_6/io_i_7_in1[7]
+ cb_2_5/io_vci cb_2_6/io_vci cb_2_5/io_vi cb_2_9/io_we_i cb_2_5/io_wo[0] cb_2_5/io_wo[10]
+ cb_2_5/io_wo[11] cb_2_5/io_wo[12] cb_2_5/io_wo[13] cb_2_5/io_wo[14] cb_2_5/io_wo[15]
+ cb_2_5/io_wo[16] cb_2_5/io_wo[17] cb_2_5/io_wo[18] cb_2_5/io_wo[19] cb_2_5/io_wo[1]
+ cb_2_5/io_wo[20] cb_2_5/io_wo[21] cb_2_5/io_wo[22] cb_2_5/io_wo[23] cb_2_5/io_wo[24]
+ cb_2_5/io_wo[25] cb_2_5/io_wo[26] cb_2_5/io_wo[27] cb_2_5/io_wo[28] cb_2_5/io_wo[29]
+ cb_2_5/io_wo[2] cb_2_5/io_wo[30] cb_2_5/io_wo[31] cb_2_5/io_wo[32] cb_2_5/io_wo[33]
+ cb_2_5/io_wo[34] cb_2_5/io_wo[35] cb_2_5/io_wo[36] cb_2_5/io_wo[37] cb_2_5/io_wo[38]
+ cb_2_5/io_wo[39] cb_2_5/io_wo[3] cb_2_5/io_wo[40] cb_2_5/io_wo[41] cb_2_5/io_wo[42]
+ cb_2_5/io_wo[43] cb_2_5/io_wo[44] cb_2_5/io_wo[45] cb_2_5/io_wo[46] cb_2_5/io_wo[47]
+ cb_2_5/io_wo[48] cb_2_5/io_wo[49] cb_2_5/io_wo[4] cb_2_5/io_wo[50] cb_2_5/io_wo[51]
+ cb_2_5/io_wo[52] cb_2_5/io_wo[53] cb_2_5/io_wo[54] cb_2_5/io_wo[55] cb_2_5/io_wo[56]
+ cb_2_5/io_wo[57] cb_2_5/io_wo[58] cb_2_5/io_wo[59] cb_2_5/io_wo[5] cb_2_5/io_wo[60]
+ cb_2_5/io_wo[61] cb_2_5/io_wo[62] cb_2_5/io_wo[63] cb_2_5/io_wo[6] cb_2_5/io_wo[7]
+ cb_2_5/io_wo[8] cb_2_5/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_0_2 cb_0_9/io_adr_i[0] cb_0_9/io_adr_i[1] cb_0_2/io_cs_i cb_0_9/io_dat_i[0] cb_0_9/io_dat_i[10]
+ cb_0_9/io_dat_i[11] cb_0_9/io_dat_i[12] cb_0_9/io_dat_i[13] cb_0_9/io_dat_i[14]
+ cb_0_9/io_dat_i[15] cb_0_9/io_dat_i[1] cb_0_9/io_dat_i[2] cb_0_9/io_dat_i[3] cb_0_9/io_dat_i[4]
+ cb_0_9/io_dat_i[5] cb_0_9/io_dat_i[6] cb_0_9/io_dat_i[7] cb_0_9/io_dat_i[8] cb_0_9/io_dat_i[9]
+ cb_0_2/io_dat_o[0] cb_0_2/io_dat_o[10] cb_0_2/io_dat_o[11] cb_0_2/io_dat_o[12] cb_0_2/io_dat_o[13]
+ cb_0_2/io_dat_o[14] cb_0_2/io_dat_o[15] cb_0_2/io_dat_o[1] cb_0_2/io_dat_o[2] cb_0_2/io_dat_o[3]
+ cb_0_2/io_dat_o[4] cb_0_2/io_dat_o[5] cb_0_2/io_dat_o[6] cb_0_2/io_dat_o[7] cb_0_2/io_dat_o[8]
+ cb_0_2/io_dat_o[9] cb_0_3/io_wo[0] cb_0_3/io_wo[10] cb_0_3/io_wo[11] cb_0_3/io_wo[12]
+ cb_0_3/io_wo[13] cb_0_3/io_wo[14] cb_0_3/io_wo[15] cb_0_3/io_wo[16] cb_0_3/io_wo[17]
+ cb_0_3/io_wo[18] cb_0_3/io_wo[19] cb_0_3/io_wo[1] cb_0_3/io_wo[20] cb_0_3/io_wo[21]
+ cb_0_3/io_wo[22] cb_0_3/io_wo[23] cb_0_3/io_wo[24] cb_0_3/io_wo[25] cb_0_3/io_wo[26]
+ cb_0_3/io_wo[27] cb_0_3/io_wo[28] cb_0_3/io_wo[29] cb_0_3/io_wo[2] cb_0_3/io_wo[30]
+ cb_0_3/io_wo[31] cb_0_3/io_wo[32] cb_0_3/io_wo[33] cb_0_3/io_wo[34] cb_0_3/io_wo[35]
+ cb_0_3/io_wo[36] cb_0_3/io_wo[37] cb_0_3/io_wo[38] cb_0_3/io_wo[39] cb_0_3/io_wo[3]
+ cb_0_3/io_wo[40] cb_0_3/io_wo[41] cb_0_3/io_wo[42] cb_0_3/io_wo[43] cb_0_3/io_wo[44]
+ cb_0_3/io_wo[45] cb_0_3/io_wo[46] cb_0_3/io_wo[47] cb_0_3/io_wo[48] cb_0_3/io_wo[49]
+ cb_0_3/io_wo[4] cb_0_3/io_wo[50] cb_0_3/io_wo[51] cb_0_3/io_wo[52] cb_0_3/io_wo[53]
+ cb_0_3/io_wo[54] cb_0_3/io_wo[55] cb_0_3/io_wo[56] cb_0_3/io_wo[57] cb_0_3/io_wo[58]
+ cb_0_3/io_wo[59] cb_0_3/io_wo[5] cb_0_3/io_wo[60] cb_0_3/io_wo[61] cb_0_3/io_wo[62]
+ cb_0_3/io_wo[63] cb_0_3/io_wo[6] cb_0_3/io_wo[7] cb_0_3/io_wo[8] cb_0_3/io_wo[9]
+ cb_0_2/io_i_0_ci cb_0_2/io_i_0_in1[0] cb_0_2/io_i_0_in1[1] cb_0_2/io_i_0_in1[2]
+ cb_0_2/io_i_0_in1[3] cb_0_2/io_i_0_in1[4] cb_0_2/io_i_0_in1[5] cb_0_2/io_i_0_in1[6]
+ cb_0_2/io_i_0_in1[7] cb_0_2/io_i_1_ci cb_0_2/io_i_1_in1[0] cb_0_2/io_i_1_in1[1]
+ cb_0_2/io_i_1_in1[2] cb_0_2/io_i_1_in1[3] cb_0_2/io_i_1_in1[4] cb_0_2/io_i_1_in1[5]
+ cb_0_2/io_i_1_in1[6] cb_0_2/io_i_1_in1[7] cb_0_2/io_i_2_ci cb_0_2/io_i_2_in1[0]
+ cb_0_2/io_i_2_in1[1] cb_0_2/io_i_2_in1[2] cb_0_2/io_i_2_in1[3] cb_0_2/io_i_2_in1[4]
+ cb_0_2/io_i_2_in1[5] cb_0_2/io_i_2_in1[6] cb_0_2/io_i_2_in1[7] cb_0_2/io_i_3_ci
+ cb_0_2/io_i_3_in1[0] cb_0_2/io_i_3_in1[1] cb_0_2/io_i_3_in1[2] cb_0_2/io_i_3_in1[3]
+ cb_0_2/io_i_3_in1[4] cb_0_2/io_i_3_in1[5] cb_0_2/io_i_3_in1[6] cb_0_2/io_i_3_in1[7]
+ cb_0_2/io_i_4_ci cb_0_2/io_i_4_in1[0] cb_0_2/io_i_4_in1[1] cb_0_2/io_i_4_in1[2]
+ cb_0_2/io_i_4_in1[3] cb_0_2/io_i_4_in1[4] cb_0_2/io_i_4_in1[5] cb_0_2/io_i_4_in1[6]
+ cb_0_2/io_i_4_in1[7] cb_0_2/io_i_5_ci cb_0_2/io_i_5_in1[0] cb_0_2/io_i_5_in1[1]
+ cb_0_2/io_i_5_in1[2] cb_0_2/io_i_5_in1[3] cb_0_2/io_i_5_in1[4] cb_0_2/io_i_5_in1[5]
+ cb_0_2/io_i_5_in1[6] cb_0_2/io_i_5_in1[7] cb_0_2/io_i_6_ci cb_0_2/io_i_6_in1[0]
+ cb_0_2/io_i_6_in1[1] cb_0_2/io_i_6_in1[2] cb_0_2/io_i_6_in1[3] cb_0_2/io_i_6_in1[4]
+ cb_0_2/io_i_6_in1[5] cb_0_2/io_i_6_in1[6] cb_0_2/io_i_6_in1[7] cb_0_2/io_i_7_ci
+ cb_0_2/io_i_7_in1[0] cb_0_2/io_i_7_in1[1] cb_0_2/io_i_7_in1[2] cb_0_2/io_i_7_in1[3]
+ cb_0_2/io_i_7_in1[4] cb_0_2/io_i_7_in1[5] cb_0_2/io_i_7_in1[6] cb_0_2/io_i_7_in1[7]
+ cb_0_3/io_i_0_ci cb_0_3/io_i_0_in1[0] cb_0_3/io_i_0_in1[1] cb_0_3/io_i_0_in1[2]
+ cb_0_3/io_i_0_in1[3] cb_0_3/io_i_0_in1[4] cb_0_3/io_i_0_in1[5] cb_0_3/io_i_0_in1[6]
+ cb_0_3/io_i_0_in1[7] cb_0_3/io_i_1_ci cb_0_3/io_i_1_in1[0] cb_0_3/io_i_1_in1[1]
+ cb_0_3/io_i_1_in1[2] cb_0_3/io_i_1_in1[3] cb_0_3/io_i_1_in1[4] cb_0_3/io_i_1_in1[5]
+ cb_0_3/io_i_1_in1[6] cb_0_3/io_i_1_in1[7] cb_0_3/io_i_2_ci cb_0_3/io_i_2_in1[0]
+ cb_0_3/io_i_2_in1[1] cb_0_3/io_i_2_in1[2] cb_0_3/io_i_2_in1[3] cb_0_3/io_i_2_in1[4]
+ cb_0_3/io_i_2_in1[5] cb_0_3/io_i_2_in1[6] cb_0_3/io_i_2_in1[7] cb_0_3/io_i_3_ci
+ cb_0_3/io_i_3_in1[0] cb_0_3/io_i_3_in1[1] cb_0_3/io_i_3_in1[2] cb_0_3/io_i_3_in1[3]
+ cb_0_3/io_i_3_in1[4] cb_0_3/io_i_3_in1[5] cb_0_3/io_i_3_in1[6] cb_0_3/io_i_3_in1[7]
+ cb_0_3/io_i_4_ci cb_0_3/io_i_4_in1[0] cb_0_3/io_i_4_in1[1] cb_0_3/io_i_4_in1[2]
+ cb_0_3/io_i_4_in1[3] cb_0_3/io_i_4_in1[4] cb_0_3/io_i_4_in1[5] cb_0_3/io_i_4_in1[6]
+ cb_0_3/io_i_4_in1[7] cb_0_3/io_i_5_ci cb_0_3/io_i_5_in1[0] cb_0_3/io_i_5_in1[1]
+ cb_0_3/io_i_5_in1[2] cb_0_3/io_i_5_in1[3] cb_0_3/io_i_5_in1[4] cb_0_3/io_i_5_in1[5]
+ cb_0_3/io_i_5_in1[6] cb_0_3/io_i_5_in1[7] cb_0_3/io_i_6_ci cb_0_3/io_i_6_in1[0]
+ cb_0_3/io_i_6_in1[1] cb_0_3/io_i_6_in1[2] cb_0_3/io_i_6_in1[3] cb_0_3/io_i_6_in1[4]
+ cb_0_3/io_i_6_in1[5] cb_0_3/io_i_6_in1[6] cb_0_3/io_i_6_in1[7] cb_0_3/io_i_7_ci
+ cb_0_3/io_i_7_in1[0] cb_0_3/io_i_7_in1[1] cb_0_3/io_i_7_in1[2] cb_0_3/io_i_7_in1[3]
+ cb_0_3/io_i_7_in1[4] cb_0_3/io_i_7_in1[5] cb_0_3/io_i_7_in1[6] cb_0_3/io_i_7_in1[7]
+ cb_0_2/io_vci cb_0_3/io_vci cb_0_2/io_vi cb_0_9/io_we_i cb_0_2/io_wo[0] cb_0_2/io_wo[10]
+ cb_0_2/io_wo[11] cb_0_2/io_wo[12] cb_0_2/io_wo[13] cb_0_2/io_wo[14] cb_0_2/io_wo[15]
+ cb_0_2/io_wo[16] cb_0_2/io_wo[17] cb_0_2/io_wo[18] cb_0_2/io_wo[19] cb_0_2/io_wo[1]
+ cb_0_2/io_wo[20] cb_0_2/io_wo[21] cb_0_2/io_wo[22] cb_0_2/io_wo[23] cb_0_2/io_wo[24]
+ cb_0_2/io_wo[25] cb_0_2/io_wo[26] cb_0_2/io_wo[27] cb_0_2/io_wo[28] cb_0_2/io_wo[29]
+ cb_0_2/io_wo[2] cb_0_2/io_wo[30] cb_0_2/io_wo[31] cb_0_2/io_wo[32] cb_0_2/io_wo[33]
+ cb_0_2/io_wo[34] cb_0_2/io_wo[35] cb_0_2/io_wo[36] cb_0_2/io_wo[37] cb_0_2/io_wo[38]
+ cb_0_2/io_wo[39] cb_0_2/io_wo[3] cb_0_2/io_wo[40] cb_0_2/io_wo[41] cb_0_2/io_wo[42]
+ cb_0_2/io_wo[43] cb_0_2/io_wo[44] cb_0_2/io_wo[45] cb_0_2/io_wo[46] cb_0_2/io_wo[47]
+ cb_0_2/io_wo[48] cb_0_2/io_wo[49] cb_0_2/io_wo[4] cb_0_2/io_wo[50] cb_0_2/io_wo[51]
+ cb_0_2/io_wo[52] cb_0_2/io_wo[53] cb_0_2/io_wo[54] cb_0_2/io_wo[55] cb_0_2/io_wo[56]
+ cb_0_2/io_wo[57] cb_0_2/io_wo[58] cb_0_2/io_wo[59] cb_0_2/io_wo[5] cb_0_2/io_wo[60]
+ cb_0_2/io_wo[61] cb_0_2/io_wo[62] cb_0_2/io_wo[63] cb_0_2/io_wo[6] cb_0_2/io_wo[7]
+ cb_0_2/io_wo[8] cb_0_2/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_4_9 cb_4_9/io_adr_i[0] cb_4_9/io_adr_i[1] cb_4_9/io_cs_i cb_4_9/io_dat_i[0] cb_4_9/io_dat_i[10]
+ cb_4_9/io_dat_i[11] cb_4_9/io_dat_i[12] cb_4_9/io_dat_i[13] cb_4_9/io_dat_i[14]
+ cb_4_9/io_dat_i[15] cb_4_9/io_dat_i[1] cb_4_9/io_dat_i[2] cb_4_9/io_dat_i[3] cb_4_9/io_dat_i[4]
+ cb_4_9/io_dat_i[5] cb_4_9/io_dat_i[6] cb_4_9/io_dat_i[7] cb_4_9/io_dat_i[8] cb_4_9/io_dat_i[9]
+ cb_4_9/io_dat_o[0] cb_4_9/io_dat_o[10] cb_4_9/io_dat_o[11] cb_4_9/io_dat_o[12] cb_4_9/io_dat_o[13]
+ cb_4_9/io_dat_o[14] cb_4_9/io_dat_o[15] cb_4_9/io_dat_o[1] cb_4_9/io_dat_o[2] cb_4_9/io_dat_o[3]
+ cb_4_9/io_dat_o[4] cb_4_9/io_dat_o[5] cb_4_9/io_dat_o[6] cb_4_9/io_dat_o[7] cb_4_9/io_dat_o[8]
+ cb_4_9/io_dat_o[9] cb_4_9/io_eo[0] cb_4_9/io_eo[10] cb_4_9/io_eo[11] cb_4_9/io_eo[12]
+ cb_4_9/io_eo[13] cb_4_9/io_eo[14] cb_4_9/io_eo[15] cb_4_9/io_eo[16] cb_4_9/io_eo[17]
+ cb_4_9/io_eo[18] cb_4_9/io_eo[19] cb_4_9/io_eo[1] cb_4_9/io_eo[20] cb_4_9/io_eo[21]
+ cb_4_9/io_eo[22] cb_4_9/io_eo[23] cb_4_9/io_eo[24] cb_4_9/io_eo[25] cb_4_9/io_eo[26]
+ cb_4_9/io_eo[27] cb_4_9/io_eo[28] cb_4_9/io_eo[29] cb_4_9/io_eo[2] cb_4_9/io_eo[30]
+ cb_4_9/io_eo[31] cb_4_9/io_eo[32] cb_4_9/io_eo[33] cb_4_9/io_eo[34] cb_4_9/io_eo[35]
+ cb_4_9/io_eo[36] cb_4_9/io_eo[37] cb_4_9/io_eo[38] cb_4_9/io_eo[39] cb_4_9/io_eo[3]
+ cb_4_9/io_eo[40] cb_4_9/io_eo[41] cb_4_9/io_eo[42] cb_4_9/io_eo[43] cb_4_9/io_eo[44]
+ cb_4_9/io_eo[45] cb_4_9/io_eo[46] cb_4_9/io_eo[47] cb_4_9/io_eo[48] cb_4_9/io_eo[49]
+ cb_4_9/io_eo[4] cb_4_9/io_eo[50] cb_4_9/io_eo[51] cb_4_9/io_eo[52] cb_4_9/io_eo[53]
+ cb_4_9/io_eo[54] cb_4_9/io_eo[55] cb_4_9/io_eo[56] cb_4_9/io_eo[57] cb_4_9/io_eo[58]
+ cb_4_9/io_eo[59] cb_4_9/io_eo[5] cb_4_9/io_eo[60] cb_4_9/io_eo[61] cb_4_9/io_eo[62]
+ cb_4_9/io_eo[63] cb_4_9/io_eo[6] cb_4_9/io_eo[7] cb_4_9/io_eo[8] cb_4_9/io_eo[9]
+ cb_4_9/io_i_0_ci cb_4_9/io_i_0_in1[0] cb_4_9/io_i_0_in1[1] cb_4_9/io_i_0_in1[2]
+ cb_4_9/io_i_0_in1[3] cb_4_9/io_i_0_in1[4] cb_4_9/io_i_0_in1[5] cb_4_9/io_i_0_in1[6]
+ cb_4_9/io_i_0_in1[7] cb_4_9/io_i_1_ci cb_4_9/io_i_1_in1[0] cb_4_9/io_i_1_in1[1]
+ cb_4_9/io_i_1_in1[2] cb_4_9/io_i_1_in1[3] cb_4_9/io_i_1_in1[4] cb_4_9/io_i_1_in1[5]
+ cb_4_9/io_i_1_in1[6] cb_4_9/io_i_1_in1[7] cb_4_9/io_i_2_ci cb_4_9/io_i_2_in1[0]
+ cb_4_9/io_i_2_in1[1] cb_4_9/io_i_2_in1[2] cb_4_9/io_i_2_in1[3] cb_4_9/io_i_2_in1[4]
+ cb_4_9/io_i_2_in1[5] cb_4_9/io_i_2_in1[6] cb_4_9/io_i_2_in1[7] cb_4_9/io_i_3_ci
+ cb_4_9/io_i_3_in1[0] cb_4_9/io_i_3_in1[1] cb_4_9/io_i_3_in1[2] cb_4_9/io_i_3_in1[3]
+ cb_4_9/io_i_3_in1[4] cb_4_9/io_i_3_in1[5] cb_4_9/io_i_3_in1[6] cb_4_9/io_i_3_in1[7]
+ cb_4_9/io_i_4_ci cb_4_9/io_i_4_in1[0] cb_4_9/io_i_4_in1[1] cb_4_9/io_i_4_in1[2]
+ cb_4_9/io_i_4_in1[3] cb_4_9/io_i_4_in1[4] cb_4_9/io_i_4_in1[5] cb_4_9/io_i_4_in1[6]
+ cb_4_9/io_i_4_in1[7] cb_4_9/io_i_5_ci cb_4_9/io_i_5_in1[0] cb_4_9/io_i_5_in1[1]
+ cb_4_9/io_i_5_in1[2] cb_4_9/io_i_5_in1[3] cb_4_9/io_i_5_in1[4] cb_4_9/io_i_5_in1[5]
+ cb_4_9/io_i_5_in1[6] cb_4_9/io_i_5_in1[7] cb_4_9/io_i_6_ci cb_4_9/io_i_6_in1[0]
+ cb_4_9/io_i_6_in1[1] cb_4_9/io_i_6_in1[2] cb_4_9/io_i_6_in1[3] cb_4_9/io_i_6_in1[4]
+ cb_4_9/io_i_6_in1[5] cb_4_9/io_i_6_in1[6] cb_4_9/io_i_6_in1[7] cb_4_9/io_i_7_ci
+ cb_4_9/io_i_7_in1[0] cb_4_9/io_i_7_in1[1] cb_4_9/io_i_7_in1[2] cb_4_9/io_i_7_in1[3]
+ cb_4_9/io_i_7_in1[4] cb_4_9/io_i_7_in1[5] cb_4_9/io_i_7_in1[6] cb_4_9/io_i_7_in1[7]
+ cb_4_9/io_o_0_co cb_4_9/io_o_0_out[0] cb_4_9/io_o_0_out[1] cb_4_9/io_o_0_out[2]
+ cb_4_9/io_o_0_out[3] cb_4_9/io_o_0_out[4] cb_4_9/io_o_0_out[5] cb_4_9/io_o_0_out[6]
+ cb_4_9/io_o_0_out[7] cb_4_9/io_o_1_co cb_4_9/io_o_1_out[0] cb_4_9/io_o_1_out[1]
+ cb_4_9/io_o_1_out[2] cb_4_9/io_o_1_out[3] cb_4_9/io_o_1_out[4] cb_4_9/io_o_1_out[5]
+ cb_4_9/io_o_1_out[6] cb_4_9/io_o_1_out[7] cb_4_9/io_o_2_co cb_4_9/io_o_2_out[0]
+ cb_4_9/io_o_2_out[1] cb_4_9/io_o_2_out[2] cb_4_9/io_o_2_out[3] cb_4_9/io_o_2_out[4]
+ cb_4_9/io_o_2_out[5] cb_4_9/io_o_2_out[6] cb_4_9/io_o_2_out[7] cb_4_9/io_o_3_co
+ cb_4_9/io_o_3_out[0] cb_4_9/io_o_3_out[1] cb_4_9/io_o_3_out[2] cb_4_9/io_o_3_out[3]
+ cb_4_9/io_o_3_out[4] cb_4_9/io_o_3_out[5] cb_4_9/io_o_3_out[6] cb_4_9/io_o_3_out[7]
+ cb_4_9/io_o_4_co cb_4_9/io_o_4_out[0] cb_4_9/io_o_4_out[1] cb_4_9/io_o_4_out[2]
+ cb_4_9/io_o_4_out[3] cb_4_9/io_o_4_out[4] cb_4_9/io_o_4_out[5] cb_4_9/io_o_4_out[6]
+ cb_4_9/io_o_4_out[7] cb_4_9/io_o_5_co cb_4_9/io_o_5_out[0] cb_4_9/io_o_5_out[1]
+ cb_4_9/io_o_5_out[2] cb_4_9/io_o_5_out[3] cb_4_9/io_o_5_out[4] cb_4_9/io_o_5_out[5]
+ cb_4_9/io_o_5_out[6] cb_4_9/io_o_5_out[7] cb_4_9/io_o_6_co cb_4_9/io_o_6_out[0]
+ cb_4_9/io_o_6_out[1] cb_4_9/io_o_6_out[2] cb_4_9/io_o_6_out[3] cb_4_9/io_o_6_out[4]
+ cb_4_9/io_o_6_out[5] cb_4_9/io_o_6_out[6] cb_4_9/io_o_6_out[7] cb_4_9/io_o_7_co
+ cb_4_9/io_o_7_out[0] cb_4_9/io_o_7_out[1] cb_4_9/io_o_7_out[2] cb_4_9/io_o_7_out[3]
+ cb_4_9/io_o_7_out[4] cb_4_9/io_o_7_out[5] cb_4_9/io_o_7_out[6] cb_4_9/io_o_7_out[7]
+ cb_4_9/io_vci cb_4_9/io_vco cb_4_9/io_vi cb_4_9/io_we_i cb_4_9/io_wo[0] cb_4_9/io_wo[10]
+ cb_4_9/io_wo[11] cb_4_9/io_wo[12] cb_4_9/io_wo[13] cb_4_9/io_wo[14] cb_4_9/io_wo[15]
+ cb_4_9/io_wo[16] cb_4_9/io_wo[17] cb_4_9/io_wo[18] cb_4_9/io_wo[19] cb_4_9/io_wo[1]
+ cb_4_9/io_wo[20] cb_4_9/io_wo[21] cb_4_9/io_wo[22] cb_4_9/io_wo[23] cb_4_9/io_wo[24]
+ cb_4_9/io_wo[25] cb_4_9/io_wo[26] cb_4_9/io_wo[27] cb_4_9/io_wo[28] cb_4_9/io_wo[29]
+ cb_4_9/io_wo[2] cb_4_9/io_wo[30] cb_4_9/io_wo[31] cb_4_9/io_wo[32] cb_4_9/io_wo[33]
+ cb_4_9/io_wo[34] cb_4_9/io_wo[35] cb_4_9/io_wo[36] cb_4_9/io_wo[37] cb_4_9/io_wo[38]
+ cb_4_9/io_wo[39] cb_4_9/io_wo[3] cb_4_9/io_wo[40] cb_4_9/io_wo[41] cb_4_9/io_wo[42]
+ cb_4_9/io_wo[43] cb_4_9/io_wo[44] cb_4_9/io_wo[45] cb_4_9/io_wo[46] cb_4_9/io_wo[47]
+ cb_4_9/io_wo[48] cb_4_9/io_wo[49] cb_4_9/io_wo[4] cb_4_9/io_wo[50] cb_4_9/io_wo[51]
+ cb_4_9/io_wo[52] cb_4_9/io_wo[53] cb_4_9/io_wo[54] cb_4_9/io_wo[55] cb_4_9/io_wo[56]
+ cb_4_9/io_wo[57] cb_4_9/io_wo[58] cb_4_9/io_wo[59] cb_4_9/io_wo[5] cb_4_9/io_wo[60]
+ cb_4_9/io_wo[61] cb_4_9/io_wo[62] cb_4_9/io_wo[63] cb_4_9/io_wo[6] cb_4_9/io_wo[7]
+ cb_4_9/io_wo[8] cb_4_9/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_2_6 cb_2_9/io_adr_i[0] cb_2_9/io_adr_i[1] cb_2_6/io_cs_i cb_2_9/io_dat_i[0] cb_2_9/io_dat_i[10]
+ cb_2_9/io_dat_i[11] cb_2_9/io_dat_i[12] cb_2_9/io_dat_i[13] cb_2_9/io_dat_i[14]
+ cb_2_9/io_dat_i[15] cb_2_9/io_dat_i[1] cb_2_9/io_dat_i[2] cb_2_9/io_dat_i[3] cb_2_9/io_dat_i[4]
+ cb_2_9/io_dat_i[5] cb_2_9/io_dat_i[6] cb_2_9/io_dat_i[7] cb_2_9/io_dat_i[8] cb_2_9/io_dat_i[9]
+ cb_2_6/io_dat_o[0] cb_2_6/io_dat_o[10] cb_2_6/io_dat_o[11] cb_2_6/io_dat_o[12] cb_2_6/io_dat_o[13]
+ cb_2_6/io_dat_o[14] cb_2_6/io_dat_o[15] cb_2_6/io_dat_o[1] cb_2_6/io_dat_o[2] cb_2_6/io_dat_o[3]
+ cb_2_6/io_dat_o[4] cb_2_6/io_dat_o[5] cb_2_6/io_dat_o[6] cb_2_6/io_dat_o[7] cb_2_6/io_dat_o[8]
+ cb_2_6/io_dat_o[9] cb_2_7/io_wo[0] cb_2_7/io_wo[10] cb_2_7/io_wo[11] cb_2_7/io_wo[12]
+ cb_2_7/io_wo[13] cb_2_7/io_wo[14] cb_2_7/io_wo[15] cb_2_7/io_wo[16] cb_2_7/io_wo[17]
+ cb_2_7/io_wo[18] cb_2_7/io_wo[19] cb_2_7/io_wo[1] cb_2_7/io_wo[20] cb_2_7/io_wo[21]
+ cb_2_7/io_wo[22] cb_2_7/io_wo[23] cb_2_7/io_wo[24] cb_2_7/io_wo[25] cb_2_7/io_wo[26]
+ cb_2_7/io_wo[27] cb_2_7/io_wo[28] cb_2_7/io_wo[29] cb_2_7/io_wo[2] cb_2_7/io_wo[30]
+ cb_2_7/io_wo[31] cb_2_7/io_wo[32] cb_2_7/io_wo[33] cb_2_7/io_wo[34] cb_2_7/io_wo[35]
+ cb_2_7/io_wo[36] cb_2_7/io_wo[37] cb_2_7/io_wo[38] cb_2_7/io_wo[39] cb_2_7/io_wo[3]
+ cb_2_7/io_wo[40] cb_2_7/io_wo[41] cb_2_7/io_wo[42] cb_2_7/io_wo[43] cb_2_7/io_wo[44]
+ cb_2_7/io_wo[45] cb_2_7/io_wo[46] cb_2_7/io_wo[47] cb_2_7/io_wo[48] cb_2_7/io_wo[49]
+ cb_2_7/io_wo[4] cb_2_7/io_wo[50] cb_2_7/io_wo[51] cb_2_7/io_wo[52] cb_2_7/io_wo[53]
+ cb_2_7/io_wo[54] cb_2_7/io_wo[55] cb_2_7/io_wo[56] cb_2_7/io_wo[57] cb_2_7/io_wo[58]
+ cb_2_7/io_wo[59] cb_2_7/io_wo[5] cb_2_7/io_wo[60] cb_2_7/io_wo[61] cb_2_7/io_wo[62]
+ cb_2_7/io_wo[63] cb_2_7/io_wo[6] cb_2_7/io_wo[7] cb_2_7/io_wo[8] cb_2_7/io_wo[9]
+ cb_2_6/io_i_0_ci cb_2_6/io_i_0_in1[0] cb_2_6/io_i_0_in1[1] cb_2_6/io_i_0_in1[2]
+ cb_2_6/io_i_0_in1[3] cb_2_6/io_i_0_in1[4] cb_2_6/io_i_0_in1[5] cb_2_6/io_i_0_in1[6]
+ cb_2_6/io_i_0_in1[7] cb_2_6/io_i_1_ci cb_2_6/io_i_1_in1[0] cb_2_6/io_i_1_in1[1]
+ cb_2_6/io_i_1_in1[2] cb_2_6/io_i_1_in1[3] cb_2_6/io_i_1_in1[4] cb_2_6/io_i_1_in1[5]
+ cb_2_6/io_i_1_in1[6] cb_2_6/io_i_1_in1[7] cb_2_6/io_i_2_ci cb_2_6/io_i_2_in1[0]
+ cb_2_6/io_i_2_in1[1] cb_2_6/io_i_2_in1[2] cb_2_6/io_i_2_in1[3] cb_2_6/io_i_2_in1[4]
+ cb_2_6/io_i_2_in1[5] cb_2_6/io_i_2_in1[6] cb_2_6/io_i_2_in1[7] cb_2_6/io_i_3_ci
+ cb_2_6/io_i_3_in1[0] cb_2_6/io_i_3_in1[1] cb_2_6/io_i_3_in1[2] cb_2_6/io_i_3_in1[3]
+ cb_2_6/io_i_3_in1[4] cb_2_6/io_i_3_in1[5] cb_2_6/io_i_3_in1[6] cb_2_6/io_i_3_in1[7]
+ cb_2_6/io_i_4_ci cb_2_6/io_i_4_in1[0] cb_2_6/io_i_4_in1[1] cb_2_6/io_i_4_in1[2]
+ cb_2_6/io_i_4_in1[3] cb_2_6/io_i_4_in1[4] cb_2_6/io_i_4_in1[5] cb_2_6/io_i_4_in1[6]
+ cb_2_6/io_i_4_in1[7] cb_2_6/io_i_5_ci cb_2_6/io_i_5_in1[0] cb_2_6/io_i_5_in1[1]
+ cb_2_6/io_i_5_in1[2] cb_2_6/io_i_5_in1[3] cb_2_6/io_i_5_in1[4] cb_2_6/io_i_5_in1[5]
+ cb_2_6/io_i_5_in1[6] cb_2_6/io_i_5_in1[7] cb_2_6/io_i_6_ci cb_2_6/io_i_6_in1[0]
+ cb_2_6/io_i_6_in1[1] cb_2_6/io_i_6_in1[2] cb_2_6/io_i_6_in1[3] cb_2_6/io_i_6_in1[4]
+ cb_2_6/io_i_6_in1[5] cb_2_6/io_i_6_in1[6] cb_2_6/io_i_6_in1[7] cb_2_6/io_i_7_ci
+ cb_2_6/io_i_7_in1[0] cb_2_6/io_i_7_in1[1] cb_2_6/io_i_7_in1[2] cb_2_6/io_i_7_in1[3]
+ cb_2_6/io_i_7_in1[4] cb_2_6/io_i_7_in1[5] cb_2_6/io_i_7_in1[6] cb_2_6/io_i_7_in1[7]
+ cb_2_7/io_i_0_ci cb_2_7/io_i_0_in1[0] cb_2_7/io_i_0_in1[1] cb_2_7/io_i_0_in1[2]
+ cb_2_7/io_i_0_in1[3] cb_2_7/io_i_0_in1[4] cb_2_7/io_i_0_in1[5] cb_2_7/io_i_0_in1[6]
+ cb_2_7/io_i_0_in1[7] cb_2_7/io_i_1_ci cb_2_7/io_i_1_in1[0] cb_2_7/io_i_1_in1[1]
+ cb_2_7/io_i_1_in1[2] cb_2_7/io_i_1_in1[3] cb_2_7/io_i_1_in1[4] cb_2_7/io_i_1_in1[5]
+ cb_2_7/io_i_1_in1[6] cb_2_7/io_i_1_in1[7] cb_2_7/io_i_2_ci cb_2_7/io_i_2_in1[0]
+ cb_2_7/io_i_2_in1[1] cb_2_7/io_i_2_in1[2] cb_2_7/io_i_2_in1[3] cb_2_7/io_i_2_in1[4]
+ cb_2_7/io_i_2_in1[5] cb_2_7/io_i_2_in1[6] cb_2_7/io_i_2_in1[7] cb_2_7/io_i_3_ci
+ cb_2_7/io_i_3_in1[0] cb_2_7/io_i_3_in1[1] cb_2_7/io_i_3_in1[2] cb_2_7/io_i_3_in1[3]
+ cb_2_7/io_i_3_in1[4] cb_2_7/io_i_3_in1[5] cb_2_7/io_i_3_in1[6] cb_2_7/io_i_3_in1[7]
+ cb_2_7/io_i_4_ci cb_2_7/io_i_4_in1[0] cb_2_7/io_i_4_in1[1] cb_2_7/io_i_4_in1[2]
+ cb_2_7/io_i_4_in1[3] cb_2_7/io_i_4_in1[4] cb_2_7/io_i_4_in1[5] cb_2_7/io_i_4_in1[6]
+ cb_2_7/io_i_4_in1[7] cb_2_7/io_i_5_ci cb_2_7/io_i_5_in1[0] cb_2_7/io_i_5_in1[1]
+ cb_2_7/io_i_5_in1[2] cb_2_7/io_i_5_in1[3] cb_2_7/io_i_5_in1[4] cb_2_7/io_i_5_in1[5]
+ cb_2_7/io_i_5_in1[6] cb_2_7/io_i_5_in1[7] cb_2_7/io_i_6_ci cb_2_7/io_i_6_in1[0]
+ cb_2_7/io_i_6_in1[1] cb_2_7/io_i_6_in1[2] cb_2_7/io_i_6_in1[3] cb_2_7/io_i_6_in1[4]
+ cb_2_7/io_i_6_in1[5] cb_2_7/io_i_6_in1[6] cb_2_7/io_i_6_in1[7] cb_2_7/io_i_7_ci
+ cb_2_7/io_i_7_in1[0] cb_2_7/io_i_7_in1[1] cb_2_7/io_i_7_in1[2] cb_2_7/io_i_7_in1[3]
+ cb_2_7/io_i_7_in1[4] cb_2_7/io_i_7_in1[5] cb_2_7/io_i_7_in1[6] cb_2_7/io_i_7_in1[7]
+ cb_2_6/io_vci cb_2_7/io_vci cb_2_6/io_vi cb_2_9/io_we_i cb_2_6/io_wo[0] cb_2_6/io_wo[10]
+ cb_2_6/io_wo[11] cb_2_6/io_wo[12] cb_2_6/io_wo[13] cb_2_6/io_wo[14] cb_2_6/io_wo[15]
+ cb_2_6/io_wo[16] cb_2_6/io_wo[17] cb_2_6/io_wo[18] cb_2_6/io_wo[19] cb_2_6/io_wo[1]
+ cb_2_6/io_wo[20] cb_2_6/io_wo[21] cb_2_6/io_wo[22] cb_2_6/io_wo[23] cb_2_6/io_wo[24]
+ cb_2_6/io_wo[25] cb_2_6/io_wo[26] cb_2_6/io_wo[27] cb_2_6/io_wo[28] cb_2_6/io_wo[29]
+ cb_2_6/io_wo[2] cb_2_6/io_wo[30] cb_2_6/io_wo[31] cb_2_6/io_wo[32] cb_2_6/io_wo[33]
+ cb_2_6/io_wo[34] cb_2_6/io_wo[35] cb_2_6/io_wo[36] cb_2_6/io_wo[37] cb_2_6/io_wo[38]
+ cb_2_6/io_wo[39] cb_2_6/io_wo[3] cb_2_6/io_wo[40] cb_2_6/io_wo[41] cb_2_6/io_wo[42]
+ cb_2_6/io_wo[43] cb_2_6/io_wo[44] cb_2_6/io_wo[45] cb_2_6/io_wo[46] cb_2_6/io_wo[47]
+ cb_2_6/io_wo[48] cb_2_6/io_wo[49] cb_2_6/io_wo[4] cb_2_6/io_wo[50] cb_2_6/io_wo[51]
+ cb_2_6/io_wo[52] cb_2_6/io_wo[53] cb_2_6/io_wo[54] cb_2_6/io_wo[55] cb_2_6/io_wo[56]
+ cb_2_6/io_wo[57] cb_2_6/io_wo[58] cb_2_6/io_wo[59] cb_2_6/io_wo[5] cb_2_6/io_wo[60]
+ cb_2_6/io_wo[61] cb_2_6/io_wo[62] cb_2_6/io_wo[63] cb_2_6/io_wo[6] cb_2_6/io_wo[7]
+ cb_2_6/io_wo[8] cb_2_6/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_0_3 cb_0_9/io_adr_i[0] cb_0_9/io_adr_i[1] cb_0_3/io_cs_i cb_0_9/io_dat_i[0] cb_0_9/io_dat_i[10]
+ cb_0_9/io_dat_i[11] cb_0_9/io_dat_i[12] cb_0_9/io_dat_i[13] cb_0_9/io_dat_i[14]
+ cb_0_9/io_dat_i[15] cb_0_9/io_dat_i[1] cb_0_9/io_dat_i[2] cb_0_9/io_dat_i[3] cb_0_9/io_dat_i[4]
+ cb_0_9/io_dat_i[5] cb_0_9/io_dat_i[6] cb_0_9/io_dat_i[7] cb_0_9/io_dat_i[8] cb_0_9/io_dat_i[9]
+ cb_0_3/io_dat_o[0] cb_0_3/io_dat_o[10] cb_0_3/io_dat_o[11] cb_0_3/io_dat_o[12] cb_0_3/io_dat_o[13]
+ cb_0_3/io_dat_o[14] cb_0_3/io_dat_o[15] cb_0_3/io_dat_o[1] cb_0_3/io_dat_o[2] cb_0_3/io_dat_o[3]
+ cb_0_3/io_dat_o[4] cb_0_3/io_dat_o[5] cb_0_3/io_dat_o[6] cb_0_3/io_dat_o[7] cb_0_3/io_dat_o[8]
+ cb_0_3/io_dat_o[9] cb_0_4/io_wo[0] cb_0_4/io_wo[10] cb_0_4/io_wo[11] cb_0_4/io_wo[12]
+ cb_0_4/io_wo[13] cb_0_4/io_wo[14] cb_0_4/io_wo[15] cb_0_4/io_wo[16] cb_0_4/io_wo[17]
+ cb_0_4/io_wo[18] cb_0_4/io_wo[19] cb_0_4/io_wo[1] cb_0_4/io_wo[20] cb_0_4/io_wo[21]
+ cb_0_4/io_wo[22] cb_0_4/io_wo[23] cb_0_4/io_wo[24] cb_0_4/io_wo[25] cb_0_4/io_wo[26]
+ cb_0_4/io_wo[27] cb_0_4/io_wo[28] cb_0_4/io_wo[29] cb_0_4/io_wo[2] cb_0_4/io_wo[30]
+ cb_0_4/io_wo[31] cb_0_4/io_wo[32] cb_0_4/io_wo[33] cb_0_4/io_wo[34] cb_0_4/io_wo[35]
+ cb_0_4/io_wo[36] cb_0_4/io_wo[37] cb_0_4/io_wo[38] cb_0_4/io_wo[39] cb_0_4/io_wo[3]
+ cb_0_4/io_wo[40] cb_0_4/io_wo[41] cb_0_4/io_wo[42] cb_0_4/io_wo[43] cb_0_4/io_wo[44]
+ cb_0_4/io_wo[45] cb_0_4/io_wo[46] cb_0_4/io_wo[47] cb_0_4/io_wo[48] cb_0_4/io_wo[49]
+ cb_0_4/io_wo[4] cb_0_4/io_wo[50] cb_0_4/io_wo[51] cb_0_4/io_wo[52] cb_0_4/io_wo[53]
+ cb_0_4/io_wo[54] cb_0_4/io_wo[55] cb_0_4/io_wo[56] cb_0_4/io_wo[57] cb_0_4/io_wo[58]
+ cb_0_4/io_wo[59] cb_0_4/io_wo[5] cb_0_4/io_wo[60] cb_0_4/io_wo[61] cb_0_4/io_wo[62]
+ cb_0_4/io_wo[63] cb_0_4/io_wo[6] cb_0_4/io_wo[7] cb_0_4/io_wo[8] cb_0_4/io_wo[9]
+ cb_0_3/io_i_0_ci cb_0_3/io_i_0_in1[0] cb_0_3/io_i_0_in1[1] cb_0_3/io_i_0_in1[2]
+ cb_0_3/io_i_0_in1[3] cb_0_3/io_i_0_in1[4] cb_0_3/io_i_0_in1[5] cb_0_3/io_i_0_in1[6]
+ cb_0_3/io_i_0_in1[7] cb_0_3/io_i_1_ci cb_0_3/io_i_1_in1[0] cb_0_3/io_i_1_in1[1]
+ cb_0_3/io_i_1_in1[2] cb_0_3/io_i_1_in1[3] cb_0_3/io_i_1_in1[4] cb_0_3/io_i_1_in1[5]
+ cb_0_3/io_i_1_in1[6] cb_0_3/io_i_1_in1[7] cb_0_3/io_i_2_ci cb_0_3/io_i_2_in1[0]
+ cb_0_3/io_i_2_in1[1] cb_0_3/io_i_2_in1[2] cb_0_3/io_i_2_in1[3] cb_0_3/io_i_2_in1[4]
+ cb_0_3/io_i_2_in1[5] cb_0_3/io_i_2_in1[6] cb_0_3/io_i_2_in1[7] cb_0_3/io_i_3_ci
+ cb_0_3/io_i_3_in1[0] cb_0_3/io_i_3_in1[1] cb_0_3/io_i_3_in1[2] cb_0_3/io_i_3_in1[3]
+ cb_0_3/io_i_3_in1[4] cb_0_3/io_i_3_in1[5] cb_0_3/io_i_3_in1[6] cb_0_3/io_i_3_in1[7]
+ cb_0_3/io_i_4_ci cb_0_3/io_i_4_in1[0] cb_0_3/io_i_4_in1[1] cb_0_3/io_i_4_in1[2]
+ cb_0_3/io_i_4_in1[3] cb_0_3/io_i_4_in1[4] cb_0_3/io_i_4_in1[5] cb_0_3/io_i_4_in1[6]
+ cb_0_3/io_i_4_in1[7] cb_0_3/io_i_5_ci cb_0_3/io_i_5_in1[0] cb_0_3/io_i_5_in1[1]
+ cb_0_3/io_i_5_in1[2] cb_0_3/io_i_5_in1[3] cb_0_3/io_i_5_in1[4] cb_0_3/io_i_5_in1[5]
+ cb_0_3/io_i_5_in1[6] cb_0_3/io_i_5_in1[7] cb_0_3/io_i_6_ci cb_0_3/io_i_6_in1[0]
+ cb_0_3/io_i_6_in1[1] cb_0_3/io_i_6_in1[2] cb_0_3/io_i_6_in1[3] cb_0_3/io_i_6_in1[4]
+ cb_0_3/io_i_6_in1[5] cb_0_3/io_i_6_in1[6] cb_0_3/io_i_6_in1[7] cb_0_3/io_i_7_ci
+ cb_0_3/io_i_7_in1[0] cb_0_3/io_i_7_in1[1] cb_0_3/io_i_7_in1[2] cb_0_3/io_i_7_in1[3]
+ cb_0_3/io_i_7_in1[4] cb_0_3/io_i_7_in1[5] cb_0_3/io_i_7_in1[6] cb_0_3/io_i_7_in1[7]
+ cb_0_4/io_i_0_ci cb_0_4/io_i_0_in1[0] cb_0_4/io_i_0_in1[1] cb_0_4/io_i_0_in1[2]
+ cb_0_4/io_i_0_in1[3] cb_0_4/io_i_0_in1[4] cb_0_4/io_i_0_in1[5] cb_0_4/io_i_0_in1[6]
+ cb_0_4/io_i_0_in1[7] cb_0_4/io_i_1_ci cb_0_4/io_i_1_in1[0] cb_0_4/io_i_1_in1[1]
+ cb_0_4/io_i_1_in1[2] cb_0_4/io_i_1_in1[3] cb_0_4/io_i_1_in1[4] cb_0_4/io_i_1_in1[5]
+ cb_0_4/io_i_1_in1[6] cb_0_4/io_i_1_in1[7] cb_0_4/io_i_2_ci cb_0_4/io_i_2_in1[0]
+ cb_0_4/io_i_2_in1[1] cb_0_4/io_i_2_in1[2] cb_0_4/io_i_2_in1[3] cb_0_4/io_i_2_in1[4]
+ cb_0_4/io_i_2_in1[5] cb_0_4/io_i_2_in1[6] cb_0_4/io_i_2_in1[7] cb_0_4/io_i_3_ci
+ cb_0_4/io_i_3_in1[0] cb_0_4/io_i_3_in1[1] cb_0_4/io_i_3_in1[2] cb_0_4/io_i_3_in1[3]
+ cb_0_4/io_i_3_in1[4] cb_0_4/io_i_3_in1[5] cb_0_4/io_i_3_in1[6] cb_0_4/io_i_3_in1[7]
+ cb_0_4/io_i_4_ci cb_0_4/io_i_4_in1[0] cb_0_4/io_i_4_in1[1] cb_0_4/io_i_4_in1[2]
+ cb_0_4/io_i_4_in1[3] cb_0_4/io_i_4_in1[4] cb_0_4/io_i_4_in1[5] cb_0_4/io_i_4_in1[6]
+ cb_0_4/io_i_4_in1[7] cb_0_4/io_i_5_ci cb_0_4/io_i_5_in1[0] cb_0_4/io_i_5_in1[1]
+ cb_0_4/io_i_5_in1[2] cb_0_4/io_i_5_in1[3] cb_0_4/io_i_5_in1[4] cb_0_4/io_i_5_in1[5]
+ cb_0_4/io_i_5_in1[6] cb_0_4/io_i_5_in1[7] cb_0_4/io_i_6_ci cb_0_4/io_i_6_in1[0]
+ cb_0_4/io_i_6_in1[1] cb_0_4/io_i_6_in1[2] cb_0_4/io_i_6_in1[3] cb_0_4/io_i_6_in1[4]
+ cb_0_4/io_i_6_in1[5] cb_0_4/io_i_6_in1[6] cb_0_4/io_i_6_in1[7] cb_0_4/io_i_7_ci
+ cb_0_4/io_i_7_in1[0] cb_0_4/io_i_7_in1[1] cb_0_4/io_i_7_in1[2] cb_0_4/io_i_7_in1[3]
+ cb_0_4/io_i_7_in1[4] cb_0_4/io_i_7_in1[5] cb_0_4/io_i_7_in1[6] cb_0_4/io_i_7_in1[7]
+ cb_0_3/io_vci cb_0_4/io_vci cb_0_3/io_vi cb_0_9/io_we_i cb_0_3/io_wo[0] cb_0_3/io_wo[10]
+ cb_0_3/io_wo[11] cb_0_3/io_wo[12] cb_0_3/io_wo[13] cb_0_3/io_wo[14] cb_0_3/io_wo[15]
+ cb_0_3/io_wo[16] cb_0_3/io_wo[17] cb_0_3/io_wo[18] cb_0_3/io_wo[19] cb_0_3/io_wo[1]
+ cb_0_3/io_wo[20] cb_0_3/io_wo[21] cb_0_3/io_wo[22] cb_0_3/io_wo[23] cb_0_3/io_wo[24]
+ cb_0_3/io_wo[25] cb_0_3/io_wo[26] cb_0_3/io_wo[27] cb_0_3/io_wo[28] cb_0_3/io_wo[29]
+ cb_0_3/io_wo[2] cb_0_3/io_wo[30] cb_0_3/io_wo[31] cb_0_3/io_wo[32] cb_0_3/io_wo[33]
+ cb_0_3/io_wo[34] cb_0_3/io_wo[35] cb_0_3/io_wo[36] cb_0_3/io_wo[37] cb_0_3/io_wo[38]
+ cb_0_3/io_wo[39] cb_0_3/io_wo[3] cb_0_3/io_wo[40] cb_0_3/io_wo[41] cb_0_3/io_wo[42]
+ cb_0_3/io_wo[43] cb_0_3/io_wo[44] cb_0_3/io_wo[45] cb_0_3/io_wo[46] cb_0_3/io_wo[47]
+ cb_0_3/io_wo[48] cb_0_3/io_wo[49] cb_0_3/io_wo[4] cb_0_3/io_wo[50] cb_0_3/io_wo[51]
+ cb_0_3/io_wo[52] cb_0_3/io_wo[53] cb_0_3/io_wo[54] cb_0_3/io_wo[55] cb_0_3/io_wo[56]
+ cb_0_3/io_wo[57] cb_0_3/io_wo[58] cb_0_3/io_wo[59] cb_0_3/io_wo[5] cb_0_3/io_wo[60]
+ cb_0_3/io_wo[61] cb_0_3/io_wo[62] cb_0_3/io_wo[63] cb_0_3/io_wo[6] cb_0_3/io_wo[7]
+ cb_0_3/io_wo[8] cb_0_3/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_2_7 cb_2_9/io_adr_i[0] cb_2_9/io_adr_i[1] cb_2_7/io_cs_i cb_2_9/io_dat_i[0] cb_2_9/io_dat_i[10]
+ cb_2_9/io_dat_i[11] cb_2_9/io_dat_i[12] cb_2_9/io_dat_i[13] cb_2_9/io_dat_i[14]
+ cb_2_9/io_dat_i[15] cb_2_9/io_dat_i[1] cb_2_9/io_dat_i[2] cb_2_9/io_dat_i[3] cb_2_9/io_dat_i[4]
+ cb_2_9/io_dat_i[5] cb_2_9/io_dat_i[6] cb_2_9/io_dat_i[7] cb_2_9/io_dat_i[8] cb_2_9/io_dat_i[9]
+ cb_2_7/io_dat_o[0] cb_2_7/io_dat_o[10] cb_2_7/io_dat_o[11] cb_2_7/io_dat_o[12] cb_2_7/io_dat_o[13]
+ cb_2_7/io_dat_o[14] cb_2_7/io_dat_o[15] cb_2_7/io_dat_o[1] cb_2_7/io_dat_o[2] cb_2_7/io_dat_o[3]
+ cb_2_7/io_dat_o[4] cb_2_7/io_dat_o[5] cb_2_7/io_dat_o[6] cb_2_7/io_dat_o[7] cb_2_7/io_dat_o[8]
+ cb_2_7/io_dat_o[9] cb_2_8/io_wo[0] cb_2_8/io_wo[10] cb_2_8/io_wo[11] cb_2_8/io_wo[12]
+ cb_2_8/io_wo[13] cb_2_8/io_wo[14] cb_2_8/io_wo[15] cb_2_8/io_wo[16] cb_2_8/io_wo[17]
+ cb_2_8/io_wo[18] cb_2_8/io_wo[19] cb_2_8/io_wo[1] cb_2_8/io_wo[20] cb_2_8/io_wo[21]
+ cb_2_8/io_wo[22] cb_2_8/io_wo[23] cb_2_8/io_wo[24] cb_2_8/io_wo[25] cb_2_8/io_wo[26]
+ cb_2_8/io_wo[27] cb_2_8/io_wo[28] cb_2_8/io_wo[29] cb_2_8/io_wo[2] cb_2_8/io_wo[30]
+ cb_2_8/io_wo[31] cb_2_8/io_wo[32] cb_2_8/io_wo[33] cb_2_8/io_wo[34] cb_2_8/io_wo[35]
+ cb_2_8/io_wo[36] cb_2_8/io_wo[37] cb_2_8/io_wo[38] cb_2_8/io_wo[39] cb_2_8/io_wo[3]
+ cb_2_8/io_wo[40] cb_2_8/io_wo[41] cb_2_8/io_wo[42] cb_2_8/io_wo[43] cb_2_8/io_wo[44]
+ cb_2_8/io_wo[45] cb_2_8/io_wo[46] cb_2_8/io_wo[47] cb_2_8/io_wo[48] cb_2_8/io_wo[49]
+ cb_2_8/io_wo[4] cb_2_8/io_wo[50] cb_2_8/io_wo[51] cb_2_8/io_wo[52] cb_2_8/io_wo[53]
+ cb_2_8/io_wo[54] cb_2_8/io_wo[55] cb_2_8/io_wo[56] cb_2_8/io_wo[57] cb_2_8/io_wo[58]
+ cb_2_8/io_wo[59] cb_2_8/io_wo[5] cb_2_8/io_wo[60] cb_2_8/io_wo[61] cb_2_8/io_wo[62]
+ cb_2_8/io_wo[63] cb_2_8/io_wo[6] cb_2_8/io_wo[7] cb_2_8/io_wo[8] cb_2_8/io_wo[9]
+ cb_2_7/io_i_0_ci cb_2_7/io_i_0_in1[0] cb_2_7/io_i_0_in1[1] cb_2_7/io_i_0_in1[2]
+ cb_2_7/io_i_0_in1[3] cb_2_7/io_i_0_in1[4] cb_2_7/io_i_0_in1[5] cb_2_7/io_i_0_in1[6]
+ cb_2_7/io_i_0_in1[7] cb_2_7/io_i_1_ci cb_2_7/io_i_1_in1[0] cb_2_7/io_i_1_in1[1]
+ cb_2_7/io_i_1_in1[2] cb_2_7/io_i_1_in1[3] cb_2_7/io_i_1_in1[4] cb_2_7/io_i_1_in1[5]
+ cb_2_7/io_i_1_in1[6] cb_2_7/io_i_1_in1[7] cb_2_7/io_i_2_ci cb_2_7/io_i_2_in1[0]
+ cb_2_7/io_i_2_in1[1] cb_2_7/io_i_2_in1[2] cb_2_7/io_i_2_in1[3] cb_2_7/io_i_2_in1[4]
+ cb_2_7/io_i_2_in1[5] cb_2_7/io_i_2_in1[6] cb_2_7/io_i_2_in1[7] cb_2_7/io_i_3_ci
+ cb_2_7/io_i_3_in1[0] cb_2_7/io_i_3_in1[1] cb_2_7/io_i_3_in1[2] cb_2_7/io_i_3_in1[3]
+ cb_2_7/io_i_3_in1[4] cb_2_7/io_i_3_in1[5] cb_2_7/io_i_3_in1[6] cb_2_7/io_i_3_in1[7]
+ cb_2_7/io_i_4_ci cb_2_7/io_i_4_in1[0] cb_2_7/io_i_4_in1[1] cb_2_7/io_i_4_in1[2]
+ cb_2_7/io_i_4_in1[3] cb_2_7/io_i_4_in1[4] cb_2_7/io_i_4_in1[5] cb_2_7/io_i_4_in1[6]
+ cb_2_7/io_i_4_in1[7] cb_2_7/io_i_5_ci cb_2_7/io_i_5_in1[0] cb_2_7/io_i_5_in1[1]
+ cb_2_7/io_i_5_in1[2] cb_2_7/io_i_5_in1[3] cb_2_7/io_i_5_in1[4] cb_2_7/io_i_5_in1[5]
+ cb_2_7/io_i_5_in1[6] cb_2_7/io_i_5_in1[7] cb_2_7/io_i_6_ci cb_2_7/io_i_6_in1[0]
+ cb_2_7/io_i_6_in1[1] cb_2_7/io_i_6_in1[2] cb_2_7/io_i_6_in1[3] cb_2_7/io_i_6_in1[4]
+ cb_2_7/io_i_6_in1[5] cb_2_7/io_i_6_in1[6] cb_2_7/io_i_6_in1[7] cb_2_7/io_i_7_ci
+ cb_2_7/io_i_7_in1[0] cb_2_7/io_i_7_in1[1] cb_2_7/io_i_7_in1[2] cb_2_7/io_i_7_in1[3]
+ cb_2_7/io_i_7_in1[4] cb_2_7/io_i_7_in1[5] cb_2_7/io_i_7_in1[6] cb_2_7/io_i_7_in1[7]
+ cb_2_8/io_i_0_ci cb_2_8/io_i_0_in1[0] cb_2_8/io_i_0_in1[1] cb_2_8/io_i_0_in1[2]
+ cb_2_8/io_i_0_in1[3] cb_2_8/io_i_0_in1[4] cb_2_8/io_i_0_in1[5] cb_2_8/io_i_0_in1[6]
+ cb_2_8/io_i_0_in1[7] cb_2_8/io_i_1_ci cb_2_8/io_i_1_in1[0] cb_2_8/io_i_1_in1[1]
+ cb_2_8/io_i_1_in1[2] cb_2_8/io_i_1_in1[3] cb_2_8/io_i_1_in1[4] cb_2_8/io_i_1_in1[5]
+ cb_2_8/io_i_1_in1[6] cb_2_8/io_i_1_in1[7] cb_2_8/io_i_2_ci cb_2_8/io_i_2_in1[0]
+ cb_2_8/io_i_2_in1[1] cb_2_8/io_i_2_in1[2] cb_2_8/io_i_2_in1[3] cb_2_8/io_i_2_in1[4]
+ cb_2_8/io_i_2_in1[5] cb_2_8/io_i_2_in1[6] cb_2_8/io_i_2_in1[7] cb_2_8/io_i_3_ci
+ cb_2_8/io_i_3_in1[0] cb_2_8/io_i_3_in1[1] cb_2_8/io_i_3_in1[2] cb_2_8/io_i_3_in1[3]
+ cb_2_8/io_i_3_in1[4] cb_2_8/io_i_3_in1[5] cb_2_8/io_i_3_in1[6] cb_2_8/io_i_3_in1[7]
+ cb_2_8/io_i_4_ci cb_2_8/io_i_4_in1[0] cb_2_8/io_i_4_in1[1] cb_2_8/io_i_4_in1[2]
+ cb_2_8/io_i_4_in1[3] cb_2_8/io_i_4_in1[4] cb_2_8/io_i_4_in1[5] cb_2_8/io_i_4_in1[6]
+ cb_2_8/io_i_4_in1[7] cb_2_8/io_i_5_ci cb_2_8/io_i_5_in1[0] cb_2_8/io_i_5_in1[1]
+ cb_2_8/io_i_5_in1[2] cb_2_8/io_i_5_in1[3] cb_2_8/io_i_5_in1[4] cb_2_8/io_i_5_in1[5]
+ cb_2_8/io_i_5_in1[6] cb_2_8/io_i_5_in1[7] cb_2_8/io_i_6_ci cb_2_8/io_i_6_in1[0]
+ cb_2_8/io_i_6_in1[1] cb_2_8/io_i_6_in1[2] cb_2_8/io_i_6_in1[3] cb_2_8/io_i_6_in1[4]
+ cb_2_8/io_i_6_in1[5] cb_2_8/io_i_6_in1[6] cb_2_8/io_i_6_in1[7] cb_2_8/io_i_7_ci
+ cb_2_8/io_i_7_in1[0] cb_2_8/io_i_7_in1[1] cb_2_8/io_i_7_in1[2] cb_2_8/io_i_7_in1[3]
+ cb_2_8/io_i_7_in1[4] cb_2_8/io_i_7_in1[5] cb_2_8/io_i_7_in1[6] cb_2_8/io_i_7_in1[7]
+ cb_2_7/io_vci cb_2_8/io_vci cb_2_7/io_vi cb_2_9/io_we_i cb_2_7/io_wo[0] cb_2_7/io_wo[10]
+ cb_2_7/io_wo[11] cb_2_7/io_wo[12] cb_2_7/io_wo[13] cb_2_7/io_wo[14] cb_2_7/io_wo[15]
+ cb_2_7/io_wo[16] cb_2_7/io_wo[17] cb_2_7/io_wo[18] cb_2_7/io_wo[19] cb_2_7/io_wo[1]
+ cb_2_7/io_wo[20] cb_2_7/io_wo[21] cb_2_7/io_wo[22] cb_2_7/io_wo[23] cb_2_7/io_wo[24]
+ cb_2_7/io_wo[25] cb_2_7/io_wo[26] cb_2_7/io_wo[27] cb_2_7/io_wo[28] cb_2_7/io_wo[29]
+ cb_2_7/io_wo[2] cb_2_7/io_wo[30] cb_2_7/io_wo[31] cb_2_7/io_wo[32] cb_2_7/io_wo[33]
+ cb_2_7/io_wo[34] cb_2_7/io_wo[35] cb_2_7/io_wo[36] cb_2_7/io_wo[37] cb_2_7/io_wo[38]
+ cb_2_7/io_wo[39] cb_2_7/io_wo[3] cb_2_7/io_wo[40] cb_2_7/io_wo[41] cb_2_7/io_wo[42]
+ cb_2_7/io_wo[43] cb_2_7/io_wo[44] cb_2_7/io_wo[45] cb_2_7/io_wo[46] cb_2_7/io_wo[47]
+ cb_2_7/io_wo[48] cb_2_7/io_wo[49] cb_2_7/io_wo[4] cb_2_7/io_wo[50] cb_2_7/io_wo[51]
+ cb_2_7/io_wo[52] cb_2_7/io_wo[53] cb_2_7/io_wo[54] cb_2_7/io_wo[55] cb_2_7/io_wo[56]
+ cb_2_7/io_wo[57] cb_2_7/io_wo[58] cb_2_7/io_wo[59] cb_2_7/io_wo[5] cb_2_7/io_wo[60]
+ cb_2_7/io_wo[61] cb_2_7/io_wo[62] cb_2_7/io_wo[63] cb_2_7/io_wo[6] cb_2_7/io_wo[7]
+ cb_2_7/io_wo[8] cb_2_7/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_0_4 cb_0_9/io_adr_i[0] cb_0_9/io_adr_i[1] cb_0_4/io_cs_i cb_0_9/io_dat_i[0] cb_0_9/io_dat_i[10]
+ cb_0_9/io_dat_i[11] cb_0_9/io_dat_i[12] cb_0_9/io_dat_i[13] cb_0_9/io_dat_i[14]
+ cb_0_9/io_dat_i[15] cb_0_9/io_dat_i[1] cb_0_9/io_dat_i[2] cb_0_9/io_dat_i[3] cb_0_9/io_dat_i[4]
+ cb_0_9/io_dat_i[5] cb_0_9/io_dat_i[6] cb_0_9/io_dat_i[7] cb_0_9/io_dat_i[8] cb_0_9/io_dat_i[9]
+ cb_0_4/io_dat_o[0] cb_0_4/io_dat_o[10] cb_0_4/io_dat_o[11] cb_0_4/io_dat_o[12] cb_0_4/io_dat_o[13]
+ cb_0_4/io_dat_o[14] cb_0_4/io_dat_o[15] cb_0_4/io_dat_o[1] cb_0_4/io_dat_o[2] cb_0_4/io_dat_o[3]
+ cb_0_4/io_dat_o[4] cb_0_4/io_dat_o[5] cb_0_4/io_dat_o[6] cb_0_4/io_dat_o[7] cb_0_4/io_dat_o[8]
+ cb_0_4/io_dat_o[9] cb_0_5/io_wo[0] cb_0_5/io_wo[10] cb_0_5/io_wo[11] cb_0_5/io_wo[12]
+ cb_0_5/io_wo[13] cb_0_5/io_wo[14] cb_0_5/io_wo[15] cb_0_5/io_wo[16] cb_0_5/io_wo[17]
+ cb_0_5/io_wo[18] cb_0_5/io_wo[19] cb_0_5/io_wo[1] cb_0_5/io_wo[20] cb_0_5/io_wo[21]
+ cb_0_5/io_wo[22] cb_0_5/io_wo[23] cb_0_5/io_wo[24] cb_0_5/io_wo[25] cb_0_5/io_wo[26]
+ cb_0_5/io_wo[27] cb_0_5/io_wo[28] cb_0_5/io_wo[29] cb_0_5/io_wo[2] cb_0_5/io_wo[30]
+ cb_0_5/io_wo[31] cb_0_5/io_wo[32] cb_0_5/io_wo[33] cb_0_5/io_wo[34] cb_0_5/io_wo[35]
+ cb_0_5/io_wo[36] cb_0_5/io_wo[37] cb_0_5/io_wo[38] cb_0_5/io_wo[39] cb_0_5/io_wo[3]
+ cb_0_5/io_wo[40] cb_0_5/io_wo[41] cb_0_5/io_wo[42] cb_0_5/io_wo[43] cb_0_5/io_wo[44]
+ cb_0_5/io_wo[45] cb_0_5/io_wo[46] cb_0_5/io_wo[47] cb_0_5/io_wo[48] cb_0_5/io_wo[49]
+ cb_0_5/io_wo[4] cb_0_5/io_wo[50] cb_0_5/io_wo[51] cb_0_5/io_wo[52] cb_0_5/io_wo[53]
+ cb_0_5/io_wo[54] cb_0_5/io_wo[55] cb_0_5/io_wo[56] cb_0_5/io_wo[57] cb_0_5/io_wo[58]
+ cb_0_5/io_wo[59] cb_0_5/io_wo[5] cb_0_5/io_wo[60] cb_0_5/io_wo[61] cb_0_5/io_wo[62]
+ cb_0_5/io_wo[63] cb_0_5/io_wo[6] cb_0_5/io_wo[7] cb_0_5/io_wo[8] cb_0_5/io_wo[9]
+ cb_0_4/io_i_0_ci cb_0_4/io_i_0_in1[0] cb_0_4/io_i_0_in1[1] cb_0_4/io_i_0_in1[2]
+ cb_0_4/io_i_0_in1[3] cb_0_4/io_i_0_in1[4] cb_0_4/io_i_0_in1[5] cb_0_4/io_i_0_in1[6]
+ cb_0_4/io_i_0_in1[7] cb_0_4/io_i_1_ci cb_0_4/io_i_1_in1[0] cb_0_4/io_i_1_in1[1]
+ cb_0_4/io_i_1_in1[2] cb_0_4/io_i_1_in1[3] cb_0_4/io_i_1_in1[4] cb_0_4/io_i_1_in1[5]
+ cb_0_4/io_i_1_in1[6] cb_0_4/io_i_1_in1[7] cb_0_4/io_i_2_ci cb_0_4/io_i_2_in1[0]
+ cb_0_4/io_i_2_in1[1] cb_0_4/io_i_2_in1[2] cb_0_4/io_i_2_in1[3] cb_0_4/io_i_2_in1[4]
+ cb_0_4/io_i_2_in1[5] cb_0_4/io_i_2_in1[6] cb_0_4/io_i_2_in1[7] cb_0_4/io_i_3_ci
+ cb_0_4/io_i_3_in1[0] cb_0_4/io_i_3_in1[1] cb_0_4/io_i_3_in1[2] cb_0_4/io_i_3_in1[3]
+ cb_0_4/io_i_3_in1[4] cb_0_4/io_i_3_in1[5] cb_0_4/io_i_3_in1[6] cb_0_4/io_i_3_in1[7]
+ cb_0_4/io_i_4_ci cb_0_4/io_i_4_in1[0] cb_0_4/io_i_4_in1[1] cb_0_4/io_i_4_in1[2]
+ cb_0_4/io_i_4_in1[3] cb_0_4/io_i_4_in1[4] cb_0_4/io_i_4_in1[5] cb_0_4/io_i_4_in1[6]
+ cb_0_4/io_i_4_in1[7] cb_0_4/io_i_5_ci cb_0_4/io_i_5_in1[0] cb_0_4/io_i_5_in1[1]
+ cb_0_4/io_i_5_in1[2] cb_0_4/io_i_5_in1[3] cb_0_4/io_i_5_in1[4] cb_0_4/io_i_5_in1[5]
+ cb_0_4/io_i_5_in1[6] cb_0_4/io_i_5_in1[7] cb_0_4/io_i_6_ci cb_0_4/io_i_6_in1[0]
+ cb_0_4/io_i_6_in1[1] cb_0_4/io_i_6_in1[2] cb_0_4/io_i_6_in1[3] cb_0_4/io_i_6_in1[4]
+ cb_0_4/io_i_6_in1[5] cb_0_4/io_i_6_in1[6] cb_0_4/io_i_6_in1[7] cb_0_4/io_i_7_ci
+ cb_0_4/io_i_7_in1[0] cb_0_4/io_i_7_in1[1] cb_0_4/io_i_7_in1[2] cb_0_4/io_i_7_in1[3]
+ cb_0_4/io_i_7_in1[4] cb_0_4/io_i_7_in1[5] cb_0_4/io_i_7_in1[6] cb_0_4/io_i_7_in1[7]
+ cb_0_5/io_i_0_ci cb_0_5/io_i_0_in1[0] cb_0_5/io_i_0_in1[1] cb_0_5/io_i_0_in1[2]
+ cb_0_5/io_i_0_in1[3] cb_0_5/io_i_0_in1[4] cb_0_5/io_i_0_in1[5] cb_0_5/io_i_0_in1[6]
+ cb_0_5/io_i_0_in1[7] cb_0_5/io_i_1_ci cb_0_5/io_i_1_in1[0] cb_0_5/io_i_1_in1[1]
+ cb_0_5/io_i_1_in1[2] cb_0_5/io_i_1_in1[3] cb_0_5/io_i_1_in1[4] cb_0_5/io_i_1_in1[5]
+ cb_0_5/io_i_1_in1[6] cb_0_5/io_i_1_in1[7] cb_0_5/io_i_2_ci cb_0_5/io_i_2_in1[0]
+ cb_0_5/io_i_2_in1[1] cb_0_5/io_i_2_in1[2] cb_0_5/io_i_2_in1[3] cb_0_5/io_i_2_in1[4]
+ cb_0_5/io_i_2_in1[5] cb_0_5/io_i_2_in1[6] cb_0_5/io_i_2_in1[7] cb_0_5/io_i_3_ci
+ cb_0_5/io_i_3_in1[0] cb_0_5/io_i_3_in1[1] cb_0_5/io_i_3_in1[2] cb_0_5/io_i_3_in1[3]
+ cb_0_5/io_i_3_in1[4] cb_0_5/io_i_3_in1[5] cb_0_5/io_i_3_in1[6] cb_0_5/io_i_3_in1[7]
+ cb_0_5/io_i_4_ci cb_0_5/io_i_4_in1[0] cb_0_5/io_i_4_in1[1] cb_0_5/io_i_4_in1[2]
+ cb_0_5/io_i_4_in1[3] cb_0_5/io_i_4_in1[4] cb_0_5/io_i_4_in1[5] cb_0_5/io_i_4_in1[6]
+ cb_0_5/io_i_4_in1[7] cb_0_5/io_i_5_ci cb_0_5/io_i_5_in1[0] cb_0_5/io_i_5_in1[1]
+ cb_0_5/io_i_5_in1[2] cb_0_5/io_i_5_in1[3] cb_0_5/io_i_5_in1[4] cb_0_5/io_i_5_in1[5]
+ cb_0_5/io_i_5_in1[6] cb_0_5/io_i_5_in1[7] cb_0_5/io_i_6_ci cb_0_5/io_i_6_in1[0]
+ cb_0_5/io_i_6_in1[1] cb_0_5/io_i_6_in1[2] cb_0_5/io_i_6_in1[3] cb_0_5/io_i_6_in1[4]
+ cb_0_5/io_i_6_in1[5] cb_0_5/io_i_6_in1[6] cb_0_5/io_i_6_in1[7] cb_0_5/io_i_7_ci
+ cb_0_5/io_i_7_in1[0] cb_0_5/io_i_7_in1[1] cb_0_5/io_i_7_in1[2] cb_0_5/io_i_7_in1[3]
+ cb_0_5/io_i_7_in1[4] cb_0_5/io_i_7_in1[5] cb_0_5/io_i_7_in1[6] cb_0_5/io_i_7_in1[7]
+ cb_0_4/io_vci cb_0_5/io_vci cb_0_4/io_vi cb_0_9/io_we_i cb_0_4/io_wo[0] cb_0_4/io_wo[10]
+ cb_0_4/io_wo[11] cb_0_4/io_wo[12] cb_0_4/io_wo[13] cb_0_4/io_wo[14] cb_0_4/io_wo[15]
+ cb_0_4/io_wo[16] cb_0_4/io_wo[17] cb_0_4/io_wo[18] cb_0_4/io_wo[19] cb_0_4/io_wo[1]
+ cb_0_4/io_wo[20] cb_0_4/io_wo[21] cb_0_4/io_wo[22] cb_0_4/io_wo[23] cb_0_4/io_wo[24]
+ cb_0_4/io_wo[25] cb_0_4/io_wo[26] cb_0_4/io_wo[27] cb_0_4/io_wo[28] cb_0_4/io_wo[29]
+ cb_0_4/io_wo[2] cb_0_4/io_wo[30] cb_0_4/io_wo[31] cb_0_4/io_wo[32] cb_0_4/io_wo[33]
+ cb_0_4/io_wo[34] cb_0_4/io_wo[35] cb_0_4/io_wo[36] cb_0_4/io_wo[37] cb_0_4/io_wo[38]
+ cb_0_4/io_wo[39] cb_0_4/io_wo[3] cb_0_4/io_wo[40] cb_0_4/io_wo[41] cb_0_4/io_wo[42]
+ cb_0_4/io_wo[43] cb_0_4/io_wo[44] cb_0_4/io_wo[45] cb_0_4/io_wo[46] cb_0_4/io_wo[47]
+ cb_0_4/io_wo[48] cb_0_4/io_wo[49] cb_0_4/io_wo[4] cb_0_4/io_wo[50] cb_0_4/io_wo[51]
+ cb_0_4/io_wo[52] cb_0_4/io_wo[53] cb_0_4/io_wo[54] cb_0_4/io_wo[55] cb_0_4/io_wo[56]
+ cb_0_4/io_wo[57] cb_0_4/io_wo[58] cb_0_4/io_wo[59] cb_0_4/io_wo[5] cb_0_4/io_wo[60]
+ cb_0_4/io_wo[61] cb_0_4/io_wo[62] cb_0_4/io_wo[63] cb_0_4/io_wo[6] cb_0_4/io_wo[7]
+ cb_0_4/io_wo[8] cb_0_4/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_2_10 cb_2_9/io_adr_i[0] cb_2_9/io_adr_i[1] cb_2_10/io_cs_i cb_2_9/io_dat_i[0]
+ cb_2_9/io_dat_i[10] cb_2_9/io_dat_i[11] cb_2_9/io_dat_i[12] cb_2_9/io_dat_i[13]
+ cb_2_9/io_dat_i[14] cb_2_9/io_dat_i[15] cb_2_9/io_dat_i[1] cb_2_9/io_dat_i[2] cb_2_9/io_dat_i[3]
+ cb_2_9/io_dat_i[4] cb_2_9/io_dat_i[5] cb_2_9/io_dat_i[6] cb_2_9/io_dat_i[7] cb_2_9/io_dat_i[8]
+ cb_2_9/io_dat_i[9] cb_2_10/io_dat_o[0] cb_2_10/io_dat_o[10] cb_2_10/io_dat_o[11]
+ cb_2_10/io_dat_o[12] cb_2_10/io_dat_o[13] cb_2_10/io_dat_o[14] cb_2_10/io_dat_o[15]
+ cb_2_10/io_dat_o[1] cb_2_10/io_dat_o[2] cb_2_10/io_dat_o[3] cb_2_10/io_dat_o[4]
+ cb_2_10/io_dat_o[5] cb_2_10/io_dat_o[6] cb_2_10/io_dat_o[7] cb_2_10/io_dat_o[8]
+ cb_2_10/io_dat_o[9] cb_2_10/io_eo[0] cb_2_10/io_eo[10] cb_2_10/io_eo[11] cb_2_10/io_eo[12]
+ cb_2_10/io_eo[13] cb_2_10/io_eo[14] cb_2_10/io_eo[15] cb_2_10/io_eo[16] cb_2_10/io_eo[17]
+ cb_2_10/io_eo[18] cb_2_10/io_eo[19] cb_2_10/io_eo[1] cb_2_10/io_eo[20] cb_2_10/io_eo[21]
+ cb_2_10/io_eo[22] cb_2_10/io_eo[23] cb_2_10/io_eo[24] cb_2_10/io_eo[25] cb_2_10/io_eo[26]
+ cb_2_10/io_eo[27] cb_2_10/io_eo[28] cb_2_10/io_eo[29] cb_2_10/io_eo[2] cb_2_10/io_eo[30]
+ cb_2_10/io_eo[31] cb_2_10/io_eo[32] cb_2_10/io_eo[33] cb_2_10/io_eo[34] cb_2_10/io_eo[35]
+ cb_2_10/io_eo[36] cb_2_10/io_eo[37] cb_2_10/io_eo[38] cb_2_10/io_eo[39] cb_2_10/io_eo[3]
+ cb_2_10/io_eo[40] cb_2_10/io_eo[41] cb_2_10/io_eo[42] cb_2_10/io_eo[43] cb_2_10/io_eo[44]
+ cb_2_10/io_eo[45] cb_2_10/io_eo[46] cb_2_10/io_eo[47] cb_2_10/io_eo[48] cb_2_10/io_eo[49]
+ cb_2_10/io_eo[4] cb_2_10/io_eo[50] cb_2_10/io_eo[51] cb_2_10/io_eo[52] cb_2_10/io_eo[53]
+ cb_2_10/io_eo[54] cb_2_10/io_eo[55] cb_2_10/io_eo[56] cb_2_10/io_eo[57] cb_2_10/io_eo[58]
+ cb_2_10/io_eo[59] cb_2_10/io_eo[5] cb_2_10/io_eo[60] cb_2_10/io_eo[61] cb_2_10/io_eo[62]
+ cb_2_10/io_eo[63] cb_2_10/io_eo[6] cb_2_10/io_eo[7] cb_2_10/io_eo[8] cb_2_10/io_eo[9]
+ cb_2_9/io_o_0_co cb_2_9/io_o_0_out[0] cb_2_9/io_o_0_out[1] cb_2_9/io_o_0_out[2]
+ cb_2_9/io_o_0_out[3] cb_2_9/io_o_0_out[4] cb_2_9/io_o_0_out[5] cb_2_9/io_o_0_out[6]
+ cb_2_9/io_o_0_out[7] cb_2_9/io_o_1_co cb_2_9/io_o_1_out[0] cb_2_9/io_o_1_out[1]
+ cb_2_9/io_o_1_out[2] cb_2_9/io_o_1_out[3] cb_2_9/io_o_1_out[4] cb_2_9/io_o_1_out[5]
+ cb_2_9/io_o_1_out[6] cb_2_9/io_o_1_out[7] cb_2_9/io_o_2_co cb_2_9/io_o_2_out[0]
+ cb_2_9/io_o_2_out[1] cb_2_9/io_o_2_out[2] cb_2_9/io_o_2_out[3] cb_2_9/io_o_2_out[4]
+ cb_2_9/io_o_2_out[5] cb_2_9/io_o_2_out[6] cb_2_9/io_o_2_out[7] cb_2_9/io_o_3_co
+ cb_2_9/io_o_3_out[0] cb_2_9/io_o_3_out[1] cb_2_9/io_o_3_out[2] cb_2_9/io_o_3_out[3]
+ cb_2_9/io_o_3_out[4] cb_2_9/io_o_3_out[5] cb_2_9/io_o_3_out[6] cb_2_9/io_o_3_out[7]
+ cb_2_9/io_o_4_co cb_2_9/io_o_4_out[0] cb_2_9/io_o_4_out[1] cb_2_9/io_o_4_out[2]
+ cb_2_9/io_o_4_out[3] cb_2_9/io_o_4_out[4] cb_2_9/io_o_4_out[5] cb_2_9/io_o_4_out[6]
+ cb_2_9/io_o_4_out[7] cb_2_9/io_o_5_co cb_2_9/io_o_5_out[0] cb_2_9/io_o_5_out[1]
+ cb_2_9/io_o_5_out[2] cb_2_9/io_o_5_out[3] cb_2_9/io_o_5_out[4] cb_2_9/io_o_5_out[5]
+ cb_2_9/io_o_5_out[6] cb_2_9/io_o_5_out[7] cb_2_9/io_o_6_co cb_2_9/io_o_6_out[0]
+ cb_2_9/io_o_6_out[1] cb_2_9/io_o_6_out[2] cb_2_9/io_o_6_out[3] cb_2_9/io_o_6_out[4]
+ cb_2_9/io_o_6_out[5] cb_2_9/io_o_6_out[6] cb_2_9/io_o_6_out[7] cb_2_9/io_o_7_co
+ cb_2_9/io_o_7_out[0] cb_2_9/io_o_7_out[1] cb_2_9/io_o_7_out[2] cb_2_9/io_o_7_out[3]
+ cb_2_9/io_o_7_out[4] cb_2_9/io_o_7_out[5] cb_2_9/io_o_7_out[6] cb_2_9/io_o_7_out[7]
+ cb_2_10/io_o_0_co cb_2_10/io_eo[0] cb_2_10/io_eo[1] cb_2_10/io_eo[2] cb_2_10/io_eo[3]
+ cb_2_10/io_eo[4] cb_2_10/io_eo[5] cb_2_10/io_eo[6] cb_2_10/io_eo[7] cb_2_10/io_o_1_co
+ cb_2_10/io_eo[8] cb_2_10/io_eo[9] cb_2_10/io_eo[10] cb_2_10/io_eo[11] cb_2_10/io_eo[12]
+ cb_2_10/io_eo[13] cb_2_10/io_eo[14] cb_2_10/io_eo[15] cb_2_10/io_o_2_co cb_2_10/io_eo[16]
+ cb_2_10/io_eo[17] cb_2_10/io_eo[18] cb_2_10/io_eo[19] cb_2_10/io_eo[20] cb_2_10/io_eo[21]
+ cb_2_10/io_eo[22] cb_2_10/io_eo[23] cb_2_10/io_o_3_co cb_2_10/io_eo[24] cb_2_10/io_eo[25]
+ cb_2_10/io_eo[26] cb_2_10/io_eo[27] cb_2_10/io_eo[28] cb_2_10/io_eo[29] cb_2_10/io_eo[30]
+ cb_2_10/io_eo[31] cb_2_10/io_o_4_co cb_2_10/io_eo[32] cb_2_10/io_eo[33] cb_2_10/io_eo[34]
+ cb_2_10/io_eo[35] cb_2_10/io_eo[36] cb_2_10/io_eo[37] cb_2_10/io_eo[38] cb_2_10/io_eo[39]
+ cb_2_10/io_o_5_co cb_2_10/io_eo[40] cb_2_10/io_eo[41] cb_2_10/io_eo[42] cb_2_10/io_eo[43]
+ cb_2_10/io_eo[44] cb_2_10/io_eo[45] cb_2_10/io_eo[46] cb_2_10/io_eo[47] cb_2_10/io_o_6_co
+ cb_2_10/io_eo[48] cb_2_10/io_eo[49] cb_2_10/io_eo[50] cb_2_10/io_eo[51] cb_2_10/io_eo[52]
+ cb_2_10/io_eo[53] cb_2_10/io_eo[54] cb_2_10/io_eo[55] cb_2_10/io_o_7_co cb_2_10/io_eo[56]
+ cb_2_10/io_eo[57] cb_2_10/io_eo[58] cb_2_10/io_eo[59] cb_2_10/io_eo[60] cb_2_10/io_eo[61]
+ cb_2_10/io_eo[62] cb_2_10/io_eo[63] cb_2_9/io_vco cb_2_10/io_vco cb_2_10/io_vi cb_2_9/io_we_i
+ cb_2_9/io_eo[0] cb_2_9/io_eo[10] cb_2_9/io_eo[11] cb_2_9/io_eo[12] cb_2_9/io_eo[13]
+ cb_2_9/io_eo[14] cb_2_9/io_eo[15] cb_2_9/io_eo[16] cb_2_9/io_eo[17] cb_2_9/io_eo[18]
+ cb_2_9/io_eo[19] cb_2_9/io_eo[1] cb_2_9/io_eo[20] cb_2_9/io_eo[21] cb_2_9/io_eo[22]
+ cb_2_9/io_eo[23] cb_2_9/io_eo[24] cb_2_9/io_eo[25] cb_2_9/io_eo[26] cb_2_9/io_eo[27]
+ cb_2_9/io_eo[28] cb_2_9/io_eo[29] cb_2_9/io_eo[2] cb_2_9/io_eo[30] cb_2_9/io_eo[31]
+ cb_2_9/io_eo[32] cb_2_9/io_eo[33] cb_2_9/io_eo[34] cb_2_9/io_eo[35] cb_2_9/io_eo[36]
+ cb_2_9/io_eo[37] cb_2_9/io_eo[38] cb_2_9/io_eo[39] cb_2_9/io_eo[3] cb_2_9/io_eo[40]
+ cb_2_9/io_eo[41] cb_2_9/io_eo[42] cb_2_9/io_eo[43] cb_2_9/io_eo[44] cb_2_9/io_eo[45]
+ cb_2_9/io_eo[46] cb_2_9/io_eo[47] cb_2_9/io_eo[48] cb_2_9/io_eo[49] cb_2_9/io_eo[4]
+ cb_2_9/io_eo[50] cb_2_9/io_eo[51] cb_2_9/io_eo[52] cb_2_9/io_eo[53] cb_2_9/io_eo[54]
+ cb_2_9/io_eo[55] cb_2_9/io_eo[56] cb_2_9/io_eo[57] cb_2_9/io_eo[58] cb_2_9/io_eo[59]
+ cb_2_9/io_eo[5] cb_2_9/io_eo[60] cb_2_9/io_eo[61] cb_2_9/io_eo[62] cb_2_9/io_eo[63]
+ cb_2_9/io_eo[6] cb_2_9/io_eo[7] cb_2_9/io_eo[8] cb_2_9/io_eo[9] mcons_3/clock mcons_3/reset
+ vccd1 vssd1 cic_block
Xcb_0_5 cb_0_9/io_adr_i[0] cb_0_9/io_adr_i[1] cb_0_5/io_cs_i cb_0_9/io_dat_i[0] cb_0_9/io_dat_i[10]
+ cb_0_9/io_dat_i[11] cb_0_9/io_dat_i[12] cb_0_9/io_dat_i[13] cb_0_9/io_dat_i[14]
+ cb_0_9/io_dat_i[15] cb_0_9/io_dat_i[1] cb_0_9/io_dat_i[2] cb_0_9/io_dat_i[3] cb_0_9/io_dat_i[4]
+ cb_0_9/io_dat_i[5] cb_0_9/io_dat_i[6] cb_0_9/io_dat_i[7] cb_0_9/io_dat_i[8] cb_0_9/io_dat_i[9]
+ cb_0_5/io_dat_o[0] cb_0_5/io_dat_o[10] cb_0_5/io_dat_o[11] cb_0_5/io_dat_o[12] cb_0_5/io_dat_o[13]
+ cb_0_5/io_dat_o[14] cb_0_5/io_dat_o[15] cb_0_5/io_dat_o[1] cb_0_5/io_dat_o[2] cb_0_5/io_dat_o[3]
+ cb_0_5/io_dat_o[4] cb_0_5/io_dat_o[5] cb_0_5/io_dat_o[6] cb_0_5/io_dat_o[7] cb_0_5/io_dat_o[8]
+ cb_0_5/io_dat_o[9] cb_0_6/io_wo[0] cb_0_6/io_wo[10] cb_0_6/io_wo[11] cb_0_6/io_wo[12]
+ cb_0_6/io_wo[13] cb_0_6/io_wo[14] cb_0_6/io_wo[15] cb_0_6/io_wo[16] cb_0_6/io_wo[17]
+ cb_0_6/io_wo[18] cb_0_6/io_wo[19] cb_0_6/io_wo[1] cb_0_6/io_wo[20] cb_0_6/io_wo[21]
+ cb_0_6/io_wo[22] cb_0_6/io_wo[23] cb_0_6/io_wo[24] cb_0_6/io_wo[25] cb_0_6/io_wo[26]
+ cb_0_6/io_wo[27] cb_0_6/io_wo[28] cb_0_6/io_wo[29] cb_0_6/io_wo[2] cb_0_6/io_wo[30]
+ cb_0_6/io_wo[31] cb_0_6/io_wo[32] cb_0_6/io_wo[33] cb_0_6/io_wo[34] cb_0_6/io_wo[35]
+ cb_0_6/io_wo[36] cb_0_6/io_wo[37] cb_0_6/io_wo[38] cb_0_6/io_wo[39] cb_0_6/io_wo[3]
+ cb_0_6/io_wo[40] cb_0_6/io_wo[41] cb_0_6/io_wo[42] cb_0_6/io_wo[43] cb_0_6/io_wo[44]
+ cb_0_6/io_wo[45] cb_0_6/io_wo[46] cb_0_6/io_wo[47] cb_0_6/io_wo[48] cb_0_6/io_wo[49]
+ cb_0_6/io_wo[4] cb_0_6/io_wo[50] cb_0_6/io_wo[51] cb_0_6/io_wo[52] cb_0_6/io_wo[53]
+ cb_0_6/io_wo[54] cb_0_6/io_wo[55] cb_0_6/io_wo[56] cb_0_6/io_wo[57] cb_0_6/io_wo[58]
+ cb_0_6/io_wo[59] cb_0_6/io_wo[5] cb_0_6/io_wo[60] cb_0_6/io_wo[61] cb_0_6/io_wo[62]
+ cb_0_6/io_wo[63] cb_0_6/io_wo[6] cb_0_6/io_wo[7] cb_0_6/io_wo[8] cb_0_6/io_wo[9]
+ cb_0_5/io_i_0_ci cb_0_5/io_i_0_in1[0] cb_0_5/io_i_0_in1[1] cb_0_5/io_i_0_in1[2]
+ cb_0_5/io_i_0_in1[3] cb_0_5/io_i_0_in1[4] cb_0_5/io_i_0_in1[5] cb_0_5/io_i_0_in1[6]
+ cb_0_5/io_i_0_in1[7] cb_0_5/io_i_1_ci cb_0_5/io_i_1_in1[0] cb_0_5/io_i_1_in1[1]
+ cb_0_5/io_i_1_in1[2] cb_0_5/io_i_1_in1[3] cb_0_5/io_i_1_in1[4] cb_0_5/io_i_1_in1[5]
+ cb_0_5/io_i_1_in1[6] cb_0_5/io_i_1_in1[7] cb_0_5/io_i_2_ci cb_0_5/io_i_2_in1[0]
+ cb_0_5/io_i_2_in1[1] cb_0_5/io_i_2_in1[2] cb_0_5/io_i_2_in1[3] cb_0_5/io_i_2_in1[4]
+ cb_0_5/io_i_2_in1[5] cb_0_5/io_i_2_in1[6] cb_0_5/io_i_2_in1[7] cb_0_5/io_i_3_ci
+ cb_0_5/io_i_3_in1[0] cb_0_5/io_i_3_in1[1] cb_0_5/io_i_3_in1[2] cb_0_5/io_i_3_in1[3]
+ cb_0_5/io_i_3_in1[4] cb_0_5/io_i_3_in1[5] cb_0_5/io_i_3_in1[6] cb_0_5/io_i_3_in1[7]
+ cb_0_5/io_i_4_ci cb_0_5/io_i_4_in1[0] cb_0_5/io_i_4_in1[1] cb_0_5/io_i_4_in1[2]
+ cb_0_5/io_i_4_in1[3] cb_0_5/io_i_4_in1[4] cb_0_5/io_i_4_in1[5] cb_0_5/io_i_4_in1[6]
+ cb_0_5/io_i_4_in1[7] cb_0_5/io_i_5_ci cb_0_5/io_i_5_in1[0] cb_0_5/io_i_5_in1[1]
+ cb_0_5/io_i_5_in1[2] cb_0_5/io_i_5_in1[3] cb_0_5/io_i_5_in1[4] cb_0_5/io_i_5_in1[5]
+ cb_0_5/io_i_5_in1[6] cb_0_5/io_i_5_in1[7] cb_0_5/io_i_6_ci cb_0_5/io_i_6_in1[0]
+ cb_0_5/io_i_6_in1[1] cb_0_5/io_i_6_in1[2] cb_0_5/io_i_6_in1[3] cb_0_5/io_i_6_in1[4]
+ cb_0_5/io_i_6_in1[5] cb_0_5/io_i_6_in1[6] cb_0_5/io_i_6_in1[7] cb_0_5/io_i_7_ci
+ cb_0_5/io_i_7_in1[0] cb_0_5/io_i_7_in1[1] cb_0_5/io_i_7_in1[2] cb_0_5/io_i_7_in1[3]
+ cb_0_5/io_i_7_in1[4] cb_0_5/io_i_7_in1[5] cb_0_5/io_i_7_in1[6] cb_0_5/io_i_7_in1[7]
+ cb_0_6/io_i_0_ci cb_0_6/io_i_0_in1[0] cb_0_6/io_i_0_in1[1] cb_0_6/io_i_0_in1[2]
+ cb_0_6/io_i_0_in1[3] cb_0_6/io_i_0_in1[4] cb_0_6/io_i_0_in1[5] cb_0_6/io_i_0_in1[6]
+ cb_0_6/io_i_0_in1[7] cb_0_6/io_i_1_ci cb_0_6/io_i_1_in1[0] cb_0_6/io_i_1_in1[1]
+ cb_0_6/io_i_1_in1[2] cb_0_6/io_i_1_in1[3] cb_0_6/io_i_1_in1[4] cb_0_6/io_i_1_in1[5]
+ cb_0_6/io_i_1_in1[6] cb_0_6/io_i_1_in1[7] cb_0_6/io_i_2_ci cb_0_6/io_i_2_in1[0]
+ cb_0_6/io_i_2_in1[1] cb_0_6/io_i_2_in1[2] cb_0_6/io_i_2_in1[3] cb_0_6/io_i_2_in1[4]
+ cb_0_6/io_i_2_in1[5] cb_0_6/io_i_2_in1[6] cb_0_6/io_i_2_in1[7] cb_0_6/io_i_3_ci
+ cb_0_6/io_i_3_in1[0] cb_0_6/io_i_3_in1[1] cb_0_6/io_i_3_in1[2] cb_0_6/io_i_3_in1[3]
+ cb_0_6/io_i_3_in1[4] cb_0_6/io_i_3_in1[5] cb_0_6/io_i_3_in1[6] cb_0_6/io_i_3_in1[7]
+ cb_0_6/io_i_4_ci cb_0_6/io_i_4_in1[0] cb_0_6/io_i_4_in1[1] cb_0_6/io_i_4_in1[2]
+ cb_0_6/io_i_4_in1[3] cb_0_6/io_i_4_in1[4] cb_0_6/io_i_4_in1[5] cb_0_6/io_i_4_in1[6]
+ cb_0_6/io_i_4_in1[7] cb_0_6/io_i_5_ci cb_0_6/io_i_5_in1[0] cb_0_6/io_i_5_in1[1]
+ cb_0_6/io_i_5_in1[2] cb_0_6/io_i_5_in1[3] cb_0_6/io_i_5_in1[4] cb_0_6/io_i_5_in1[5]
+ cb_0_6/io_i_5_in1[6] cb_0_6/io_i_5_in1[7] cb_0_6/io_i_6_ci cb_0_6/io_i_6_in1[0]
+ cb_0_6/io_i_6_in1[1] cb_0_6/io_i_6_in1[2] cb_0_6/io_i_6_in1[3] cb_0_6/io_i_6_in1[4]
+ cb_0_6/io_i_6_in1[5] cb_0_6/io_i_6_in1[6] cb_0_6/io_i_6_in1[7] cb_0_6/io_i_7_ci
+ cb_0_6/io_i_7_in1[0] cb_0_6/io_i_7_in1[1] cb_0_6/io_i_7_in1[2] cb_0_6/io_i_7_in1[3]
+ cb_0_6/io_i_7_in1[4] cb_0_6/io_i_7_in1[5] cb_0_6/io_i_7_in1[6] cb_0_6/io_i_7_in1[7]
+ cb_0_5/io_vci cb_0_6/io_vci cb_0_5/io_vi cb_0_9/io_we_i cb_0_5/io_wo[0] cb_0_5/io_wo[10]
+ cb_0_5/io_wo[11] cb_0_5/io_wo[12] cb_0_5/io_wo[13] cb_0_5/io_wo[14] cb_0_5/io_wo[15]
+ cb_0_5/io_wo[16] cb_0_5/io_wo[17] cb_0_5/io_wo[18] cb_0_5/io_wo[19] cb_0_5/io_wo[1]
+ cb_0_5/io_wo[20] cb_0_5/io_wo[21] cb_0_5/io_wo[22] cb_0_5/io_wo[23] cb_0_5/io_wo[24]
+ cb_0_5/io_wo[25] cb_0_5/io_wo[26] cb_0_5/io_wo[27] cb_0_5/io_wo[28] cb_0_5/io_wo[29]
+ cb_0_5/io_wo[2] cb_0_5/io_wo[30] cb_0_5/io_wo[31] cb_0_5/io_wo[32] cb_0_5/io_wo[33]
+ cb_0_5/io_wo[34] cb_0_5/io_wo[35] cb_0_5/io_wo[36] cb_0_5/io_wo[37] cb_0_5/io_wo[38]
+ cb_0_5/io_wo[39] cb_0_5/io_wo[3] cb_0_5/io_wo[40] cb_0_5/io_wo[41] cb_0_5/io_wo[42]
+ cb_0_5/io_wo[43] cb_0_5/io_wo[44] cb_0_5/io_wo[45] cb_0_5/io_wo[46] cb_0_5/io_wo[47]
+ cb_0_5/io_wo[48] cb_0_5/io_wo[49] cb_0_5/io_wo[4] cb_0_5/io_wo[50] cb_0_5/io_wo[51]
+ cb_0_5/io_wo[52] cb_0_5/io_wo[53] cb_0_5/io_wo[54] cb_0_5/io_wo[55] cb_0_5/io_wo[56]
+ cb_0_5/io_wo[57] cb_0_5/io_wo[58] cb_0_5/io_wo[59] cb_0_5/io_wo[5] cb_0_5/io_wo[60]
+ cb_0_5/io_wo[61] cb_0_5/io_wo[62] cb_0_5/io_wo[63] cb_0_5/io_wo[6] cb_0_5/io_wo[7]
+ cb_0_5/io_wo[8] cb_0_5/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_2_8 cb_2_9/io_adr_i[0] cb_2_9/io_adr_i[1] cb_2_8/io_cs_i cb_2_9/io_dat_i[0] cb_2_9/io_dat_i[10]
+ cb_2_9/io_dat_i[11] cb_2_9/io_dat_i[12] cb_2_9/io_dat_i[13] cb_2_9/io_dat_i[14]
+ cb_2_9/io_dat_i[15] cb_2_9/io_dat_i[1] cb_2_9/io_dat_i[2] cb_2_9/io_dat_i[3] cb_2_9/io_dat_i[4]
+ cb_2_9/io_dat_i[5] cb_2_9/io_dat_i[6] cb_2_9/io_dat_i[7] cb_2_9/io_dat_i[8] cb_2_9/io_dat_i[9]
+ cb_2_8/io_dat_o[0] cb_2_8/io_dat_o[10] cb_2_8/io_dat_o[11] cb_2_8/io_dat_o[12] cb_2_8/io_dat_o[13]
+ cb_2_8/io_dat_o[14] cb_2_8/io_dat_o[15] cb_2_8/io_dat_o[1] cb_2_8/io_dat_o[2] cb_2_8/io_dat_o[3]
+ cb_2_8/io_dat_o[4] cb_2_8/io_dat_o[5] cb_2_8/io_dat_o[6] cb_2_8/io_dat_o[7] cb_2_8/io_dat_o[8]
+ cb_2_8/io_dat_o[9] cb_2_9/io_wo[0] cb_2_9/io_wo[10] cb_2_9/io_wo[11] cb_2_9/io_wo[12]
+ cb_2_9/io_wo[13] cb_2_9/io_wo[14] cb_2_9/io_wo[15] cb_2_9/io_wo[16] cb_2_9/io_wo[17]
+ cb_2_9/io_wo[18] cb_2_9/io_wo[19] cb_2_9/io_wo[1] cb_2_9/io_wo[20] cb_2_9/io_wo[21]
+ cb_2_9/io_wo[22] cb_2_9/io_wo[23] cb_2_9/io_wo[24] cb_2_9/io_wo[25] cb_2_9/io_wo[26]
+ cb_2_9/io_wo[27] cb_2_9/io_wo[28] cb_2_9/io_wo[29] cb_2_9/io_wo[2] cb_2_9/io_wo[30]
+ cb_2_9/io_wo[31] cb_2_9/io_wo[32] cb_2_9/io_wo[33] cb_2_9/io_wo[34] cb_2_9/io_wo[35]
+ cb_2_9/io_wo[36] cb_2_9/io_wo[37] cb_2_9/io_wo[38] cb_2_9/io_wo[39] cb_2_9/io_wo[3]
+ cb_2_9/io_wo[40] cb_2_9/io_wo[41] cb_2_9/io_wo[42] cb_2_9/io_wo[43] cb_2_9/io_wo[44]
+ cb_2_9/io_wo[45] cb_2_9/io_wo[46] cb_2_9/io_wo[47] cb_2_9/io_wo[48] cb_2_9/io_wo[49]
+ cb_2_9/io_wo[4] cb_2_9/io_wo[50] cb_2_9/io_wo[51] cb_2_9/io_wo[52] cb_2_9/io_wo[53]
+ cb_2_9/io_wo[54] cb_2_9/io_wo[55] cb_2_9/io_wo[56] cb_2_9/io_wo[57] cb_2_9/io_wo[58]
+ cb_2_9/io_wo[59] cb_2_9/io_wo[5] cb_2_9/io_wo[60] cb_2_9/io_wo[61] cb_2_9/io_wo[62]
+ cb_2_9/io_wo[63] cb_2_9/io_wo[6] cb_2_9/io_wo[7] cb_2_9/io_wo[8] cb_2_9/io_wo[9]
+ cb_2_8/io_i_0_ci cb_2_8/io_i_0_in1[0] cb_2_8/io_i_0_in1[1] cb_2_8/io_i_0_in1[2]
+ cb_2_8/io_i_0_in1[3] cb_2_8/io_i_0_in1[4] cb_2_8/io_i_0_in1[5] cb_2_8/io_i_0_in1[6]
+ cb_2_8/io_i_0_in1[7] cb_2_8/io_i_1_ci cb_2_8/io_i_1_in1[0] cb_2_8/io_i_1_in1[1]
+ cb_2_8/io_i_1_in1[2] cb_2_8/io_i_1_in1[3] cb_2_8/io_i_1_in1[4] cb_2_8/io_i_1_in1[5]
+ cb_2_8/io_i_1_in1[6] cb_2_8/io_i_1_in1[7] cb_2_8/io_i_2_ci cb_2_8/io_i_2_in1[0]
+ cb_2_8/io_i_2_in1[1] cb_2_8/io_i_2_in1[2] cb_2_8/io_i_2_in1[3] cb_2_8/io_i_2_in1[4]
+ cb_2_8/io_i_2_in1[5] cb_2_8/io_i_2_in1[6] cb_2_8/io_i_2_in1[7] cb_2_8/io_i_3_ci
+ cb_2_8/io_i_3_in1[0] cb_2_8/io_i_3_in1[1] cb_2_8/io_i_3_in1[2] cb_2_8/io_i_3_in1[3]
+ cb_2_8/io_i_3_in1[4] cb_2_8/io_i_3_in1[5] cb_2_8/io_i_3_in1[6] cb_2_8/io_i_3_in1[7]
+ cb_2_8/io_i_4_ci cb_2_8/io_i_4_in1[0] cb_2_8/io_i_4_in1[1] cb_2_8/io_i_4_in1[2]
+ cb_2_8/io_i_4_in1[3] cb_2_8/io_i_4_in1[4] cb_2_8/io_i_4_in1[5] cb_2_8/io_i_4_in1[6]
+ cb_2_8/io_i_4_in1[7] cb_2_8/io_i_5_ci cb_2_8/io_i_5_in1[0] cb_2_8/io_i_5_in1[1]
+ cb_2_8/io_i_5_in1[2] cb_2_8/io_i_5_in1[3] cb_2_8/io_i_5_in1[4] cb_2_8/io_i_5_in1[5]
+ cb_2_8/io_i_5_in1[6] cb_2_8/io_i_5_in1[7] cb_2_8/io_i_6_ci cb_2_8/io_i_6_in1[0]
+ cb_2_8/io_i_6_in1[1] cb_2_8/io_i_6_in1[2] cb_2_8/io_i_6_in1[3] cb_2_8/io_i_6_in1[4]
+ cb_2_8/io_i_6_in1[5] cb_2_8/io_i_6_in1[6] cb_2_8/io_i_6_in1[7] cb_2_8/io_i_7_ci
+ cb_2_8/io_i_7_in1[0] cb_2_8/io_i_7_in1[1] cb_2_8/io_i_7_in1[2] cb_2_8/io_i_7_in1[3]
+ cb_2_8/io_i_7_in1[4] cb_2_8/io_i_7_in1[5] cb_2_8/io_i_7_in1[6] cb_2_8/io_i_7_in1[7]
+ cb_2_9/io_i_0_ci cb_2_9/io_i_0_in1[0] cb_2_9/io_i_0_in1[1] cb_2_9/io_i_0_in1[2]
+ cb_2_9/io_i_0_in1[3] cb_2_9/io_i_0_in1[4] cb_2_9/io_i_0_in1[5] cb_2_9/io_i_0_in1[6]
+ cb_2_9/io_i_0_in1[7] cb_2_9/io_i_1_ci cb_2_9/io_i_1_in1[0] cb_2_9/io_i_1_in1[1]
+ cb_2_9/io_i_1_in1[2] cb_2_9/io_i_1_in1[3] cb_2_9/io_i_1_in1[4] cb_2_9/io_i_1_in1[5]
+ cb_2_9/io_i_1_in1[6] cb_2_9/io_i_1_in1[7] cb_2_9/io_i_2_ci cb_2_9/io_i_2_in1[0]
+ cb_2_9/io_i_2_in1[1] cb_2_9/io_i_2_in1[2] cb_2_9/io_i_2_in1[3] cb_2_9/io_i_2_in1[4]
+ cb_2_9/io_i_2_in1[5] cb_2_9/io_i_2_in1[6] cb_2_9/io_i_2_in1[7] cb_2_9/io_i_3_ci
+ cb_2_9/io_i_3_in1[0] cb_2_9/io_i_3_in1[1] cb_2_9/io_i_3_in1[2] cb_2_9/io_i_3_in1[3]
+ cb_2_9/io_i_3_in1[4] cb_2_9/io_i_3_in1[5] cb_2_9/io_i_3_in1[6] cb_2_9/io_i_3_in1[7]
+ cb_2_9/io_i_4_ci cb_2_9/io_i_4_in1[0] cb_2_9/io_i_4_in1[1] cb_2_9/io_i_4_in1[2]
+ cb_2_9/io_i_4_in1[3] cb_2_9/io_i_4_in1[4] cb_2_9/io_i_4_in1[5] cb_2_9/io_i_4_in1[6]
+ cb_2_9/io_i_4_in1[7] cb_2_9/io_i_5_ci cb_2_9/io_i_5_in1[0] cb_2_9/io_i_5_in1[1]
+ cb_2_9/io_i_5_in1[2] cb_2_9/io_i_5_in1[3] cb_2_9/io_i_5_in1[4] cb_2_9/io_i_5_in1[5]
+ cb_2_9/io_i_5_in1[6] cb_2_9/io_i_5_in1[7] cb_2_9/io_i_6_ci cb_2_9/io_i_6_in1[0]
+ cb_2_9/io_i_6_in1[1] cb_2_9/io_i_6_in1[2] cb_2_9/io_i_6_in1[3] cb_2_9/io_i_6_in1[4]
+ cb_2_9/io_i_6_in1[5] cb_2_9/io_i_6_in1[6] cb_2_9/io_i_6_in1[7] cb_2_9/io_i_7_ci
+ cb_2_9/io_i_7_in1[0] cb_2_9/io_i_7_in1[1] cb_2_9/io_i_7_in1[2] cb_2_9/io_i_7_in1[3]
+ cb_2_9/io_i_7_in1[4] cb_2_9/io_i_7_in1[5] cb_2_9/io_i_7_in1[6] cb_2_9/io_i_7_in1[7]
+ cb_2_8/io_vci cb_2_9/io_vci cb_2_8/io_vi cb_2_9/io_we_i cb_2_8/io_wo[0] cb_2_8/io_wo[10]
+ cb_2_8/io_wo[11] cb_2_8/io_wo[12] cb_2_8/io_wo[13] cb_2_8/io_wo[14] cb_2_8/io_wo[15]
+ cb_2_8/io_wo[16] cb_2_8/io_wo[17] cb_2_8/io_wo[18] cb_2_8/io_wo[19] cb_2_8/io_wo[1]
+ cb_2_8/io_wo[20] cb_2_8/io_wo[21] cb_2_8/io_wo[22] cb_2_8/io_wo[23] cb_2_8/io_wo[24]
+ cb_2_8/io_wo[25] cb_2_8/io_wo[26] cb_2_8/io_wo[27] cb_2_8/io_wo[28] cb_2_8/io_wo[29]
+ cb_2_8/io_wo[2] cb_2_8/io_wo[30] cb_2_8/io_wo[31] cb_2_8/io_wo[32] cb_2_8/io_wo[33]
+ cb_2_8/io_wo[34] cb_2_8/io_wo[35] cb_2_8/io_wo[36] cb_2_8/io_wo[37] cb_2_8/io_wo[38]
+ cb_2_8/io_wo[39] cb_2_8/io_wo[3] cb_2_8/io_wo[40] cb_2_8/io_wo[41] cb_2_8/io_wo[42]
+ cb_2_8/io_wo[43] cb_2_8/io_wo[44] cb_2_8/io_wo[45] cb_2_8/io_wo[46] cb_2_8/io_wo[47]
+ cb_2_8/io_wo[48] cb_2_8/io_wo[49] cb_2_8/io_wo[4] cb_2_8/io_wo[50] cb_2_8/io_wo[51]
+ cb_2_8/io_wo[52] cb_2_8/io_wo[53] cb_2_8/io_wo[54] cb_2_8/io_wo[55] cb_2_8/io_wo[56]
+ cb_2_8/io_wo[57] cb_2_8/io_wo[58] cb_2_8/io_wo[59] cb_2_8/io_wo[5] cb_2_8/io_wo[60]
+ cb_2_8/io_wo[61] cb_2_8/io_wo[62] cb_2_8/io_wo[63] cb_2_8/io_wo[6] cb_2_8/io_wo[7]
+ cb_2_8/io_wo[8] cb_2_8/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_5_10 cb_5_9/io_adr_i[0] cb_5_9/io_adr_i[1] cb_5_10/io_cs_i cb_5_9/io_dat_i[0]
+ cb_5_9/io_dat_i[10] cb_5_9/io_dat_i[11] cb_5_9/io_dat_i[12] cb_5_9/io_dat_i[13]
+ cb_5_9/io_dat_i[14] cb_5_9/io_dat_i[15] cb_5_9/io_dat_i[1] cb_5_9/io_dat_i[2] cb_5_9/io_dat_i[3]
+ cb_5_9/io_dat_i[4] cb_5_9/io_dat_i[5] cb_5_9/io_dat_i[6] cb_5_9/io_dat_i[7] cb_5_9/io_dat_i[8]
+ cb_5_9/io_dat_i[9] cb_5_10/io_dat_o[0] cb_5_10/io_dat_o[10] cb_5_10/io_dat_o[11]
+ cb_5_10/io_dat_o[12] cb_5_10/io_dat_o[13] cb_5_10/io_dat_o[14] cb_5_10/io_dat_o[15]
+ cb_5_10/io_dat_o[1] cb_5_10/io_dat_o[2] cb_5_10/io_dat_o[3] cb_5_10/io_dat_o[4]
+ cb_5_10/io_dat_o[5] cb_5_10/io_dat_o[6] cb_5_10/io_dat_o[7] cb_5_10/io_dat_o[8]
+ cb_5_10/io_dat_o[9] cb_5_10/io_eo[0] cb_5_10/io_eo[10] cb_5_10/io_eo[11] cb_5_10/io_eo[12]
+ cb_5_10/io_eo[13] cb_5_10/io_eo[14] cb_5_10/io_eo[15] cb_5_10/io_eo[16] cb_5_10/io_eo[17]
+ cb_5_10/io_eo[18] cb_5_10/io_eo[19] cb_5_10/io_eo[1] cb_5_10/io_eo[20] cb_5_10/io_eo[21]
+ cb_5_10/io_eo[22] cb_5_10/io_eo[23] cb_5_10/io_eo[24] cb_5_10/io_eo[25] cb_5_10/io_eo[26]
+ cb_5_10/io_eo[27] cb_5_10/io_eo[28] cb_5_10/io_eo[29] cb_5_10/io_eo[2] cb_5_10/io_eo[30]
+ cb_5_10/io_eo[31] cb_5_10/io_eo[32] cb_5_10/io_eo[33] cb_5_10/io_eo[34] cb_5_10/io_eo[35]
+ cb_5_10/io_eo[36] cb_5_10/io_eo[37] cb_5_10/io_eo[38] cb_5_10/io_eo[39] cb_5_10/io_eo[3]
+ cb_5_10/io_eo[40] cb_5_10/io_eo[41] cb_5_10/io_eo[42] cb_5_10/io_eo[43] cb_5_10/io_eo[44]
+ cb_5_10/io_eo[45] cb_5_10/io_eo[46] cb_5_10/io_eo[47] cb_5_10/io_eo[48] cb_5_10/io_eo[49]
+ cb_5_10/io_eo[4] cb_5_10/io_eo[50] cb_5_10/io_eo[51] cb_5_10/io_eo[52] cb_5_10/io_eo[53]
+ cb_5_10/io_eo[54] cb_5_10/io_eo[55] cb_5_10/io_eo[56] cb_5_10/io_eo[57] cb_5_10/io_eo[58]
+ cb_5_10/io_eo[59] cb_5_10/io_eo[5] cb_5_10/io_eo[60] cb_5_10/io_eo[61] cb_5_10/io_eo[62]
+ cb_5_10/io_eo[63] cb_5_10/io_eo[6] cb_5_10/io_eo[7] cb_5_10/io_eo[8] cb_5_10/io_eo[9]
+ cb_5_9/io_o_0_co cb_5_9/io_o_0_out[0] cb_5_9/io_o_0_out[1] cb_5_9/io_o_0_out[2]
+ cb_5_9/io_o_0_out[3] cb_5_9/io_o_0_out[4] cb_5_9/io_o_0_out[5] cb_5_9/io_o_0_out[6]
+ cb_5_9/io_o_0_out[7] cb_5_9/io_o_1_co cb_5_9/io_o_1_out[0] cb_5_9/io_o_1_out[1]
+ cb_5_9/io_o_1_out[2] cb_5_9/io_o_1_out[3] cb_5_9/io_o_1_out[4] cb_5_9/io_o_1_out[5]
+ cb_5_9/io_o_1_out[6] cb_5_9/io_o_1_out[7] cb_5_9/io_o_2_co cb_5_9/io_o_2_out[0]
+ cb_5_9/io_o_2_out[1] cb_5_9/io_o_2_out[2] cb_5_9/io_o_2_out[3] cb_5_9/io_o_2_out[4]
+ cb_5_9/io_o_2_out[5] cb_5_9/io_o_2_out[6] cb_5_9/io_o_2_out[7] cb_5_9/io_o_3_co
+ cb_5_9/io_o_3_out[0] cb_5_9/io_o_3_out[1] cb_5_9/io_o_3_out[2] cb_5_9/io_o_3_out[3]
+ cb_5_9/io_o_3_out[4] cb_5_9/io_o_3_out[5] cb_5_9/io_o_3_out[6] cb_5_9/io_o_3_out[7]
+ cb_5_9/io_o_4_co cb_5_9/io_o_4_out[0] cb_5_9/io_o_4_out[1] cb_5_9/io_o_4_out[2]
+ cb_5_9/io_o_4_out[3] cb_5_9/io_o_4_out[4] cb_5_9/io_o_4_out[5] cb_5_9/io_o_4_out[6]
+ cb_5_9/io_o_4_out[7] cb_5_9/io_o_5_co cb_5_9/io_o_5_out[0] cb_5_9/io_o_5_out[1]
+ cb_5_9/io_o_5_out[2] cb_5_9/io_o_5_out[3] cb_5_9/io_o_5_out[4] cb_5_9/io_o_5_out[5]
+ cb_5_9/io_o_5_out[6] cb_5_9/io_o_5_out[7] cb_5_9/io_o_6_co cb_5_9/io_o_6_out[0]
+ cb_5_9/io_o_6_out[1] cb_5_9/io_o_6_out[2] cb_5_9/io_o_6_out[3] cb_5_9/io_o_6_out[4]
+ cb_5_9/io_o_6_out[5] cb_5_9/io_o_6_out[6] cb_5_9/io_o_6_out[7] cb_5_9/io_o_7_co
+ cb_5_9/io_o_7_out[0] cb_5_9/io_o_7_out[1] cb_5_9/io_o_7_out[2] cb_5_9/io_o_7_out[3]
+ cb_5_9/io_o_7_out[4] cb_5_9/io_o_7_out[5] cb_5_9/io_o_7_out[6] cb_5_9/io_o_7_out[7]
+ cb_5_10/io_o_0_co cb_5_10/io_eo[0] cb_5_10/io_eo[1] cb_5_10/io_eo[2] cb_5_10/io_eo[3]
+ cb_5_10/io_eo[4] cb_5_10/io_eo[5] cb_5_10/io_eo[6] cb_5_10/io_eo[7] cb_5_10/io_o_1_co
+ cb_5_10/io_eo[8] cb_5_10/io_eo[9] cb_5_10/io_eo[10] cb_5_10/io_eo[11] cb_5_10/io_eo[12]
+ cb_5_10/io_eo[13] cb_5_10/io_eo[14] cb_5_10/io_eo[15] cb_5_10/io_o_2_co cb_5_10/io_eo[16]
+ cb_5_10/io_eo[17] cb_5_10/io_eo[18] cb_5_10/io_eo[19] cb_5_10/io_eo[20] cb_5_10/io_eo[21]
+ cb_5_10/io_eo[22] cb_5_10/io_eo[23] cb_5_10/io_o_3_co cb_5_10/io_eo[24] cb_5_10/io_eo[25]
+ cb_5_10/io_eo[26] cb_5_10/io_eo[27] cb_5_10/io_eo[28] cb_5_10/io_eo[29] cb_5_10/io_eo[30]
+ cb_5_10/io_eo[31] cb_5_10/io_o_4_co cb_5_10/io_eo[32] cb_5_10/io_eo[33] cb_5_10/io_eo[34]
+ cb_5_10/io_eo[35] cb_5_10/io_eo[36] cb_5_10/io_eo[37] cb_5_10/io_eo[38] cb_5_10/io_eo[39]
+ cb_5_10/io_o_5_co cb_5_10/io_eo[40] cb_5_10/io_eo[41] cb_5_10/io_eo[42] cb_5_10/io_eo[43]
+ cb_5_10/io_eo[44] cb_5_10/io_eo[45] cb_5_10/io_eo[46] cb_5_10/io_eo[47] cb_5_10/io_o_6_co
+ cb_5_10/io_eo[48] cb_5_10/io_eo[49] cb_5_10/io_eo[50] cb_5_10/io_eo[51] cb_5_10/io_eo[52]
+ cb_5_10/io_eo[53] cb_5_10/io_eo[54] cb_5_10/io_eo[55] cb_5_10/io_o_7_co cb_5_10/io_eo[56]
+ cb_5_10/io_eo[57] cb_5_10/io_eo[58] cb_5_10/io_eo[59] cb_5_10/io_eo[60] cb_5_10/io_eo[61]
+ cb_5_10/io_eo[62] cb_5_10/io_eo[63] cb_5_9/io_vco cb_5_10/io_vco cb_5_10/io_vi cb_5_9/io_we_i
+ cb_5_9/io_eo[0] cb_5_9/io_eo[10] cb_5_9/io_eo[11] cb_5_9/io_eo[12] cb_5_9/io_eo[13]
+ cb_5_9/io_eo[14] cb_5_9/io_eo[15] cb_5_9/io_eo[16] cb_5_9/io_eo[17] cb_5_9/io_eo[18]
+ cb_5_9/io_eo[19] cb_5_9/io_eo[1] cb_5_9/io_eo[20] cb_5_9/io_eo[21] cb_5_9/io_eo[22]
+ cb_5_9/io_eo[23] cb_5_9/io_eo[24] cb_5_9/io_eo[25] cb_5_9/io_eo[26] cb_5_9/io_eo[27]
+ cb_5_9/io_eo[28] cb_5_9/io_eo[29] cb_5_9/io_eo[2] cb_5_9/io_eo[30] cb_5_9/io_eo[31]
+ cb_5_9/io_eo[32] cb_5_9/io_eo[33] cb_5_9/io_eo[34] cb_5_9/io_eo[35] cb_5_9/io_eo[36]
+ cb_5_9/io_eo[37] cb_5_9/io_eo[38] cb_5_9/io_eo[39] cb_5_9/io_eo[3] cb_5_9/io_eo[40]
+ cb_5_9/io_eo[41] cb_5_9/io_eo[42] cb_5_9/io_eo[43] cb_5_9/io_eo[44] cb_5_9/io_eo[45]
+ cb_5_9/io_eo[46] cb_5_9/io_eo[47] cb_5_9/io_eo[48] cb_5_9/io_eo[49] cb_5_9/io_eo[4]
+ cb_5_9/io_eo[50] cb_5_9/io_eo[51] cb_5_9/io_eo[52] cb_5_9/io_eo[53] cb_5_9/io_eo[54]
+ cb_5_9/io_eo[55] cb_5_9/io_eo[56] cb_5_9/io_eo[57] cb_5_9/io_eo[58] cb_5_9/io_eo[59]
+ cb_5_9/io_eo[5] cb_5_9/io_eo[60] cb_5_9/io_eo[61] cb_5_9/io_eo[62] cb_5_9/io_eo[63]
+ cb_5_9/io_eo[6] cb_5_9/io_eo[7] cb_5_9/io_eo[8] cb_5_9/io_eo[9] mcons_3/clock mcons_3/reset
+ vccd1 vssd1 cic_block
Xcb_2_9 cb_2_9/io_adr_i[0] cb_2_9/io_adr_i[1] cb_2_9/io_cs_i cb_2_9/io_dat_i[0] cb_2_9/io_dat_i[10]
+ cb_2_9/io_dat_i[11] cb_2_9/io_dat_i[12] cb_2_9/io_dat_i[13] cb_2_9/io_dat_i[14]
+ cb_2_9/io_dat_i[15] cb_2_9/io_dat_i[1] cb_2_9/io_dat_i[2] cb_2_9/io_dat_i[3] cb_2_9/io_dat_i[4]
+ cb_2_9/io_dat_i[5] cb_2_9/io_dat_i[6] cb_2_9/io_dat_i[7] cb_2_9/io_dat_i[8] cb_2_9/io_dat_i[9]
+ cb_2_9/io_dat_o[0] cb_2_9/io_dat_o[10] cb_2_9/io_dat_o[11] cb_2_9/io_dat_o[12] cb_2_9/io_dat_o[13]
+ cb_2_9/io_dat_o[14] cb_2_9/io_dat_o[15] cb_2_9/io_dat_o[1] cb_2_9/io_dat_o[2] cb_2_9/io_dat_o[3]
+ cb_2_9/io_dat_o[4] cb_2_9/io_dat_o[5] cb_2_9/io_dat_o[6] cb_2_9/io_dat_o[7] cb_2_9/io_dat_o[8]
+ cb_2_9/io_dat_o[9] cb_2_9/io_eo[0] cb_2_9/io_eo[10] cb_2_9/io_eo[11] cb_2_9/io_eo[12]
+ cb_2_9/io_eo[13] cb_2_9/io_eo[14] cb_2_9/io_eo[15] cb_2_9/io_eo[16] cb_2_9/io_eo[17]
+ cb_2_9/io_eo[18] cb_2_9/io_eo[19] cb_2_9/io_eo[1] cb_2_9/io_eo[20] cb_2_9/io_eo[21]
+ cb_2_9/io_eo[22] cb_2_9/io_eo[23] cb_2_9/io_eo[24] cb_2_9/io_eo[25] cb_2_9/io_eo[26]
+ cb_2_9/io_eo[27] cb_2_9/io_eo[28] cb_2_9/io_eo[29] cb_2_9/io_eo[2] cb_2_9/io_eo[30]
+ cb_2_9/io_eo[31] cb_2_9/io_eo[32] cb_2_9/io_eo[33] cb_2_9/io_eo[34] cb_2_9/io_eo[35]
+ cb_2_9/io_eo[36] cb_2_9/io_eo[37] cb_2_9/io_eo[38] cb_2_9/io_eo[39] cb_2_9/io_eo[3]
+ cb_2_9/io_eo[40] cb_2_9/io_eo[41] cb_2_9/io_eo[42] cb_2_9/io_eo[43] cb_2_9/io_eo[44]
+ cb_2_9/io_eo[45] cb_2_9/io_eo[46] cb_2_9/io_eo[47] cb_2_9/io_eo[48] cb_2_9/io_eo[49]
+ cb_2_9/io_eo[4] cb_2_9/io_eo[50] cb_2_9/io_eo[51] cb_2_9/io_eo[52] cb_2_9/io_eo[53]
+ cb_2_9/io_eo[54] cb_2_9/io_eo[55] cb_2_9/io_eo[56] cb_2_9/io_eo[57] cb_2_9/io_eo[58]
+ cb_2_9/io_eo[59] cb_2_9/io_eo[5] cb_2_9/io_eo[60] cb_2_9/io_eo[61] cb_2_9/io_eo[62]
+ cb_2_9/io_eo[63] cb_2_9/io_eo[6] cb_2_9/io_eo[7] cb_2_9/io_eo[8] cb_2_9/io_eo[9]
+ cb_2_9/io_i_0_ci cb_2_9/io_i_0_in1[0] cb_2_9/io_i_0_in1[1] cb_2_9/io_i_0_in1[2]
+ cb_2_9/io_i_0_in1[3] cb_2_9/io_i_0_in1[4] cb_2_9/io_i_0_in1[5] cb_2_9/io_i_0_in1[6]
+ cb_2_9/io_i_0_in1[7] cb_2_9/io_i_1_ci cb_2_9/io_i_1_in1[0] cb_2_9/io_i_1_in1[1]
+ cb_2_9/io_i_1_in1[2] cb_2_9/io_i_1_in1[3] cb_2_9/io_i_1_in1[4] cb_2_9/io_i_1_in1[5]
+ cb_2_9/io_i_1_in1[6] cb_2_9/io_i_1_in1[7] cb_2_9/io_i_2_ci cb_2_9/io_i_2_in1[0]
+ cb_2_9/io_i_2_in1[1] cb_2_9/io_i_2_in1[2] cb_2_9/io_i_2_in1[3] cb_2_9/io_i_2_in1[4]
+ cb_2_9/io_i_2_in1[5] cb_2_9/io_i_2_in1[6] cb_2_9/io_i_2_in1[7] cb_2_9/io_i_3_ci
+ cb_2_9/io_i_3_in1[0] cb_2_9/io_i_3_in1[1] cb_2_9/io_i_3_in1[2] cb_2_9/io_i_3_in1[3]
+ cb_2_9/io_i_3_in1[4] cb_2_9/io_i_3_in1[5] cb_2_9/io_i_3_in1[6] cb_2_9/io_i_3_in1[7]
+ cb_2_9/io_i_4_ci cb_2_9/io_i_4_in1[0] cb_2_9/io_i_4_in1[1] cb_2_9/io_i_4_in1[2]
+ cb_2_9/io_i_4_in1[3] cb_2_9/io_i_4_in1[4] cb_2_9/io_i_4_in1[5] cb_2_9/io_i_4_in1[6]
+ cb_2_9/io_i_4_in1[7] cb_2_9/io_i_5_ci cb_2_9/io_i_5_in1[0] cb_2_9/io_i_5_in1[1]
+ cb_2_9/io_i_5_in1[2] cb_2_9/io_i_5_in1[3] cb_2_9/io_i_5_in1[4] cb_2_9/io_i_5_in1[5]
+ cb_2_9/io_i_5_in1[6] cb_2_9/io_i_5_in1[7] cb_2_9/io_i_6_ci cb_2_9/io_i_6_in1[0]
+ cb_2_9/io_i_6_in1[1] cb_2_9/io_i_6_in1[2] cb_2_9/io_i_6_in1[3] cb_2_9/io_i_6_in1[4]
+ cb_2_9/io_i_6_in1[5] cb_2_9/io_i_6_in1[6] cb_2_9/io_i_6_in1[7] cb_2_9/io_i_7_ci
+ cb_2_9/io_i_7_in1[0] cb_2_9/io_i_7_in1[1] cb_2_9/io_i_7_in1[2] cb_2_9/io_i_7_in1[3]
+ cb_2_9/io_i_7_in1[4] cb_2_9/io_i_7_in1[5] cb_2_9/io_i_7_in1[6] cb_2_9/io_i_7_in1[7]
+ cb_2_9/io_o_0_co cb_2_9/io_o_0_out[0] cb_2_9/io_o_0_out[1] cb_2_9/io_o_0_out[2]
+ cb_2_9/io_o_0_out[3] cb_2_9/io_o_0_out[4] cb_2_9/io_o_0_out[5] cb_2_9/io_o_0_out[6]
+ cb_2_9/io_o_0_out[7] cb_2_9/io_o_1_co cb_2_9/io_o_1_out[0] cb_2_9/io_o_1_out[1]
+ cb_2_9/io_o_1_out[2] cb_2_9/io_o_1_out[3] cb_2_9/io_o_1_out[4] cb_2_9/io_o_1_out[5]
+ cb_2_9/io_o_1_out[6] cb_2_9/io_o_1_out[7] cb_2_9/io_o_2_co cb_2_9/io_o_2_out[0]
+ cb_2_9/io_o_2_out[1] cb_2_9/io_o_2_out[2] cb_2_9/io_o_2_out[3] cb_2_9/io_o_2_out[4]
+ cb_2_9/io_o_2_out[5] cb_2_9/io_o_2_out[6] cb_2_9/io_o_2_out[7] cb_2_9/io_o_3_co
+ cb_2_9/io_o_3_out[0] cb_2_9/io_o_3_out[1] cb_2_9/io_o_3_out[2] cb_2_9/io_o_3_out[3]
+ cb_2_9/io_o_3_out[4] cb_2_9/io_o_3_out[5] cb_2_9/io_o_3_out[6] cb_2_9/io_o_3_out[7]
+ cb_2_9/io_o_4_co cb_2_9/io_o_4_out[0] cb_2_9/io_o_4_out[1] cb_2_9/io_o_4_out[2]
+ cb_2_9/io_o_4_out[3] cb_2_9/io_o_4_out[4] cb_2_9/io_o_4_out[5] cb_2_9/io_o_4_out[6]
+ cb_2_9/io_o_4_out[7] cb_2_9/io_o_5_co cb_2_9/io_o_5_out[0] cb_2_9/io_o_5_out[1]
+ cb_2_9/io_o_5_out[2] cb_2_9/io_o_5_out[3] cb_2_9/io_o_5_out[4] cb_2_9/io_o_5_out[5]
+ cb_2_9/io_o_5_out[6] cb_2_9/io_o_5_out[7] cb_2_9/io_o_6_co cb_2_9/io_o_6_out[0]
+ cb_2_9/io_o_6_out[1] cb_2_9/io_o_6_out[2] cb_2_9/io_o_6_out[3] cb_2_9/io_o_6_out[4]
+ cb_2_9/io_o_6_out[5] cb_2_9/io_o_6_out[6] cb_2_9/io_o_6_out[7] cb_2_9/io_o_7_co
+ cb_2_9/io_o_7_out[0] cb_2_9/io_o_7_out[1] cb_2_9/io_o_7_out[2] cb_2_9/io_o_7_out[3]
+ cb_2_9/io_o_7_out[4] cb_2_9/io_o_7_out[5] cb_2_9/io_o_7_out[6] cb_2_9/io_o_7_out[7]
+ cb_2_9/io_vci cb_2_9/io_vco cb_2_9/io_vi cb_2_9/io_we_i cb_2_9/io_wo[0] cb_2_9/io_wo[10]
+ cb_2_9/io_wo[11] cb_2_9/io_wo[12] cb_2_9/io_wo[13] cb_2_9/io_wo[14] cb_2_9/io_wo[15]
+ cb_2_9/io_wo[16] cb_2_9/io_wo[17] cb_2_9/io_wo[18] cb_2_9/io_wo[19] cb_2_9/io_wo[1]
+ cb_2_9/io_wo[20] cb_2_9/io_wo[21] cb_2_9/io_wo[22] cb_2_9/io_wo[23] cb_2_9/io_wo[24]
+ cb_2_9/io_wo[25] cb_2_9/io_wo[26] cb_2_9/io_wo[27] cb_2_9/io_wo[28] cb_2_9/io_wo[29]
+ cb_2_9/io_wo[2] cb_2_9/io_wo[30] cb_2_9/io_wo[31] cb_2_9/io_wo[32] cb_2_9/io_wo[33]
+ cb_2_9/io_wo[34] cb_2_9/io_wo[35] cb_2_9/io_wo[36] cb_2_9/io_wo[37] cb_2_9/io_wo[38]
+ cb_2_9/io_wo[39] cb_2_9/io_wo[3] cb_2_9/io_wo[40] cb_2_9/io_wo[41] cb_2_9/io_wo[42]
+ cb_2_9/io_wo[43] cb_2_9/io_wo[44] cb_2_9/io_wo[45] cb_2_9/io_wo[46] cb_2_9/io_wo[47]
+ cb_2_9/io_wo[48] cb_2_9/io_wo[49] cb_2_9/io_wo[4] cb_2_9/io_wo[50] cb_2_9/io_wo[51]
+ cb_2_9/io_wo[52] cb_2_9/io_wo[53] cb_2_9/io_wo[54] cb_2_9/io_wo[55] cb_2_9/io_wo[56]
+ cb_2_9/io_wo[57] cb_2_9/io_wo[58] cb_2_9/io_wo[59] cb_2_9/io_wo[5] cb_2_9/io_wo[60]
+ cb_2_9/io_wo[61] cb_2_9/io_wo[62] cb_2_9/io_wo[63] cb_2_9/io_wo[6] cb_2_9/io_wo[7]
+ cb_2_9/io_wo[8] cb_2_9/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_0_6 cb_0_9/io_adr_i[0] cb_0_9/io_adr_i[1] cb_0_6/io_cs_i cb_0_9/io_dat_i[0] cb_0_9/io_dat_i[10]
+ cb_0_9/io_dat_i[11] cb_0_9/io_dat_i[12] cb_0_9/io_dat_i[13] cb_0_9/io_dat_i[14]
+ cb_0_9/io_dat_i[15] cb_0_9/io_dat_i[1] cb_0_9/io_dat_i[2] cb_0_9/io_dat_i[3] cb_0_9/io_dat_i[4]
+ cb_0_9/io_dat_i[5] cb_0_9/io_dat_i[6] cb_0_9/io_dat_i[7] cb_0_9/io_dat_i[8] cb_0_9/io_dat_i[9]
+ cb_0_6/io_dat_o[0] cb_0_6/io_dat_o[10] cb_0_6/io_dat_o[11] cb_0_6/io_dat_o[12] cb_0_6/io_dat_o[13]
+ cb_0_6/io_dat_o[14] cb_0_6/io_dat_o[15] cb_0_6/io_dat_o[1] cb_0_6/io_dat_o[2] cb_0_6/io_dat_o[3]
+ cb_0_6/io_dat_o[4] cb_0_6/io_dat_o[5] cb_0_6/io_dat_o[6] cb_0_6/io_dat_o[7] cb_0_6/io_dat_o[8]
+ cb_0_6/io_dat_o[9] cb_0_7/io_wo[0] cb_0_7/io_wo[10] cb_0_7/io_wo[11] cb_0_7/io_wo[12]
+ cb_0_7/io_wo[13] cb_0_7/io_wo[14] cb_0_7/io_wo[15] cb_0_7/io_wo[16] cb_0_7/io_wo[17]
+ cb_0_7/io_wo[18] cb_0_7/io_wo[19] cb_0_7/io_wo[1] cb_0_7/io_wo[20] cb_0_7/io_wo[21]
+ cb_0_7/io_wo[22] cb_0_7/io_wo[23] cb_0_7/io_wo[24] cb_0_7/io_wo[25] cb_0_7/io_wo[26]
+ cb_0_7/io_wo[27] cb_0_7/io_wo[28] cb_0_7/io_wo[29] cb_0_7/io_wo[2] cb_0_7/io_wo[30]
+ cb_0_7/io_wo[31] cb_0_7/io_wo[32] cb_0_7/io_wo[33] cb_0_7/io_wo[34] cb_0_7/io_wo[35]
+ cb_0_7/io_wo[36] cb_0_7/io_wo[37] cb_0_7/io_wo[38] cb_0_7/io_wo[39] cb_0_7/io_wo[3]
+ cb_0_7/io_wo[40] cb_0_7/io_wo[41] cb_0_7/io_wo[42] cb_0_7/io_wo[43] cb_0_7/io_wo[44]
+ cb_0_7/io_wo[45] cb_0_7/io_wo[46] cb_0_7/io_wo[47] cb_0_7/io_wo[48] cb_0_7/io_wo[49]
+ cb_0_7/io_wo[4] cb_0_7/io_wo[50] cb_0_7/io_wo[51] cb_0_7/io_wo[52] cb_0_7/io_wo[53]
+ cb_0_7/io_wo[54] cb_0_7/io_wo[55] cb_0_7/io_wo[56] cb_0_7/io_wo[57] cb_0_7/io_wo[58]
+ cb_0_7/io_wo[59] cb_0_7/io_wo[5] cb_0_7/io_wo[60] cb_0_7/io_wo[61] cb_0_7/io_wo[62]
+ cb_0_7/io_wo[63] cb_0_7/io_wo[6] cb_0_7/io_wo[7] cb_0_7/io_wo[8] cb_0_7/io_wo[9]
+ cb_0_6/io_i_0_ci cb_0_6/io_i_0_in1[0] cb_0_6/io_i_0_in1[1] cb_0_6/io_i_0_in1[2]
+ cb_0_6/io_i_0_in1[3] cb_0_6/io_i_0_in1[4] cb_0_6/io_i_0_in1[5] cb_0_6/io_i_0_in1[6]
+ cb_0_6/io_i_0_in1[7] cb_0_6/io_i_1_ci cb_0_6/io_i_1_in1[0] cb_0_6/io_i_1_in1[1]
+ cb_0_6/io_i_1_in1[2] cb_0_6/io_i_1_in1[3] cb_0_6/io_i_1_in1[4] cb_0_6/io_i_1_in1[5]
+ cb_0_6/io_i_1_in1[6] cb_0_6/io_i_1_in1[7] cb_0_6/io_i_2_ci cb_0_6/io_i_2_in1[0]
+ cb_0_6/io_i_2_in1[1] cb_0_6/io_i_2_in1[2] cb_0_6/io_i_2_in1[3] cb_0_6/io_i_2_in1[4]
+ cb_0_6/io_i_2_in1[5] cb_0_6/io_i_2_in1[6] cb_0_6/io_i_2_in1[7] cb_0_6/io_i_3_ci
+ cb_0_6/io_i_3_in1[0] cb_0_6/io_i_3_in1[1] cb_0_6/io_i_3_in1[2] cb_0_6/io_i_3_in1[3]
+ cb_0_6/io_i_3_in1[4] cb_0_6/io_i_3_in1[5] cb_0_6/io_i_3_in1[6] cb_0_6/io_i_3_in1[7]
+ cb_0_6/io_i_4_ci cb_0_6/io_i_4_in1[0] cb_0_6/io_i_4_in1[1] cb_0_6/io_i_4_in1[2]
+ cb_0_6/io_i_4_in1[3] cb_0_6/io_i_4_in1[4] cb_0_6/io_i_4_in1[5] cb_0_6/io_i_4_in1[6]
+ cb_0_6/io_i_4_in1[7] cb_0_6/io_i_5_ci cb_0_6/io_i_5_in1[0] cb_0_6/io_i_5_in1[1]
+ cb_0_6/io_i_5_in1[2] cb_0_6/io_i_5_in1[3] cb_0_6/io_i_5_in1[4] cb_0_6/io_i_5_in1[5]
+ cb_0_6/io_i_5_in1[6] cb_0_6/io_i_5_in1[7] cb_0_6/io_i_6_ci cb_0_6/io_i_6_in1[0]
+ cb_0_6/io_i_6_in1[1] cb_0_6/io_i_6_in1[2] cb_0_6/io_i_6_in1[3] cb_0_6/io_i_6_in1[4]
+ cb_0_6/io_i_6_in1[5] cb_0_6/io_i_6_in1[6] cb_0_6/io_i_6_in1[7] cb_0_6/io_i_7_ci
+ cb_0_6/io_i_7_in1[0] cb_0_6/io_i_7_in1[1] cb_0_6/io_i_7_in1[2] cb_0_6/io_i_7_in1[3]
+ cb_0_6/io_i_7_in1[4] cb_0_6/io_i_7_in1[5] cb_0_6/io_i_7_in1[6] cb_0_6/io_i_7_in1[7]
+ cb_0_7/io_i_0_ci cb_0_7/io_i_0_in1[0] cb_0_7/io_i_0_in1[1] cb_0_7/io_i_0_in1[2]
+ cb_0_7/io_i_0_in1[3] cb_0_7/io_i_0_in1[4] cb_0_7/io_i_0_in1[5] cb_0_7/io_i_0_in1[6]
+ cb_0_7/io_i_0_in1[7] cb_0_7/io_i_1_ci cb_0_7/io_i_1_in1[0] cb_0_7/io_i_1_in1[1]
+ cb_0_7/io_i_1_in1[2] cb_0_7/io_i_1_in1[3] cb_0_7/io_i_1_in1[4] cb_0_7/io_i_1_in1[5]
+ cb_0_7/io_i_1_in1[6] cb_0_7/io_i_1_in1[7] cb_0_7/io_i_2_ci cb_0_7/io_i_2_in1[0]
+ cb_0_7/io_i_2_in1[1] cb_0_7/io_i_2_in1[2] cb_0_7/io_i_2_in1[3] cb_0_7/io_i_2_in1[4]
+ cb_0_7/io_i_2_in1[5] cb_0_7/io_i_2_in1[6] cb_0_7/io_i_2_in1[7] cb_0_7/io_i_3_ci
+ cb_0_7/io_i_3_in1[0] cb_0_7/io_i_3_in1[1] cb_0_7/io_i_3_in1[2] cb_0_7/io_i_3_in1[3]
+ cb_0_7/io_i_3_in1[4] cb_0_7/io_i_3_in1[5] cb_0_7/io_i_3_in1[6] cb_0_7/io_i_3_in1[7]
+ cb_0_7/io_i_4_ci cb_0_7/io_i_4_in1[0] cb_0_7/io_i_4_in1[1] cb_0_7/io_i_4_in1[2]
+ cb_0_7/io_i_4_in1[3] cb_0_7/io_i_4_in1[4] cb_0_7/io_i_4_in1[5] cb_0_7/io_i_4_in1[6]
+ cb_0_7/io_i_4_in1[7] cb_0_7/io_i_5_ci cb_0_7/io_i_5_in1[0] cb_0_7/io_i_5_in1[1]
+ cb_0_7/io_i_5_in1[2] cb_0_7/io_i_5_in1[3] cb_0_7/io_i_5_in1[4] cb_0_7/io_i_5_in1[5]
+ cb_0_7/io_i_5_in1[6] cb_0_7/io_i_5_in1[7] cb_0_7/io_i_6_ci cb_0_7/io_i_6_in1[0]
+ cb_0_7/io_i_6_in1[1] cb_0_7/io_i_6_in1[2] cb_0_7/io_i_6_in1[3] cb_0_7/io_i_6_in1[4]
+ cb_0_7/io_i_6_in1[5] cb_0_7/io_i_6_in1[6] cb_0_7/io_i_6_in1[7] cb_0_7/io_i_7_ci
+ cb_0_7/io_i_7_in1[0] cb_0_7/io_i_7_in1[1] cb_0_7/io_i_7_in1[2] cb_0_7/io_i_7_in1[3]
+ cb_0_7/io_i_7_in1[4] cb_0_7/io_i_7_in1[5] cb_0_7/io_i_7_in1[6] cb_0_7/io_i_7_in1[7]
+ cb_0_6/io_vci cb_0_7/io_vci cb_0_6/io_vi cb_0_9/io_we_i cb_0_6/io_wo[0] cb_0_6/io_wo[10]
+ cb_0_6/io_wo[11] cb_0_6/io_wo[12] cb_0_6/io_wo[13] cb_0_6/io_wo[14] cb_0_6/io_wo[15]
+ cb_0_6/io_wo[16] cb_0_6/io_wo[17] cb_0_6/io_wo[18] cb_0_6/io_wo[19] cb_0_6/io_wo[1]
+ cb_0_6/io_wo[20] cb_0_6/io_wo[21] cb_0_6/io_wo[22] cb_0_6/io_wo[23] cb_0_6/io_wo[24]
+ cb_0_6/io_wo[25] cb_0_6/io_wo[26] cb_0_6/io_wo[27] cb_0_6/io_wo[28] cb_0_6/io_wo[29]
+ cb_0_6/io_wo[2] cb_0_6/io_wo[30] cb_0_6/io_wo[31] cb_0_6/io_wo[32] cb_0_6/io_wo[33]
+ cb_0_6/io_wo[34] cb_0_6/io_wo[35] cb_0_6/io_wo[36] cb_0_6/io_wo[37] cb_0_6/io_wo[38]
+ cb_0_6/io_wo[39] cb_0_6/io_wo[3] cb_0_6/io_wo[40] cb_0_6/io_wo[41] cb_0_6/io_wo[42]
+ cb_0_6/io_wo[43] cb_0_6/io_wo[44] cb_0_6/io_wo[45] cb_0_6/io_wo[46] cb_0_6/io_wo[47]
+ cb_0_6/io_wo[48] cb_0_6/io_wo[49] cb_0_6/io_wo[4] cb_0_6/io_wo[50] cb_0_6/io_wo[51]
+ cb_0_6/io_wo[52] cb_0_6/io_wo[53] cb_0_6/io_wo[54] cb_0_6/io_wo[55] cb_0_6/io_wo[56]
+ cb_0_6/io_wo[57] cb_0_6/io_wo[58] cb_0_6/io_wo[59] cb_0_6/io_wo[5] cb_0_6/io_wo[60]
+ cb_0_6/io_wo[61] cb_0_6/io_wo[62] cb_0_6/io_wo[63] cb_0_6/io_wo[6] cb_0_6/io_wo[7]
+ cb_0_6/io_wo[8] cb_0_6/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_0_7 cb_0_9/io_adr_i[0] cb_0_9/io_adr_i[1] cb_0_7/io_cs_i cb_0_9/io_dat_i[0] cb_0_9/io_dat_i[10]
+ cb_0_9/io_dat_i[11] cb_0_9/io_dat_i[12] cb_0_9/io_dat_i[13] cb_0_9/io_dat_i[14]
+ cb_0_9/io_dat_i[15] cb_0_9/io_dat_i[1] cb_0_9/io_dat_i[2] cb_0_9/io_dat_i[3] cb_0_9/io_dat_i[4]
+ cb_0_9/io_dat_i[5] cb_0_9/io_dat_i[6] cb_0_9/io_dat_i[7] cb_0_9/io_dat_i[8] cb_0_9/io_dat_i[9]
+ cb_0_7/io_dat_o[0] cb_0_7/io_dat_o[10] cb_0_7/io_dat_o[11] cb_0_7/io_dat_o[12] cb_0_7/io_dat_o[13]
+ cb_0_7/io_dat_o[14] cb_0_7/io_dat_o[15] cb_0_7/io_dat_o[1] cb_0_7/io_dat_o[2] cb_0_7/io_dat_o[3]
+ cb_0_7/io_dat_o[4] cb_0_7/io_dat_o[5] cb_0_7/io_dat_o[6] cb_0_7/io_dat_o[7] cb_0_7/io_dat_o[8]
+ cb_0_7/io_dat_o[9] cb_0_8/io_wo[0] cb_0_8/io_wo[10] cb_0_8/io_wo[11] cb_0_8/io_wo[12]
+ cb_0_8/io_wo[13] cb_0_8/io_wo[14] cb_0_8/io_wo[15] cb_0_8/io_wo[16] cb_0_8/io_wo[17]
+ cb_0_8/io_wo[18] cb_0_8/io_wo[19] cb_0_8/io_wo[1] cb_0_8/io_wo[20] cb_0_8/io_wo[21]
+ cb_0_8/io_wo[22] cb_0_8/io_wo[23] cb_0_8/io_wo[24] cb_0_8/io_wo[25] cb_0_8/io_wo[26]
+ cb_0_8/io_wo[27] cb_0_8/io_wo[28] cb_0_8/io_wo[29] cb_0_8/io_wo[2] cb_0_8/io_wo[30]
+ cb_0_8/io_wo[31] cb_0_8/io_wo[32] cb_0_8/io_wo[33] cb_0_8/io_wo[34] cb_0_8/io_wo[35]
+ cb_0_8/io_wo[36] cb_0_8/io_wo[37] cb_0_8/io_wo[38] cb_0_8/io_wo[39] cb_0_8/io_wo[3]
+ cb_0_8/io_wo[40] cb_0_8/io_wo[41] cb_0_8/io_wo[42] cb_0_8/io_wo[43] cb_0_8/io_wo[44]
+ cb_0_8/io_wo[45] cb_0_8/io_wo[46] cb_0_8/io_wo[47] cb_0_8/io_wo[48] cb_0_8/io_wo[49]
+ cb_0_8/io_wo[4] cb_0_8/io_wo[50] cb_0_8/io_wo[51] cb_0_8/io_wo[52] cb_0_8/io_wo[53]
+ cb_0_8/io_wo[54] cb_0_8/io_wo[55] cb_0_8/io_wo[56] cb_0_8/io_wo[57] cb_0_8/io_wo[58]
+ cb_0_8/io_wo[59] cb_0_8/io_wo[5] cb_0_8/io_wo[60] cb_0_8/io_wo[61] cb_0_8/io_wo[62]
+ cb_0_8/io_wo[63] cb_0_8/io_wo[6] cb_0_8/io_wo[7] cb_0_8/io_wo[8] cb_0_8/io_wo[9]
+ cb_0_7/io_i_0_ci cb_0_7/io_i_0_in1[0] cb_0_7/io_i_0_in1[1] cb_0_7/io_i_0_in1[2]
+ cb_0_7/io_i_0_in1[3] cb_0_7/io_i_0_in1[4] cb_0_7/io_i_0_in1[5] cb_0_7/io_i_0_in1[6]
+ cb_0_7/io_i_0_in1[7] cb_0_7/io_i_1_ci cb_0_7/io_i_1_in1[0] cb_0_7/io_i_1_in1[1]
+ cb_0_7/io_i_1_in1[2] cb_0_7/io_i_1_in1[3] cb_0_7/io_i_1_in1[4] cb_0_7/io_i_1_in1[5]
+ cb_0_7/io_i_1_in1[6] cb_0_7/io_i_1_in1[7] cb_0_7/io_i_2_ci cb_0_7/io_i_2_in1[0]
+ cb_0_7/io_i_2_in1[1] cb_0_7/io_i_2_in1[2] cb_0_7/io_i_2_in1[3] cb_0_7/io_i_2_in1[4]
+ cb_0_7/io_i_2_in1[5] cb_0_7/io_i_2_in1[6] cb_0_7/io_i_2_in1[7] cb_0_7/io_i_3_ci
+ cb_0_7/io_i_3_in1[0] cb_0_7/io_i_3_in1[1] cb_0_7/io_i_3_in1[2] cb_0_7/io_i_3_in1[3]
+ cb_0_7/io_i_3_in1[4] cb_0_7/io_i_3_in1[5] cb_0_7/io_i_3_in1[6] cb_0_7/io_i_3_in1[7]
+ cb_0_7/io_i_4_ci cb_0_7/io_i_4_in1[0] cb_0_7/io_i_4_in1[1] cb_0_7/io_i_4_in1[2]
+ cb_0_7/io_i_4_in1[3] cb_0_7/io_i_4_in1[4] cb_0_7/io_i_4_in1[5] cb_0_7/io_i_4_in1[6]
+ cb_0_7/io_i_4_in1[7] cb_0_7/io_i_5_ci cb_0_7/io_i_5_in1[0] cb_0_7/io_i_5_in1[1]
+ cb_0_7/io_i_5_in1[2] cb_0_7/io_i_5_in1[3] cb_0_7/io_i_5_in1[4] cb_0_7/io_i_5_in1[5]
+ cb_0_7/io_i_5_in1[6] cb_0_7/io_i_5_in1[7] cb_0_7/io_i_6_ci cb_0_7/io_i_6_in1[0]
+ cb_0_7/io_i_6_in1[1] cb_0_7/io_i_6_in1[2] cb_0_7/io_i_6_in1[3] cb_0_7/io_i_6_in1[4]
+ cb_0_7/io_i_6_in1[5] cb_0_7/io_i_6_in1[6] cb_0_7/io_i_6_in1[7] cb_0_7/io_i_7_ci
+ cb_0_7/io_i_7_in1[0] cb_0_7/io_i_7_in1[1] cb_0_7/io_i_7_in1[2] cb_0_7/io_i_7_in1[3]
+ cb_0_7/io_i_7_in1[4] cb_0_7/io_i_7_in1[5] cb_0_7/io_i_7_in1[6] cb_0_7/io_i_7_in1[7]
+ cb_0_8/io_i_0_ci cb_0_8/io_i_0_in1[0] cb_0_8/io_i_0_in1[1] cb_0_8/io_i_0_in1[2]
+ cb_0_8/io_i_0_in1[3] cb_0_8/io_i_0_in1[4] cb_0_8/io_i_0_in1[5] cb_0_8/io_i_0_in1[6]
+ cb_0_8/io_i_0_in1[7] cb_0_8/io_i_1_ci cb_0_8/io_i_1_in1[0] cb_0_8/io_i_1_in1[1]
+ cb_0_8/io_i_1_in1[2] cb_0_8/io_i_1_in1[3] cb_0_8/io_i_1_in1[4] cb_0_8/io_i_1_in1[5]
+ cb_0_8/io_i_1_in1[6] cb_0_8/io_i_1_in1[7] cb_0_8/io_i_2_ci cb_0_8/io_i_2_in1[0]
+ cb_0_8/io_i_2_in1[1] cb_0_8/io_i_2_in1[2] cb_0_8/io_i_2_in1[3] cb_0_8/io_i_2_in1[4]
+ cb_0_8/io_i_2_in1[5] cb_0_8/io_i_2_in1[6] cb_0_8/io_i_2_in1[7] cb_0_8/io_i_3_ci
+ cb_0_8/io_i_3_in1[0] cb_0_8/io_i_3_in1[1] cb_0_8/io_i_3_in1[2] cb_0_8/io_i_3_in1[3]
+ cb_0_8/io_i_3_in1[4] cb_0_8/io_i_3_in1[5] cb_0_8/io_i_3_in1[6] cb_0_8/io_i_3_in1[7]
+ cb_0_8/io_i_4_ci cb_0_8/io_i_4_in1[0] cb_0_8/io_i_4_in1[1] cb_0_8/io_i_4_in1[2]
+ cb_0_8/io_i_4_in1[3] cb_0_8/io_i_4_in1[4] cb_0_8/io_i_4_in1[5] cb_0_8/io_i_4_in1[6]
+ cb_0_8/io_i_4_in1[7] cb_0_8/io_i_5_ci cb_0_8/io_i_5_in1[0] cb_0_8/io_i_5_in1[1]
+ cb_0_8/io_i_5_in1[2] cb_0_8/io_i_5_in1[3] cb_0_8/io_i_5_in1[4] cb_0_8/io_i_5_in1[5]
+ cb_0_8/io_i_5_in1[6] cb_0_8/io_i_5_in1[7] cb_0_8/io_i_6_ci cb_0_8/io_i_6_in1[0]
+ cb_0_8/io_i_6_in1[1] cb_0_8/io_i_6_in1[2] cb_0_8/io_i_6_in1[3] cb_0_8/io_i_6_in1[4]
+ cb_0_8/io_i_6_in1[5] cb_0_8/io_i_6_in1[6] cb_0_8/io_i_6_in1[7] cb_0_8/io_i_7_ci
+ cb_0_8/io_i_7_in1[0] cb_0_8/io_i_7_in1[1] cb_0_8/io_i_7_in1[2] cb_0_8/io_i_7_in1[3]
+ cb_0_8/io_i_7_in1[4] cb_0_8/io_i_7_in1[5] cb_0_8/io_i_7_in1[6] cb_0_8/io_i_7_in1[7]
+ cb_0_7/io_vci cb_0_8/io_vci cb_0_7/io_vi cb_0_9/io_we_i cb_0_7/io_wo[0] cb_0_7/io_wo[10]
+ cb_0_7/io_wo[11] cb_0_7/io_wo[12] cb_0_7/io_wo[13] cb_0_7/io_wo[14] cb_0_7/io_wo[15]
+ cb_0_7/io_wo[16] cb_0_7/io_wo[17] cb_0_7/io_wo[18] cb_0_7/io_wo[19] cb_0_7/io_wo[1]
+ cb_0_7/io_wo[20] cb_0_7/io_wo[21] cb_0_7/io_wo[22] cb_0_7/io_wo[23] cb_0_7/io_wo[24]
+ cb_0_7/io_wo[25] cb_0_7/io_wo[26] cb_0_7/io_wo[27] cb_0_7/io_wo[28] cb_0_7/io_wo[29]
+ cb_0_7/io_wo[2] cb_0_7/io_wo[30] cb_0_7/io_wo[31] cb_0_7/io_wo[32] cb_0_7/io_wo[33]
+ cb_0_7/io_wo[34] cb_0_7/io_wo[35] cb_0_7/io_wo[36] cb_0_7/io_wo[37] cb_0_7/io_wo[38]
+ cb_0_7/io_wo[39] cb_0_7/io_wo[3] cb_0_7/io_wo[40] cb_0_7/io_wo[41] cb_0_7/io_wo[42]
+ cb_0_7/io_wo[43] cb_0_7/io_wo[44] cb_0_7/io_wo[45] cb_0_7/io_wo[46] cb_0_7/io_wo[47]
+ cb_0_7/io_wo[48] cb_0_7/io_wo[49] cb_0_7/io_wo[4] cb_0_7/io_wo[50] cb_0_7/io_wo[51]
+ cb_0_7/io_wo[52] cb_0_7/io_wo[53] cb_0_7/io_wo[54] cb_0_7/io_wo[55] cb_0_7/io_wo[56]
+ cb_0_7/io_wo[57] cb_0_7/io_wo[58] cb_0_7/io_wo[59] cb_0_7/io_wo[5] cb_0_7/io_wo[60]
+ cb_0_7/io_wo[61] cb_0_7/io_wo[62] cb_0_7/io_wo[63] cb_0_7/io_wo[6] cb_0_7/io_wo[7]
+ cb_0_7/io_wo[8] cb_0_7/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_7_0 cb_7_9/io_adr_i[0] cb_7_9/io_adr_i[1] cb_7_0/io_cs_i cb_7_9/io_dat_i[0] cb_7_9/io_dat_i[10]
+ cb_7_9/io_dat_i[11] cb_7_9/io_dat_i[12] cb_7_9/io_dat_i[13] cb_7_9/io_dat_i[14]
+ cb_7_9/io_dat_i[15] cb_7_9/io_dat_i[1] cb_7_9/io_dat_i[2] cb_7_9/io_dat_i[3] cb_7_9/io_dat_i[4]
+ cb_7_9/io_dat_i[5] cb_7_9/io_dat_i[6] cb_7_9/io_dat_i[7] cb_7_9/io_dat_i[8] cb_7_9/io_dat_i[9]
+ cb_7_0/io_dat_o[0] cb_7_0/io_dat_o[10] cb_7_0/io_dat_o[11] cb_7_0/io_dat_o[12] cb_7_0/io_dat_o[13]
+ cb_7_0/io_dat_o[14] cb_7_0/io_dat_o[15] cb_7_0/io_dat_o[1] cb_7_0/io_dat_o[2] cb_7_0/io_dat_o[3]
+ cb_7_0/io_dat_o[4] cb_7_0/io_dat_o[5] cb_7_0/io_dat_o[6] cb_7_0/io_dat_o[7] cb_7_0/io_dat_o[8]
+ cb_7_0/io_dat_o[9] cb_7_1/io_wo[0] cb_7_1/io_wo[10] cb_7_1/io_wo[11] cb_7_1/io_wo[12]
+ cb_7_1/io_wo[13] cb_7_1/io_wo[14] cb_7_1/io_wo[15] cb_7_1/io_wo[16] cb_7_1/io_wo[17]
+ cb_7_1/io_wo[18] cb_7_1/io_wo[19] cb_7_1/io_wo[1] cb_7_1/io_wo[20] cb_7_1/io_wo[21]
+ cb_7_1/io_wo[22] cb_7_1/io_wo[23] cb_7_1/io_wo[24] cb_7_1/io_wo[25] cb_7_1/io_wo[26]
+ cb_7_1/io_wo[27] cb_7_1/io_wo[28] cb_7_1/io_wo[29] cb_7_1/io_wo[2] cb_7_1/io_wo[30]
+ cb_7_1/io_wo[31] cb_7_1/io_wo[32] cb_7_1/io_wo[33] cb_7_1/io_wo[34] cb_7_1/io_wo[35]
+ cb_7_1/io_wo[36] cb_7_1/io_wo[37] cb_7_1/io_wo[38] cb_7_1/io_wo[39] cb_7_1/io_wo[3]
+ cb_7_1/io_wo[40] cb_7_1/io_wo[41] cb_7_1/io_wo[42] cb_7_1/io_wo[43] cb_7_1/io_wo[44]
+ cb_7_1/io_wo[45] cb_7_1/io_wo[46] cb_7_1/io_wo[47] cb_7_1/io_wo[48] cb_7_1/io_wo[49]
+ cb_7_1/io_wo[4] cb_7_1/io_wo[50] cb_7_1/io_wo[51] cb_7_1/io_wo[52] cb_7_1/io_wo[53]
+ cb_7_1/io_wo[54] cb_7_1/io_wo[55] cb_7_1/io_wo[56] cb_7_1/io_wo[57] cb_7_1/io_wo[58]
+ cb_7_1/io_wo[59] cb_7_1/io_wo[5] cb_7_1/io_wo[60] cb_7_1/io_wo[61] cb_7_1/io_wo[62]
+ cb_7_1/io_wo[63] cb_7_1/io_wo[6] cb_7_1/io_wo[7] cb_7_1/io_wo[8] cb_7_1/io_wo[9]
+ ccon_7/io_dsi_o cb_7_0/io_i_0_in1[0] cb_7_0/io_i_0_in1[1] cb_7_0/io_i_0_in1[2] cb_7_0/io_i_0_in1[3]
+ cb_7_0/io_i_0_in1[4] cb_7_0/io_i_0_in1[5] cb_7_0/io_i_0_in1[6] cb_7_0/io_i_0_in1[7]
+ cb_7_0/io_i_1_ci cb_7_0/io_i_1_in1[0] cb_7_0/io_i_1_in1[1] cb_7_0/io_i_1_in1[2]
+ cb_7_0/io_i_1_in1[3] cb_7_0/io_i_1_in1[4] cb_7_0/io_i_1_in1[5] cb_7_0/io_i_1_in1[6]
+ cb_7_0/io_i_1_in1[7] cb_7_0/io_i_2_ci cb_7_0/io_i_2_in1[0] cb_7_0/io_i_2_in1[1]
+ cb_7_0/io_i_2_in1[2] cb_7_0/io_i_2_in1[3] cb_7_0/io_i_2_in1[4] cb_7_0/io_i_2_in1[5]
+ cb_7_0/io_i_2_in1[6] cb_7_0/io_i_2_in1[7] cb_7_0/io_i_3_ci cb_7_0/io_i_3_in1[0]
+ cb_7_0/io_i_3_in1[1] cb_7_0/io_i_3_in1[2] cb_7_0/io_i_3_in1[3] cb_7_0/io_i_3_in1[4]
+ cb_7_0/io_i_3_in1[5] cb_7_0/io_i_3_in1[6] cb_7_0/io_i_3_in1[7] cb_7_0/io_i_4_ci
+ cb_7_0/io_i_4_in1[0] cb_7_0/io_i_4_in1[1] cb_7_0/io_i_4_in1[2] cb_7_0/io_i_4_in1[3]
+ cb_7_0/io_i_4_in1[4] cb_7_0/io_i_4_in1[5] cb_7_0/io_i_4_in1[6] cb_7_0/io_i_4_in1[7]
+ cb_7_0/io_i_5_ci cb_7_0/io_i_5_in1[0] cb_7_0/io_i_5_in1[1] cb_7_0/io_i_5_in1[2]
+ cb_7_0/io_i_5_in1[3] cb_7_0/io_i_5_in1[4] cb_7_0/io_i_5_in1[5] cb_7_0/io_i_5_in1[6]
+ cb_7_0/io_i_5_in1[7] cb_7_0/io_i_6_ci cb_7_0/io_i_6_in1[0] cb_7_0/io_i_6_in1[1]
+ cb_7_0/io_i_6_in1[2] cb_7_0/io_i_6_in1[3] cb_7_0/io_i_6_in1[4] cb_7_0/io_i_6_in1[5]
+ cb_7_0/io_i_6_in1[6] cb_7_0/io_i_6_in1[7] cb_7_0/io_i_7_ci cb_7_0/io_i_7_in1[0]
+ cb_7_0/io_i_7_in1[1] cb_7_0/io_i_7_in1[2] cb_7_0/io_i_7_in1[3] cb_7_0/io_i_7_in1[4]
+ cb_7_0/io_i_7_in1[5] cb_7_0/io_i_7_in1[6] cb_7_0/io_i_7_in1[7] cb_7_1/io_i_0_ci
+ cb_7_1/io_i_0_in1[0] cb_7_1/io_i_0_in1[1] cb_7_1/io_i_0_in1[2] cb_7_1/io_i_0_in1[3]
+ cb_7_1/io_i_0_in1[4] cb_7_1/io_i_0_in1[5] cb_7_1/io_i_0_in1[6] cb_7_1/io_i_0_in1[7]
+ cb_7_1/io_i_1_ci cb_7_1/io_i_1_in1[0] cb_7_1/io_i_1_in1[1] cb_7_1/io_i_1_in1[2]
+ cb_7_1/io_i_1_in1[3] cb_7_1/io_i_1_in1[4] cb_7_1/io_i_1_in1[5] cb_7_1/io_i_1_in1[6]
+ cb_7_1/io_i_1_in1[7] cb_7_1/io_i_2_ci cb_7_1/io_i_2_in1[0] cb_7_1/io_i_2_in1[1]
+ cb_7_1/io_i_2_in1[2] cb_7_1/io_i_2_in1[3] cb_7_1/io_i_2_in1[4] cb_7_1/io_i_2_in1[5]
+ cb_7_1/io_i_2_in1[6] cb_7_1/io_i_2_in1[7] cb_7_1/io_i_3_ci cb_7_1/io_i_3_in1[0]
+ cb_7_1/io_i_3_in1[1] cb_7_1/io_i_3_in1[2] cb_7_1/io_i_3_in1[3] cb_7_1/io_i_3_in1[4]
+ cb_7_1/io_i_3_in1[5] cb_7_1/io_i_3_in1[6] cb_7_1/io_i_3_in1[7] cb_7_1/io_i_4_ci
+ cb_7_1/io_i_4_in1[0] cb_7_1/io_i_4_in1[1] cb_7_1/io_i_4_in1[2] cb_7_1/io_i_4_in1[3]
+ cb_7_1/io_i_4_in1[4] cb_7_1/io_i_4_in1[5] cb_7_1/io_i_4_in1[6] cb_7_1/io_i_4_in1[7]
+ cb_7_1/io_i_5_ci cb_7_1/io_i_5_in1[0] cb_7_1/io_i_5_in1[1] cb_7_1/io_i_5_in1[2]
+ cb_7_1/io_i_5_in1[3] cb_7_1/io_i_5_in1[4] cb_7_1/io_i_5_in1[5] cb_7_1/io_i_5_in1[6]
+ cb_7_1/io_i_5_in1[7] cb_7_1/io_i_6_ci cb_7_1/io_i_6_in1[0] cb_7_1/io_i_6_in1[1]
+ cb_7_1/io_i_6_in1[2] cb_7_1/io_i_6_in1[3] cb_7_1/io_i_6_in1[4] cb_7_1/io_i_6_in1[5]
+ cb_7_1/io_i_6_in1[6] cb_7_1/io_i_6_in1[7] cb_7_1/io_i_7_ci cb_7_1/io_i_7_in1[0]
+ cb_7_1/io_i_7_in1[1] cb_7_1/io_i_7_in1[2] cb_7_1/io_i_7_in1[3] cb_7_1/io_i_7_in1[4]
+ cb_7_1/io_i_7_in1[5] cb_7_1/io_i_7_in1[6] cb_7_1/io_i_7_in1[7] cb_7_0/io_vci cb_7_1/io_vci
+ cb_7_0/io_vi cb_7_9/io_we_i cb_7_0/io_wo[0] cb_7_0/io_wo[10] cb_7_0/io_wo[11] cb_7_0/io_wo[12]
+ cb_7_0/io_wo[13] cb_7_0/io_wo[14] cb_7_0/io_wo[15] cb_7_0/io_wo[16] cb_7_0/io_wo[17]
+ cb_7_0/io_wo[18] cb_7_0/io_wo[19] cb_7_0/io_wo[1] cb_7_0/io_wo[20] cb_7_0/io_wo[21]
+ cb_7_0/io_wo[22] cb_7_0/io_wo[23] cb_7_0/io_wo[24] cb_7_0/io_wo[25] cb_7_0/io_wo[26]
+ cb_7_0/io_wo[27] cb_7_0/io_wo[28] cb_7_0/io_wo[29] cb_7_0/io_wo[2] cb_7_0/io_wo[30]
+ cb_7_0/io_wo[31] cb_7_0/io_wo[32] cb_7_0/io_wo[33] cb_7_0/io_wo[34] cb_7_0/io_wo[35]
+ cb_7_0/io_wo[36] cb_7_0/io_wo[37] cb_7_0/io_wo[38] cb_7_0/io_wo[39] cb_7_0/io_wo[3]
+ cb_7_0/io_wo[40] cb_7_0/io_wo[41] cb_7_0/io_wo[42] cb_7_0/io_wo[43] cb_7_0/io_wo[44]
+ cb_7_0/io_wo[45] cb_7_0/io_wo[46] cb_7_0/io_wo[47] cb_7_0/io_wo[48] cb_7_0/io_wo[49]
+ cb_7_0/io_wo[4] cb_7_0/io_wo[50] cb_7_0/io_wo[51] cb_7_0/io_wo[52] cb_7_0/io_wo[53]
+ cb_7_0/io_wo[54] cb_7_0/io_wo[55] cb_7_0/io_wo[56] cb_7_0/io_wo[57] cb_7_0/io_wo[58]
+ cb_7_0/io_wo[59] cb_7_0/io_wo[5] cb_7_0/io_wo[60] cb_7_0/io_wo[61] cb_7_0/io_wo[62]
+ cb_7_0/io_wo[63] cb_7_0/io_wo[6] cb_7_0/io_wo[7] cb_7_0/io_wo[8] cb_7_0/io_wo[9]
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_7_1 cb_7_9/io_adr_i[0] cb_7_9/io_adr_i[1] cb_7_1/io_cs_i cb_7_9/io_dat_i[0] cb_7_9/io_dat_i[10]
+ cb_7_9/io_dat_i[11] cb_7_9/io_dat_i[12] cb_7_9/io_dat_i[13] cb_7_9/io_dat_i[14]
+ cb_7_9/io_dat_i[15] cb_7_9/io_dat_i[1] cb_7_9/io_dat_i[2] cb_7_9/io_dat_i[3] cb_7_9/io_dat_i[4]
+ cb_7_9/io_dat_i[5] cb_7_9/io_dat_i[6] cb_7_9/io_dat_i[7] cb_7_9/io_dat_i[8] cb_7_9/io_dat_i[9]
+ cb_7_1/io_dat_o[0] cb_7_1/io_dat_o[10] cb_7_1/io_dat_o[11] cb_7_1/io_dat_o[12] cb_7_1/io_dat_o[13]
+ cb_7_1/io_dat_o[14] cb_7_1/io_dat_o[15] cb_7_1/io_dat_o[1] cb_7_1/io_dat_o[2] cb_7_1/io_dat_o[3]
+ cb_7_1/io_dat_o[4] cb_7_1/io_dat_o[5] cb_7_1/io_dat_o[6] cb_7_1/io_dat_o[7] cb_7_1/io_dat_o[8]
+ cb_7_1/io_dat_o[9] cb_7_2/io_wo[0] cb_7_2/io_wo[10] cb_7_2/io_wo[11] cb_7_2/io_wo[12]
+ cb_7_2/io_wo[13] cb_7_2/io_wo[14] cb_7_2/io_wo[15] cb_7_2/io_wo[16] cb_7_2/io_wo[17]
+ cb_7_2/io_wo[18] cb_7_2/io_wo[19] cb_7_2/io_wo[1] cb_7_2/io_wo[20] cb_7_2/io_wo[21]
+ cb_7_2/io_wo[22] cb_7_2/io_wo[23] cb_7_2/io_wo[24] cb_7_2/io_wo[25] cb_7_2/io_wo[26]
+ cb_7_2/io_wo[27] cb_7_2/io_wo[28] cb_7_2/io_wo[29] cb_7_2/io_wo[2] cb_7_2/io_wo[30]
+ cb_7_2/io_wo[31] cb_7_2/io_wo[32] cb_7_2/io_wo[33] cb_7_2/io_wo[34] cb_7_2/io_wo[35]
+ cb_7_2/io_wo[36] cb_7_2/io_wo[37] cb_7_2/io_wo[38] cb_7_2/io_wo[39] cb_7_2/io_wo[3]
+ cb_7_2/io_wo[40] cb_7_2/io_wo[41] cb_7_2/io_wo[42] cb_7_2/io_wo[43] cb_7_2/io_wo[44]
+ cb_7_2/io_wo[45] cb_7_2/io_wo[46] cb_7_2/io_wo[47] cb_7_2/io_wo[48] cb_7_2/io_wo[49]
+ cb_7_2/io_wo[4] cb_7_2/io_wo[50] cb_7_2/io_wo[51] cb_7_2/io_wo[52] cb_7_2/io_wo[53]
+ cb_7_2/io_wo[54] cb_7_2/io_wo[55] cb_7_2/io_wo[56] cb_7_2/io_wo[57] cb_7_2/io_wo[58]
+ cb_7_2/io_wo[59] cb_7_2/io_wo[5] cb_7_2/io_wo[60] cb_7_2/io_wo[61] cb_7_2/io_wo[62]
+ cb_7_2/io_wo[63] cb_7_2/io_wo[6] cb_7_2/io_wo[7] cb_7_2/io_wo[8] cb_7_2/io_wo[9]
+ cb_7_1/io_i_0_ci cb_7_1/io_i_0_in1[0] cb_7_1/io_i_0_in1[1] cb_7_1/io_i_0_in1[2]
+ cb_7_1/io_i_0_in1[3] cb_7_1/io_i_0_in1[4] cb_7_1/io_i_0_in1[5] cb_7_1/io_i_0_in1[6]
+ cb_7_1/io_i_0_in1[7] cb_7_1/io_i_1_ci cb_7_1/io_i_1_in1[0] cb_7_1/io_i_1_in1[1]
+ cb_7_1/io_i_1_in1[2] cb_7_1/io_i_1_in1[3] cb_7_1/io_i_1_in1[4] cb_7_1/io_i_1_in1[5]
+ cb_7_1/io_i_1_in1[6] cb_7_1/io_i_1_in1[7] cb_7_1/io_i_2_ci cb_7_1/io_i_2_in1[0]
+ cb_7_1/io_i_2_in1[1] cb_7_1/io_i_2_in1[2] cb_7_1/io_i_2_in1[3] cb_7_1/io_i_2_in1[4]
+ cb_7_1/io_i_2_in1[5] cb_7_1/io_i_2_in1[6] cb_7_1/io_i_2_in1[7] cb_7_1/io_i_3_ci
+ cb_7_1/io_i_3_in1[0] cb_7_1/io_i_3_in1[1] cb_7_1/io_i_3_in1[2] cb_7_1/io_i_3_in1[3]
+ cb_7_1/io_i_3_in1[4] cb_7_1/io_i_3_in1[5] cb_7_1/io_i_3_in1[6] cb_7_1/io_i_3_in1[7]
+ cb_7_1/io_i_4_ci cb_7_1/io_i_4_in1[0] cb_7_1/io_i_4_in1[1] cb_7_1/io_i_4_in1[2]
+ cb_7_1/io_i_4_in1[3] cb_7_1/io_i_4_in1[4] cb_7_1/io_i_4_in1[5] cb_7_1/io_i_4_in1[6]
+ cb_7_1/io_i_4_in1[7] cb_7_1/io_i_5_ci cb_7_1/io_i_5_in1[0] cb_7_1/io_i_5_in1[1]
+ cb_7_1/io_i_5_in1[2] cb_7_1/io_i_5_in1[3] cb_7_1/io_i_5_in1[4] cb_7_1/io_i_5_in1[5]
+ cb_7_1/io_i_5_in1[6] cb_7_1/io_i_5_in1[7] cb_7_1/io_i_6_ci cb_7_1/io_i_6_in1[0]
+ cb_7_1/io_i_6_in1[1] cb_7_1/io_i_6_in1[2] cb_7_1/io_i_6_in1[3] cb_7_1/io_i_6_in1[4]
+ cb_7_1/io_i_6_in1[5] cb_7_1/io_i_6_in1[6] cb_7_1/io_i_6_in1[7] cb_7_1/io_i_7_ci
+ cb_7_1/io_i_7_in1[0] cb_7_1/io_i_7_in1[1] cb_7_1/io_i_7_in1[2] cb_7_1/io_i_7_in1[3]
+ cb_7_1/io_i_7_in1[4] cb_7_1/io_i_7_in1[5] cb_7_1/io_i_7_in1[6] cb_7_1/io_i_7_in1[7]
+ cb_7_2/io_i_0_ci cb_7_2/io_i_0_in1[0] cb_7_2/io_i_0_in1[1] cb_7_2/io_i_0_in1[2]
+ cb_7_2/io_i_0_in1[3] cb_7_2/io_i_0_in1[4] cb_7_2/io_i_0_in1[5] cb_7_2/io_i_0_in1[6]
+ cb_7_2/io_i_0_in1[7] cb_7_2/io_i_1_ci cb_7_2/io_i_1_in1[0] cb_7_2/io_i_1_in1[1]
+ cb_7_2/io_i_1_in1[2] cb_7_2/io_i_1_in1[3] cb_7_2/io_i_1_in1[4] cb_7_2/io_i_1_in1[5]
+ cb_7_2/io_i_1_in1[6] cb_7_2/io_i_1_in1[7] cb_7_2/io_i_2_ci cb_7_2/io_i_2_in1[0]
+ cb_7_2/io_i_2_in1[1] cb_7_2/io_i_2_in1[2] cb_7_2/io_i_2_in1[3] cb_7_2/io_i_2_in1[4]
+ cb_7_2/io_i_2_in1[5] cb_7_2/io_i_2_in1[6] cb_7_2/io_i_2_in1[7] cb_7_2/io_i_3_ci
+ cb_7_2/io_i_3_in1[0] cb_7_2/io_i_3_in1[1] cb_7_2/io_i_3_in1[2] cb_7_2/io_i_3_in1[3]
+ cb_7_2/io_i_3_in1[4] cb_7_2/io_i_3_in1[5] cb_7_2/io_i_3_in1[6] cb_7_2/io_i_3_in1[7]
+ cb_7_2/io_i_4_ci cb_7_2/io_i_4_in1[0] cb_7_2/io_i_4_in1[1] cb_7_2/io_i_4_in1[2]
+ cb_7_2/io_i_4_in1[3] cb_7_2/io_i_4_in1[4] cb_7_2/io_i_4_in1[5] cb_7_2/io_i_4_in1[6]
+ cb_7_2/io_i_4_in1[7] cb_7_2/io_i_5_ci cb_7_2/io_i_5_in1[0] cb_7_2/io_i_5_in1[1]
+ cb_7_2/io_i_5_in1[2] cb_7_2/io_i_5_in1[3] cb_7_2/io_i_5_in1[4] cb_7_2/io_i_5_in1[5]
+ cb_7_2/io_i_5_in1[6] cb_7_2/io_i_5_in1[7] cb_7_2/io_i_6_ci cb_7_2/io_i_6_in1[0]
+ cb_7_2/io_i_6_in1[1] cb_7_2/io_i_6_in1[2] cb_7_2/io_i_6_in1[3] cb_7_2/io_i_6_in1[4]
+ cb_7_2/io_i_6_in1[5] cb_7_2/io_i_6_in1[6] cb_7_2/io_i_6_in1[7] cb_7_2/io_i_7_ci
+ cb_7_2/io_i_7_in1[0] cb_7_2/io_i_7_in1[1] cb_7_2/io_i_7_in1[2] cb_7_2/io_i_7_in1[3]
+ cb_7_2/io_i_7_in1[4] cb_7_2/io_i_7_in1[5] cb_7_2/io_i_7_in1[6] cb_7_2/io_i_7_in1[7]
+ cb_7_1/io_vci cb_7_2/io_vci cb_7_1/io_vi cb_7_9/io_we_i cb_7_1/io_wo[0] cb_7_1/io_wo[10]
+ cb_7_1/io_wo[11] cb_7_1/io_wo[12] cb_7_1/io_wo[13] cb_7_1/io_wo[14] cb_7_1/io_wo[15]
+ cb_7_1/io_wo[16] cb_7_1/io_wo[17] cb_7_1/io_wo[18] cb_7_1/io_wo[19] cb_7_1/io_wo[1]
+ cb_7_1/io_wo[20] cb_7_1/io_wo[21] cb_7_1/io_wo[22] cb_7_1/io_wo[23] cb_7_1/io_wo[24]
+ cb_7_1/io_wo[25] cb_7_1/io_wo[26] cb_7_1/io_wo[27] cb_7_1/io_wo[28] cb_7_1/io_wo[29]
+ cb_7_1/io_wo[2] cb_7_1/io_wo[30] cb_7_1/io_wo[31] cb_7_1/io_wo[32] cb_7_1/io_wo[33]
+ cb_7_1/io_wo[34] cb_7_1/io_wo[35] cb_7_1/io_wo[36] cb_7_1/io_wo[37] cb_7_1/io_wo[38]
+ cb_7_1/io_wo[39] cb_7_1/io_wo[3] cb_7_1/io_wo[40] cb_7_1/io_wo[41] cb_7_1/io_wo[42]
+ cb_7_1/io_wo[43] cb_7_1/io_wo[44] cb_7_1/io_wo[45] cb_7_1/io_wo[46] cb_7_1/io_wo[47]
+ cb_7_1/io_wo[48] cb_7_1/io_wo[49] cb_7_1/io_wo[4] cb_7_1/io_wo[50] cb_7_1/io_wo[51]
+ cb_7_1/io_wo[52] cb_7_1/io_wo[53] cb_7_1/io_wo[54] cb_7_1/io_wo[55] cb_7_1/io_wo[56]
+ cb_7_1/io_wo[57] cb_7_1/io_wo[58] cb_7_1/io_wo[59] cb_7_1/io_wo[5] cb_7_1/io_wo[60]
+ cb_7_1/io_wo[61] cb_7_1/io_wo[62] cb_7_1/io_wo[63] cb_7_1/io_wo[6] cb_7_1/io_wo[7]
+ cb_7_1/io_wo[8] cb_7_1/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_0_8 cb_0_9/io_adr_i[0] cb_0_9/io_adr_i[1] cb_0_8/io_cs_i cb_0_9/io_dat_i[0] cb_0_9/io_dat_i[10]
+ cb_0_9/io_dat_i[11] cb_0_9/io_dat_i[12] cb_0_9/io_dat_i[13] cb_0_9/io_dat_i[14]
+ cb_0_9/io_dat_i[15] cb_0_9/io_dat_i[1] cb_0_9/io_dat_i[2] cb_0_9/io_dat_i[3] cb_0_9/io_dat_i[4]
+ cb_0_9/io_dat_i[5] cb_0_9/io_dat_i[6] cb_0_9/io_dat_i[7] cb_0_9/io_dat_i[8] cb_0_9/io_dat_i[9]
+ cb_0_8/io_dat_o[0] cb_0_8/io_dat_o[10] cb_0_8/io_dat_o[11] cb_0_8/io_dat_o[12] cb_0_8/io_dat_o[13]
+ cb_0_8/io_dat_o[14] cb_0_8/io_dat_o[15] cb_0_8/io_dat_o[1] cb_0_8/io_dat_o[2] cb_0_8/io_dat_o[3]
+ cb_0_8/io_dat_o[4] cb_0_8/io_dat_o[5] cb_0_8/io_dat_o[6] cb_0_8/io_dat_o[7] cb_0_8/io_dat_o[8]
+ cb_0_8/io_dat_o[9] cb_0_9/io_wo[0] cb_0_9/io_wo[10] cb_0_9/io_wo[11] cb_0_9/io_wo[12]
+ cb_0_9/io_wo[13] cb_0_9/io_wo[14] cb_0_9/io_wo[15] cb_0_9/io_wo[16] cb_0_9/io_wo[17]
+ cb_0_9/io_wo[18] cb_0_9/io_wo[19] cb_0_9/io_wo[1] cb_0_9/io_wo[20] cb_0_9/io_wo[21]
+ cb_0_9/io_wo[22] cb_0_9/io_wo[23] cb_0_9/io_wo[24] cb_0_9/io_wo[25] cb_0_9/io_wo[26]
+ cb_0_9/io_wo[27] cb_0_9/io_wo[28] cb_0_9/io_wo[29] cb_0_9/io_wo[2] cb_0_9/io_wo[30]
+ cb_0_9/io_wo[31] cb_0_9/io_wo[32] cb_0_9/io_wo[33] cb_0_9/io_wo[34] cb_0_9/io_wo[35]
+ cb_0_9/io_wo[36] cb_0_9/io_wo[37] cb_0_9/io_wo[38] cb_0_9/io_wo[39] cb_0_9/io_wo[3]
+ cb_0_9/io_wo[40] cb_0_9/io_wo[41] cb_0_9/io_wo[42] cb_0_9/io_wo[43] cb_0_9/io_wo[44]
+ cb_0_9/io_wo[45] cb_0_9/io_wo[46] cb_0_9/io_wo[47] cb_0_9/io_wo[48] cb_0_9/io_wo[49]
+ cb_0_9/io_wo[4] cb_0_9/io_wo[50] cb_0_9/io_wo[51] cb_0_9/io_wo[52] cb_0_9/io_wo[53]
+ cb_0_9/io_wo[54] cb_0_9/io_wo[55] cb_0_9/io_wo[56] cb_0_9/io_wo[57] cb_0_9/io_wo[58]
+ cb_0_9/io_wo[59] cb_0_9/io_wo[5] cb_0_9/io_wo[60] cb_0_9/io_wo[61] cb_0_9/io_wo[62]
+ cb_0_9/io_wo[63] cb_0_9/io_wo[6] cb_0_9/io_wo[7] cb_0_9/io_wo[8] cb_0_9/io_wo[9]
+ cb_0_8/io_i_0_ci cb_0_8/io_i_0_in1[0] cb_0_8/io_i_0_in1[1] cb_0_8/io_i_0_in1[2]
+ cb_0_8/io_i_0_in1[3] cb_0_8/io_i_0_in1[4] cb_0_8/io_i_0_in1[5] cb_0_8/io_i_0_in1[6]
+ cb_0_8/io_i_0_in1[7] cb_0_8/io_i_1_ci cb_0_8/io_i_1_in1[0] cb_0_8/io_i_1_in1[1]
+ cb_0_8/io_i_1_in1[2] cb_0_8/io_i_1_in1[3] cb_0_8/io_i_1_in1[4] cb_0_8/io_i_1_in1[5]
+ cb_0_8/io_i_1_in1[6] cb_0_8/io_i_1_in1[7] cb_0_8/io_i_2_ci cb_0_8/io_i_2_in1[0]
+ cb_0_8/io_i_2_in1[1] cb_0_8/io_i_2_in1[2] cb_0_8/io_i_2_in1[3] cb_0_8/io_i_2_in1[4]
+ cb_0_8/io_i_2_in1[5] cb_0_8/io_i_2_in1[6] cb_0_8/io_i_2_in1[7] cb_0_8/io_i_3_ci
+ cb_0_8/io_i_3_in1[0] cb_0_8/io_i_3_in1[1] cb_0_8/io_i_3_in1[2] cb_0_8/io_i_3_in1[3]
+ cb_0_8/io_i_3_in1[4] cb_0_8/io_i_3_in1[5] cb_0_8/io_i_3_in1[6] cb_0_8/io_i_3_in1[7]
+ cb_0_8/io_i_4_ci cb_0_8/io_i_4_in1[0] cb_0_8/io_i_4_in1[1] cb_0_8/io_i_4_in1[2]
+ cb_0_8/io_i_4_in1[3] cb_0_8/io_i_4_in1[4] cb_0_8/io_i_4_in1[5] cb_0_8/io_i_4_in1[6]
+ cb_0_8/io_i_4_in1[7] cb_0_8/io_i_5_ci cb_0_8/io_i_5_in1[0] cb_0_8/io_i_5_in1[1]
+ cb_0_8/io_i_5_in1[2] cb_0_8/io_i_5_in1[3] cb_0_8/io_i_5_in1[4] cb_0_8/io_i_5_in1[5]
+ cb_0_8/io_i_5_in1[6] cb_0_8/io_i_5_in1[7] cb_0_8/io_i_6_ci cb_0_8/io_i_6_in1[0]
+ cb_0_8/io_i_6_in1[1] cb_0_8/io_i_6_in1[2] cb_0_8/io_i_6_in1[3] cb_0_8/io_i_6_in1[4]
+ cb_0_8/io_i_6_in1[5] cb_0_8/io_i_6_in1[6] cb_0_8/io_i_6_in1[7] cb_0_8/io_i_7_ci
+ cb_0_8/io_i_7_in1[0] cb_0_8/io_i_7_in1[1] cb_0_8/io_i_7_in1[2] cb_0_8/io_i_7_in1[3]
+ cb_0_8/io_i_7_in1[4] cb_0_8/io_i_7_in1[5] cb_0_8/io_i_7_in1[6] cb_0_8/io_i_7_in1[7]
+ cb_0_9/io_i_0_ci cb_0_9/io_i_0_in1[0] cb_0_9/io_i_0_in1[1] cb_0_9/io_i_0_in1[2]
+ cb_0_9/io_i_0_in1[3] cb_0_9/io_i_0_in1[4] cb_0_9/io_i_0_in1[5] cb_0_9/io_i_0_in1[6]
+ cb_0_9/io_i_0_in1[7] cb_0_9/io_i_1_ci cb_0_9/io_i_1_in1[0] cb_0_9/io_i_1_in1[1]
+ cb_0_9/io_i_1_in1[2] cb_0_9/io_i_1_in1[3] cb_0_9/io_i_1_in1[4] cb_0_9/io_i_1_in1[5]
+ cb_0_9/io_i_1_in1[6] cb_0_9/io_i_1_in1[7] cb_0_9/io_i_2_ci cb_0_9/io_i_2_in1[0]
+ cb_0_9/io_i_2_in1[1] cb_0_9/io_i_2_in1[2] cb_0_9/io_i_2_in1[3] cb_0_9/io_i_2_in1[4]
+ cb_0_9/io_i_2_in1[5] cb_0_9/io_i_2_in1[6] cb_0_9/io_i_2_in1[7] cb_0_9/io_i_3_ci
+ cb_0_9/io_i_3_in1[0] cb_0_9/io_i_3_in1[1] cb_0_9/io_i_3_in1[2] cb_0_9/io_i_3_in1[3]
+ cb_0_9/io_i_3_in1[4] cb_0_9/io_i_3_in1[5] cb_0_9/io_i_3_in1[6] cb_0_9/io_i_3_in1[7]
+ cb_0_9/io_i_4_ci cb_0_9/io_i_4_in1[0] cb_0_9/io_i_4_in1[1] cb_0_9/io_i_4_in1[2]
+ cb_0_9/io_i_4_in1[3] cb_0_9/io_i_4_in1[4] cb_0_9/io_i_4_in1[5] cb_0_9/io_i_4_in1[6]
+ cb_0_9/io_i_4_in1[7] cb_0_9/io_i_5_ci cb_0_9/io_i_5_in1[0] cb_0_9/io_i_5_in1[1]
+ cb_0_9/io_i_5_in1[2] cb_0_9/io_i_5_in1[3] cb_0_9/io_i_5_in1[4] cb_0_9/io_i_5_in1[5]
+ cb_0_9/io_i_5_in1[6] cb_0_9/io_i_5_in1[7] cb_0_9/io_i_6_ci cb_0_9/io_i_6_in1[0]
+ cb_0_9/io_i_6_in1[1] cb_0_9/io_i_6_in1[2] cb_0_9/io_i_6_in1[3] cb_0_9/io_i_6_in1[4]
+ cb_0_9/io_i_6_in1[5] cb_0_9/io_i_6_in1[6] cb_0_9/io_i_6_in1[7] cb_0_9/io_i_7_ci
+ cb_0_9/io_i_7_in1[0] cb_0_9/io_i_7_in1[1] cb_0_9/io_i_7_in1[2] cb_0_9/io_i_7_in1[3]
+ cb_0_9/io_i_7_in1[4] cb_0_9/io_i_7_in1[5] cb_0_9/io_i_7_in1[6] cb_0_9/io_i_7_in1[7]
+ cb_0_8/io_vci cb_0_9/io_vci cb_0_8/io_vi cb_0_9/io_we_i cb_0_8/io_wo[0] cb_0_8/io_wo[10]
+ cb_0_8/io_wo[11] cb_0_8/io_wo[12] cb_0_8/io_wo[13] cb_0_8/io_wo[14] cb_0_8/io_wo[15]
+ cb_0_8/io_wo[16] cb_0_8/io_wo[17] cb_0_8/io_wo[18] cb_0_8/io_wo[19] cb_0_8/io_wo[1]
+ cb_0_8/io_wo[20] cb_0_8/io_wo[21] cb_0_8/io_wo[22] cb_0_8/io_wo[23] cb_0_8/io_wo[24]
+ cb_0_8/io_wo[25] cb_0_8/io_wo[26] cb_0_8/io_wo[27] cb_0_8/io_wo[28] cb_0_8/io_wo[29]
+ cb_0_8/io_wo[2] cb_0_8/io_wo[30] cb_0_8/io_wo[31] cb_0_8/io_wo[32] cb_0_8/io_wo[33]
+ cb_0_8/io_wo[34] cb_0_8/io_wo[35] cb_0_8/io_wo[36] cb_0_8/io_wo[37] cb_0_8/io_wo[38]
+ cb_0_8/io_wo[39] cb_0_8/io_wo[3] cb_0_8/io_wo[40] cb_0_8/io_wo[41] cb_0_8/io_wo[42]
+ cb_0_8/io_wo[43] cb_0_8/io_wo[44] cb_0_8/io_wo[45] cb_0_8/io_wo[46] cb_0_8/io_wo[47]
+ cb_0_8/io_wo[48] cb_0_8/io_wo[49] cb_0_8/io_wo[4] cb_0_8/io_wo[50] cb_0_8/io_wo[51]
+ cb_0_8/io_wo[52] cb_0_8/io_wo[53] cb_0_8/io_wo[54] cb_0_8/io_wo[55] cb_0_8/io_wo[56]
+ cb_0_8/io_wo[57] cb_0_8/io_wo[58] cb_0_8/io_wo[59] cb_0_8/io_wo[5] cb_0_8/io_wo[60]
+ cb_0_8/io_wo[61] cb_0_8/io_wo[62] cb_0_8/io_wo[63] cb_0_8/io_wo[6] cb_0_8/io_wo[7]
+ cb_0_8/io_wo[8] cb_0_8/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_0_9 cb_0_9/io_adr_i[0] cb_0_9/io_adr_i[1] cb_0_9/io_cs_i cb_0_9/io_dat_i[0] cb_0_9/io_dat_i[10]
+ cb_0_9/io_dat_i[11] cb_0_9/io_dat_i[12] cb_0_9/io_dat_i[13] cb_0_9/io_dat_i[14]
+ cb_0_9/io_dat_i[15] cb_0_9/io_dat_i[1] cb_0_9/io_dat_i[2] cb_0_9/io_dat_i[3] cb_0_9/io_dat_i[4]
+ cb_0_9/io_dat_i[5] cb_0_9/io_dat_i[6] cb_0_9/io_dat_i[7] cb_0_9/io_dat_i[8] cb_0_9/io_dat_i[9]
+ cb_0_9/io_dat_o[0] cb_0_9/io_dat_o[10] cb_0_9/io_dat_o[11] cb_0_9/io_dat_o[12] cb_0_9/io_dat_o[13]
+ cb_0_9/io_dat_o[14] cb_0_9/io_dat_o[15] cb_0_9/io_dat_o[1] cb_0_9/io_dat_o[2] cb_0_9/io_dat_o[3]
+ cb_0_9/io_dat_o[4] cb_0_9/io_dat_o[5] cb_0_9/io_dat_o[6] cb_0_9/io_dat_o[7] cb_0_9/io_dat_o[8]
+ cb_0_9/io_dat_o[9] cb_0_9/io_eo[0] cb_0_9/io_eo[10] cb_0_9/io_eo[11] cb_0_9/io_eo[12]
+ cb_0_9/io_eo[13] cb_0_9/io_eo[14] cb_0_9/io_eo[15] cb_0_9/io_eo[16] cb_0_9/io_eo[17]
+ cb_0_9/io_eo[18] cb_0_9/io_eo[19] cb_0_9/io_eo[1] cb_0_9/io_eo[20] cb_0_9/io_eo[21]
+ cb_0_9/io_eo[22] cb_0_9/io_eo[23] cb_0_9/io_eo[24] cb_0_9/io_eo[25] cb_0_9/io_eo[26]
+ cb_0_9/io_eo[27] cb_0_9/io_eo[28] cb_0_9/io_eo[29] cb_0_9/io_eo[2] cb_0_9/io_eo[30]
+ cb_0_9/io_eo[31] cb_0_9/io_eo[32] cb_0_9/io_eo[33] cb_0_9/io_eo[34] cb_0_9/io_eo[35]
+ cb_0_9/io_eo[36] cb_0_9/io_eo[37] cb_0_9/io_eo[38] cb_0_9/io_eo[39] cb_0_9/io_eo[3]
+ cb_0_9/io_eo[40] cb_0_9/io_eo[41] cb_0_9/io_eo[42] cb_0_9/io_eo[43] cb_0_9/io_eo[44]
+ cb_0_9/io_eo[45] cb_0_9/io_eo[46] cb_0_9/io_eo[47] cb_0_9/io_eo[48] cb_0_9/io_eo[49]
+ cb_0_9/io_eo[4] cb_0_9/io_eo[50] cb_0_9/io_eo[51] cb_0_9/io_eo[52] cb_0_9/io_eo[53]
+ cb_0_9/io_eo[54] cb_0_9/io_eo[55] cb_0_9/io_eo[56] cb_0_9/io_eo[57] cb_0_9/io_eo[58]
+ cb_0_9/io_eo[59] cb_0_9/io_eo[5] cb_0_9/io_eo[60] cb_0_9/io_eo[61] cb_0_9/io_eo[62]
+ cb_0_9/io_eo[63] cb_0_9/io_eo[6] cb_0_9/io_eo[7] cb_0_9/io_eo[8] cb_0_9/io_eo[9]
+ cb_0_9/io_i_0_ci cb_0_9/io_i_0_in1[0] cb_0_9/io_i_0_in1[1] cb_0_9/io_i_0_in1[2]
+ cb_0_9/io_i_0_in1[3] cb_0_9/io_i_0_in1[4] cb_0_9/io_i_0_in1[5] cb_0_9/io_i_0_in1[6]
+ cb_0_9/io_i_0_in1[7] cb_0_9/io_i_1_ci cb_0_9/io_i_1_in1[0] cb_0_9/io_i_1_in1[1]
+ cb_0_9/io_i_1_in1[2] cb_0_9/io_i_1_in1[3] cb_0_9/io_i_1_in1[4] cb_0_9/io_i_1_in1[5]
+ cb_0_9/io_i_1_in1[6] cb_0_9/io_i_1_in1[7] cb_0_9/io_i_2_ci cb_0_9/io_i_2_in1[0]
+ cb_0_9/io_i_2_in1[1] cb_0_9/io_i_2_in1[2] cb_0_9/io_i_2_in1[3] cb_0_9/io_i_2_in1[4]
+ cb_0_9/io_i_2_in1[5] cb_0_9/io_i_2_in1[6] cb_0_9/io_i_2_in1[7] cb_0_9/io_i_3_ci
+ cb_0_9/io_i_3_in1[0] cb_0_9/io_i_3_in1[1] cb_0_9/io_i_3_in1[2] cb_0_9/io_i_3_in1[3]
+ cb_0_9/io_i_3_in1[4] cb_0_9/io_i_3_in1[5] cb_0_9/io_i_3_in1[6] cb_0_9/io_i_3_in1[7]
+ cb_0_9/io_i_4_ci cb_0_9/io_i_4_in1[0] cb_0_9/io_i_4_in1[1] cb_0_9/io_i_4_in1[2]
+ cb_0_9/io_i_4_in1[3] cb_0_9/io_i_4_in1[4] cb_0_9/io_i_4_in1[5] cb_0_9/io_i_4_in1[6]
+ cb_0_9/io_i_4_in1[7] cb_0_9/io_i_5_ci cb_0_9/io_i_5_in1[0] cb_0_9/io_i_5_in1[1]
+ cb_0_9/io_i_5_in1[2] cb_0_9/io_i_5_in1[3] cb_0_9/io_i_5_in1[4] cb_0_9/io_i_5_in1[5]
+ cb_0_9/io_i_5_in1[6] cb_0_9/io_i_5_in1[7] cb_0_9/io_i_6_ci cb_0_9/io_i_6_in1[0]
+ cb_0_9/io_i_6_in1[1] cb_0_9/io_i_6_in1[2] cb_0_9/io_i_6_in1[3] cb_0_9/io_i_6_in1[4]
+ cb_0_9/io_i_6_in1[5] cb_0_9/io_i_6_in1[6] cb_0_9/io_i_6_in1[7] cb_0_9/io_i_7_ci
+ cb_0_9/io_i_7_in1[0] cb_0_9/io_i_7_in1[1] cb_0_9/io_i_7_in1[2] cb_0_9/io_i_7_in1[3]
+ cb_0_9/io_i_7_in1[4] cb_0_9/io_i_7_in1[5] cb_0_9/io_i_7_in1[6] cb_0_9/io_i_7_in1[7]
+ cb_0_9/io_o_0_co cb_0_9/io_o_0_out[0] cb_0_9/io_o_0_out[1] cb_0_9/io_o_0_out[2]
+ cb_0_9/io_o_0_out[3] cb_0_9/io_o_0_out[4] cb_0_9/io_o_0_out[5] cb_0_9/io_o_0_out[6]
+ cb_0_9/io_o_0_out[7] cb_0_9/io_o_1_co cb_0_9/io_o_1_out[0] cb_0_9/io_o_1_out[1]
+ cb_0_9/io_o_1_out[2] cb_0_9/io_o_1_out[3] cb_0_9/io_o_1_out[4] cb_0_9/io_o_1_out[5]
+ cb_0_9/io_o_1_out[6] cb_0_9/io_o_1_out[7] cb_0_9/io_o_2_co cb_0_9/io_o_2_out[0]
+ cb_0_9/io_o_2_out[1] cb_0_9/io_o_2_out[2] cb_0_9/io_o_2_out[3] cb_0_9/io_o_2_out[4]
+ cb_0_9/io_o_2_out[5] cb_0_9/io_o_2_out[6] cb_0_9/io_o_2_out[7] cb_0_9/io_o_3_co
+ cb_0_9/io_o_3_out[0] cb_0_9/io_o_3_out[1] cb_0_9/io_o_3_out[2] cb_0_9/io_o_3_out[3]
+ cb_0_9/io_o_3_out[4] cb_0_9/io_o_3_out[5] cb_0_9/io_o_3_out[6] cb_0_9/io_o_3_out[7]
+ cb_0_9/io_o_4_co cb_0_9/io_o_4_out[0] cb_0_9/io_o_4_out[1] cb_0_9/io_o_4_out[2]
+ cb_0_9/io_o_4_out[3] cb_0_9/io_o_4_out[4] cb_0_9/io_o_4_out[5] cb_0_9/io_o_4_out[6]
+ cb_0_9/io_o_4_out[7] cb_0_9/io_o_5_co cb_0_9/io_o_5_out[0] cb_0_9/io_o_5_out[1]
+ cb_0_9/io_o_5_out[2] cb_0_9/io_o_5_out[3] cb_0_9/io_o_5_out[4] cb_0_9/io_o_5_out[5]
+ cb_0_9/io_o_5_out[6] cb_0_9/io_o_5_out[7] cb_0_9/io_o_6_co cb_0_9/io_o_6_out[0]
+ cb_0_9/io_o_6_out[1] cb_0_9/io_o_6_out[2] cb_0_9/io_o_6_out[3] cb_0_9/io_o_6_out[4]
+ cb_0_9/io_o_6_out[5] cb_0_9/io_o_6_out[6] cb_0_9/io_o_6_out[7] cb_0_9/io_o_7_co
+ cb_0_9/io_o_7_out[0] cb_0_9/io_o_7_out[1] cb_0_9/io_o_7_out[2] cb_0_9/io_o_7_out[3]
+ cb_0_9/io_o_7_out[4] cb_0_9/io_o_7_out[5] cb_0_9/io_o_7_out[6] cb_0_9/io_o_7_out[7]
+ cb_0_9/io_vci cb_0_9/io_vco cb_0_9/io_vi cb_0_9/io_we_i cb_0_9/io_wo[0] cb_0_9/io_wo[10]
+ cb_0_9/io_wo[11] cb_0_9/io_wo[12] cb_0_9/io_wo[13] cb_0_9/io_wo[14] cb_0_9/io_wo[15]
+ cb_0_9/io_wo[16] cb_0_9/io_wo[17] cb_0_9/io_wo[18] cb_0_9/io_wo[19] cb_0_9/io_wo[1]
+ cb_0_9/io_wo[20] cb_0_9/io_wo[21] cb_0_9/io_wo[22] cb_0_9/io_wo[23] cb_0_9/io_wo[24]
+ cb_0_9/io_wo[25] cb_0_9/io_wo[26] cb_0_9/io_wo[27] cb_0_9/io_wo[28] cb_0_9/io_wo[29]
+ cb_0_9/io_wo[2] cb_0_9/io_wo[30] cb_0_9/io_wo[31] cb_0_9/io_wo[32] cb_0_9/io_wo[33]
+ cb_0_9/io_wo[34] cb_0_9/io_wo[35] cb_0_9/io_wo[36] cb_0_9/io_wo[37] cb_0_9/io_wo[38]
+ cb_0_9/io_wo[39] cb_0_9/io_wo[3] cb_0_9/io_wo[40] cb_0_9/io_wo[41] cb_0_9/io_wo[42]
+ cb_0_9/io_wo[43] cb_0_9/io_wo[44] cb_0_9/io_wo[45] cb_0_9/io_wo[46] cb_0_9/io_wo[47]
+ cb_0_9/io_wo[48] cb_0_9/io_wo[49] cb_0_9/io_wo[4] cb_0_9/io_wo[50] cb_0_9/io_wo[51]
+ cb_0_9/io_wo[52] cb_0_9/io_wo[53] cb_0_9/io_wo[54] cb_0_9/io_wo[55] cb_0_9/io_wo[56]
+ cb_0_9/io_wo[57] cb_0_9/io_wo[58] cb_0_9/io_wo[59] cb_0_9/io_wo[5] cb_0_9/io_wo[60]
+ cb_0_9/io_wo[61] cb_0_9/io_wo[62] cb_0_9/io_wo[63] cb_0_9/io_wo[6] cb_0_9/io_wo[7]
+ cb_0_9/io_wo[8] cb_0_9/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_7_2 cb_7_9/io_adr_i[0] cb_7_9/io_adr_i[1] cb_7_2/io_cs_i cb_7_9/io_dat_i[0] cb_7_9/io_dat_i[10]
+ cb_7_9/io_dat_i[11] cb_7_9/io_dat_i[12] cb_7_9/io_dat_i[13] cb_7_9/io_dat_i[14]
+ cb_7_9/io_dat_i[15] cb_7_9/io_dat_i[1] cb_7_9/io_dat_i[2] cb_7_9/io_dat_i[3] cb_7_9/io_dat_i[4]
+ cb_7_9/io_dat_i[5] cb_7_9/io_dat_i[6] cb_7_9/io_dat_i[7] cb_7_9/io_dat_i[8] cb_7_9/io_dat_i[9]
+ cb_7_2/io_dat_o[0] cb_7_2/io_dat_o[10] cb_7_2/io_dat_o[11] cb_7_2/io_dat_o[12] cb_7_2/io_dat_o[13]
+ cb_7_2/io_dat_o[14] cb_7_2/io_dat_o[15] cb_7_2/io_dat_o[1] cb_7_2/io_dat_o[2] cb_7_2/io_dat_o[3]
+ cb_7_2/io_dat_o[4] cb_7_2/io_dat_o[5] cb_7_2/io_dat_o[6] cb_7_2/io_dat_o[7] cb_7_2/io_dat_o[8]
+ cb_7_2/io_dat_o[9] cb_7_3/io_wo[0] cb_7_3/io_wo[10] cb_7_3/io_wo[11] cb_7_3/io_wo[12]
+ cb_7_3/io_wo[13] cb_7_3/io_wo[14] cb_7_3/io_wo[15] cb_7_3/io_wo[16] cb_7_3/io_wo[17]
+ cb_7_3/io_wo[18] cb_7_3/io_wo[19] cb_7_3/io_wo[1] cb_7_3/io_wo[20] cb_7_3/io_wo[21]
+ cb_7_3/io_wo[22] cb_7_3/io_wo[23] cb_7_3/io_wo[24] cb_7_3/io_wo[25] cb_7_3/io_wo[26]
+ cb_7_3/io_wo[27] cb_7_3/io_wo[28] cb_7_3/io_wo[29] cb_7_3/io_wo[2] cb_7_3/io_wo[30]
+ cb_7_3/io_wo[31] cb_7_3/io_wo[32] cb_7_3/io_wo[33] cb_7_3/io_wo[34] cb_7_3/io_wo[35]
+ cb_7_3/io_wo[36] cb_7_3/io_wo[37] cb_7_3/io_wo[38] cb_7_3/io_wo[39] cb_7_3/io_wo[3]
+ cb_7_3/io_wo[40] cb_7_3/io_wo[41] cb_7_3/io_wo[42] cb_7_3/io_wo[43] cb_7_3/io_wo[44]
+ cb_7_3/io_wo[45] cb_7_3/io_wo[46] cb_7_3/io_wo[47] cb_7_3/io_wo[48] cb_7_3/io_wo[49]
+ cb_7_3/io_wo[4] cb_7_3/io_wo[50] cb_7_3/io_wo[51] cb_7_3/io_wo[52] cb_7_3/io_wo[53]
+ cb_7_3/io_wo[54] cb_7_3/io_wo[55] cb_7_3/io_wo[56] cb_7_3/io_wo[57] cb_7_3/io_wo[58]
+ cb_7_3/io_wo[59] cb_7_3/io_wo[5] cb_7_3/io_wo[60] cb_7_3/io_wo[61] cb_7_3/io_wo[62]
+ cb_7_3/io_wo[63] cb_7_3/io_wo[6] cb_7_3/io_wo[7] cb_7_3/io_wo[8] cb_7_3/io_wo[9]
+ cb_7_2/io_i_0_ci cb_7_2/io_i_0_in1[0] cb_7_2/io_i_0_in1[1] cb_7_2/io_i_0_in1[2]
+ cb_7_2/io_i_0_in1[3] cb_7_2/io_i_0_in1[4] cb_7_2/io_i_0_in1[5] cb_7_2/io_i_0_in1[6]
+ cb_7_2/io_i_0_in1[7] cb_7_2/io_i_1_ci cb_7_2/io_i_1_in1[0] cb_7_2/io_i_1_in1[1]
+ cb_7_2/io_i_1_in1[2] cb_7_2/io_i_1_in1[3] cb_7_2/io_i_1_in1[4] cb_7_2/io_i_1_in1[5]
+ cb_7_2/io_i_1_in1[6] cb_7_2/io_i_1_in1[7] cb_7_2/io_i_2_ci cb_7_2/io_i_2_in1[0]
+ cb_7_2/io_i_2_in1[1] cb_7_2/io_i_2_in1[2] cb_7_2/io_i_2_in1[3] cb_7_2/io_i_2_in1[4]
+ cb_7_2/io_i_2_in1[5] cb_7_2/io_i_2_in1[6] cb_7_2/io_i_2_in1[7] cb_7_2/io_i_3_ci
+ cb_7_2/io_i_3_in1[0] cb_7_2/io_i_3_in1[1] cb_7_2/io_i_3_in1[2] cb_7_2/io_i_3_in1[3]
+ cb_7_2/io_i_3_in1[4] cb_7_2/io_i_3_in1[5] cb_7_2/io_i_3_in1[6] cb_7_2/io_i_3_in1[7]
+ cb_7_2/io_i_4_ci cb_7_2/io_i_4_in1[0] cb_7_2/io_i_4_in1[1] cb_7_2/io_i_4_in1[2]
+ cb_7_2/io_i_4_in1[3] cb_7_2/io_i_4_in1[4] cb_7_2/io_i_4_in1[5] cb_7_2/io_i_4_in1[6]
+ cb_7_2/io_i_4_in1[7] cb_7_2/io_i_5_ci cb_7_2/io_i_5_in1[0] cb_7_2/io_i_5_in1[1]
+ cb_7_2/io_i_5_in1[2] cb_7_2/io_i_5_in1[3] cb_7_2/io_i_5_in1[4] cb_7_2/io_i_5_in1[5]
+ cb_7_2/io_i_5_in1[6] cb_7_2/io_i_5_in1[7] cb_7_2/io_i_6_ci cb_7_2/io_i_6_in1[0]
+ cb_7_2/io_i_6_in1[1] cb_7_2/io_i_6_in1[2] cb_7_2/io_i_6_in1[3] cb_7_2/io_i_6_in1[4]
+ cb_7_2/io_i_6_in1[5] cb_7_2/io_i_6_in1[6] cb_7_2/io_i_6_in1[7] cb_7_2/io_i_7_ci
+ cb_7_2/io_i_7_in1[0] cb_7_2/io_i_7_in1[1] cb_7_2/io_i_7_in1[2] cb_7_2/io_i_7_in1[3]
+ cb_7_2/io_i_7_in1[4] cb_7_2/io_i_7_in1[5] cb_7_2/io_i_7_in1[6] cb_7_2/io_i_7_in1[7]
+ cb_7_3/io_i_0_ci cb_7_3/io_i_0_in1[0] cb_7_3/io_i_0_in1[1] cb_7_3/io_i_0_in1[2]
+ cb_7_3/io_i_0_in1[3] cb_7_3/io_i_0_in1[4] cb_7_3/io_i_0_in1[5] cb_7_3/io_i_0_in1[6]
+ cb_7_3/io_i_0_in1[7] cb_7_3/io_i_1_ci cb_7_3/io_i_1_in1[0] cb_7_3/io_i_1_in1[1]
+ cb_7_3/io_i_1_in1[2] cb_7_3/io_i_1_in1[3] cb_7_3/io_i_1_in1[4] cb_7_3/io_i_1_in1[5]
+ cb_7_3/io_i_1_in1[6] cb_7_3/io_i_1_in1[7] cb_7_3/io_i_2_ci cb_7_3/io_i_2_in1[0]
+ cb_7_3/io_i_2_in1[1] cb_7_3/io_i_2_in1[2] cb_7_3/io_i_2_in1[3] cb_7_3/io_i_2_in1[4]
+ cb_7_3/io_i_2_in1[5] cb_7_3/io_i_2_in1[6] cb_7_3/io_i_2_in1[7] cb_7_3/io_i_3_ci
+ cb_7_3/io_i_3_in1[0] cb_7_3/io_i_3_in1[1] cb_7_3/io_i_3_in1[2] cb_7_3/io_i_3_in1[3]
+ cb_7_3/io_i_3_in1[4] cb_7_3/io_i_3_in1[5] cb_7_3/io_i_3_in1[6] cb_7_3/io_i_3_in1[7]
+ cb_7_3/io_i_4_ci cb_7_3/io_i_4_in1[0] cb_7_3/io_i_4_in1[1] cb_7_3/io_i_4_in1[2]
+ cb_7_3/io_i_4_in1[3] cb_7_3/io_i_4_in1[4] cb_7_3/io_i_4_in1[5] cb_7_3/io_i_4_in1[6]
+ cb_7_3/io_i_4_in1[7] cb_7_3/io_i_5_ci cb_7_3/io_i_5_in1[0] cb_7_3/io_i_5_in1[1]
+ cb_7_3/io_i_5_in1[2] cb_7_3/io_i_5_in1[3] cb_7_3/io_i_5_in1[4] cb_7_3/io_i_5_in1[5]
+ cb_7_3/io_i_5_in1[6] cb_7_3/io_i_5_in1[7] cb_7_3/io_i_6_ci cb_7_3/io_i_6_in1[0]
+ cb_7_3/io_i_6_in1[1] cb_7_3/io_i_6_in1[2] cb_7_3/io_i_6_in1[3] cb_7_3/io_i_6_in1[4]
+ cb_7_3/io_i_6_in1[5] cb_7_3/io_i_6_in1[6] cb_7_3/io_i_6_in1[7] cb_7_3/io_i_7_ci
+ cb_7_3/io_i_7_in1[0] cb_7_3/io_i_7_in1[1] cb_7_3/io_i_7_in1[2] cb_7_3/io_i_7_in1[3]
+ cb_7_3/io_i_7_in1[4] cb_7_3/io_i_7_in1[5] cb_7_3/io_i_7_in1[6] cb_7_3/io_i_7_in1[7]
+ cb_7_2/io_vci cb_7_3/io_vci cb_7_2/io_vi cb_7_9/io_we_i cb_7_2/io_wo[0] cb_7_2/io_wo[10]
+ cb_7_2/io_wo[11] cb_7_2/io_wo[12] cb_7_2/io_wo[13] cb_7_2/io_wo[14] cb_7_2/io_wo[15]
+ cb_7_2/io_wo[16] cb_7_2/io_wo[17] cb_7_2/io_wo[18] cb_7_2/io_wo[19] cb_7_2/io_wo[1]
+ cb_7_2/io_wo[20] cb_7_2/io_wo[21] cb_7_2/io_wo[22] cb_7_2/io_wo[23] cb_7_2/io_wo[24]
+ cb_7_2/io_wo[25] cb_7_2/io_wo[26] cb_7_2/io_wo[27] cb_7_2/io_wo[28] cb_7_2/io_wo[29]
+ cb_7_2/io_wo[2] cb_7_2/io_wo[30] cb_7_2/io_wo[31] cb_7_2/io_wo[32] cb_7_2/io_wo[33]
+ cb_7_2/io_wo[34] cb_7_2/io_wo[35] cb_7_2/io_wo[36] cb_7_2/io_wo[37] cb_7_2/io_wo[38]
+ cb_7_2/io_wo[39] cb_7_2/io_wo[3] cb_7_2/io_wo[40] cb_7_2/io_wo[41] cb_7_2/io_wo[42]
+ cb_7_2/io_wo[43] cb_7_2/io_wo[44] cb_7_2/io_wo[45] cb_7_2/io_wo[46] cb_7_2/io_wo[47]
+ cb_7_2/io_wo[48] cb_7_2/io_wo[49] cb_7_2/io_wo[4] cb_7_2/io_wo[50] cb_7_2/io_wo[51]
+ cb_7_2/io_wo[52] cb_7_2/io_wo[53] cb_7_2/io_wo[54] cb_7_2/io_wo[55] cb_7_2/io_wo[56]
+ cb_7_2/io_wo[57] cb_7_2/io_wo[58] cb_7_2/io_wo[59] cb_7_2/io_wo[5] cb_7_2/io_wo[60]
+ cb_7_2/io_wo[61] cb_7_2/io_wo[62] cb_7_2/io_wo[63] cb_7_2/io_wo[6] cb_7_2/io_wo[7]
+ cb_7_2/io_wo[8] cb_7_2/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_7_3 cb_7_9/io_adr_i[0] cb_7_9/io_adr_i[1] cb_7_3/io_cs_i cb_7_9/io_dat_i[0] cb_7_9/io_dat_i[10]
+ cb_7_9/io_dat_i[11] cb_7_9/io_dat_i[12] cb_7_9/io_dat_i[13] cb_7_9/io_dat_i[14]
+ cb_7_9/io_dat_i[15] cb_7_9/io_dat_i[1] cb_7_9/io_dat_i[2] cb_7_9/io_dat_i[3] cb_7_9/io_dat_i[4]
+ cb_7_9/io_dat_i[5] cb_7_9/io_dat_i[6] cb_7_9/io_dat_i[7] cb_7_9/io_dat_i[8] cb_7_9/io_dat_i[9]
+ cb_7_3/io_dat_o[0] cb_7_3/io_dat_o[10] cb_7_3/io_dat_o[11] cb_7_3/io_dat_o[12] cb_7_3/io_dat_o[13]
+ cb_7_3/io_dat_o[14] cb_7_3/io_dat_o[15] cb_7_3/io_dat_o[1] cb_7_3/io_dat_o[2] cb_7_3/io_dat_o[3]
+ cb_7_3/io_dat_o[4] cb_7_3/io_dat_o[5] cb_7_3/io_dat_o[6] cb_7_3/io_dat_o[7] cb_7_3/io_dat_o[8]
+ cb_7_3/io_dat_o[9] cb_7_4/io_wo[0] cb_7_4/io_wo[10] cb_7_4/io_wo[11] cb_7_4/io_wo[12]
+ cb_7_4/io_wo[13] cb_7_4/io_wo[14] cb_7_4/io_wo[15] cb_7_4/io_wo[16] cb_7_4/io_wo[17]
+ cb_7_4/io_wo[18] cb_7_4/io_wo[19] cb_7_4/io_wo[1] cb_7_4/io_wo[20] cb_7_4/io_wo[21]
+ cb_7_4/io_wo[22] cb_7_4/io_wo[23] cb_7_4/io_wo[24] cb_7_4/io_wo[25] cb_7_4/io_wo[26]
+ cb_7_4/io_wo[27] cb_7_4/io_wo[28] cb_7_4/io_wo[29] cb_7_4/io_wo[2] cb_7_4/io_wo[30]
+ cb_7_4/io_wo[31] cb_7_4/io_wo[32] cb_7_4/io_wo[33] cb_7_4/io_wo[34] cb_7_4/io_wo[35]
+ cb_7_4/io_wo[36] cb_7_4/io_wo[37] cb_7_4/io_wo[38] cb_7_4/io_wo[39] cb_7_4/io_wo[3]
+ cb_7_4/io_wo[40] cb_7_4/io_wo[41] cb_7_4/io_wo[42] cb_7_4/io_wo[43] cb_7_4/io_wo[44]
+ cb_7_4/io_wo[45] cb_7_4/io_wo[46] cb_7_4/io_wo[47] cb_7_4/io_wo[48] cb_7_4/io_wo[49]
+ cb_7_4/io_wo[4] cb_7_4/io_wo[50] cb_7_4/io_wo[51] cb_7_4/io_wo[52] cb_7_4/io_wo[53]
+ cb_7_4/io_wo[54] cb_7_4/io_wo[55] cb_7_4/io_wo[56] cb_7_4/io_wo[57] cb_7_4/io_wo[58]
+ cb_7_4/io_wo[59] cb_7_4/io_wo[5] cb_7_4/io_wo[60] cb_7_4/io_wo[61] cb_7_4/io_wo[62]
+ cb_7_4/io_wo[63] cb_7_4/io_wo[6] cb_7_4/io_wo[7] cb_7_4/io_wo[8] cb_7_4/io_wo[9]
+ cb_7_3/io_i_0_ci cb_7_3/io_i_0_in1[0] cb_7_3/io_i_0_in1[1] cb_7_3/io_i_0_in1[2]
+ cb_7_3/io_i_0_in1[3] cb_7_3/io_i_0_in1[4] cb_7_3/io_i_0_in1[5] cb_7_3/io_i_0_in1[6]
+ cb_7_3/io_i_0_in1[7] cb_7_3/io_i_1_ci cb_7_3/io_i_1_in1[0] cb_7_3/io_i_1_in1[1]
+ cb_7_3/io_i_1_in1[2] cb_7_3/io_i_1_in1[3] cb_7_3/io_i_1_in1[4] cb_7_3/io_i_1_in1[5]
+ cb_7_3/io_i_1_in1[6] cb_7_3/io_i_1_in1[7] cb_7_3/io_i_2_ci cb_7_3/io_i_2_in1[0]
+ cb_7_3/io_i_2_in1[1] cb_7_3/io_i_2_in1[2] cb_7_3/io_i_2_in1[3] cb_7_3/io_i_2_in1[4]
+ cb_7_3/io_i_2_in1[5] cb_7_3/io_i_2_in1[6] cb_7_3/io_i_2_in1[7] cb_7_3/io_i_3_ci
+ cb_7_3/io_i_3_in1[0] cb_7_3/io_i_3_in1[1] cb_7_3/io_i_3_in1[2] cb_7_3/io_i_3_in1[3]
+ cb_7_3/io_i_3_in1[4] cb_7_3/io_i_3_in1[5] cb_7_3/io_i_3_in1[6] cb_7_3/io_i_3_in1[7]
+ cb_7_3/io_i_4_ci cb_7_3/io_i_4_in1[0] cb_7_3/io_i_4_in1[1] cb_7_3/io_i_4_in1[2]
+ cb_7_3/io_i_4_in1[3] cb_7_3/io_i_4_in1[4] cb_7_3/io_i_4_in1[5] cb_7_3/io_i_4_in1[6]
+ cb_7_3/io_i_4_in1[7] cb_7_3/io_i_5_ci cb_7_3/io_i_5_in1[0] cb_7_3/io_i_5_in1[1]
+ cb_7_3/io_i_5_in1[2] cb_7_3/io_i_5_in1[3] cb_7_3/io_i_5_in1[4] cb_7_3/io_i_5_in1[5]
+ cb_7_3/io_i_5_in1[6] cb_7_3/io_i_5_in1[7] cb_7_3/io_i_6_ci cb_7_3/io_i_6_in1[0]
+ cb_7_3/io_i_6_in1[1] cb_7_3/io_i_6_in1[2] cb_7_3/io_i_6_in1[3] cb_7_3/io_i_6_in1[4]
+ cb_7_3/io_i_6_in1[5] cb_7_3/io_i_6_in1[6] cb_7_3/io_i_6_in1[7] cb_7_3/io_i_7_ci
+ cb_7_3/io_i_7_in1[0] cb_7_3/io_i_7_in1[1] cb_7_3/io_i_7_in1[2] cb_7_3/io_i_7_in1[3]
+ cb_7_3/io_i_7_in1[4] cb_7_3/io_i_7_in1[5] cb_7_3/io_i_7_in1[6] cb_7_3/io_i_7_in1[7]
+ cb_7_4/io_i_0_ci cb_7_4/io_i_0_in1[0] cb_7_4/io_i_0_in1[1] cb_7_4/io_i_0_in1[2]
+ cb_7_4/io_i_0_in1[3] cb_7_4/io_i_0_in1[4] cb_7_4/io_i_0_in1[5] cb_7_4/io_i_0_in1[6]
+ cb_7_4/io_i_0_in1[7] cb_7_4/io_i_1_ci cb_7_4/io_i_1_in1[0] cb_7_4/io_i_1_in1[1]
+ cb_7_4/io_i_1_in1[2] cb_7_4/io_i_1_in1[3] cb_7_4/io_i_1_in1[4] cb_7_4/io_i_1_in1[5]
+ cb_7_4/io_i_1_in1[6] cb_7_4/io_i_1_in1[7] cb_7_4/io_i_2_ci cb_7_4/io_i_2_in1[0]
+ cb_7_4/io_i_2_in1[1] cb_7_4/io_i_2_in1[2] cb_7_4/io_i_2_in1[3] cb_7_4/io_i_2_in1[4]
+ cb_7_4/io_i_2_in1[5] cb_7_4/io_i_2_in1[6] cb_7_4/io_i_2_in1[7] cb_7_4/io_i_3_ci
+ cb_7_4/io_i_3_in1[0] cb_7_4/io_i_3_in1[1] cb_7_4/io_i_3_in1[2] cb_7_4/io_i_3_in1[3]
+ cb_7_4/io_i_3_in1[4] cb_7_4/io_i_3_in1[5] cb_7_4/io_i_3_in1[6] cb_7_4/io_i_3_in1[7]
+ cb_7_4/io_i_4_ci cb_7_4/io_i_4_in1[0] cb_7_4/io_i_4_in1[1] cb_7_4/io_i_4_in1[2]
+ cb_7_4/io_i_4_in1[3] cb_7_4/io_i_4_in1[4] cb_7_4/io_i_4_in1[5] cb_7_4/io_i_4_in1[6]
+ cb_7_4/io_i_4_in1[7] cb_7_4/io_i_5_ci cb_7_4/io_i_5_in1[0] cb_7_4/io_i_5_in1[1]
+ cb_7_4/io_i_5_in1[2] cb_7_4/io_i_5_in1[3] cb_7_4/io_i_5_in1[4] cb_7_4/io_i_5_in1[5]
+ cb_7_4/io_i_5_in1[6] cb_7_4/io_i_5_in1[7] cb_7_4/io_i_6_ci cb_7_4/io_i_6_in1[0]
+ cb_7_4/io_i_6_in1[1] cb_7_4/io_i_6_in1[2] cb_7_4/io_i_6_in1[3] cb_7_4/io_i_6_in1[4]
+ cb_7_4/io_i_6_in1[5] cb_7_4/io_i_6_in1[6] cb_7_4/io_i_6_in1[7] cb_7_4/io_i_7_ci
+ cb_7_4/io_i_7_in1[0] cb_7_4/io_i_7_in1[1] cb_7_4/io_i_7_in1[2] cb_7_4/io_i_7_in1[3]
+ cb_7_4/io_i_7_in1[4] cb_7_4/io_i_7_in1[5] cb_7_4/io_i_7_in1[6] cb_7_4/io_i_7_in1[7]
+ cb_7_3/io_vci cb_7_4/io_vci cb_7_3/io_vi cb_7_9/io_we_i cb_7_3/io_wo[0] cb_7_3/io_wo[10]
+ cb_7_3/io_wo[11] cb_7_3/io_wo[12] cb_7_3/io_wo[13] cb_7_3/io_wo[14] cb_7_3/io_wo[15]
+ cb_7_3/io_wo[16] cb_7_3/io_wo[17] cb_7_3/io_wo[18] cb_7_3/io_wo[19] cb_7_3/io_wo[1]
+ cb_7_3/io_wo[20] cb_7_3/io_wo[21] cb_7_3/io_wo[22] cb_7_3/io_wo[23] cb_7_3/io_wo[24]
+ cb_7_3/io_wo[25] cb_7_3/io_wo[26] cb_7_3/io_wo[27] cb_7_3/io_wo[28] cb_7_3/io_wo[29]
+ cb_7_3/io_wo[2] cb_7_3/io_wo[30] cb_7_3/io_wo[31] cb_7_3/io_wo[32] cb_7_3/io_wo[33]
+ cb_7_3/io_wo[34] cb_7_3/io_wo[35] cb_7_3/io_wo[36] cb_7_3/io_wo[37] cb_7_3/io_wo[38]
+ cb_7_3/io_wo[39] cb_7_3/io_wo[3] cb_7_3/io_wo[40] cb_7_3/io_wo[41] cb_7_3/io_wo[42]
+ cb_7_3/io_wo[43] cb_7_3/io_wo[44] cb_7_3/io_wo[45] cb_7_3/io_wo[46] cb_7_3/io_wo[47]
+ cb_7_3/io_wo[48] cb_7_3/io_wo[49] cb_7_3/io_wo[4] cb_7_3/io_wo[50] cb_7_3/io_wo[51]
+ cb_7_3/io_wo[52] cb_7_3/io_wo[53] cb_7_3/io_wo[54] cb_7_3/io_wo[55] cb_7_3/io_wo[56]
+ cb_7_3/io_wo[57] cb_7_3/io_wo[58] cb_7_3/io_wo[59] cb_7_3/io_wo[5] cb_7_3/io_wo[60]
+ cb_7_3/io_wo[61] cb_7_3/io_wo[62] cb_7_3/io_wo[63] cb_7_3/io_wo[6] cb_7_3/io_wo[7]
+ cb_7_3/io_wo[8] cb_7_3/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_5_0 cb_5_9/io_adr_i[0] cb_5_9/io_adr_i[1] cb_5_0/io_cs_i cb_5_9/io_dat_i[0] cb_5_9/io_dat_i[10]
+ cb_5_9/io_dat_i[11] cb_5_9/io_dat_i[12] cb_5_9/io_dat_i[13] cb_5_9/io_dat_i[14]
+ cb_5_9/io_dat_i[15] cb_5_9/io_dat_i[1] cb_5_9/io_dat_i[2] cb_5_9/io_dat_i[3] cb_5_9/io_dat_i[4]
+ cb_5_9/io_dat_i[5] cb_5_9/io_dat_i[6] cb_5_9/io_dat_i[7] cb_5_9/io_dat_i[8] cb_5_9/io_dat_i[9]
+ cb_5_0/io_dat_o[0] cb_5_0/io_dat_o[10] cb_5_0/io_dat_o[11] cb_5_0/io_dat_o[12] cb_5_0/io_dat_o[13]
+ cb_5_0/io_dat_o[14] cb_5_0/io_dat_o[15] cb_5_0/io_dat_o[1] cb_5_0/io_dat_o[2] cb_5_0/io_dat_o[3]
+ cb_5_0/io_dat_o[4] cb_5_0/io_dat_o[5] cb_5_0/io_dat_o[6] cb_5_0/io_dat_o[7] cb_5_0/io_dat_o[8]
+ cb_5_0/io_dat_o[9] cb_5_1/io_wo[0] cb_5_1/io_wo[10] cb_5_1/io_wo[11] cb_5_1/io_wo[12]
+ cb_5_1/io_wo[13] cb_5_1/io_wo[14] cb_5_1/io_wo[15] cb_5_1/io_wo[16] cb_5_1/io_wo[17]
+ cb_5_1/io_wo[18] cb_5_1/io_wo[19] cb_5_1/io_wo[1] cb_5_1/io_wo[20] cb_5_1/io_wo[21]
+ cb_5_1/io_wo[22] cb_5_1/io_wo[23] cb_5_1/io_wo[24] cb_5_1/io_wo[25] cb_5_1/io_wo[26]
+ cb_5_1/io_wo[27] cb_5_1/io_wo[28] cb_5_1/io_wo[29] cb_5_1/io_wo[2] cb_5_1/io_wo[30]
+ cb_5_1/io_wo[31] cb_5_1/io_wo[32] cb_5_1/io_wo[33] cb_5_1/io_wo[34] cb_5_1/io_wo[35]
+ cb_5_1/io_wo[36] cb_5_1/io_wo[37] cb_5_1/io_wo[38] cb_5_1/io_wo[39] cb_5_1/io_wo[3]
+ cb_5_1/io_wo[40] cb_5_1/io_wo[41] cb_5_1/io_wo[42] cb_5_1/io_wo[43] cb_5_1/io_wo[44]
+ cb_5_1/io_wo[45] cb_5_1/io_wo[46] cb_5_1/io_wo[47] cb_5_1/io_wo[48] cb_5_1/io_wo[49]
+ cb_5_1/io_wo[4] cb_5_1/io_wo[50] cb_5_1/io_wo[51] cb_5_1/io_wo[52] cb_5_1/io_wo[53]
+ cb_5_1/io_wo[54] cb_5_1/io_wo[55] cb_5_1/io_wo[56] cb_5_1/io_wo[57] cb_5_1/io_wo[58]
+ cb_5_1/io_wo[59] cb_5_1/io_wo[5] cb_5_1/io_wo[60] cb_5_1/io_wo[61] cb_5_1/io_wo[62]
+ cb_5_1/io_wo[63] cb_5_1/io_wo[6] cb_5_1/io_wo[7] cb_5_1/io_wo[8] cb_5_1/io_wo[9]
+ ccon_5/io_dsi_o cb_5_0/io_i_0_in1[0] cb_5_0/io_i_0_in1[1] cb_5_0/io_i_0_in1[2] cb_5_0/io_i_0_in1[3]
+ cb_5_0/io_i_0_in1[4] cb_5_0/io_i_0_in1[5] cb_5_0/io_i_0_in1[6] cb_5_0/io_i_0_in1[7]
+ cb_5_0/io_i_1_ci cb_5_0/io_i_1_in1[0] cb_5_0/io_i_1_in1[1] cb_5_0/io_i_1_in1[2]
+ cb_5_0/io_i_1_in1[3] cb_5_0/io_i_1_in1[4] cb_5_0/io_i_1_in1[5] cb_5_0/io_i_1_in1[6]
+ cb_5_0/io_i_1_in1[7] cb_5_0/io_i_2_ci cb_5_0/io_i_2_in1[0] cb_5_0/io_i_2_in1[1]
+ cb_5_0/io_i_2_in1[2] cb_5_0/io_i_2_in1[3] cb_5_0/io_i_2_in1[4] cb_5_0/io_i_2_in1[5]
+ cb_5_0/io_i_2_in1[6] cb_5_0/io_i_2_in1[7] cb_5_0/io_i_3_ci cb_5_0/io_i_3_in1[0]
+ cb_5_0/io_i_3_in1[1] cb_5_0/io_i_3_in1[2] cb_5_0/io_i_3_in1[3] cb_5_0/io_i_3_in1[4]
+ cb_5_0/io_i_3_in1[5] cb_5_0/io_i_3_in1[6] cb_5_0/io_i_3_in1[7] cb_5_0/io_i_4_ci
+ cb_5_0/io_i_4_in1[0] cb_5_0/io_i_4_in1[1] cb_5_0/io_i_4_in1[2] cb_5_0/io_i_4_in1[3]
+ cb_5_0/io_i_4_in1[4] cb_5_0/io_i_4_in1[5] cb_5_0/io_i_4_in1[6] cb_5_0/io_i_4_in1[7]
+ cb_5_0/io_i_5_ci cb_5_0/io_i_5_in1[0] cb_5_0/io_i_5_in1[1] cb_5_0/io_i_5_in1[2]
+ cb_5_0/io_i_5_in1[3] cb_5_0/io_i_5_in1[4] cb_5_0/io_i_5_in1[5] cb_5_0/io_i_5_in1[6]
+ cb_5_0/io_i_5_in1[7] cb_5_0/io_i_6_ci cb_5_0/io_i_6_in1[0] cb_5_0/io_i_6_in1[1]
+ cb_5_0/io_i_6_in1[2] cb_5_0/io_i_6_in1[3] cb_5_0/io_i_6_in1[4] cb_5_0/io_i_6_in1[5]
+ cb_5_0/io_i_6_in1[6] cb_5_0/io_i_6_in1[7] cb_5_0/io_i_7_ci cb_5_0/io_i_7_in1[0]
+ cb_5_0/io_i_7_in1[1] cb_5_0/io_i_7_in1[2] cb_5_0/io_i_7_in1[3] cb_5_0/io_i_7_in1[4]
+ cb_5_0/io_i_7_in1[5] cb_5_0/io_i_7_in1[6] cb_5_0/io_i_7_in1[7] cb_5_1/io_i_0_ci
+ cb_5_1/io_i_0_in1[0] cb_5_1/io_i_0_in1[1] cb_5_1/io_i_0_in1[2] cb_5_1/io_i_0_in1[3]
+ cb_5_1/io_i_0_in1[4] cb_5_1/io_i_0_in1[5] cb_5_1/io_i_0_in1[6] cb_5_1/io_i_0_in1[7]
+ cb_5_1/io_i_1_ci cb_5_1/io_i_1_in1[0] cb_5_1/io_i_1_in1[1] cb_5_1/io_i_1_in1[2]
+ cb_5_1/io_i_1_in1[3] cb_5_1/io_i_1_in1[4] cb_5_1/io_i_1_in1[5] cb_5_1/io_i_1_in1[6]
+ cb_5_1/io_i_1_in1[7] cb_5_1/io_i_2_ci cb_5_1/io_i_2_in1[0] cb_5_1/io_i_2_in1[1]
+ cb_5_1/io_i_2_in1[2] cb_5_1/io_i_2_in1[3] cb_5_1/io_i_2_in1[4] cb_5_1/io_i_2_in1[5]
+ cb_5_1/io_i_2_in1[6] cb_5_1/io_i_2_in1[7] cb_5_1/io_i_3_ci cb_5_1/io_i_3_in1[0]
+ cb_5_1/io_i_3_in1[1] cb_5_1/io_i_3_in1[2] cb_5_1/io_i_3_in1[3] cb_5_1/io_i_3_in1[4]
+ cb_5_1/io_i_3_in1[5] cb_5_1/io_i_3_in1[6] cb_5_1/io_i_3_in1[7] cb_5_1/io_i_4_ci
+ cb_5_1/io_i_4_in1[0] cb_5_1/io_i_4_in1[1] cb_5_1/io_i_4_in1[2] cb_5_1/io_i_4_in1[3]
+ cb_5_1/io_i_4_in1[4] cb_5_1/io_i_4_in1[5] cb_5_1/io_i_4_in1[6] cb_5_1/io_i_4_in1[7]
+ cb_5_1/io_i_5_ci cb_5_1/io_i_5_in1[0] cb_5_1/io_i_5_in1[1] cb_5_1/io_i_5_in1[2]
+ cb_5_1/io_i_5_in1[3] cb_5_1/io_i_5_in1[4] cb_5_1/io_i_5_in1[5] cb_5_1/io_i_5_in1[6]
+ cb_5_1/io_i_5_in1[7] cb_5_1/io_i_6_ci cb_5_1/io_i_6_in1[0] cb_5_1/io_i_6_in1[1]
+ cb_5_1/io_i_6_in1[2] cb_5_1/io_i_6_in1[3] cb_5_1/io_i_6_in1[4] cb_5_1/io_i_6_in1[5]
+ cb_5_1/io_i_6_in1[6] cb_5_1/io_i_6_in1[7] cb_5_1/io_i_7_ci cb_5_1/io_i_7_in1[0]
+ cb_5_1/io_i_7_in1[1] cb_5_1/io_i_7_in1[2] cb_5_1/io_i_7_in1[3] cb_5_1/io_i_7_in1[4]
+ cb_5_1/io_i_7_in1[5] cb_5_1/io_i_7_in1[6] cb_5_1/io_i_7_in1[7] cb_5_0/io_vci cb_5_1/io_vci
+ cb_5_0/io_vi cb_5_9/io_we_i cb_5_0/io_wo[0] cb_5_0/io_wo[10] cb_5_0/io_wo[11] cb_5_0/io_wo[12]
+ cb_5_0/io_wo[13] cb_5_0/io_wo[14] cb_5_0/io_wo[15] cb_5_0/io_wo[16] cb_5_0/io_wo[17]
+ cb_5_0/io_wo[18] cb_5_0/io_wo[19] cb_5_0/io_wo[1] cb_5_0/io_wo[20] cb_5_0/io_wo[21]
+ cb_5_0/io_wo[22] cb_5_0/io_wo[23] cb_5_0/io_wo[24] cb_5_0/io_wo[25] cb_5_0/io_wo[26]
+ cb_5_0/io_wo[27] cb_5_0/io_wo[28] cb_5_0/io_wo[29] cb_5_0/io_wo[2] cb_5_0/io_wo[30]
+ cb_5_0/io_wo[31] cb_5_0/io_wo[32] cb_5_0/io_wo[33] cb_5_0/io_wo[34] cb_5_0/io_wo[35]
+ cb_5_0/io_wo[36] cb_5_0/io_wo[37] cb_5_0/io_wo[38] cb_5_0/io_wo[39] cb_5_0/io_wo[3]
+ cb_5_0/io_wo[40] cb_5_0/io_wo[41] cb_5_0/io_wo[42] cb_5_0/io_wo[43] cb_5_0/io_wo[44]
+ cb_5_0/io_wo[45] cb_5_0/io_wo[46] cb_5_0/io_wo[47] cb_5_0/io_wo[48] cb_5_0/io_wo[49]
+ cb_5_0/io_wo[4] cb_5_0/io_wo[50] cb_5_0/io_wo[51] cb_5_0/io_wo[52] cb_5_0/io_wo[53]
+ cb_5_0/io_wo[54] cb_5_0/io_wo[55] cb_5_0/io_wo[56] cb_5_0/io_wo[57] cb_5_0/io_wo[58]
+ cb_5_0/io_wo[59] cb_5_0/io_wo[5] cb_5_0/io_wo[60] cb_5_0/io_wo[61] cb_5_0/io_wo[62]
+ cb_5_0/io_wo[63] cb_5_0/io_wo[6] cb_5_0/io_wo[7] cb_5_0/io_wo[8] cb_5_0/io_wo[9]
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcordic cordic/ao_reg[0] cordic/ao_reg[10] cordic/ao_reg[11] cordic/ao_reg[12] cordic/ao_reg[13]
+ cordic/ao_reg[14] cordic/ao_reg[15] cordic/ao_reg[16] cordic/ao_reg[17] cordic/ao_reg[18]
+ cordic/ao_reg[19] cordic/ao_reg[1] cordic/ao_reg[20] cordic/ao_reg[21] cordic/ao_reg[22]
+ cordic/ao_reg[23] cordic/ao_reg[24] cordic/ao_reg[25] cordic/ao_reg[26] cordic/ao_reg[27]
+ cordic/ao_reg[28] cordic/ao_reg[29] cordic/ao_reg[2] cordic/ao_reg[30] cordic/ao_reg[31]
+ cordic/ao_reg[3] cordic/ao_reg[4] cordic/ao_reg[5] cordic/ao_reg[6] cordic/ao_reg[7]
+ cordic/ao_reg[8] cordic/ao_reg[9] cordic/asel cordic/bo_reg[0] cordic/bo_reg[10]
+ cordic/bo_reg[11] cordic/bo_reg[12] cordic/bo_reg[13] cordic/bo_reg[14] cordic/bo_reg[15]
+ cordic/bo_reg[16] cordic/bo_reg[17] cordic/bo_reg[18] cordic/bo_reg[19] cordic/bo_reg[1]
+ cordic/bo_reg[20] cordic/bo_reg[21] cordic/bo_reg[22] cordic/bo_reg[23] cordic/bo_reg[24]
+ cordic/bo_reg[25] cordic/bo_reg[26] cordic/bo_reg[27] cordic/bo_reg[28] cordic/bo_reg[29]
+ cordic/bo_reg[2] cordic/bo_reg[30] cordic/bo_reg[31] cordic/bo_reg[3] cordic/bo_reg[4]
+ cordic/bo_reg[5] cordic/bo_reg[6] cordic/bo_reg[7] cordic/bo_reg[8] cordic/bo_reg[9]
+ cordic/clk la_data_in[96] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[97] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[98] la_data_in[126] la_data_in[127] la_data_in[99] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_out[96] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[97] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[98] la_data_out[126] la_data_out[127]
+ la_data_out[99] la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103]
+ la_data_out[104] la_data_out[105] la_data_in[64] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[80] la_data_in[81] la_data_in[82]
+ la_data_in[83] la_data_in[65] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93]
+ la_data_in[66] la_data_in[94] la_data_in[95] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_out[64] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[65]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[66] la_data_out[94] la_data_out[95] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_in[32] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[50] la_data_in[51] la_data_in[33]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[60] la_data_in[61] la_data_in[34] la_data_in[62]
+ la_data_in[63] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[40] la_data_in[41] la_data_out[32] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[50] la_data_out[51] la_data_out[33] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[60] la_data_out[61] la_data_out[34] la_data_out[62]
+ la_data_out[63] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[40] la_data_out[41] la_data_in[0] la_data_in[10] la_data_in[11]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22]
+ la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28]
+ la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[3] la_data_in[4]
+ la_data_in[5] la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0]
+ la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[3] la_data_out[4] la_data_out[5]
+ la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9] vccd1 vssd1 sin3
Xcb_7_4 cb_7_9/io_adr_i[0] cb_7_9/io_adr_i[1] cb_7_4/io_cs_i cb_7_9/io_dat_i[0] cb_7_9/io_dat_i[10]
+ cb_7_9/io_dat_i[11] cb_7_9/io_dat_i[12] cb_7_9/io_dat_i[13] cb_7_9/io_dat_i[14]
+ cb_7_9/io_dat_i[15] cb_7_9/io_dat_i[1] cb_7_9/io_dat_i[2] cb_7_9/io_dat_i[3] cb_7_9/io_dat_i[4]
+ cb_7_9/io_dat_i[5] cb_7_9/io_dat_i[6] cb_7_9/io_dat_i[7] cb_7_9/io_dat_i[8] cb_7_9/io_dat_i[9]
+ cb_7_4/io_dat_o[0] cb_7_4/io_dat_o[10] cb_7_4/io_dat_o[11] cb_7_4/io_dat_o[12] cb_7_4/io_dat_o[13]
+ cb_7_4/io_dat_o[14] cb_7_4/io_dat_o[15] cb_7_4/io_dat_o[1] cb_7_4/io_dat_o[2] cb_7_4/io_dat_o[3]
+ cb_7_4/io_dat_o[4] cb_7_4/io_dat_o[5] cb_7_4/io_dat_o[6] cb_7_4/io_dat_o[7] cb_7_4/io_dat_o[8]
+ cb_7_4/io_dat_o[9] cb_7_5/io_wo[0] cb_7_5/io_wo[10] cb_7_5/io_wo[11] cb_7_5/io_wo[12]
+ cb_7_5/io_wo[13] cb_7_5/io_wo[14] cb_7_5/io_wo[15] cb_7_5/io_wo[16] cb_7_5/io_wo[17]
+ cb_7_5/io_wo[18] cb_7_5/io_wo[19] cb_7_5/io_wo[1] cb_7_5/io_wo[20] cb_7_5/io_wo[21]
+ cb_7_5/io_wo[22] cb_7_5/io_wo[23] cb_7_5/io_wo[24] cb_7_5/io_wo[25] cb_7_5/io_wo[26]
+ cb_7_5/io_wo[27] cb_7_5/io_wo[28] cb_7_5/io_wo[29] cb_7_5/io_wo[2] cb_7_5/io_wo[30]
+ cb_7_5/io_wo[31] cb_7_5/io_wo[32] cb_7_5/io_wo[33] cb_7_5/io_wo[34] cb_7_5/io_wo[35]
+ cb_7_5/io_wo[36] cb_7_5/io_wo[37] cb_7_5/io_wo[38] cb_7_5/io_wo[39] cb_7_5/io_wo[3]
+ cb_7_5/io_wo[40] cb_7_5/io_wo[41] cb_7_5/io_wo[42] cb_7_5/io_wo[43] cb_7_5/io_wo[44]
+ cb_7_5/io_wo[45] cb_7_5/io_wo[46] cb_7_5/io_wo[47] cb_7_5/io_wo[48] cb_7_5/io_wo[49]
+ cb_7_5/io_wo[4] cb_7_5/io_wo[50] cb_7_5/io_wo[51] cb_7_5/io_wo[52] cb_7_5/io_wo[53]
+ cb_7_5/io_wo[54] cb_7_5/io_wo[55] cb_7_5/io_wo[56] cb_7_5/io_wo[57] cb_7_5/io_wo[58]
+ cb_7_5/io_wo[59] cb_7_5/io_wo[5] cb_7_5/io_wo[60] cb_7_5/io_wo[61] cb_7_5/io_wo[62]
+ cb_7_5/io_wo[63] cb_7_5/io_wo[6] cb_7_5/io_wo[7] cb_7_5/io_wo[8] cb_7_5/io_wo[9]
+ cb_7_4/io_i_0_ci cb_7_4/io_i_0_in1[0] cb_7_4/io_i_0_in1[1] cb_7_4/io_i_0_in1[2]
+ cb_7_4/io_i_0_in1[3] cb_7_4/io_i_0_in1[4] cb_7_4/io_i_0_in1[5] cb_7_4/io_i_0_in1[6]
+ cb_7_4/io_i_0_in1[7] cb_7_4/io_i_1_ci cb_7_4/io_i_1_in1[0] cb_7_4/io_i_1_in1[1]
+ cb_7_4/io_i_1_in1[2] cb_7_4/io_i_1_in1[3] cb_7_4/io_i_1_in1[4] cb_7_4/io_i_1_in1[5]
+ cb_7_4/io_i_1_in1[6] cb_7_4/io_i_1_in1[7] cb_7_4/io_i_2_ci cb_7_4/io_i_2_in1[0]
+ cb_7_4/io_i_2_in1[1] cb_7_4/io_i_2_in1[2] cb_7_4/io_i_2_in1[3] cb_7_4/io_i_2_in1[4]
+ cb_7_4/io_i_2_in1[5] cb_7_4/io_i_2_in1[6] cb_7_4/io_i_2_in1[7] cb_7_4/io_i_3_ci
+ cb_7_4/io_i_3_in1[0] cb_7_4/io_i_3_in1[1] cb_7_4/io_i_3_in1[2] cb_7_4/io_i_3_in1[3]
+ cb_7_4/io_i_3_in1[4] cb_7_4/io_i_3_in1[5] cb_7_4/io_i_3_in1[6] cb_7_4/io_i_3_in1[7]
+ cb_7_4/io_i_4_ci cb_7_4/io_i_4_in1[0] cb_7_4/io_i_4_in1[1] cb_7_4/io_i_4_in1[2]
+ cb_7_4/io_i_4_in1[3] cb_7_4/io_i_4_in1[4] cb_7_4/io_i_4_in1[5] cb_7_4/io_i_4_in1[6]
+ cb_7_4/io_i_4_in1[7] cb_7_4/io_i_5_ci cb_7_4/io_i_5_in1[0] cb_7_4/io_i_5_in1[1]
+ cb_7_4/io_i_5_in1[2] cb_7_4/io_i_5_in1[3] cb_7_4/io_i_5_in1[4] cb_7_4/io_i_5_in1[5]
+ cb_7_4/io_i_5_in1[6] cb_7_4/io_i_5_in1[7] cb_7_4/io_i_6_ci cb_7_4/io_i_6_in1[0]
+ cb_7_4/io_i_6_in1[1] cb_7_4/io_i_6_in1[2] cb_7_4/io_i_6_in1[3] cb_7_4/io_i_6_in1[4]
+ cb_7_4/io_i_6_in1[5] cb_7_4/io_i_6_in1[6] cb_7_4/io_i_6_in1[7] cb_7_4/io_i_7_ci
+ cb_7_4/io_i_7_in1[0] cb_7_4/io_i_7_in1[1] cb_7_4/io_i_7_in1[2] cb_7_4/io_i_7_in1[3]
+ cb_7_4/io_i_7_in1[4] cb_7_4/io_i_7_in1[5] cb_7_4/io_i_7_in1[6] cb_7_4/io_i_7_in1[7]
+ cb_7_5/io_i_0_ci cb_7_5/io_i_0_in1[0] cb_7_5/io_i_0_in1[1] cb_7_5/io_i_0_in1[2]
+ cb_7_5/io_i_0_in1[3] cb_7_5/io_i_0_in1[4] cb_7_5/io_i_0_in1[5] cb_7_5/io_i_0_in1[6]
+ cb_7_5/io_i_0_in1[7] cb_7_5/io_i_1_ci cb_7_5/io_i_1_in1[0] cb_7_5/io_i_1_in1[1]
+ cb_7_5/io_i_1_in1[2] cb_7_5/io_i_1_in1[3] cb_7_5/io_i_1_in1[4] cb_7_5/io_i_1_in1[5]
+ cb_7_5/io_i_1_in1[6] cb_7_5/io_i_1_in1[7] cb_7_5/io_i_2_ci cb_7_5/io_i_2_in1[0]
+ cb_7_5/io_i_2_in1[1] cb_7_5/io_i_2_in1[2] cb_7_5/io_i_2_in1[3] cb_7_5/io_i_2_in1[4]
+ cb_7_5/io_i_2_in1[5] cb_7_5/io_i_2_in1[6] cb_7_5/io_i_2_in1[7] cb_7_5/io_i_3_ci
+ cb_7_5/io_i_3_in1[0] cb_7_5/io_i_3_in1[1] cb_7_5/io_i_3_in1[2] cb_7_5/io_i_3_in1[3]
+ cb_7_5/io_i_3_in1[4] cb_7_5/io_i_3_in1[5] cb_7_5/io_i_3_in1[6] cb_7_5/io_i_3_in1[7]
+ cb_7_5/io_i_4_ci cb_7_5/io_i_4_in1[0] cb_7_5/io_i_4_in1[1] cb_7_5/io_i_4_in1[2]
+ cb_7_5/io_i_4_in1[3] cb_7_5/io_i_4_in1[4] cb_7_5/io_i_4_in1[5] cb_7_5/io_i_4_in1[6]
+ cb_7_5/io_i_4_in1[7] cb_7_5/io_i_5_ci cb_7_5/io_i_5_in1[0] cb_7_5/io_i_5_in1[1]
+ cb_7_5/io_i_5_in1[2] cb_7_5/io_i_5_in1[3] cb_7_5/io_i_5_in1[4] cb_7_5/io_i_5_in1[5]
+ cb_7_5/io_i_5_in1[6] cb_7_5/io_i_5_in1[7] cb_7_5/io_i_6_ci cb_7_5/io_i_6_in1[0]
+ cb_7_5/io_i_6_in1[1] cb_7_5/io_i_6_in1[2] cb_7_5/io_i_6_in1[3] cb_7_5/io_i_6_in1[4]
+ cb_7_5/io_i_6_in1[5] cb_7_5/io_i_6_in1[6] cb_7_5/io_i_6_in1[7] cb_7_5/io_i_7_ci
+ cb_7_5/io_i_7_in1[0] cb_7_5/io_i_7_in1[1] cb_7_5/io_i_7_in1[2] cb_7_5/io_i_7_in1[3]
+ cb_7_5/io_i_7_in1[4] cb_7_5/io_i_7_in1[5] cb_7_5/io_i_7_in1[6] cb_7_5/io_i_7_in1[7]
+ cb_7_4/io_vci cb_7_5/io_vci cb_7_4/io_vi cb_7_9/io_we_i cb_7_4/io_wo[0] cb_7_4/io_wo[10]
+ cb_7_4/io_wo[11] cb_7_4/io_wo[12] cb_7_4/io_wo[13] cb_7_4/io_wo[14] cb_7_4/io_wo[15]
+ cb_7_4/io_wo[16] cb_7_4/io_wo[17] cb_7_4/io_wo[18] cb_7_4/io_wo[19] cb_7_4/io_wo[1]
+ cb_7_4/io_wo[20] cb_7_4/io_wo[21] cb_7_4/io_wo[22] cb_7_4/io_wo[23] cb_7_4/io_wo[24]
+ cb_7_4/io_wo[25] cb_7_4/io_wo[26] cb_7_4/io_wo[27] cb_7_4/io_wo[28] cb_7_4/io_wo[29]
+ cb_7_4/io_wo[2] cb_7_4/io_wo[30] cb_7_4/io_wo[31] cb_7_4/io_wo[32] cb_7_4/io_wo[33]
+ cb_7_4/io_wo[34] cb_7_4/io_wo[35] cb_7_4/io_wo[36] cb_7_4/io_wo[37] cb_7_4/io_wo[38]
+ cb_7_4/io_wo[39] cb_7_4/io_wo[3] cb_7_4/io_wo[40] cb_7_4/io_wo[41] cb_7_4/io_wo[42]
+ cb_7_4/io_wo[43] cb_7_4/io_wo[44] cb_7_4/io_wo[45] cb_7_4/io_wo[46] cb_7_4/io_wo[47]
+ cb_7_4/io_wo[48] cb_7_4/io_wo[49] cb_7_4/io_wo[4] cb_7_4/io_wo[50] cb_7_4/io_wo[51]
+ cb_7_4/io_wo[52] cb_7_4/io_wo[53] cb_7_4/io_wo[54] cb_7_4/io_wo[55] cb_7_4/io_wo[56]
+ cb_7_4/io_wo[57] cb_7_4/io_wo[58] cb_7_4/io_wo[59] cb_7_4/io_wo[5] cb_7_4/io_wo[60]
+ cb_7_4/io_wo[61] cb_7_4/io_wo[62] cb_7_4/io_wo[63] cb_7_4/io_wo[6] cb_7_4/io_wo[7]
+ cb_7_4/io_wo[8] cb_7_4/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_5_1 cb_5_9/io_adr_i[0] cb_5_9/io_adr_i[1] cb_5_1/io_cs_i cb_5_9/io_dat_i[0] cb_5_9/io_dat_i[10]
+ cb_5_9/io_dat_i[11] cb_5_9/io_dat_i[12] cb_5_9/io_dat_i[13] cb_5_9/io_dat_i[14]
+ cb_5_9/io_dat_i[15] cb_5_9/io_dat_i[1] cb_5_9/io_dat_i[2] cb_5_9/io_dat_i[3] cb_5_9/io_dat_i[4]
+ cb_5_9/io_dat_i[5] cb_5_9/io_dat_i[6] cb_5_9/io_dat_i[7] cb_5_9/io_dat_i[8] cb_5_9/io_dat_i[9]
+ cb_5_1/io_dat_o[0] cb_5_1/io_dat_o[10] cb_5_1/io_dat_o[11] cb_5_1/io_dat_o[12] cb_5_1/io_dat_o[13]
+ cb_5_1/io_dat_o[14] cb_5_1/io_dat_o[15] cb_5_1/io_dat_o[1] cb_5_1/io_dat_o[2] cb_5_1/io_dat_o[3]
+ cb_5_1/io_dat_o[4] cb_5_1/io_dat_o[5] cb_5_1/io_dat_o[6] cb_5_1/io_dat_o[7] cb_5_1/io_dat_o[8]
+ cb_5_1/io_dat_o[9] cb_5_2/io_wo[0] cb_5_2/io_wo[10] cb_5_2/io_wo[11] cb_5_2/io_wo[12]
+ cb_5_2/io_wo[13] cb_5_2/io_wo[14] cb_5_2/io_wo[15] cb_5_2/io_wo[16] cb_5_2/io_wo[17]
+ cb_5_2/io_wo[18] cb_5_2/io_wo[19] cb_5_2/io_wo[1] cb_5_2/io_wo[20] cb_5_2/io_wo[21]
+ cb_5_2/io_wo[22] cb_5_2/io_wo[23] cb_5_2/io_wo[24] cb_5_2/io_wo[25] cb_5_2/io_wo[26]
+ cb_5_2/io_wo[27] cb_5_2/io_wo[28] cb_5_2/io_wo[29] cb_5_2/io_wo[2] cb_5_2/io_wo[30]
+ cb_5_2/io_wo[31] cb_5_2/io_wo[32] cb_5_2/io_wo[33] cb_5_2/io_wo[34] cb_5_2/io_wo[35]
+ cb_5_2/io_wo[36] cb_5_2/io_wo[37] cb_5_2/io_wo[38] cb_5_2/io_wo[39] cb_5_2/io_wo[3]
+ cb_5_2/io_wo[40] cb_5_2/io_wo[41] cb_5_2/io_wo[42] cb_5_2/io_wo[43] cb_5_2/io_wo[44]
+ cb_5_2/io_wo[45] cb_5_2/io_wo[46] cb_5_2/io_wo[47] cb_5_2/io_wo[48] cb_5_2/io_wo[49]
+ cb_5_2/io_wo[4] cb_5_2/io_wo[50] cb_5_2/io_wo[51] cb_5_2/io_wo[52] cb_5_2/io_wo[53]
+ cb_5_2/io_wo[54] cb_5_2/io_wo[55] cb_5_2/io_wo[56] cb_5_2/io_wo[57] cb_5_2/io_wo[58]
+ cb_5_2/io_wo[59] cb_5_2/io_wo[5] cb_5_2/io_wo[60] cb_5_2/io_wo[61] cb_5_2/io_wo[62]
+ cb_5_2/io_wo[63] cb_5_2/io_wo[6] cb_5_2/io_wo[7] cb_5_2/io_wo[8] cb_5_2/io_wo[9]
+ cb_5_1/io_i_0_ci cb_5_1/io_i_0_in1[0] cb_5_1/io_i_0_in1[1] cb_5_1/io_i_0_in1[2]
+ cb_5_1/io_i_0_in1[3] cb_5_1/io_i_0_in1[4] cb_5_1/io_i_0_in1[5] cb_5_1/io_i_0_in1[6]
+ cb_5_1/io_i_0_in1[7] cb_5_1/io_i_1_ci cb_5_1/io_i_1_in1[0] cb_5_1/io_i_1_in1[1]
+ cb_5_1/io_i_1_in1[2] cb_5_1/io_i_1_in1[3] cb_5_1/io_i_1_in1[4] cb_5_1/io_i_1_in1[5]
+ cb_5_1/io_i_1_in1[6] cb_5_1/io_i_1_in1[7] cb_5_1/io_i_2_ci cb_5_1/io_i_2_in1[0]
+ cb_5_1/io_i_2_in1[1] cb_5_1/io_i_2_in1[2] cb_5_1/io_i_2_in1[3] cb_5_1/io_i_2_in1[4]
+ cb_5_1/io_i_2_in1[5] cb_5_1/io_i_2_in1[6] cb_5_1/io_i_2_in1[7] cb_5_1/io_i_3_ci
+ cb_5_1/io_i_3_in1[0] cb_5_1/io_i_3_in1[1] cb_5_1/io_i_3_in1[2] cb_5_1/io_i_3_in1[3]
+ cb_5_1/io_i_3_in1[4] cb_5_1/io_i_3_in1[5] cb_5_1/io_i_3_in1[6] cb_5_1/io_i_3_in1[7]
+ cb_5_1/io_i_4_ci cb_5_1/io_i_4_in1[0] cb_5_1/io_i_4_in1[1] cb_5_1/io_i_4_in1[2]
+ cb_5_1/io_i_4_in1[3] cb_5_1/io_i_4_in1[4] cb_5_1/io_i_4_in1[5] cb_5_1/io_i_4_in1[6]
+ cb_5_1/io_i_4_in1[7] cb_5_1/io_i_5_ci cb_5_1/io_i_5_in1[0] cb_5_1/io_i_5_in1[1]
+ cb_5_1/io_i_5_in1[2] cb_5_1/io_i_5_in1[3] cb_5_1/io_i_5_in1[4] cb_5_1/io_i_5_in1[5]
+ cb_5_1/io_i_5_in1[6] cb_5_1/io_i_5_in1[7] cb_5_1/io_i_6_ci cb_5_1/io_i_6_in1[0]
+ cb_5_1/io_i_6_in1[1] cb_5_1/io_i_6_in1[2] cb_5_1/io_i_6_in1[3] cb_5_1/io_i_6_in1[4]
+ cb_5_1/io_i_6_in1[5] cb_5_1/io_i_6_in1[6] cb_5_1/io_i_6_in1[7] cb_5_1/io_i_7_ci
+ cb_5_1/io_i_7_in1[0] cb_5_1/io_i_7_in1[1] cb_5_1/io_i_7_in1[2] cb_5_1/io_i_7_in1[3]
+ cb_5_1/io_i_7_in1[4] cb_5_1/io_i_7_in1[5] cb_5_1/io_i_7_in1[6] cb_5_1/io_i_7_in1[7]
+ cb_5_2/io_i_0_ci cb_5_2/io_i_0_in1[0] cb_5_2/io_i_0_in1[1] cb_5_2/io_i_0_in1[2]
+ cb_5_2/io_i_0_in1[3] cb_5_2/io_i_0_in1[4] cb_5_2/io_i_0_in1[5] cb_5_2/io_i_0_in1[6]
+ cb_5_2/io_i_0_in1[7] cb_5_2/io_i_1_ci cb_5_2/io_i_1_in1[0] cb_5_2/io_i_1_in1[1]
+ cb_5_2/io_i_1_in1[2] cb_5_2/io_i_1_in1[3] cb_5_2/io_i_1_in1[4] cb_5_2/io_i_1_in1[5]
+ cb_5_2/io_i_1_in1[6] cb_5_2/io_i_1_in1[7] cb_5_2/io_i_2_ci cb_5_2/io_i_2_in1[0]
+ cb_5_2/io_i_2_in1[1] cb_5_2/io_i_2_in1[2] cb_5_2/io_i_2_in1[3] cb_5_2/io_i_2_in1[4]
+ cb_5_2/io_i_2_in1[5] cb_5_2/io_i_2_in1[6] cb_5_2/io_i_2_in1[7] cb_5_2/io_i_3_ci
+ cb_5_2/io_i_3_in1[0] cb_5_2/io_i_3_in1[1] cb_5_2/io_i_3_in1[2] cb_5_2/io_i_3_in1[3]
+ cb_5_2/io_i_3_in1[4] cb_5_2/io_i_3_in1[5] cb_5_2/io_i_3_in1[6] cb_5_2/io_i_3_in1[7]
+ cb_5_2/io_i_4_ci cb_5_2/io_i_4_in1[0] cb_5_2/io_i_4_in1[1] cb_5_2/io_i_4_in1[2]
+ cb_5_2/io_i_4_in1[3] cb_5_2/io_i_4_in1[4] cb_5_2/io_i_4_in1[5] cb_5_2/io_i_4_in1[6]
+ cb_5_2/io_i_4_in1[7] cb_5_2/io_i_5_ci cb_5_2/io_i_5_in1[0] cb_5_2/io_i_5_in1[1]
+ cb_5_2/io_i_5_in1[2] cb_5_2/io_i_5_in1[3] cb_5_2/io_i_5_in1[4] cb_5_2/io_i_5_in1[5]
+ cb_5_2/io_i_5_in1[6] cb_5_2/io_i_5_in1[7] cb_5_2/io_i_6_ci cb_5_2/io_i_6_in1[0]
+ cb_5_2/io_i_6_in1[1] cb_5_2/io_i_6_in1[2] cb_5_2/io_i_6_in1[3] cb_5_2/io_i_6_in1[4]
+ cb_5_2/io_i_6_in1[5] cb_5_2/io_i_6_in1[6] cb_5_2/io_i_6_in1[7] cb_5_2/io_i_7_ci
+ cb_5_2/io_i_7_in1[0] cb_5_2/io_i_7_in1[1] cb_5_2/io_i_7_in1[2] cb_5_2/io_i_7_in1[3]
+ cb_5_2/io_i_7_in1[4] cb_5_2/io_i_7_in1[5] cb_5_2/io_i_7_in1[6] cb_5_2/io_i_7_in1[7]
+ cb_5_1/io_vci cb_5_2/io_vci cb_5_1/io_vi cb_5_9/io_we_i cb_5_1/io_wo[0] cb_5_1/io_wo[10]
+ cb_5_1/io_wo[11] cb_5_1/io_wo[12] cb_5_1/io_wo[13] cb_5_1/io_wo[14] cb_5_1/io_wo[15]
+ cb_5_1/io_wo[16] cb_5_1/io_wo[17] cb_5_1/io_wo[18] cb_5_1/io_wo[19] cb_5_1/io_wo[1]
+ cb_5_1/io_wo[20] cb_5_1/io_wo[21] cb_5_1/io_wo[22] cb_5_1/io_wo[23] cb_5_1/io_wo[24]
+ cb_5_1/io_wo[25] cb_5_1/io_wo[26] cb_5_1/io_wo[27] cb_5_1/io_wo[28] cb_5_1/io_wo[29]
+ cb_5_1/io_wo[2] cb_5_1/io_wo[30] cb_5_1/io_wo[31] cb_5_1/io_wo[32] cb_5_1/io_wo[33]
+ cb_5_1/io_wo[34] cb_5_1/io_wo[35] cb_5_1/io_wo[36] cb_5_1/io_wo[37] cb_5_1/io_wo[38]
+ cb_5_1/io_wo[39] cb_5_1/io_wo[3] cb_5_1/io_wo[40] cb_5_1/io_wo[41] cb_5_1/io_wo[42]
+ cb_5_1/io_wo[43] cb_5_1/io_wo[44] cb_5_1/io_wo[45] cb_5_1/io_wo[46] cb_5_1/io_wo[47]
+ cb_5_1/io_wo[48] cb_5_1/io_wo[49] cb_5_1/io_wo[4] cb_5_1/io_wo[50] cb_5_1/io_wo[51]
+ cb_5_1/io_wo[52] cb_5_1/io_wo[53] cb_5_1/io_wo[54] cb_5_1/io_wo[55] cb_5_1/io_wo[56]
+ cb_5_1/io_wo[57] cb_5_1/io_wo[58] cb_5_1/io_wo[59] cb_5_1/io_wo[5] cb_5_1/io_wo[60]
+ cb_5_1/io_wo[61] cb_5_1/io_wo[62] cb_5_1/io_wo[63] cb_5_1/io_wo[6] cb_5_1/io_wo[7]
+ cb_5_1/io_wo[8] cb_5_1/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_7_5 cb_7_9/io_adr_i[0] cb_7_9/io_adr_i[1] cb_7_5/io_cs_i cb_7_9/io_dat_i[0] cb_7_9/io_dat_i[10]
+ cb_7_9/io_dat_i[11] cb_7_9/io_dat_i[12] cb_7_9/io_dat_i[13] cb_7_9/io_dat_i[14]
+ cb_7_9/io_dat_i[15] cb_7_9/io_dat_i[1] cb_7_9/io_dat_i[2] cb_7_9/io_dat_i[3] cb_7_9/io_dat_i[4]
+ cb_7_9/io_dat_i[5] cb_7_9/io_dat_i[6] cb_7_9/io_dat_i[7] cb_7_9/io_dat_i[8] cb_7_9/io_dat_i[9]
+ cb_7_5/io_dat_o[0] cb_7_5/io_dat_o[10] cb_7_5/io_dat_o[11] cb_7_5/io_dat_o[12] cb_7_5/io_dat_o[13]
+ cb_7_5/io_dat_o[14] cb_7_5/io_dat_o[15] cb_7_5/io_dat_o[1] cb_7_5/io_dat_o[2] cb_7_5/io_dat_o[3]
+ cb_7_5/io_dat_o[4] cb_7_5/io_dat_o[5] cb_7_5/io_dat_o[6] cb_7_5/io_dat_o[7] cb_7_5/io_dat_o[8]
+ cb_7_5/io_dat_o[9] cb_7_6/io_wo[0] cb_7_6/io_wo[10] cb_7_6/io_wo[11] cb_7_6/io_wo[12]
+ cb_7_6/io_wo[13] cb_7_6/io_wo[14] cb_7_6/io_wo[15] cb_7_6/io_wo[16] cb_7_6/io_wo[17]
+ cb_7_6/io_wo[18] cb_7_6/io_wo[19] cb_7_6/io_wo[1] cb_7_6/io_wo[20] cb_7_6/io_wo[21]
+ cb_7_6/io_wo[22] cb_7_6/io_wo[23] cb_7_6/io_wo[24] cb_7_6/io_wo[25] cb_7_6/io_wo[26]
+ cb_7_6/io_wo[27] cb_7_6/io_wo[28] cb_7_6/io_wo[29] cb_7_6/io_wo[2] cb_7_6/io_wo[30]
+ cb_7_6/io_wo[31] cb_7_6/io_wo[32] cb_7_6/io_wo[33] cb_7_6/io_wo[34] cb_7_6/io_wo[35]
+ cb_7_6/io_wo[36] cb_7_6/io_wo[37] cb_7_6/io_wo[38] cb_7_6/io_wo[39] cb_7_6/io_wo[3]
+ cb_7_6/io_wo[40] cb_7_6/io_wo[41] cb_7_6/io_wo[42] cb_7_6/io_wo[43] cb_7_6/io_wo[44]
+ cb_7_6/io_wo[45] cb_7_6/io_wo[46] cb_7_6/io_wo[47] cb_7_6/io_wo[48] cb_7_6/io_wo[49]
+ cb_7_6/io_wo[4] cb_7_6/io_wo[50] cb_7_6/io_wo[51] cb_7_6/io_wo[52] cb_7_6/io_wo[53]
+ cb_7_6/io_wo[54] cb_7_6/io_wo[55] cb_7_6/io_wo[56] cb_7_6/io_wo[57] cb_7_6/io_wo[58]
+ cb_7_6/io_wo[59] cb_7_6/io_wo[5] cb_7_6/io_wo[60] cb_7_6/io_wo[61] cb_7_6/io_wo[62]
+ cb_7_6/io_wo[63] cb_7_6/io_wo[6] cb_7_6/io_wo[7] cb_7_6/io_wo[8] cb_7_6/io_wo[9]
+ cb_7_5/io_i_0_ci cb_7_5/io_i_0_in1[0] cb_7_5/io_i_0_in1[1] cb_7_5/io_i_0_in1[2]
+ cb_7_5/io_i_0_in1[3] cb_7_5/io_i_0_in1[4] cb_7_5/io_i_0_in1[5] cb_7_5/io_i_0_in1[6]
+ cb_7_5/io_i_0_in1[7] cb_7_5/io_i_1_ci cb_7_5/io_i_1_in1[0] cb_7_5/io_i_1_in1[1]
+ cb_7_5/io_i_1_in1[2] cb_7_5/io_i_1_in1[3] cb_7_5/io_i_1_in1[4] cb_7_5/io_i_1_in1[5]
+ cb_7_5/io_i_1_in1[6] cb_7_5/io_i_1_in1[7] cb_7_5/io_i_2_ci cb_7_5/io_i_2_in1[0]
+ cb_7_5/io_i_2_in1[1] cb_7_5/io_i_2_in1[2] cb_7_5/io_i_2_in1[3] cb_7_5/io_i_2_in1[4]
+ cb_7_5/io_i_2_in1[5] cb_7_5/io_i_2_in1[6] cb_7_5/io_i_2_in1[7] cb_7_5/io_i_3_ci
+ cb_7_5/io_i_3_in1[0] cb_7_5/io_i_3_in1[1] cb_7_5/io_i_3_in1[2] cb_7_5/io_i_3_in1[3]
+ cb_7_5/io_i_3_in1[4] cb_7_5/io_i_3_in1[5] cb_7_5/io_i_3_in1[6] cb_7_5/io_i_3_in1[7]
+ cb_7_5/io_i_4_ci cb_7_5/io_i_4_in1[0] cb_7_5/io_i_4_in1[1] cb_7_5/io_i_4_in1[2]
+ cb_7_5/io_i_4_in1[3] cb_7_5/io_i_4_in1[4] cb_7_5/io_i_4_in1[5] cb_7_5/io_i_4_in1[6]
+ cb_7_5/io_i_4_in1[7] cb_7_5/io_i_5_ci cb_7_5/io_i_5_in1[0] cb_7_5/io_i_5_in1[1]
+ cb_7_5/io_i_5_in1[2] cb_7_5/io_i_5_in1[3] cb_7_5/io_i_5_in1[4] cb_7_5/io_i_5_in1[5]
+ cb_7_5/io_i_5_in1[6] cb_7_5/io_i_5_in1[7] cb_7_5/io_i_6_ci cb_7_5/io_i_6_in1[0]
+ cb_7_5/io_i_6_in1[1] cb_7_5/io_i_6_in1[2] cb_7_5/io_i_6_in1[3] cb_7_5/io_i_6_in1[4]
+ cb_7_5/io_i_6_in1[5] cb_7_5/io_i_6_in1[6] cb_7_5/io_i_6_in1[7] cb_7_5/io_i_7_ci
+ cb_7_5/io_i_7_in1[0] cb_7_5/io_i_7_in1[1] cb_7_5/io_i_7_in1[2] cb_7_5/io_i_7_in1[3]
+ cb_7_5/io_i_7_in1[4] cb_7_5/io_i_7_in1[5] cb_7_5/io_i_7_in1[6] cb_7_5/io_i_7_in1[7]
+ cb_7_6/io_i_0_ci cb_7_6/io_i_0_in1[0] cb_7_6/io_i_0_in1[1] cb_7_6/io_i_0_in1[2]
+ cb_7_6/io_i_0_in1[3] cb_7_6/io_i_0_in1[4] cb_7_6/io_i_0_in1[5] cb_7_6/io_i_0_in1[6]
+ cb_7_6/io_i_0_in1[7] cb_7_6/io_i_1_ci cb_7_6/io_i_1_in1[0] cb_7_6/io_i_1_in1[1]
+ cb_7_6/io_i_1_in1[2] cb_7_6/io_i_1_in1[3] cb_7_6/io_i_1_in1[4] cb_7_6/io_i_1_in1[5]
+ cb_7_6/io_i_1_in1[6] cb_7_6/io_i_1_in1[7] cb_7_6/io_i_2_ci cb_7_6/io_i_2_in1[0]
+ cb_7_6/io_i_2_in1[1] cb_7_6/io_i_2_in1[2] cb_7_6/io_i_2_in1[3] cb_7_6/io_i_2_in1[4]
+ cb_7_6/io_i_2_in1[5] cb_7_6/io_i_2_in1[6] cb_7_6/io_i_2_in1[7] cb_7_6/io_i_3_ci
+ cb_7_6/io_i_3_in1[0] cb_7_6/io_i_3_in1[1] cb_7_6/io_i_3_in1[2] cb_7_6/io_i_3_in1[3]
+ cb_7_6/io_i_3_in1[4] cb_7_6/io_i_3_in1[5] cb_7_6/io_i_3_in1[6] cb_7_6/io_i_3_in1[7]
+ cb_7_6/io_i_4_ci cb_7_6/io_i_4_in1[0] cb_7_6/io_i_4_in1[1] cb_7_6/io_i_4_in1[2]
+ cb_7_6/io_i_4_in1[3] cb_7_6/io_i_4_in1[4] cb_7_6/io_i_4_in1[5] cb_7_6/io_i_4_in1[6]
+ cb_7_6/io_i_4_in1[7] cb_7_6/io_i_5_ci cb_7_6/io_i_5_in1[0] cb_7_6/io_i_5_in1[1]
+ cb_7_6/io_i_5_in1[2] cb_7_6/io_i_5_in1[3] cb_7_6/io_i_5_in1[4] cb_7_6/io_i_5_in1[5]
+ cb_7_6/io_i_5_in1[6] cb_7_6/io_i_5_in1[7] cb_7_6/io_i_6_ci cb_7_6/io_i_6_in1[0]
+ cb_7_6/io_i_6_in1[1] cb_7_6/io_i_6_in1[2] cb_7_6/io_i_6_in1[3] cb_7_6/io_i_6_in1[4]
+ cb_7_6/io_i_6_in1[5] cb_7_6/io_i_6_in1[6] cb_7_6/io_i_6_in1[7] cb_7_6/io_i_7_ci
+ cb_7_6/io_i_7_in1[0] cb_7_6/io_i_7_in1[1] cb_7_6/io_i_7_in1[2] cb_7_6/io_i_7_in1[3]
+ cb_7_6/io_i_7_in1[4] cb_7_6/io_i_7_in1[5] cb_7_6/io_i_7_in1[6] cb_7_6/io_i_7_in1[7]
+ cb_7_5/io_vci cb_7_6/io_vci cb_7_5/io_vi cb_7_9/io_we_i cb_7_5/io_wo[0] cb_7_5/io_wo[10]
+ cb_7_5/io_wo[11] cb_7_5/io_wo[12] cb_7_5/io_wo[13] cb_7_5/io_wo[14] cb_7_5/io_wo[15]
+ cb_7_5/io_wo[16] cb_7_5/io_wo[17] cb_7_5/io_wo[18] cb_7_5/io_wo[19] cb_7_5/io_wo[1]
+ cb_7_5/io_wo[20] cb_7_5/io_wo[21] cb_7_5/io_wo[22] cb_7_5/io_wo[23] cb_7_5/io_wo[24]
+ cb_7_5/io_wo[25] cb_7_5/io_wo[26] cb_7_5/io_wo[27] cb_7_5/io_wo[28] cb_7_5/io_wo[29]
+ cb_7_5/io_wo[2] cb_7_5/io_wo[30] cb_7_5/io_wo[31] cb_7_5/io_wo[32] cb_7_5/io_wo[33]
+ cb_7_5/io_wo[34] cb_7_5/io_wo[35] cb_7_5/io_wo[36] cb_7_5/io_wo[37] cb_7_5/io_wo[38]
+ cb_7_5/io_wo[39] cb_7_5/io_wo[3] cb_7_5/io_wo[40] cb_7_5/io_wo[41] cb_7_5/io_wo[42]
+ cb_7_5/io_wo[43] cb_7_5/io_wo[44] cb_7_5/io_wo[45] cb_7_5/io_wo[46] cb_7_5/io_wo[47]
+ cb_7_5/io_wo[48] cb_7_5/io_wo[49] cb_7_5/io_wo[4] cb_7_5/io_wo[50] cb_7_5/io_wo[51]
+ cb_7_5/io_wo[52] cb_7_5/io_wo[53] cb_7_5/io_wo[54] cb_7_5/io_wo[55] cb_7_5/io_wo[56]
+ cb_7_5/io_wo[57] cb_7_5/io_wo[58] cb_7_5/io_wo[59] cb_7_5/io_wo[5] cb_7_5/io_wo[60]
+ cb_7_5/io_wo[61] cb_7_5/io_wo[62] cb_7_5/io_wo[63] cb_7_5/io_wo[6] cb_7_5/io_wo[7]
+ cb_7_5/io_wo[8] cb_7_5/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_5_2 cb_5_9/io_adr_i[0] cb_5_9/io_adr_i[1] cb_5_2/io_cs_i cb_5_9/io_dat_i[0] cb_5_9/io_dat_i[10]
+ cb_5_9/io_dat_i[11] cb_5_9/io_dat_i[12] cb_5_9/io_dat_i[13] cb_5_9/io_dat_i[14]
+ cb_5_9/io_dat_i[15] cb_5_9/io_dat_i[1] cb_5_9/io_dat_i[2] cb_5_9/io_dat_i[3] cb_5_9/io_dat_i[4]
+ cb_5_9/io_dat_i[5] cb_5_9/io_dat_i[6] cb_5_9/io_dat_i[7] cb_5_9/io_dat_i[8] cb_5_9/io_dat_i[9]
+ cb_5_2/io_dat_o[0] cb_5_2/io_dat_o[10] cb_5_2/io_dat_o[11] cb_5_2/io_dat_o[12] cb_5_2/io_dat_o[13]
+ cb_5_2/io_dat_o[14] cb_5_2/io_dat_o[15] cb_5_2/io_dat_o[1] cb_5_2/io_dat_o[2] cb_5_2/io_dat_o[3]
+ cb_5_2/io_dat_o[4] cb_5_2/io_dat_o[5] cb_5_2/io_dat_o[6] cb_5_2/io_dat_o[7] cb_5_2/io_dat_o[8]
+ cb_5_2/io_dat_o[9] cb_5_3/io_wo[0] cb_5_3/io_wo[10] cb_5_3/io_wo[11] cb_5_3/io_wo[12]
+ cb_5_3/io_wo[13] cb_5_3/io_wo[14] cb_5_3/io_wo[15] cb_5_3/io_wo[16] cb_5_3/io_wo[17]
+ cb_5_3/io_wo[18] cb_5_3/io_wo[19] cb_5_3/io_wo[1] cb_5_3/io_wo[20] cb_5_3/io_wo[21]
+ cb_5_3/io_wo[22] cb_5_3/io_wo[23] cb_5_3/io_wo[24] cb_5_3/io_wo[25] cb_5_3/io_wo[26]
+ cb_5_3/io_wo[27] cb_5_3/io_wo[28] cb_5_3/io_wo[29] cb_5_3/io_wo[2] cb_5_3/io_wo[30]
+ cb_5_3/io_wo[31] cb_5_3/io_wo[32] cb_5_3/io_wo[33] cb_5_3/io_wo[34] cb_5_3/io_wo[35]
+ cb_5_3/io_wo[36] cb_5_3/io_wo[37] cb_5_3/io_wo[38] cb_5_3/io_wo[39] cb_5_3/io_wo[3]
+ cb_5_3/io_wo[40] cb_5_3/io_wo[41] cb_5_3/io_wo[42] cb_5_3/io_wo[43] cb_5_3/io_wo[44]
+ cb_5_3/io_wo[45] cb_5_3/io_wo[46] cb_5_3/io_wo[47] cb_5_3/io_wo[48] cb_5_3/io_wo[49]
+ cb_5_3/io_wo[4] cb_5_3/io_wo[50] cb_5_3/io_wo[51] cb_5_3/io_wo[52] cb_5_3/io_wo[53]
+ cb_5_3/io_wo[54] cb_5_3/io_wo[55] cb_5_3/io_wo[56] cb_5_3/io_wo[57] cb_5_3/io_wo[58]
+ cb_5_3/io_wo[59] cb_5_3/io_wo[5] cb_5_3/io_wo[60] cb_5_3/io_wo[61] cb_5_3/io_wo[62]
+ cb_5_3/io_wo[63] cb_5_3/io_wo[6] cb_5_3/io_wo[7] cb_5_3/io_wo[8] cb_5_3/io_wo[9]
+ cb_5_2/io_i_0_ci cb_5_2/io_i_0_in1[0] cb_5_2/io_i_0_in1[1] cb_5_2/io_i_0_in1[2]
+ cb_5_2/io_i_0_in1[3] cb_5_2/io_i_0_in1[4] cb_5_2/io_i_0_in1[5] cb_5_2/io_i_0_in1[6]
+ cb_5_2/io_i_0_in1[7] cb_5_2/io_i_1_ci cb_5_2/io_i_1_in1[0] cb_5_2/io_i_1_in1[1]
+ cb_5_2/io_i_1_in1[2] cb_5_2/io_i_1_in1[3] cb_5_2/io_i_1_in1[4] cb_5_2/io_i_1_in1[5]
+ cb_5_2/io_i_1_in1[6] cb_5_2/io_i_1_in1[7] cb_5_2/io_i_2_ci cb_5_2/io_i_2_in1[0]
+ cb_5_2/io_i_2_in1[1] cb_5_2/io_i_2_in1[2] cb_5_2/io_i_2_in1[3] cb_5_2/io_i_2_in1[4]
+ cb_5_2/io_i_2_in1[5] cb_5_2/io_i_2_in1[6] cb_5_2/io_i_2_in1[7] cb_5_2/io_i_3_ci
+ cb_5_2/io_i_3_in1[0] cb_5_2/io_i_3_in1[1] cb_5_2/io_i_3_in1[2] cb_5_2/io_i_3_in1[3]
+ cb_5_2/io_i_3_in1[4] cb_5_2/io_i_3_in1[5] cb_5_2/io_i_3_in1[6] cb_5_2/io_i_3_in1[7]
+ cb_5_2/io_i_4_ci cb_5_2/io_i_4_in1[0] cb_5_2/io_i_4_in1[1] cb_5_2/io_i_4_in1[2]
+ cb_5_2/io_i_4_in1[3] cb_5_2/io_i_4_in1[4] cb_5_2/io_i_4_in1[5] cb_5_2/io_i_4_in1[6]
+ cb_5_2/io_i_4_in1[7] cb_5_2/io_i_5_ci cb_5_2/io_i_5_in1[0] cb_5_2/io_i_5_in1[1]
+ cb_5_2/io_i_5_in1[2] cb_5_2/io_i_5_in1[3] cb_5_2/io_i_5_in1[4] cb_5_2/io_i_5_in1[5]
+ cb_5_2/io_i_5_in1[6] cb_5_2/io_i_5_in1[7] cb_5_2/io_i_6_ci cb_5_2/io_i_6_in1[0]
+ cb_5_2/io_i_6_in1[1] cb_5_2/io_i_6_in1[2] cb_5_2/io_i_6_in1[3] cb_5_2/io_i_6_in1[4]
+ cb_5_2/io_i_6_in1[5] cb_5_2/io_i_6_in1[6] cb_5_2/io_i_6_in1[7] cb_5_2/io_i_7_ci
+ cb_5_2/io_i_7_in1[0] cb_5_2/io_i_7_in1[1] cb_5_2/io_i_7_in1[2] cb_5_2/io_i_7_in1[3]
+ cb_5_2/io_i_7_in1[4] cb_5_2/io_i_7_in1[5] cb_5_2/io_i_7_in1[6] cb_5_2/io_i_7_in1[7]
+ cb_5_3/io_i_0_ci cb_5_3/io_i_0_in1[0] cb_5_3/io_i_0_in1[1] cb_5_3/io_i_0_in1[2]
+ cb_5_3/io_i_0_in1[3] cb_5_3/io_i_0_in1[4] cb_5_3/io_i_0_in1[5] cb_5_3/io_i_0_in1[6]
+ cb_5_3/io_i_0_in1[7] cb_5_3/io_i_1_ci cb_5_3/io_i_1_in1[0] cb_5_3/io_i_1_in1[1]
+ cb_5_3/io_i_1_in1[2] cb_5_3/io_i_1_in1[3] cb_5_3/io_i_1_in1[4] cb_5_3/io_i_1_in1[5]
+ cb_5_3/io_i_1_in1[6] cb_5_3/io_i_1_in1[7] cb_5_3/io_i_2_ci cb_5_3/io_i_2_in1[0]
+ cb_5_3/io_i_2_in1[1] cb_5_3/io_i_2_in1[2] cb_5_3/io_i_2_in1[3] cb_5_3/io_i_2_in1[4]
+ cb_5_3/io_i_2_in1[5] cb_5_3/io_i_2_in1[6] cb_5_3/io_i_2_in1[7] cb_5_3/io_i_3_ci
+ cb_5_3/io_i_3_in1[0] cb_5_3/io_i_3_in1[1] cb_5_3/io_i_3_in1[2] cb_5_3/io_i_3_in1[3]
+ cb_5_3/io_i_3_in1[4] cb_5_3/io_i_3_in1[5] cb_5_3/io_i_3_in1[6] cb_5_3/io_i_3_in1[7]
+ cb_5_3/io_i_4_ci cb_5_3/io_i_4_in1[0] cb_5_3/io_i_4_in1[1] cb_5_3/io_i_4_in1[2]
+ cb_5_3/io_i_4_in1[3] cb_5_3/io_i_4_in1[4] cb_5_3/io_i_4_in1[5] cb_5_3/io_i_4_in1[6]
+ cb_5_3/io_i_4_in1[7] cb_5_3/io_i_5_ci cb_5_3/io_i_5_in1[0] cb_5_3/io_i_5_in1[1]
+ cb_5_3/io_i_5_in1[2] cb_5_3/io_i_5_in1[3] cb_5_3/io_i_5_in1[4] cb_5_3/io_i_5_in1[5]
+ cb_5_3/io_i_5_in1[6] cb_5_3/io_i_5_in1[7] cb_5_3/io_i_6_ci cb_5_3/io_i_6_in1[0]
+ cb_5_3/io_i_6_in1[1] cb_5_3/io_i_6_in1[2] cb_5_3/io_i_6_in1[3] cb_5_3/io_i_6_in1[4]
+ cb_5_3/io_i_6_in1[5] cb_5_3/io_i_6_in1[6] cb_5_3/io_i_6_in1[7] cb_5_3/io_i_7_ci
+ cb_5_3/io_i_7_in1[0] cb_5_3/io_i_7_in1[1] cb_5_3/io_i_7_in1[2] cb_5_3/io_i_7_in1[3]
+ cb_5_3/io_i_7_in1[4] cb_5_3/io_i_7_in1[5] cb_5_3/io_i_7_in1[6] cb_5_3/io_i_7_in1[7]
+ cb_5_2/io_vci cb_5_3/io_vci cb_5_2/io_vi cb_5_9/io_we_i cb_5_2/io_wo[0] cb_5_2/io_wo[10]
+ cb_5_2/io_wo[11] cb_5_2/io_wo[12] cb_5_2/io_wo[13] cb_5_2/io_wo[14] cb_5_2/io_wo[15]
+ cb_5_2/io_wo[16] cb_5_2/io_wo[17] cb_5_2/io_wo[18] cb_5_2/io_wo[19] cb_5_2/io_wo[1]
+ cb_5_2/io_wo[20] cb_5_2/io_wo[21] cb_5_2/io_wo[22] cb_5_2/io_wo[23] cb_5_2/io_wo[24]
+ cb_5_2/io_wo[25] cb_5_2/io_wo[26] cb_5_2/io_wo[27] cb_5_2/io_wo[28] cb_5_2/io_wo[29]
+ cb_5_2/io_wo[2] cb_5_2/io_wo[30] cb_5_2/io_wo[31] cb_5_2/io_wo[32] cb_5_2/io_wo[33]
+ cb_5_2/io_wo[34] cb_5_2/io_wo[35] cb_5_2/io_wo[36] cb_5_2/io_wo[37] cb_5_2/io_wo[38]
+ cb_5_2/io_wo[39] cb_5_2/io_wo[3] cb_5_2/io_wo[40] cb_5_2/io_wo[41] cb_5_2/io_wo[42]
+ cb_5_2/io_wo[43] cb_5_2/io_wo[44] cb_5_2/io_wo[45] cb_5_2/io_wo[46] cb_5_2/io_wo[47]
+ cb_5_2/io_wo[48] cb_5_2/io_wo[49] cb_5_2/io_wo[4] cb_5_2/io_wo[50] cb_5_2/io_wo[51]
+ cb_5_2/io_wo[52] cb_5_2/io_wo[53] cb_5_2/io_wo[54] cb_5_2/io_wo[55] cb_5_2/io_wo[56]
+ cb_5_2/io_wo[57] cb_5_2/io_wo[58] cb_5_2/io_wo[59] cb_5_2/io_wo[5] cb_5_2/io_wo[60]
+ cb_5_2/io_wo[61] cb_5_2/io_wo[62] cb_5_2/io_wo[63] cb_5_2/io_wo[6] cb_5_2/io_wo[7]
+ cb_5_2/io_wo[8] cb_5_2/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_7_6 cb_7_9/io_adr_i[0] cb_7_9/io_adr_i[1] cb_7_6/io_cs_i cb_7_9/io_dat_i[0] cb_7_9/io_dat_i[10]
+ cb_7_9/io_dat_i[11] cb_7_9/io_dat_i[12] cb_7_9/io_dat_i[13] cb_7_9/io_dat_i[14]
+ cb_7_9/io_dat_i[15] cb_7_9/io_dat_i[1] cb_7_9/io_dat_i[2] cb_7_9/io_dat_i[3] cb_7_9/io_dat_i[4]
+ cb_7_9/io_dat_i[5] cb_7_9/io_dat_i[6] cb_7_9/io_dat_i[7] cb_7_9/io_dat_i[8] cb_7_9/io_dat_i[9]
+ cb_7_6/io_dat_o[0] cb_7_6/io_dat_o[10] cb_7_6/io_dat_o[11] cb_7_6/io_dat_o[12] cb_7_6/io_dat_o[13]
+ cb_7_6/io_dat_o[14] cb_7_6/io_dat_o[15] cb_7_6/io_dat_o[1] cb_7_6/io_dat_o[2] cb_7_6/io_dat_o[3]
+ cb_7_6/io_dat_o[4] cb_7_6/io_dat_o[5] cb_7_6/io_dat_o[6] cb_7_6/io_dat_o[7] cb_7_6/io_dat_o[8]
+ cb_7_6/io_dat_o[9] cb_7_7/io_wo[0] cb_7_7/io_wo[10] cb_7_7/io_wo[11] cb_7_7/io_wo[12]
+ cb_7_7/io_wo[13] cb_7_7/io_wo[14] cb_7_7/io_wo[15] cb_7_7/io_wo[16] cb_7_7/io_wo[17]
+ cb_7_7/io_wo[18] cb_7_7/io_wo[19] cb_7_7/io_wo[1] cb_7_7/io_wo[20] cb_7_7/io_wo[21]
+ cb_7_7/io_wo[22] cb_7_7/io_wo[23] cb_7_7/io_wo[24] cb_7_7/io_wo[25] cb_7_7/io_wo[26]
+ cb_7_7/io_wo[27] cb_7_7/io_wo[28] cb_7_7/io_wo[29] cb_7_7/io_wo[2] cb_7_7/io_wo[30]
+ cb_7_7/io_wo[31] cb_7_7/io_wo[32] cb_7_7/io_wo[33] cb_7_7/io_wo[34] cb_7_7/io_wo[35]
+ cb_7_7/io_wo[36] cb_7_7/io_wo[37] cb_7_7/io_wo[38] cb_7_7/io_wo[39] cb_7_7/io_wo[3]
+ cb_7_7/io_wo[40] cb_7_7/io_wo[41] cb_7_7/io_wo[42] cb_7_7/io_wo[43] cb_7_7/io_wo[44]
+ cb_7_7/io_wo[45] cb_7_7/io_wo[46] cb_7_7/io_wo[47] cb_7_7/io_wo[48] cb_7_7/io_wo[49]
+ cb_7_7/io_wo[4] cb_7_7/io_wo[50] cb_7_7/io_wo[51] cb_7_7/io_wo[52] cb_7_7/io_wo[53]
+ cb_7_7/io_wo[54] cb_7_7/io_wo[55] cb_7_7/io_wo[56] cb_7_7/io_wo[57] cb_7_7/io_wo[58]
+ cb_7_7/io_wo[59] cb_7_7/io_wo[5] cb_7_7/io_wo[60] cb_7_7/io_wo[61] cb_7_7/io_wo[62]
+ cb_7_7/io_wo[63] cb_7_7/io_wo[6] cb_7_7/io_wo[7] cb_7_7/io_wo[8] cb_7_7/io_wo[9]
+ cb_7_6/io_i_0_ci cb_7_6/io_i_0_in1[0] cb_7_6/io_i_0_in1[1] cb_7_6/io_i_0_in1[2]
+ cb_7_6/io_i_0_in1[3] cb_7_6/io_i_0_in1[4] cb_7_6/io_i_0_in1[5] cb_7_6/io_i_0_in1[6]
+ cb_7_6/io_i_0_in1[7] cb_7_6/io_i_1_ci cb_7_6/io_i_1_in1[0] cb_7_6/io_i_1_in1[1]
+ cb_7_6/io_i_1_in1[2] cb_7_6/io_i_1_in1[3] cb_7_6/io_i_1_in1[4] cb_7_6/io_i_1_in1[5]
+ cb_7_6/io_i_1_in1[6] cb_7_6/io_i_1_in1[7] cb_7_6/io_i_2_ci cb_7_6/io_i_2_in1[0]
+ cb_7_6/io_i_2_in1[1] cb_7_6/io_i_2_in1[2] cb_7_6/io_i_2_in1[3] cb_7_6/io_i_2_in1[4]
+ cb_7_6/io_i_2_in1[5] cb_7_6/io_i_2_in1[6] cb_7_6/io_i_2_in1[7] cb_7_6/io_i_3_ci
+ cb_7_6/io_i_3_in1[0] cb_7_6/io_i_3_in1[1] cb_7_6/io_i_3_in1[2] cb_7_6/io_i_3_in1[3]
+ cb_7_6/io_i_3_in1[4] cb_7_6/io_i_3_in1[5] cb_7_6/io_i_3_in1[6] cb_7_6/io_i_3_in1[7]
+ cb_7_6/io_i_4_ci cb_7_6/io_i_4_in1[0] cb_7_6/io_i_4_in1[1] cb_7_6/io_i_4_in1[2]
+ cb_7_6/io_i_4_in1[3] cb_7_6/io_i_4_in1[4] cb_7_6/io_i_4_in1[5] cb_7_6/io_i_4_in1[6]
+ cb_7_6/io_i_4_in1[7] cb_7_6/io_i_5_ci cb_7_6/io_i_5_in1[0] cb_7_6/io_i_5_in1[1]
+ cb_7_6/io_i_5_in1[2] cb_7_6/io_i_5_in1[3] cb_7_6/io_i_5_in1[4] cb_7_6/io_i_5_in1[5]
+ cb_7_6/io_i_5_in1[6] cb_7_6/io_i_5_in1[7] cb_7_6/io_i_6_ci cb_7_6/io_i_6_in1[0]
+ cb_7_6/io_i_6_in1[1] cb_7_6/io_i_6_in1[2] cb_7_6/io_i_6_in1[3] cb_7_6/io_i_6_in1[4]
+ cb_7_6/io_i_6_in1[5] cb_7_6/io_i_6_in1[6] cb_7_6/io_i_6_in1[7] cb_7_6/io_i_7_ci
+ cb_7_6/io_i_7_in1[0] cb_7_6/io_i_7_in1[1] cb_7_6/io_i_7_in1[2] cb_7_6/io_i_7_in1[3]
+ cb_7_6/io_i_7_in1[4] cb_7_6/io_i_7_in1[5] cb_7_6/io_i_7_in1[6] cb_7_6/io_i_7_in1[7]
+ cb_7_7/io_i_0_ci cb_7_7/io_i_0_in1[0] cb_7_7/io_i_0_in1[1] cb_7_7/io_i_0_in1[2]
+ cb_7_7/io_i_0_in1[3] cb_7_7/io_i_0_in1[4] cb_7_7/io_i_0_in1[5] cb_7_7/io_i_0_in1[6]
+ cb_7_7/io_i_0_in1[7] cb_7_7/io_i_1_ci cb_7_7/io_i_1_in1[0] cb_7_7/io_i_1_in1[1]
+ cb_7_7/io_i_1_in1[2] cb_7_7/io_i_1_in1[3] cb_7_7/io_i_1_in1[4] cb_7_7/io_i_1_in1[5]
+ cb_7_7/io_i_1_in1[6] cb_7_7/io_i_1_in1[7] cb_7_7/io_i_2_ci cb_7_7/io_i_2_in1[0]
+ cb_7_7/io_i_2_in1[1] cb_7_7/io_i_2_in1[2] cb_7_7/io_i_2_in1[3] cb_7_7/io_i_2_in1[4]
+ cb_7_7/io_i_2_in1[5] cb_7_7/io_i_2_in1[6] cb_7_7/io_i_2_in1[7] cb_7_7/io_i_3_ci
+ cb_7_7/io_i_3_in1[0] cb_7_7/io_i_3_in1[1] cb_7_7/io_i_3_in1[2] cb_7_7/io_i_3_in1[3]
+ cb_7_7/io_i_3_in1[4] cb_7_7/io_i_3_in1[5] cb_7_7/io_i_3_in1[6] cb_7_7/io_i_3_in1[7]
+ cb_7_7/io_i_4_ci cb_7_7/io_i_4_in1[0] cb_7_7/io_i_4_in1[1] cb_7_7/io_i_4_in1[2]
+ cb_7_7/io_i_4_in1[3] cb_7_7/io_i_4_in1[4] cb_7_7/io_i_4_in1[5] cb_7_7/io_i_4_in1[6]
+ cb_7_7/io_i_4_in1[7] cb_7_7/io_i_5_ci cb_7_7/io_i_5_in1[0] cb_7_7/io_i_5_in1[1]
+ cb_7_7/io_i_5_in1[2] cb_7_7/io_i_5_in1[3] cb_7_7/io_i_5_in1[4] cb_7_7/io_i_5_in1[5]
+ cb_7_7/io_i_5_in1[6] cb_7_7/io_i_5_in1[7] cb_7_7/io_i_6_ci cb_7_7/io_i_6_in1[0]
+ cb_7_7/io_i_6_in1[1] cb_7_7/io_i_6_in1[2] cb_7_7/io_i_6_in1[3] cb_7_7/io_i_6_in1[4]
+ cb_7_7/io_i_6_in1[5] cb_7_7/io_i_6_in1[6] cb_7_7/io_i_6_in1[7] cb_7_7/io_i_7_ci
+ cb_7_7/io_i_7_in1[0] cb_7_7/io_i_7_in1[1] cb_7_7/io_i_7_in1[2] cb_7_7/io_i_7_in1[3]
+ cb_7_7/io_i_7_in1[4] cb_7_7/io_i_7_in1[5] cb_7_7/io_i_7_in1[6] cb_7_7/io_i_7_in1[7]
+ cb_7_6/io_vci cb_7_7/io_vci cb_7_6/io_vi cb_7_9/io_we_i cb_7_6/io_wo[0] cb_7_6/io_wo[10]
+ cb_7_6/io_wo[11] cb_7_6/io_wo[12] cb_7_6/io_wo[13] cb_7_6/io_wo[14] cb_7_6/io_wo[15]
+ cb_7_6/io_wo[16] cb_7_6/io_wo[17] cb_7_6/io_wo[18] cb_7_6/io_wo[19] cb_7_6/io_wo[1]
+ cb_7_6/io_wo[20] cb_7_6/io_wo[21] cb_7_6/io_wo[22] cb_7_6/io_wo[23] cb_7_6/io_wo[24]
+ cb_7_6/io_wo[25] cb_7_6/io_wo[26] cb_7_6/io_wo[27] cb_7_6/io_wo[28] cb_7_6/io_wo[29]
+ cb_7_6/io_wo[2] cb_7_6/io_wo[30] cb_7_6/io_wo[31] cb_7_6/io_wo[32] cb_7_6/io_wo[33]
+ cb_7_6/io_wo[34] cb_7_6/io_wo[35] cb_7_6/io_wo[36] cb_7_6/io_wo[37] cb_7_6/io_wo[38]
+ cb_7_6/io_wo[39] cb_7_6/io_wo[3] cb_7_6/io_wo[40] cb_7_6/io_wo[41] cb_7_6/io_wo[42]
+ cb_7_6/io_wo[43] cb_7_6/io_wo[44] cb_7_6/io_wo[45] cb_7_6/io_wo[46] cb_7_6/io_wo[47]
+ cb_7_6/io_wo[48] cb_7_6/io_wo[49] cb_7_6/io_wo[4] cb_7_6/io_wo[50] cb_7_6/io_wo[51]
+ cb_7_6/io_wo[52] cb_7_6/io_wo[53] cb_7_6/io_wo[54] cb_7_6/io_wo[55] cb_7_6/io_wo[56]
+ cb_7_6/io_wo[57] cb_7_6/io_wo[58] cb_7_6/io_wo[59] cb_7_6/io_wo[5] cb_7_6/io_wo[60]
+ cb_7_6/io_wo[61] cb_7_6/io_wo[62] cb_7_6/io_wo[63] cb_7_6/io_wo[6] cb_7_6/io_wo[7]
+ cb_7_6/io_wo[8] cb_7_6/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_5_3 cb_5_9/io_adr_i[0] cb_5_9/io_adr_i[1] cb_5_3/io_cs_i cb_5_9/io_dat_i[0] cb_5_9/io_dat_i[10]
+ cb_5_9/io_dat_i[11] cb_5_9/io_dat_i[12] cb_5_9/io_dat_i[13] cb_5_9/io_dat_i[14]
+ cb_5_9/io_dat_i[15] cb_5_9/io_dat_i[1] cb_5_9/io_dat_i[2] cb_5_9/io_dat_i[3] cb_5_9/io_dat_i[4]
+ cb_5_9/io_dat_i[5] cb_5_9/io_dat_i[6] cb_5_9/io_dat_i[7] cb_5_9/io_dat_i[8] cb_5_9/io_dat_i[9]
+ cb_5_3/io_dat_o[0] cb_5_3/io_dat_o[10] cb_5_3/io_dat_o[11] cb_5_3/io_dat_o[12] cb_5_3/io_dat_o[13]
+ cb_5_3/io_dat_o[14] cb_5_3/io_dat_o[15] cb_5_3/io_dat_o[1] cb_5_3/io_dat_o[2] cb_5_3/io_dat_o[3]
+ cb_5_3/io_dat_o[4] cb_5_3/io_dat_o[5] cb_5_3/io_dat_o[6] cb_5_3/io_dat_o[7] cb_5_3/io_dat_o[8]
+ cb_5_3/io_dat_o[9] cb_5_4/io_wo[0] cb_5_4/io_wo[10] cb_5_4/io_wo[11] cb_5_4/io_wo[12]
+ cb_5_4/io_wo[13] cb_5_4/io_wo[14] cb_5_4/io_wo[15] cb_5_4/io_wo[16] cb_5_4/io_wo[17]
+ cb_5_4/io_wo[18] cb_5_4/io_wo[19] cb_5_4/io_wo[1] cb_5_4/io_wo[20] cb_5_4/io_wo[21]
+ cb_5_4/io_wo[22] cb_5_4/io_wo[23] cb_5_4/io_wo[24] cb_5_4/io_wo[25] cb_5_4/io_wo[26]
+ cb_5_4/io_wo[27] cb_5_4/io_wo[28] cb_5_4/io_wo[29] cb_5_4/io_wo[2] cb_5_4/io_wo[30]
+ cb_5_4/io_wo[31] cb_5_4/io_wo[32] cb_5_4/io_wo[33] cb_5_4/io_wo[34] cb_5_4/io_wo[35]
+ cb_5_4/io_wo[36] cb_5_4/io_wo[37] cb_5_4/io_wo[38] cb_5_4/io_wo[39] cb_5_4/io_wo[3]
+ cb_5_4/io_wo[40] cb_5_4/io_wo[41] cb_5_4/io_wo[42] cb_5_4/io_wo[43] cb_5_4/io_wo[44]
+ cb_5_4/io_wo[45] cb_5_4/io_wo[46] cb_5_4/io_wo[47] cb_5_4/io_wo[48] cb_5_4/io_wo[49]
+ cb_5_4/io_wo[4] cb_5_4/io_wo[50] cb_5_4/io_wo[51] cb_5_4/io_wo[52] cb_5_4/io_wo[53]
+ cb_5_4/io_wo[54] cb_5_4/io_wo[55] cb_5_4/io_wo[56] cb_5_4/io_wo[57] cb_5_4/io_wo[58]
+ cb_5_4/io_wo[59] cb_5_4/io_wo[5] cb_5_4/io_wo[60] cb_5_4/io_wo[61] cb_5_4/io_wo[62]
+ cb_5_4/io_wo[63] cb_5_4/io_wo[6] cb_5_4/io_wo[7] cb_5_4/io_wo[8] cb_5_4/io_wo[9]
+ cb_5_3/io_i_0_ci cb_5_3/io_i_0_in1[0] cb_5_3/io_i_0_in1[1] cb_5_3/io_i_0_in1[2]
+ cb_5_3/io_i_0_in1[3] cb_5_3/io_i_0_in1[4] cb_5_3/io_i_0_in1[5] cb_5_3/io_i_0_in1[6]
+ cb_5_3/io_i_0_in1[7] cb_5_3/io_i_1_ci cb_5_3/io_i_1_in1[0] cb_5_3/io_i_1_in1[1]
+ cb_5_3/io_i_1_in1[2] cb_5_3/io_i_1_in1[3] cb_5_3/io_i_1_in1[4] cb_5_3/io_i_1_in1[5]
+ cb_5_3/io_i_1_in1[6] cb_5_3/io_i_1_in1[7] cb_5_3/io_i_2_ci cb_5_3/io_i_2_in1[0]
+ cb_5_3/io_i_2_in1[1] cb_5_3/io_i_2_in1[2] cb_5_3/io_i_2_in1[3] cb_5_3/io_i_2_in1[4]
+ cb_5_3/io_i_2_in1[5] cb_5_3/io_i_2_in1[6] cb_5_3/io_i_2_in1[7] cb_5_3/io_i_3_ci
+ cb_5_3/io_i_3_in1[0] cb_5_3/io_i_3_in1[1] cb_5_3/io_i_3_in1[2] cb_5_3/io_i_3_in1[3]
+ cb_5_3/io_i_3_in1[4] cb_5_3/io_i_3_in1[5] cb_5_3/io_i_3_in1[6] cb_5_3/io_i_3_in1[7]
+ cb_5_3/io_i_4_ci cb_5_3/io_i_4_in1[0] cb_5_3/io_i_4_in1[1] cb_5_3/io_i_4_in1[2]
+ cb_5_3/io_i_4_in1[3] cb_5_3/io_i_4_in1[4] cb_5_3/io_i_4_in1[5] cb_5_3/io_i_4_in1[6]
+ cb_5_3/io_i_4_in1[7] cb_5_3/io_i_5_ci cb_5_3/io_i_5_in1[0] cb_5_3/io_i_5_in1[1]
+ cb_5_3/io_i_5_in1[2] cb_5_3/io_i_5_in1[3] cb_5_3/io_i_5_in1[4] cb_5_3/io_i_5_in1[5]
+ cb_5_3/io_i_5_in1[6] cb_5_3/io_i_5_in1[7] cb_5_3/io_i_6_ci cb_5_3/io_i_6_in1[0]
+ cb_5_3/io_i_6_in1[1] cb_5_3/io_i_6_in1[2] cb_5_3/io_i_6_in1[3] cb_5_3/io_i_6_in1[4]
+ cb_5_3/io_i_6_in1[5] cb_5_3/io_i_6_in1[6] cb_5_3/io_i_6_in1[7] cb_5_3/io_i_7_ci
+ cb_5_3/io_i_7_in1[0] cb_5_3/io_i_7_in1[1] cb_5_3/io_i_7_in1[2] cb_5_3/io_i_7_in1[3]
+ cb_5_3/io_i_7_in1[4] cb_5_3/io_i_7_in1[5] cb_5_3/io_i_7_in1[6] cb_5_3/io_i_7_in1[7]
+ cb_5_4/io_i_0_ci cb_5_4/io_i_0_in1[0] cb_5_4/io_i_0_in1[1] cb_5_4/io_i_0_in1[2]
+ cb_5_4/io_i_0_in1[3] cb_5_4/io_i_0_in1[4] cb_5_4/io_i_0_in1[5] cb_5_4/io_i_0_in1[6]
+ cb_5_4/io_i_0_in1[7] cb_5_4/io_i_1_ci cb_5_4/io_i_1_in1[0] cb_5_4/io_i_1_in1[1]
+ cb_5_4/io_i_1_in1[2] cb_5_4/io_i_1_in1[3] cb_5_4/io_i_1_in1[4] cb_5_4/io_i_1_in1[5]
+ cb_5_4/io_i_1_in1[6] cb_5_4/io_i_1_in1[7] cb_5_4/io_i_2_ci cb_5_4/io_i_2_in1[0]
+ cb_5_4/io_i_2_in1[1] cb_5_4/io_i_2_in1[2] cb_5_4/io_i_2_in1[3] cb_5_4/io_i_2_in1[4]
+ cb_5_4/io_i_2_in1[5] cb_5_4/io_i_2_in1[6] cb_5_4/io_i_2_in1[7] cb_5_4/io_i_3_ci
+ cb_5_4/io_i_3_in1[0] cb_5_4/io_i_3_in1[1] cb_5_4/io_i_3_in1[2] cb_5_4/io_i_3_in1[3]
+ cb_5_4/io_i_3_in1[4] cb_5_4/io_i_3_in1[5] cb_5_4/io_i_3_in1[6] cb_5_4/io_i_3_in1[7]
+ cb_5_4/io_i_4_ci cb_5_4/io_i_4_in1[0] cb_5_4/io_i_4_in1[1] cb_5_4/io_i_4_in1[2]
+ cb_5_4/io_i_4_in1[3] cb_5_4/io_i_4_in1[4] cb_5_4/io_i_4_in1[5] cb_5_4/io_i_4_in1[6]
+ cb_5_4/io_i_4_in1[7] cb_5_4/io_i_5_ci cb_5_4/io_i_5_in1[0] cb_5_4/io_i_5_in1[1]
+ cb_5_4/io_i_5_in1[2] cb_5_4/io_i_5_in1[3] cb_5_4/io_i_5_in1[4] cb_5_4/io_i_5_in1[5]
+ cb_5_4/io_i_5_in1[6] cb_5_4/io_i_5_in1[7] cb_5_4/io_i_6_ci cb_5_4/io_i_6_in1[0]
+ cb_5_4/io_i_6_in1[1] cb_5_4/io_i_6_in1[2] cb_5_4/io_i_6_in1[3] cb_5_4/io_i_6_in1[4]
+ cb_5_4/io_i_6_in1[5] cb_5_4/io_i_6_in1[6] cb_5_4/io_i_6_in1[7] cb_5_4/io_i_7_ci
+ cb_5_4/io_i_7_in1[0] cb_5_4/io_i_7_in1[1] cb_5_4/io_i_7_in1[2] cb_5_4/io_i_7_in1[3]
+ cb_5_4/io_i_7_in1[4] cb_5_4/io_i_7_in1[5] cb_5_4/io_i_7_in1[6] cb_5_4/io_i_7_in1[7]
+ cb_5_3/io_vci cb_5_4/io_vci cb_5_3/io_vi cb_5_9/io_we_i cb_5_3/io_wo[0] cb_5_3/io_wo[10]
+ cb_5_3/io_wo[11] cb_5_3/io_wo[12] cb_5_3/io_wo[13] cb_5_3/io_wo[14] cb_5_3/io_wo[15]
+ cb_5_3/io_wo[16] cb_5_3/io_wo[17] cb_5_3/io_wo[18] cb_5_3/io_wo[19] cb_5_3/io_wo[1]
+ cb_5_3/io_wo[20] cb_5_3/io_wo[21] cb_5_3/io_wo[22] cb_5_3/io_wo[23] cb_5_3/io_wo[24]
+ cb_5_3/io_wo[25] cb_5_3/io_wo[26] cb_5_3/io_wo[27] cb_5_3/io_wo[28] cb_5_3/io_wo[29]
+ cb_5_3/io_wo[2] cb_5_3/io_wo[30] cb_5_3/io_wo[31] cb_5_3/io_wo[32] cb_5_3/io_wo[33]
+ cb_5_3/io_wo[34] cb_5_3/io_wo[35] cb_5_3/io_wo[36] cb_5_3/io_wo[37] cb_5_3/io_wo[38]
+ cb_5_3/io_wo[39] cb_5_3/io_wo[3] cb_5_3/io_wo[40] cb_5_3/io_wo[41] cb_5_3/io_wo[42]
+ cb_5_3/io_wo[43] cb_5_3/io_wo[44] cb_5_3/io_wo[45] cb_5_3/io_wo[46] cb_5_3/io_wo[47]
+ cb_5_3/io_wo[48] cb_5_3/io_wo[49] cb_5_3/io_wo[4] cb_5_3/io_wo[50] cb_5_3/io_wo[51]
+ cb_5_3/io_wo[52] cb_5_3/io_wo[53] cb_5_3/io_wo[54] cb_5_3/io_wo[55] cb_5_3/io_wo[56]
+ cb_5_3/io_wo[57] cb_5_3/io_wo[58] cb_5_3/io_wo[59] cb_5_3/io_wo[5] cb_5_3/io_wo[60]
+ cb_5_3/io_wo[61] cb_5_3/io_wo[62] cb_5_3/io_wo[63] cb_5_3/io_wo[6] cb_5_3/io_wo[7]
+ cb_5_3/io_wo[8] cb_5_3/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_3_0 cb_3_9/io_adr_i[0] cb_3_9/io_adr_i[1] cb_3_0/io_cs_i cb_3_9/io_dat_i[0] cb_3_9/io_dat_i[10]
+ cb_3_9/io_dat_i[11] cb_3_9/io_dat_i[12] cb_3_9/io_dat_i[13] cb_3_9/io_dat_i[14]
+ cb_3_9/io_dat_i[15] cb_3_9/io_dat_i[1] cb_3_9/io_dat_i[2] cb_3_9/io_dat_i[3] cb_3_9/io_dat_i[4]
+ cb_3_9/io_dat_i[5] cb_3_9/io_dat_i[6] cb_3_9/io_dat_i[7] cb_3_9/io_dat_i[8] cb_3_9/io_dat_i[9]
+ cb_3_0/io_dat_o[0] cb_3_0/io_dat_o[10] cb_3_0/io_dat_o[11] cb_3_0/io_dat_o[12] cb_3_0/io_dat_o[13]
+ cb_3_0/io_dat_o[14] cb_3_0/io_dat_o[15] cb_3_0/io_dat_o[1] cb_3_0/io_dat_o[2] cb_3_0/io_dat_o[3]
+ cb_3_0/io_dat_o[4] cb_3_0/io_dat_o[5] cb_3_0/io_dat_o[6] cb_3_0/io_dat_o[7] cb_3_0/io_dat_o[8]
+ cb_3_0/io_dat_o[9] cb_3_1/io_wo[0] cb_3_1/io_wo[10] cb_3_1/io_wo[11] cb_3_1/io_wo[12]
+ cb_3_1/io_wo[13] cb_3_1/io_wo[14] cb_3_1/io_wo[15] cb_3_1/io_wo[16] cb_3_1/io_wo[17]
+ cb_3_1/io_wo[18] cb_3_1/io_wo[19] cb_3_1/io_wo[1] cb_3_1/io_wo[20] cb_3_1/io_wo[21]
+ cb_3_1/io_wo[22] cb_3_1/io_wo[23] cb_3_1/io_wo[24] cb_3_1/io_wo[25] cb_3_1/io_wo[26]
+ cb_3_1/io_wo[27] cb_3_1/io_wo[28] cb_3_1/io_wo[29] cb_3_1/io_wo[2] cb_3_1/io_wo[30]
+ cb_3_1/io_wo[31] cb_3_1/io_wo[32] cb_3_1/io_wo[33] cb_3_1/io_wo[34] cb_3_1/io_wo[35]
+ cb_3_1/io_wo[36] cb_3_1/io_wo[37] cb_3_1/io_wo[38] cb_3_1/io_wo[39] cb_3_1/io_wo[3]
+ cb_3_1/io_wo[40] cb_3_1/io_wo[41] cb_3_1/io_wo[42] cb_3_1/io_wo[43] cb_3_1/io_wo[44]
+ cb_3_1/io_wo[45] cb_3_1/io_wo[46] cb_3_1/io_wo[47] cb_3_1/io_wo[48] cb_3_1/io_wo[49]
+ cb_3_1/io_wo[4] cb_3_1/io_wo[50] cb_3_1/io_wo[51] cb_3_1/io_wo[52] cb_3_1/io_wo[53]
+ cb_3_1/io_wo[54] cb_3_1/io_wo[55] cb_3_1/io_wo[56] cb_3_1/io_wo[57] cb_3_1/io_wo[58]
+ cb_3_1/io_wo[59] cb_3_1/io_wo[5] cb_3_1/io_wo[60] cb_3_1/io_wo[61] cb_3_1/io_wo[62]
+ cb_3_1/io_wo[63] cb_3_1/io_wo[6] cb_3_1/io_wo[7] cb_3_1/io_wo[8] cb_3_1/io_wo[9]
+ ccon_3/io_dsi_o cb_3_0/io_i_0_in1[0] cb_3_0/io_i_0_in1[1] cb_3_0/io_i_0_in1[2] cb_3_0/io_i_0_in1[3]
+ cb_3_0/io_i_0_in1[4] cb_3_0/io_i_0_in1[5] cb_3_0/io_i_0_in1[6] cb_3_0/io_i_0_in1[7]
+ cb_3_0/io_i_1_ci cb_3_0/io_i_1_in1[0] cb_3_0/io_i_1_in1[1] cb_3_0/io_i_1_in1[2]
+ cb_3_0/io_i_1_in1[3] cb_3_0/io_i_1_in1[4] cb_3_0/io_i_1_in1[5] cb_3_0/io_i_1_in1[6]
+ cb_3_0/io_i_1_in1[7] cb_3_0/io_i_2_ci cb_3_0/io_i_2_in1[0] cb_3_0/io_i_2_in1[1]
+ cb_3_0/io_i_2_in1[2] cb_3_0/io_i_2_in1[3] cb_3_0/io_i_2_in1[4] cb_3_0/io_i_2_in1[5]
+ cb_3_0/io_i_2_in1[6] cb_3_0/io_i_2_in1[7] cb_3_0/io_i_3_ci cb_3_0/io_i_3_in1[0]
+ cb_3_0/io_i_3_in1[1] cb_3_0/io_i_3_in1[2] cb_3_0/io_i_3_in1[3] cb_3_0/io_i_3_in1[4]
+ cb_3_0/io_i_3_in1[5] cb_3_0/io_i_3_in1[6] cb_3_0/io_i_3_in1[7] cb_3_0/io_i_4_ci
+ cb_3_0/io_i_4_in1[0] cb_3_0/io_i_4_in1[1] cb_3_0/io_i_4_in1[2] cb_3_0/io_i_4_in1[3]
+ cb_3_0/io_i_4_in1[4] cb_3_0/io_i_4_in1[5] cb_3_0/io_i_4_in1[6] cb_3_0/io_i_4_in1[7]
+ cb_3_0/io_i_5_ci cb_3_0/io_i_5_in1[0] cb_3_0/io_i_5_in1[1] cb_3_0/io_i_5_in1[2]
+ cb_3_0/io_i_5_in1[3] cb_3_0/io_i_5_in1[4] cb_3_0/io_i_5_in1[5] cb_3_0/io_i_5_in1[6]
+ cb_3_0/io_i_5_in1[7] cb_3_0/io_i_6_ci cb_3_0/io_i_6_in1[0] cb_3_0/io_i_6_in1[1]
+ cb_3_0/io_i_6_in1[2] cb_3_0/io_i_6_in1[3] cb_3_0/io_i_6_in1[4] cb_3_0/io_i_6_in1[5]
+ cb_3_0/io_i_6_in1[6] cb_3_0/io_i_6_in1[7] cb_3_0/io_i_7_ci cb_3_0/io_i_7_in1[0]
+ cb_3_0/io_i_7_in1[1] cb_3_0/io_i_7_in1[2] cb_3_0/io_i_7_in1[3] cb_3_0/io_i_7_in1[4]
+ cb_3_0/io_i_7_in1[5] cb_3_0/io_i_7_in1[6] cb_3_0/io_i_7_in1[7] cb_3_1/io_i_0_ci
+ cb_3_1/io_i_0_in1[0] cb_3_1/io_i_0_in1[1] cb_3_1/io_i_0_in1[2] cb_3_1/io_i_0_in1[3]
+ cb_3_1/io_i_0_in1[4] cb_3_1/io_i_0_in1[5] cb_3_1/io_i_0_in1[6] cb_3_1/io_i_0_in1[7]
+ cb_3_1/io_i_1_ci cb_3_1/io_i_1_in1[0] cb_3_1/io_i_1_in1[1] cb_3_1/io_i_1_in1[2]
+ cb_3_1/io_i_1_in1[3] cb_3_1/io_i_1_in1[4] cb_3_1/io_i_1_in1[5] cb_3_1/io_i_1_in1[6]
+ cb_3_1/io_i_1_in1[7] cb_3_1/io_i_2_ci cb_3_1/io_i_2_in1[0] cb_3_1/io_i_2_in1[1]
+ cb_3_1/io_i_2_in1[2] cb_3_1/io_i_2_in1[3] cb_3_1/io_i_2_in1[4] cb_3_1/io_i_2_in1[5]
+ cb_3_1/io_i_2_in1[6] cb_3_1/io_i_2_in1[7] cb_3_1/io_i_3_ci cb_3_1/io_i_3_in1[0]
+ cb_3_1/io_i_3_in1[1] cb_3_1/io_i_3_in1[2] cb_3_1/io_i_3_in1[3] cb_3_1/io_i_3_in1[4]
+ cb_3_1/io_i_3_in1[5] cb_3_1/io_i_3_in1[6] cb_3_1/io_i_3_in1[7] cb_3_1/io_i_4_ci
+ cb_3_1/io_i_4_in1[0] cb_3_1/io_i_4_in1[1] cb_3_1/io_i_4_in1[2] cb_3_1/io_i_4_in1[3]
+ cb_3_1/io_i_4_in1[4] cb_3_1/io_i_4_in1[5] cb_3_1/io_i_4_in1[6] cb_3_1/io_i_4_in1[7]
+ cb_3_1/io_i_5_ci cb_3_1/io_i_5_in1[0] cb_3_1/io_i_5_in1[1] cb_3_1/io_i_5_in1[2]
+ cb_3_1/io_i_5_in1[3] cb_3_1/io_i_5_in1[4] cb_3_1/io_i_5_in1[5] cb_3_1/io_i_5_in1[6]
+ cb_3_1/io_i_5_in1[7] cb_3_1/io_i_6_ci cb_3_1/io_i_6_in1[0] cb_3_1/io_i_6_in1[1]
+ cb_3_1/io_i_6_in1[2] cb_3_1/io_i_6_in1[3] cb_3_1/io_i_6_in1[4] cb_3_1/io_i_6_in1[5]
+ cb_3_1/io_i_6_in1[6] cb_3_1/io_i_6_in1[7] cb_3_1/io_i_7_ci cb_3_1/io_i_7_in1[0]
+ cb_3_1/io_i_7_in1[1] cb_3_1/io_i_7_in1[2] cb_3_1/io_i_7_in1[3] cb_3_1/io_i_7_in1[4]
+ cb_3_1/io_i_7_in1[5] cb_3_1/io_i_7_in1[6] cb_3_1/io_i_7_in1[7] cb_3_0/io_vci cb_3_1/io_vci
+ cb_3_0/io_vi cb_3_9/io_we_i cb_3_0/io_wo[0] cb_3_0/io_wo[10] cb_3_0/io_wo[11] cb_3_0/io_wo[12]
+ cb_3_0/io_wo[13] cb_3_0/io_wo[14] cb_3_0/io_wo[15] cb_3_0/io_wo[16] cb_3_0/io_wo[17]
+ cb_3_0/io_wo[18] cb_3_0/io_wo[19] cb_3_0/io_wo[1] cb_3_0/io_wo[20] cb_3_0/io_wo[21]
+ cb_3_0/io_wo[22] cb_3_0/io_wo[23] cb_3_0/io_wo[24] cb_3_0/io_wo[25] cb_3_0/io_wo[26]
+ cb_3_0/io_wo[27] cb_3_0/io_wo[28] cb_3_0/io_wo[29] cb_3_0/io_wo[2] cb_3_0/io_wo[30]
+ cb_3_0/io_wo[31] cb_3_0/io_wo[32] cb_3_0/io_wo[33] cb_3_0/io_wo[34] cb_3_0/io_wo[35]
+ cb_3_0/io_wo[36] cb_3_0/io_wo[37] cb_3_0/io_wo[38] cb_3_0/io_wo[39] cb_3_0/io_wo[3]
+ cb_3_0/io_wo[40] cb_3_0/io_wo[41] cb_3_0/io_wo[42] cb_3_0/io_wo[43] cb_3_0/io_wo[44]
+ cb_3_0/io_wo[45] cb_3_0/io_wo[46] cb_3_0/io_wo[47] cb_3_0/io_wo[48] cb_3_0/io_wo[49]
+ cb_3_0/io_wo[4] cb_3_0/io_wo[50] cb_3_0/io_wo[51] cb_3_0/io_wo[52] cb_3_0/io_wo[53]
+ cb_3_0/io_wo[54] cb_3_0/io_wo[55] cb_3_0/io_wo[56] cb_3_0/io_wo[57] cb_3_0/io_wo[58]
+ cb_3_0/io_wo[59] cb_3_0/io_wo[5] cb_3_0/io_wo[60] cb_3_0/io_wo[61] cb_3_0/io_wo[62]
+ cb_3_0/io_wo[63] cb_3_0/io_wo[6] cb_3_0/io_wo[7] cb_3_0/io_wo[8] cb_3_0/io_wo[9]
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_7_7 cb_7_9/io_adr_i[0] cb_7_9/io_adr_i[1] cb_7_7/io_cs_i cb_7_9/io_dat_i[0] cb_7_9/io_dat_i[10]
+ cb_7_9/io_dat_i[11] cb_7_9/io_dat_i[12] cb_7_9/io_dat_i[13] cb_7_9/io_dat_i[14]
+ cb_7_9/io_dat_i[15] cb_7_9/io_dat_i[1] cb_7_9/io_dat_i[2] cb_7_9/io_dat_i[3] cb_7_9/io_dat_i[4]
+ cb_7_9/io_dat_i[5] cb_7_9/io_dat_i[6] cb_7_9/io_dat_i[7] cb_7_9/io_dat_i[8] cb_7_9/io_dat_i[9]
+ cb_7_7/io_dat_o[0] cb_7_7/io_dat_o[10] cb_7_7/io_dat_o[11] cb_7_7/io_dat_o[12] cb_7_7/io_dat_o[13]
+ cb_7_7/io_dat_o[14] cb_7_7/io_dat_o[15] cb_7_7/io_dat_o[1] cb_7_7/io_dat_o[2] cb_7_7/io_dat_o[3]
+ cb_7_7/io_dat_o[4] cb_7_7/io_dat_o[5] cb_7_7/io_dat_o[6] cb_7_7/io_dat_o[7] cb_7_7/io_dat_o[8]
+ cb_7_7/io_dat_o[9] cb_7_8/io_wo[0] cb_7_8/io_wo[10] cb_7_8/io_wo[11] cb_7_8/io_wo[12]
+ cb_7_8/io_wo[13] cb_7_8/io_wo[14] cb_7_8/io_wo[15] cb_7_8/io_wo[16] cb_7_8/io_wo[17]
+ cb_7_8/io_wo[18] cb_7_8/io_wo[19] cb_7_8/io_wo[1] cb_7_8/io_wo[20] cb_7_8/io_wo[21]
+ cb_7_8/io_wo[22] cb_7_8/io_wo[23] cb_7_8/io_wo[24] cb_7_8/io_wo[25] cb_7_8/io_wo[26]
+ cb_7_8/io_wo[27] cb_7_8/io_wo[28] cb_7_8/io_wo[29] cb_7_8/io_wo[2] cb_7_8/io_wo[30]
+ cb_7_8/io_wo[31] cb_7_8/io_wo[32] cb_7_8/io_wo[33] cb_7_8/io_wo[34] cb_7_8/io_wo[35]
+ cb_7_8/io_wo[36] cb_7_8/io_wo[37] cb_7_8/io_wo[38] cb_7_8/io_wo[39] cb_7_8/io_wo[3]
+ cb_7_8/io_wo[40] cb_7_8/io_wo[41] cb_7_8/io_wo[42] cb_7_8/io_wo[43] cb_7_8/io_wo[44]
+ cb_7_8/io_wo[45] cb_7_8/io_wo[46] cb_7_8/io_wo[47] cb_7_8/io_wo[48] cb_7_8/io_wo[49]
+ cb_7_8/io_wo[4] cb_7_8/io_wo[50] cb_7_8/io_wo[51] cb_7_8/io_wo[52] cb_7_8/io_wo[53]
+ cb_7_8/io_wo[54] cb_7_8/io_wo[55] cb_7_8/io_wo[56] cb_7_8/io_wo[57] cb_7_8/io_wo[58]
+ cb_7_8/io_wo[59] cb_7_8/io_wo[5] cb_7_8/io_wo[60] cb_7_8/io_wo[61] cb_7_8/io_wo[62]
+ cb_7_8/io_wo[63] cb_7_8/io_wo[6] cb_7_8/io_wo[7] cb_7_8/io_wo[8] cb_7_8/io_wo[9]
+ cb_7_7/io_i_0_ci cb_7_7/io_i_0_in1[0] cb_7_7/io_i_0_in1[1] cb_7_7/io_i_0_in1[2]
+ cb_7_7/io_i_0_in1[3] cb_7_7/io_i_0_in1[4] cb_7_7/io_i_0_in1[5] cb_7_7/io_i_0_in1[6]
+ cb_7_7/io_i_0_in1[7] cb_7_7/io_i_1_ci cb_7_7/io_i_1_in1[0] cb_7_7/io_i_1_in1[1]
+ cb_7_7/io_i_1_in1[2] cb_7_7/io_i_1_in1[3] cb_7_7/io_i_1_in1[4] cb_7_7/io_i_1_in1[5]
+ cb_7_7/io_i_1_in1[6] cb_7_7/io_i_1_in1[7] cb_7_7/io_i_2_ci cb_7_7/io_i_2_in1[0]
+ cb_7_7/io_i_2_in1[1] cb_7_7/io_i_2_in1[2] cb_7_7/io_i_2_in1[3] cb_7_7/io_i_2_in1[4]
+ cb_7_7/io_i_2_in1[5] cb_7_7/io_i_2_in1[6] cb_7_7/io_i_2_in1[7] cb_7_7/io_i_3_ci
+ cb_7_7/io_i_3_in1[0] cb_7_7/io_i_3_in1[1] cb_7_7/io_i_3_in1[2] cb_7_7/io_i_3_in1[3]
+ cb_7_7/io_i_3_in1[4] cb_7_7/io_i_3_in1[5] cb_7_7/io_i_3_in1[6] cb_7_7/io_i_3_in1[7]
+ cb_7_7/io_i_4_ci cb_7_7/io_i_4_in1[0] cb_7_7/io_i_4_in1[1] cb_7_7/io_i_4_in1[2]
+ cb_7_7/io_i_4_in1[3] cb_7_7/io_i_4_in1[4] cb_7_7/io_i_4_in1[5] cb_7_7/io_i_4_in1[6]
+ cb_7_7/io_i_4_in1[7] cb_7_7/io_i_5_ci cb_7_7/io_i_5_in1[0] cb_7_7/io_i_5_in1[1]
+ cb_7_7/io_i_5_in1[2] cb_7_7/io_i_5_in1[3] cb_7_7/io_i_5_in1[4] cb_7_7/io_i_5_in1[5]
+ cb_7_7/io_i_5_in1[6] cb_7_7/io_i_5_in1[7] cb_7_7/io_i_6_ci cb_7_7/io_i_6_in1[0]
+ cb_7_7/io_i_6_in1[1] cb_7_7/io_i_6_in1[2] cb_7_7/io_i_6_in1[3] cb_7_7/io_i_6_in1[4]
+ cb_7_7/io_i_6_in1[5] cb_7_7/io_i_6_in1[6] cb_7_7/io_i_6_in1[7] cb_7_7/io_i_7_ci
+ cb_7_7/io_i_7_in1[0] cb_7_7/io_i_7_in1[1] cb_7_7/io_i_7_in1[2] cb_7_7/io_i_7_in1[3]
+ cb_7_7/io_i_7_in1[4] cb_7_7/io_i_7_in1[5] cb_7_7/io_i_7_in1[6] cb_7_7/io_i_7_in1[7]
+ cb_7_8/io_i_0_ci cb_7_8/io_i_0_in1[0] cb_7_8/io_i_0_in1[1] cb_7_8/io_i_0_in1[2]
+ cb_7_8/io_i_0_in1[3] cb_7_8/io_i_0_in1[4] cb_7_8/io_i_0_in1[5] cb_7_8/io_i_0_in1[6]
+ cb_7_8/io_i_0_in1[7] cb_7_8/io_i_1_ci cb_7_8/io_i_1_in1[0] cb_7_8/io_i_1_in1[1]
+ cb_7_8/io_i_1_in1[2] cb_7_8/io_i_1_in1[3] cb_7_8/io_i_1_in1[4] cb_7_8/io_i_1_in1[5]
+ cb_7_8/io_i_1_in1[6] cb_7_8/io_i_1_in1[7] cb_7_8/io_i_2_ci cb_7_8/io_i_2_in1[0]
+ cb_7_8/io_i_2_in1[1] cb_7_8/io_i_2_in1[2] cb_7_8/io_i_2_in1[3] cb_7_8/io_i_2_in1[4]
+ cb_7_8/io_i_2_in1[5] cb_7_8/io_i_2_in1[6] cb_7_8/io_i_2_in1[7] cb_7_8/io_i_3_ci
+ cb_7_8/io_i_3_in1[0] cb_7_8/io_i_3_in1[1] cb_7_8/io_i_3_in1[2] cb_7_8/io_i_3_in1[3]
+ cb_7_8/io_i_3_in1[4] cb_7_8/io_i_3_in1[5] cb_7_8/io_i_3_in1[6] cb_7_8/io_i_3_in1[7]
+ cb_7_8/io_i_4_ci cb_7_8/io_i_4_in1[0] cb_7_8/io_i_4_in1[1] cb_7_8/io_i_4_in1[2]
+ cb_7_8/io_i_4_in1[3] cb_7_8/io_i_4_in1[4] cb_7_8/io_i_4_in1[5] cb_7_8/io_i_4_in1[6]
+ cb_7_8/io_i_4_in1[7] cb_7_8/io_i_5_ci cb_7_8/io_i_5_in1[0] cb_7_8/io_i_5_in1[1]
+ cb_7_8/io_i_5_in1[2] cb_7_8/io_i_5_in1[3] cb_7_8/io_i_5_in1[4] cb_7_8/io_i_5_in1[5]
+ cb_7_8/io_i_5_in1[6] cb_7_8/io_i_5_in1[7] cb_7_8/io_i_6_ci cb_7_8/io_i_6_in1[0]
+ cb_7_8/io_i_6_in1[1] cb_7_8/io_i_6_in1[2] cb_7_8/io_i_6_in1[3] cb_7_8/io_i_6_in1[4]
+ cb_7_8/io_i_6_in1[5] cb_7_8/io_i_6_in1[6] cb_7_8/io_i_6_in1[7] cb_7_8/io_i_7_ci
+ cb_7_8/io_i_7_in1[0] cb_7_8/io_i_7_in1[1] cb_7_8/io_i_7_in1[2] cb_7_8/io_i_7_in1[3]
+ cb_7_8/io_i_7_in1[4] cb_7_8/io_i_7_in1[5] cb_7_8/io_i_7_in1[6] cb_7_8/io_i_7_in1[7]
+ cb_7_7/io_vci cb_7_8/io_vci cb_7_7/io_vi cb_7_9/io_we_i cb_7_7/io_wo[0] cb_7_7/io_wo[10]
+ cb_7_7/io_wo[11] cb_7_7/io_wo[12] cb_7_7/io_wo[13] cb_7_7/io_wo[14] cb_7_7/io_wo[15]
+ cb_7_7/io_wo[16] cb_7_7/io_wo[17] cb_7_7/io_wo[18] cb_7_7/io_wo[19] cb_7_7/io_wo[1]
+ cb_7_7/io_wo[20] cb_7_7/io_wo[21] cb_7_7/io_wo[22] cb_7_7/io_wo[23] cb_7_7/io_wo[24]
+ cb_7_7/io_wo[25] cb_7_7/io_wo[26] cb_7_7/io_wo[27] cb_7_7/io_wo[28] cb_7_7/io_wo[29]
+ cb_7_7/io_wo[2] cb_7_7/io_wo[30] cb_7_7/io_wo[31] cb_7_7/io_wo[32] cb_7_7/io_wo[33]
+ cb_7_7/io_wo[34] cb_7_7/io_wo[35] cb_7_7/io_wo[36] cb_7_7/io_wo[37] cb_7_7/io_wo[38]
+ cb_7_7/io_wo[39] cb_7_7/io_wo[3] cb_7_7/io_wo[40] cb_7_7/io_wo[41] cb_7_7/io_wo[42]
+ cb_7_7/io_wo[43] cb_7_7/io_wo[44] cb_7_7/io_wo[45] cb_7_7/io_wo[46] cb_7_7/io_wo[47]
+ cb_7_7/io_wo[48] cb_7_7/io_wo[49] cb_7_7/io_wo[4] cb_7_7/io_wo[50] cb_7_7/io_wo[51]
+ cb_7_7/io_wo[52] cb_7_7/io_wo[53] cb_7_7/io_wo[54] cb_7_7/io_wo[55] cb_7_7/io_wo[56]
+ cb_7_7/io_wo[57] cb_7_7/io_wo[58] cb_7_7/io_wo[59] cb_7_7/io_wo[5] cb_7_7/io_wo[60]
+ cb_7_7/io_wo[61] cb_7_7/io_wo[62] cb_7_7/io_wo[63] cb_7_7/io_wo[6] cb_7_7/io_wo[7]
+ cb_7_7/io_wo[8] cb_7_7/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_5_4 cb_5_9/io_adr_i[0] cb_5_9/io_adr_i[1] cb_5_4/io_cs_i cb_5_9/io_dat_i[0] cb_5_9/io_dat_i[10]
+ cb_5_9/io_dat_i[11] cb_5_9/io_dat_i[12] cb_5_9/io_dat_i[13] cb_5_9/io_dat_i[14]
+ cb_5_9/io_dat_i[15] cb_5_9/io_dat_i[1] cb_5_9/io_dat_i[2] cb_5_9/io_dat_i[3] cb_5_9/io_dat_i[4]
+ cb_5_9/io_dat_i[5] cb_5_9/io_dat_i[6] cb_5_9/io_dat_i[7] cb_5_9/io_dat_i[8] cb_5_9/io_dat_i[9]
+ cb_5_4/io_dat_o[0] cb_5_4/io_dat_o[10] cb_5_4/io_dat_o[11] cb_5_4/io_dat_o[12] cb_5_4/io_dat_o[13]
+ cb_5_4/io_dat_o[14] cb_5_4/io_dat_o[15] cb_5_4/io_dat_o[1] cb_5_4/io_dat_o[2] cb_5_4/io_dat_o[3]
+ cb_5_4/io_dat_o[4] cb_5_4/io_dat_o[5] cb_5_4/io_dat_o[6] cb_5_4/io_dat_o[7] cb_5_4/io_dat_o[8]
+ cb_5_4/io_dat_o[9] cb_5_5/io_wo[0] cb_5_5/io_wo[10] cb_5_5/io_wo[11] cb_5_5/io_wo[12]
+ cb_5_5/io_wo[13] cb_5_5/io_wo[14] cb_5_5/io_wo[15] cb_5_5/io_wo[16] cb_5_5/io_wo[17]
+ cb_5_5/io_wo[18] cb_5_5/io_wo[19] cb_5_5/io_wo[1] cb_5_5/io_wo[20] cb_5_5/io_wo[21]
+ cb_5_5/io_wo[22] cb_5_5/io_wo[23] cb_5_5/io_wo[24] cb_5_5/io_wo[25] cb_5_5/io_wo[26]
+ cb_5_5/io_wo[27] cb_5_5/io_wo[28] cb_5_5/io_wo[29] cb_5_5/io_wo[2] cb_5_5/io_wo[30]
+ cb_5_5/io_wo[31] cb_5_5/io_wo[32] cb_5_5/io_wo[33] cb_5_5/io_wo[34] cb_5_5/io_wo[35]
+ cb_5_5/io_wo[36] cb_5_5/io_wo[37] cb_5_5/io_wo[38] cb_5_5/io_wo[39] cb_5_5/io_wo[3]
+ cb_5_5/io_wo[40] cb_5_5/io_wo[41] cb_5_5/io_wo[42] cb_5_5/io_wo[43] cb_5_5/io_wo[44]
+ cb_5_5/io_wo[45] cb_5_5/io_wo[46] cb_5_5/io_wo[47] cb_5_5/io_wo[48] cb_5_5/io_wo[49]
+ cb_5_5/io_wo[4] cb_5_5/io_wo[50] cb_5_5/io_wo[51] cb_5_5/io_wo[52] cb_5_5/io_wo[53]
+ cb_5_5/io_wo[54] cb_5_5/io_wo[55] cb_5_5/io_wo[56] cb_5_5/io_wo[57] cb_5_5/io_wo[58]
+ cb_5_5/io_wo[59] cb_5_5/io_wo[5] cb_5_5/io_wo[60] cb_5_5/io_wo[61] cb_5_5/io_wo[62]
+ cb_5_5/io_wo[63] cb_5_5/io_wo[6] cb_5_5/io_wo[7] cb_5_5/io_wo[8] cb_5_5/io_wo[9]
+ cb_5_4/io_i_0_ci cb_5_4/io_i_0_in1[0] cb_5_4/io_i_0_in1[1] cb_5_4/io_i_0_in1[2]
+ cb_5_4/io_i_0_in1[3] cb_5_4/io_i_0_in1[4] cb_5_4/io_i_0_in1[5] cb_5_4/io_i_0_in1[6]
+ cb_5_4/io_i_0_in1[7] cb_5_4/io_i_1_ci cb_5_4/io_i_1_in1[0] cb_5_4/io_i_1_in1[1]
+ cb_5_4/io_i_1_in1[2] cb_5_4/io_i_1_in1[3] cb_5_4/io_i_1_in1[4] cb_5_4/io_i_1_in1[5]
+ cb_5_4/io_i_1_in1[6] cb_5_4/io_i_1_in1[7] cb_5_4/io_i_2_ci cb_5_4/io_i_2_in1[0]
+ cb_5_4/io_i_2_in1[1] cb_5_4/io_i_2_in1[2] cb_5_4/io_i_2_in1[3] cb_5_4/io_i_2_in1[4]
+ cb_5_4/io_i_2_in1[5] cb_5_4/io_i_2_in1[6] cb_5_4/io_i_2_in1[7] cb_5_4/io_i_3_ci
+ cb_5_4/io_i_3_in1[0] cb_5_4/io_i_3_in1[1] cb_5_4/io_i_3_in1[2] cb_5_4/io_i_3_in1[3]
+ cb_5_4/io_i_3_in1[4] cb_5_4/io_i_3_in1[5] cb_5_4/io_i_3_in1[6] cb_5_4/io_i_3_in1[7]
+ cb_5_4/io_i_4_ci cb_5_4/io_i_4_in1[0] cb_5_4/io_i_4_in1[1] cb_5_4/io_i_4_in1[2]
+ cb_5_4/io_i_4_in1[3] cb_5_4/io_i_4_in1[4] cb_5_4/io_i_4_in1[5] cb_5_4/io_i_4_in1[6]
+ cb_5_4/io_i_4_in1[7] cb_5_4/io_i_5_ci cb_5_4/io_i_5_in1[0] cb_5_4/io_i_5_in1[1]
+ cb_5_4/io_i_5_in1[2] cb_5_4/io_i_5_in1[3] cb_5_4/io_i_5_in1[4] cb_5_4/io_i_5_in1[5]
+ cb_5_4/io_i_5_in1[6] cb_5_4/io_i_5_in1[7] cb_5_4/io_i_6_ci cb_5_4/io_i_6_in1[0]
+ cb_5_4/io_i_6_in1[1] cb_5_4/io_i_6_in1[2] cb_5_4/io_i_6_in1[3] cb_5_4/io_i_6_in1[4]
+ cb_5_4/io_i_6_in1[5] cb_5_4/io_i_6_in1[6] cb_5_4/io_i_6_in1[7] cb_5_4/io_i_7_ci
+ cb_5_4/io_i_7_in1[0] cb_5_4/io_i_7_in1[1] cb_5_4/io_i_7_in1[2] cb_5_4/io_i_7_in1[3]
+ cb_5_4/io_i_7_in1[4] cb_5_4/io_i_7_in1[5] cb_5_4/io_i_7_in1[6] cb_5_4/io_i_7_in1[7]
+ cb_5_5/io_i_0_ci cb_5_5/io_i_0_in1[0] cb_5_5/io_i_0_in1[1] cb_5_5/io_i_0_in1[2]
+ cb_5_5/io_i_0_in1[3] cb_5_5/io_i_0_in1[4] cb_5_5/io_i_0_in1[5] cb_5_5/io_i_0_in1[6]
+ cb_5_5/io_i_0_in1[7] cb_5_5/io_i_1_ci cb_5_5/io_i_1_in1[0] cb_5_5/io_i_1_in1[1]
+ cb_5_5/io_i_1_in1[2] cb_5_5/io_i_1_in1[3] cb_5_5/io_i_1_in1[4] cb_5_5/io_i_1_in1[5]
+ cb_5_5/io_i_1_in1[6] cb_5_5/io_i_1_in1[7] cb_5_5/io_i_2_ci cb_5_5/io_i_2_in1[0]
+ cb_5_5/io_i_2_in1[1] cb_5_5/io_i_2_in1[2] cb_5_5/io_i_2_in1[3] cb_5_5/io_i_2_in1[4]
+ cb_5_5/io_i_2_in1[5] cb_5_5/io_i_2_in1[6] cb_5_5/io_i_2_in1[7] cb_5_5/io_i_3_ci
+ cb_5_5/io_i_3_in1[0] cb_5_5/io_i_3_in1[1] cb_5_5/io_i_3_in1[2] cb_5_5/io_i_3_in1[3]
+ cb_5_5/io_i_3_in1[4] cb_5_5/io_i_3_in1[5] cb_5_5/io_i_3_in1[6] cb_5_5/io_i_3_in1[7]
+ cb_5_5/io_i_4_ci cb_5_5/io_i_4_in1[0] cb_5_5/io_i_4_in1[1] cb_5_5/io_i_4_in1[2]
+ cb_5_5/io_i_4_in1[3] cb_5_5/io_i_4_in1[4] cb_5_5/io_i_4_in1[5] cb_5_5/io_i_4_in1[6]
+ cb_5_5/io_i_4_in1[7] cb_5_5/io_i_5_ci cb_5_5/io_i_5_in1[0] cb_5_5/io_i_5_in1[1]
+ cb_5_5/io_i_5_in1[2] cb_5_5/io_i_5_in1[3] cb_5_5/io_i_5_in1[4] cb_5_5/io_i_5_in1[5]
+ cb_5_5/io_i_5_in1[6] cb_5_5/io_i_5_in1[7] cb_5_5/io_i_6_ci cb_5_5/io_i_6_in1[0]
+ cb_5_5/io_i_6_in1[1] cb_5_5/io_i_6_in1[2] cb_5_5/io_i_6_in1[3] cb_5_5/io_i_6_in1[4]
+ cb_5_5/io_i_6_in1[5] cb_5_5/io_i_6_in1[6] cb_5_5/io_i_6_in1[7] cb_5_5/io_i_7_ci
+ cb_5_5/io_i_7_in1[0] cb_5_5/io_i_7_in1[1] cb_5_5/io_i_7_in1[2] cb_5_5/io_i_7_in1[3]
+ cb_5_5/io_i_7_in1[4] cb_5_5/io_i_7_in1[5] cb_5_5/io_i_7_in1[6] cb_5_5/io_i_7_in1[7]
+ cb_5_4/io_vci cb_5_5/io_vci cb_5_4/io_vi cb_5_9/io_we_i cb_5_4/io_wo[0] cb_5_4/io_wo[10]
+ cb_5_4/io_wo[11] cb_5_4/io_wo[12] cb_5_4/io_wo[13] cb_5_4/io_wo[14] cb_5_4/io_wo[15]
+ cb_5_4/io_wo[16] cb_5_4/io_wo[17] cb_5_4/io_wo[18] cb_5_4/io_wo[19] cb_5_4/io_wo[1]
+ cb_5_4/io_wo[20] cb_5_4/io_wo[21] cb_5_4/io_wo[22] cb_5_4/io_wo[23] cb_5_4/io_wo[24]
+ cb_5_4/io_wo[25] cb_5_4/io_wo[26] cb_5_4/io_wo[27] cb_5_4/io_wo[28] cb_5_4/io_wo[29]
+ cb_5_4/io_wo[2] cb_5_4/io_wo[30] cb_5_4/io_wo[31] cb_5_4/io_wo[32] cb_5_4/io_wo[33]
+ cb_5_4/io_wo[34] cb_5_4/io_wo[35] cb_5_4/io_wo[36] cb_5_4/io_wo[37] cb_5_4/io_wo[38]
+ cb_5_4/io_wo[39] cb_5_4/io_wo[3] cb_5_4/io_wo[40] cb_5_4/io_wo[41] cb_5_4/io_wo[42]
+ cb_5_4/io_wo[43] cb_5_4/io_wo[44] cb_5_4/io_wo[45] cb_5_4/io_wo[46] cb_5_4/io_wo[47]
+ cb_5_4/io_wo[48] cb_5_4/io_wo[49] cb_5_4/io_wo[4] cb_5_4/io_wo[50] cb_5_4/io_wo[51]
+ cb_5_4/io_wo[52] cb_5_4/io_wo[53] cb_5_4/io_wo[54] cb_5_4/io_wo[55] cb_5_4/io_wo[56]
+ cb_5_4/io_wo[57] cb_5_4/io_wo[58] cb_5_4/io_wo[59] cb_5_4/io_wo[5] cb_5_4/io_wo[60]
+ cb_5_4/io_wo[61] cb_5_4/io_wo[62] cb_5_4/io_wo[63] cb_5_4/io_wo[6] cb_5_4/io_wo[7]
+ cb_5_4/io_wo[8] cb_5_4/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xccon_0 ccon_0/io_ack_o ccon_7/io_adr_i[0] ccon_7/io_adr_i[10] ccon_7/io_adr_i[11]
+ ccon_7/io_adr_i[1] ccon_7/io_adr_i[2] ccon_7/io_adr_i[3] ccon_7/io_adr_i[4] ccon_7/io_adr_i[5]
+ ccon_7/io_adr_i[6] ccon_7/io_adr_i[7] ccon_7/io_adr_i[8] ccon_7/io_adr_i[9] cb_0_9/io_adr_i[0]
+ cb_0_9/io_adr_i[1] cb_0_0/io_cs_i cb_0_1/io_cs_i cb_0_10/io_cs_i cb_0_2/io_cs_i
+ cb_0_3/io_cs_i cb_0_4/io_cs_i cb_0_5/io_cs_i cb_0_6/io_cs_i cb_0_7/io_cs_i cb_0_8/io_cs_i
+ cb_0_9/io_cs_i cb_0_9/io_dat_i[0] cb_0_9/io_dat_i[10] cb_0_9/io_dat_i[11] cb_0_9/io_dat_i[12]
+ cb_0_9/io_dat_i[13] cb_0_9/io_dat_i[14] cb_0_9/io_dat_i[15] cb_0_9/io_dat_i[1] cb_0_9/io_dat_i[2]
+ cb_0_9/io_dat_i[3] cb_0_9/io_dat_i[4] cb_0_9/io_dat_i[5] cb_0_9/io_dat_i[6] cb_0_9/io_dat_i[7]
+ cb_0_9/io_dat_i[8] cb_0_9/io_dat_i[9] cb_0_0/io_dat_o[0] cb_0_0/io_dat_o[10] cb_0_0/io_dat_o[11]
+ cb_0_0/io_dat_o[12] cb_0_0/io_dat_o[13] cb_0_0/io_dat_o[14] cb_0_0/io_dat_o[15]
+ cb_0_0/io_dat_o[1] cb_0_0/io_dat_o[2] cb_0_0/io_dat_o[3] cb_0_0/io_dat_o[4] cb_0_0/io_dat_o[5]
+ cb_0_0/io_dat_o[6] cb_0_0/io_dat_o[7] cb_0_0/io_dat_o[8] cb_0_0/io_dat_o[9] cb_0_10/io_dat_o[0]
+ cb_0_10/io_dat_o[10] cb_0_10/io_dat_o[11] cb_0_10/io_dat_o[12] cb_0_10/io_dat_o[13]
+ cb_0_10/io_dat_o[14] cb_0_10/io_dat_o[15] cb_0_10/io_dat_o[1] cb_0_10/io_dat_o[2]
+ cb_0_10/io_dat_o[3] cb_0_10/io_dat_o[4] cb_0_10/io_dat_o[5] cb_0_10/io_dat_o[6]
+ cb_0_10/io_dat_o[7] cb_0_10/io_dat_o[8] cb_0_10/io_dat_o[9] cb_0_1/io_dat_o[0] cb_0_1/io_dat_o[10]
+ cb_0_1/io_dat_o[11] cb_0_1/io_dat_o[12] cb_0_1/io_dat_o[13] cb_0_1/io_dat_o[14]
+ cb_0_1/io_dat_o[15] cb_0_1/io_dat_o[1] cb_0_1/io_dat_o[2] cb_0_1/io_dat_o[3] cb_0_1/io_dat_o[4]
+ cb_0_1/io_dat_o[5] cb_0_1/io_dat_o[6] cb_0_1/io_dat_o[7] cb_0_1/io_dat_o[8] cb_0_1/io_dat_o[9]
+ cb_0_2/io_dat_o[0] cb_0_2/io_dat_o[10] cb_0_2/io_dat_o[11] cb_0_2/io_dat_o[12] cb_0_2/io_dat_o[13]
+ cb_0_2/io_dat_o[14] cb_0_2/io_dat_o[15] cb_0_2/io_dat_o[1] cb_0_2/io_dat_o[2] cb_0_2/io_dat_o[3]
+ cb_0_2/io_dat_o[4] cb_0_2/io_dat_o[5] cb_0_2/io_dat_o[6] cb_0_2/io_dat_o[7] cb_0_2/io_dat_o[8]
+ cb_0_2/io_dat_o[9] cb_0_3/io_dat_o[0] cb_0_3/io_dat_o[10] cb_0_3/io_dat_o[11] cb_0_3/io_dat_o[12]
+ cb_0_3/io_dat_o[13] cb_0_3/io_dat_o[14] cb_0_3/io_dat_o[15] cb_0_3/io_dat_o[1] cb_0_3/io_dat_o[2]
+ cb_0_3/io_dat_o[3] cb_0_3/io_dat_o[4] cb_0_3/io_dat_o[5] cb_0_3/io_dat_o[6] cb_0_3/io_dat_o[7]
+ cb_0_3/io_dat_o[8] cb_0_3/io_dat_o[9] cb_0_4/io_dat_o[0] cb_0_4/io_dat_o[10] cb_0_4/io_dat_o[11]
+ cb_0_4/io_dat_o[12] cb_0_4/io_dat_o[13] cb_0_4/io_dat_o[14] cb_0_4/io_dat_o[15]
+ cb_0_4/io_dat_o[1] cb_0_4/io_dat_o[2] cb_0_4/io_dat_o[3] cb_0_4/io_dat_o[4] cb_0_4/io_dat_o[5]
+ cb_0_4/io_dat_o[6] cb_0_4/io_dat_o[7] cb_0_4/io_dat_o[8] cb_0_4/io_dat_o[9] cb_0_5/io_dat_o[0]
+ cb_0_5/io_dat_o[10] cb_0_5/io_dat_o[11] cb_0_5/io_dat_o[12] cb_0_5/io_dat_o[13]
+ cb_0_5/io_dat_o[14] cb_0_5/io_dat_o[15] cb_0_5/io_dat_o[1] cb_0_5/io_dat_o[2] cb_0_5/io_dat_o[3]
+ cb_0_5/io_dat_o[4] cb_0_5/io_dat_o[5] cb_0_5/io_dat_o[6] cb_0_5/io_dat_o[7] cb_0_5/io_dat_o[8]
+ cb_0_5/io_dat_o[9] cb_0_6/io_dat_o[0] cb_0_6/io_dat_o[10] cb_0_6/io_dat_o[11] cb_0_6/io_dat_o[12]
+ cb_0_6/io_dat_o[13] cb_0_6/io_dat_o[14] cb_0_6/io_dat_o[15] cb_0_6/io_dat_o[1] cb_0_6/io_dat_o[2]
+ cb_0_6/io_dat_o[3] cb_0_6/io_dat_o[4] cb_0_6/io_dat_o[5] cb_0_6/io_dat_o[6] cb_0_6/io_dat_o[7]
+ cb_0_6/io_dat_o[8] cb_0_6/io_dat_o[9] cb_0_7/io_dat_o[0] cb_0_7/io_dat_o[10] cb_0_7/io_dat_o[11]
+ cb_0_7/io_dat_o[12] cb_0_7/io_dat_o[13] cb_0_7/io_dat_o[14] cb_0_7/io_dat_o[15]
+ cb_0_7/io_dat_o[1] cb_0_7/io_dat_o[2] cb_0_7/io_dat_o[3] cb_0_7/io_dat_o[4] cb_0_7/io_dat_o[5]
+ cb_0_7/io_dat_o[6] cb_0_7/io_dat_o[7] cb_0_7/io_dat_o[8] cb_0_7/io_dat_o[9] cb_0_8/io_dat_o[0]
+ cb_0_8/io_dat_o[10] cb_0_8/io_dat_o[11] cb_0_8/io_dat_o[12] cb_0_8/io_dat_o[13]
+ cb_0_8/io_dat_o[14] cb_0_8/io_dat_o[15] cb_0_8/io_dat_o[1] cb_0_8/io_dat_o[2] cb_0_8/io_dat_o[3]
+ cb_0_8/io_dat_o[4] cb_0_8/io_dat_o[5] cb_0_8/io_dat_o[6] cb_0_8/io_dat_o[7] cb_0_8/io_dat_o[8]
+ cb_0_8/io_dat_o[9] cb_0_9/io_dat_o[0] cb_0_9/io_dat_o[10] cb_0_9/io_dat_o[11] cb_0_9/io_dat_o[12]
+ cb_0_9/io_dat_o[13] cb_0_9/io_dat_o[14] cb_0_9/io_dat_o[15] cb_0_9/io_dat_o[1] cb_0_9/io_dat_o[2]
+ cb_0_9/io_dat_o[3] cb_0_9/io_dat_o[4] cb_0_9/io_dat_o[5] cb_0_9/io_dat_o[6] cb_0_9/io_dat_o[7]
+ cb_0_9/io_dat_o[8] cb_0_9/io_dat_o[9] cb_0_9/io_we_i ccon_0/io_cs_i ccon_7/io_dat_i[0]
+ ccon_7/io_dat_i[10] ccon_7/io_dat_i[11] ccon_7/io_dat_i[12] ccon_7/io_dat_i[13]
+ ccon_7/io_dat_i[14] ccon_7/io_dat_i[15] ccon_7/io_dat_i[16] ccon_7/io_dat_i[17]
+ ccon_7/io_dat_i[18] ccon_7/io_dat_i[19] ccon_7/io_dat_i[1] ccon_7/io_dat_i[20] ccon_7/io_dat_i[21]
+ ccon_7/io_dat_i[22] ccon_7/io_dat_i[23] ccon_7/io_dat_i[24] ccon_7/io_dat_i[25]
+ ccon_7/io_dat_i[26] ccon_7/io_dat_i[27] ccon_7/io_dat_i[28] ccon_7/io_dat_i[29]
+ ccon_7/io_dat_i[2] ccon_7/io_dat_i[30] ccon_7/io_dat_i[31] ccon_7/io_dat_i[3] ccon_7/io_dat_i[4]
+ ccon_7/io_dat_i[5] ccon_7/io_dat_i[6] ccon_7/io_dat_i[7] ccon_7/io_dat_i[8] ccon_7/io_dat_i[9]
+ ccon_0/io_dat_o[0] ccon_0/io_dat_o[10] ccon_0/io_dat_o[11] ccon_0/io_dat_o[12] ccon_0/io_dat_o[13]
+ ccon_0/io_dat_o[14] ccon_0/io_dat_o[15] ccon_0/io_dat_o[16] ccon_0/io_dat_o[17]
+ ccon_0/io_dat_o[18] ccon_0/io_dat_o[19] ccon_0/io_dat_o[1] ccon_0/io_dat_o[20] ccon_0/io_dat_o[21]
+ ccon_0/io_dat_o[22] ccon_0/io_dat_o[23] ccon_0/io_dat_o[24] ccon_0/io_dat_o[25]
+ ccon_0/io_dat_o[26] ccon_0/io_dat_o[27] ccon_0/io_dat_o[28] ccon_0/io_dat_o[29]
+ ccon_0/io_dat_o[2] ccon_0/io_dat_o[30] ccon_0/io_dat_o[31] ccon_0/io_dat_o[3] ccon_0/io_dat_o[4]
+ ccon_0/io_dat_o[5] ccon_0/io_dat_o[6] ccon_0/io_dat_o[7] ccon_0/io_dat_o[8] ccon_0/io_dat_o[9]
+ cb_0_0/io_wo[0] cb_0_0/io_wo[10] cb_0_0/io_wo[11] cb_0_0/io_wo[12] cb_0_0/io_wo[13]
+ cb_0_0/io_wo[14] cb_0_0/io_wo[15] cb_0_0/io_wo[16] cb_0_0/io_wo[17] cb_0_0/io_wo[18]
+ cb_0_0/io_wo[19] cb_0_0/io_wo[1] cb_0_0/io_wo[20] cb_0_0/io_wo[21] cb_0_0/io_wo[22]
+ cb_0_0/io_wo[23] cb_0_0/io_wo[24] cb_0_0/io_wo[25] cb_0_0/io_wo[26] cb_0_0/io_wo[27]
+ cb_0_0/io_wo[28] cb_0_0/io_wo[29] cb_0_0/io_wo[2] cb_0_0/io_wo[30] cb_0_0/io_wo[31]
+ cb_0_0/io_wo[32] cb_0_0/io_wo[33] cb_0_0/io_wo[34] cb_0_0/io_wo[35] cb_0_0/io_wo[36]
+ cb_0_0/io_wo[37] cb_0_0/io_wo[38] cb_0_0/io_wo[39] cb_0_0/io_wo[3] cb_0_0/io_wo[40]
+ cb_0_0/io_wo[41] cb_0_0/io_wo[42] cb_0_0/io_wo[43] cb_0_0/io_wo[44] cb_0_0/io_wo[45]
+ cb_0_0/io_wo[46] cb_0_0/io_wo[47] cb_0_0/io_wo[48] cb_0_0/io_wo[49] cb_0_0/io_wo[4]
+ cb_0_0/io_wo[50] cb_0_0/io_wo[51] cb_0_0/io_wo[52] cb_0_0/io_wo[53] cb_0_0/io_wo[54]
+ cb_0_0/io_wo[55] cb_0_0/io_wo[56] cb_0_0/io_wo[57] cb_0_0/io_wo[58] cb_0_0/io_wo[59]
+ cb_0_0/io_wo[5] cb_0_0/io_wo[60] cb_0_0/io_wo[61] cb_0_0/io_wo[62] cb_0_0/io_wo[63]
+ cb_0_0/io_wo[6] cb_0_0/io_wo[7] cb_0_0/io_wo[8] cb_0_0/io_wo[9] icon/dsi[0] icon/dsi[1]
+ icon/dsi[2] icon/dsi[3] icon/dsi[4] icon/dsi[5] icon/dsi[6] icon/dsi[7] ccon_0/io_dsi_o
+ ccon_0/io_irq cb_0_0/io_vi cb_0_10/io_vi cb_0_1/io_vi cb_0_2/io_vi cb_0_3/io_vi
+ cb_0_4/io_vi cb_0_5/io_vi cb_0_6/io_vi cb_0_7/io_vi cb_0_8/io_vi cb_0_9/io_vi ccon_7/io_we_i
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_con
Xcb_3_1 cb_3_9/io_adr_i[0] cb_3_9/io_adr_i[1] cb_3_1/io_cs_i cb_3_9/io_dat_i[0] cb_3_9/io_dat_i[10]
+ cb_3_9/io_dat_i[11] cb_3_9/io_dat_i[12] cb_3_9/io_dat_i[13] cb_3_9/io_dat_i[14]
+ cb_3_9/io_dat_i[15] cb_3_9/io_dat_i[1] cb_3_9/io_dat_i[2] cb_3_9/io_dat_i[3] cb_3_9/io_dat_i[4]
+ cb_3_9/io_dat_i[5] cb_3_9/io_dat_i[6] cb_3_9/io_dat_i[7] cb_3_9/io_dat_i[8] cb_3_9/io_dat_i[9]
+ cb_3_1/io_dat_o[0] cb_3_1/io_dat_o[10] cb_3_1/io_dat_o[11] cb_3_1/io_dat_o[12] cb_3_1/io_dat_o[13]
+ cb_3_1/io_dat_o[14] cb_3_1/io_dat_o[15] cb_3_1/io_dat_o[1] cb_3_1/io_dat_o[2] cb_3_1/io_dat_o[3]
+ cb_3_1/io_dat_o[4] cb_3_1/io_dat_o[5] cb_3_1/io_dat_o[6] cb_3_1/io_dat_o[7] cb_3_1/io_dat_o[8]
+ cb_3_1/io_dat_o[9] cb_3_2/io_wo[0] cb_3_2/io_wo[10] cb_3_2/io_wo[11] cb_3_2/io_wo[12]
+ cb_3_2/io_wo[13] cb_3_2/io_wo[14] cb_3_2/io_wo[15] cb_3_2/io_wo[16] cb_3_2/io_wo[17]
+ cb_3_2/io_wo[18] cb_3_2/io_wo[19] cb_3_2/io_wo[1] cb_3_2/io_wo[20] cb_3_2/io_wo[21]
+ cb_3_2/io_wo[22] cb_3_2/io_wo[23] cb_3_2/io_wo[24] cb_3_2/io_wo[25] cb_3_2/io_wo[26]
+ cb_3_2/io_wo[27] cb_3_2/io_wo[28] cb_3_2/io_wo[29] cb_3_2/io_wo[2] cb_3_2/io_wo[30]
+ cb_3_2/io_wo[31] cb_3_2/io_wo[32] cb_3_2/io_wo[33] cb_3_2/io_wo[34] cb_3_2/io_wo[35]
+ cb_3_2/io_wo[36] cb_3_2/io_wo[37] cb_3_2/io_wo[38] cb_3_2/io_wo[39] cb_3_2/io_wo[3]
+ cb_3_2/io_wo[40] cb_3_2/io_wo[41] cb_3_2/io_wo[42] cb_3_2/io_wo[43] cb_3_2/io_wo[44]
+ cb_3_2/io_wo[45] cb_3_2/io_wo[46] cb_3_2/io_wo[47] cb_3_2/io_wo[48] cb_3_2/io_wo[49]
+ cb_3_2/io_wo[4] cb_3_2/io_wo[50] cb_3_2/io_wo[51] cb_3_2/io_wo[52] cb_3_2/io_wo[53]
+ cb_3_2/io_wo[54] cb_3_2/io_wo[55] cb_3_2/io_wo[56] cb_3_2/io_wo[57] cb_3_2/io_wo[58]
+ cb_3_2/io_wo[59] cb_3_2/io_wo[5] cb_3_2/io_wo[60] cb_3_2/io_wo[61] cb_3_2/io_wo[62]
+ cb_3_2/io_wo[63] cb_3_2/io_wo[6] cb_3_2/io_wo[7] cb_3_2/io_wo[8] cb_3_2/io_wo[9]
+ cb_3_1/io_i_0_ci cb_3_1/io_i_0_in1[0] cb_3_1/io_i_0_in1[1] cb_3_1/io_i_0_in1[2]
+ cb_3_1/io_i_0_in1[3] cb_3_1/io_i_0_in1[4] cb_3_1/io_i_0_in1[5] cb_3_1/io_i_0_in1[6]
+ cb_3_1/io_i_0_in1[7] cb_3_1/io_i_1_ci cb_3_1/io_i_1_in1[0] cb_3_1/io_i_1_in1[1]
+ cb_3_1/io_i_1_in1[2] cb_3_1/io_i_1_in1[3] cb_3_1/io_i_1_in1[4] cb_3_1/io_i_1_in1[5]
+ cb_3_1/io_i_1_in1[6] cb_3_1/io_i_1_in1[7] cb_3_1/io_i_2_ci cb_3_1/io_i_2_in1[0]
+ cb_3_1/io_i_2_in1[1] cb_3_1/io_i_2_in1[2] cb_3_1/io_i_2_in1[3] cb_3_1/io_i_2_in1[4]
+ cb_3_1/io_i_2_in1[5] cb_3_1/io_i_2_in1[6] cb_3_1/io_i_2_in1[7] cb_3_1/io_i_3_ci
+ cb_3_1/io_i_3_in1[0] cb_3_1/io_i_3_in1[1] cb_3_1/io_i_3_in1[2] cb_3_1/io_i_3_in1[3]
+ cb_3_1/io_i_3_in1[4] cb_3_1/io_i_3_in1[5] cb_3_1/io_i_3_in1[6] cb_3_1/io_i_3_in1[7]
+ cb_3_1/io_i_4_ci cb_3_1/io_i_4_in1[0] cb_3_1/io_i_4_in1[1] cb_3_1/io_i_4_in1[2]
+ cb_3_1/io_i_4_in1[3] cb_3_1/io_i_4_in1[4] cb_3_1/io_i_4_in1[5] cb_3_1/io_i_4_in1[6]
+ cb_3_1/io_i_4_in1[7] cb_3_1/io_i_5_ci cb_3_1/io_i_5_in1[0] cb_3_1/io_i_5_in1[1]
+ cb_3_1/io_i_5_in1[2] cb_3_1/io_i_5_in1[3] cb_3_1/io_i_5_in1[4] cb_3_1/io_i_5_in1[5]
+ cb_3_1/io_i_5_in1[6] cb_3_1/io_i_5_in1[7] cb_3_1/io_i_6_ci cb_3_1/io_i_6_in1[0]
+ cb_3_1/io_i_6_in1[1] cb_3_1/io_i_6_in1[2] cb_3_1/io_i_6_in1[3] cb_3_1/io_i_6_in1[4]
+ cb_3_1/io_i_6_in1[5] cb_3_1/io_i_6_in1[6] cb_3_1/io_i_6_in1[7] cb_3_1/io_i_7_ci
+ cb_3_1/io_i_7_in1[0] cb_3_1/io_i_7_in1[1] cb_3_1/io_i_7_in1[2] cb_3_1/io_i_7_in1[3]
+ cb_3_1/io_i_7_in1[4] cb_3_1/io_i_7_in1[5] cb_3_1/io_i_7_in1[6] cb_3_1/io_i_7_in1[7]
+ cb_3_2/io_i_0_ci cb_3_2/io_i_0_in1[0] cb_3_2/io_i_0_in1[1] cb_3_2/io_i_0_in1[2]
+ cb_3_2/io_i_0_in1[3] cb_3_2/io_i_0_in1[4] cb_3_2/io_i_0_in1[5] cb_3_2/io_i_0_in1[6]
+ cb_3_2/io_i_0_in1[7] cb_3_2/io_i_1_ci cb_3_2/io_i_1_in1[0] cb_3_2/io_i_1_in1[1]
+ cb_3_2/io_i_1_in1[2] cb_3_2/io_i_1_in1[3] cb_3_2/io_i_1_in1[4] cb_3_2/io_i_1_in1[5]
+ cb_3_2/io_i_1_in1[6] cb_3_2/io_i_1_in1[7] cb_3_2/io_i_2_ci cb_3_2/io_i_2_in1[0]
+ cb_3_2/io_i_2_in1[1] cb_3_2/io_i_2_in1[2] cb_3_2/io_i_2_in1[3] cb_3_2/io_i_2_in1[4]
+ cb_3_2/io_i_2_in1[5] cb_3_2/io_i_2_in1[6] cb_3_2/io_i_2_in1[7] cb_3_2/io_i_3_ci
+ cb_3_2/io_i_3_in1[0] cb_3_2/io_i_3_in1[1] cb_3_2/io_i_3_in1[2] cb_3_2/io_i_3_in1[3]
+ cb_3_2/io_i_3_in1[4] cb_3_2/io_i_3_in1[5] cb_3_2/io_i_3_in1[6] cb_3_2/io_i_3_in1[7]
+ cb_3_2/io_i_4_ci cb_3_2/io_i_4_in1[0] cb_3_2/io_i_4_in1[1] cb_3_2/io_i_4_in1[2]
+ cb_3_2/io_i_4_in1[3] cb_3_2/io_i_4_in1[4] cb_3_2/io_i_4_in1[5] cb_3_2/io_i_4_in1[6]
+ cb_3_2/io_i_4_in1[7] cb_3_2/io_i_5_ci cb_3_2/io_i_5_in1[0] cb_3_2/io_i_5_in1[1]
+ cb_3_2/io_i_5_in1[2] cb_3_2/io_i_5_in1[3] cb_3_2/io_i_5_in1[4] cb_3_2/io_i_5_in1[5]
+ cb_3_2/io_i_5_in1[6] cb_3_2/io_i_5_in1[7] cb_3_2/io_i_6_ci cb_3_2/io_i_6_in1[0]
+ cb_3_2/io_i_6_in1[1] cb_3_2/io_i_6_in1[2] cb_3_2/io_i_6_in1[3] cb_3_2/io_i_6_in1[4]
+ cb_3_2/io_i_6_in1[5] cb_3_2/io_i_6_in1[6] cb_3_2/io_i_6_in1[7] cb_3_2/io_i_7_ci
+ cb_3_2/io_i_7_in1[0] cb_3_2/io_i_7_in1[1] cb_3_2/io_i_7_in1[2] cb_3_2/io_i_7_in1[3]
+ cb_3_2/io_i_7_in1[4] cb_3_2/io_i_7_in1[5] cb_3_2/io_i_7_in1[6] cb_3_2/io_i_7_in1[7]
+ cb_3_1/io_vci cb_3_2/io_vci cb_3_1/io_vi cb_3_9/io_we_i cb_3_1/io_wo[0] cb_3_1/io_wo[10]
+ cb_3_1/io_wo[11] cb_3_1/io_wo[12] cb_3_1/io_wo[13] cb_3_1/io_wo[14] cb_3_1/io_wo[15]
+ cb_3_1/io_wo[16] cb_3_1/io_wo[17] cb_3_1/io_wo[18] cb_3_1/io_wo[19] cb_3_1/io_wo[1]
+ cb_3_1/io_wo[20] cb_3_1/io_wo[21] cb_3_1/io_wo[22] cb_3_1/io_wo[23] cb_3_1/io_wo[24]
+ cb_3_1/io_wo[25] cb_3_1/io_wo[26] cb_3_1/io_wo[27] cb_3_1/io_wo[28] cb_3_1/io_wo[29]
+ cb_3_1/io_wo[2] cb_3_1/io_wo[30] cb_3_1/io_wo[31] cb_3_1/io_wo[32] cb_3_1/io_wo[33]
+ cb_3_1/io_wo[34] cb_3_1/io_wo[35] cb_3_1/io_wo[36] cb_3_1/io_wo[37] cb_3_1/io_wo[38]
+ cb_3_1/io_wo[39] cb_3_1/io_wo[3] cb_3_1/io_wo[40] cb_3_1/io_wo[41] cb_3_1/io_wo[42]
+ cb_3_1/io_wo[43] cb_3_1/io_wo[44] cb_3_1/io_wo[45] cb_3_1/io_wo[46] cb_3_1/io_wo[47]
+ cb_3_1/io_wo[48] cb_3_1/io_wo[49] cb_3_1/io_wo[4] cb_3_1/io_wo[50] cb_3_1/io_wo[51]
+ cb_3_1/io_wo[52] cb_3_1/io_wo[53] cb_3_1/io_wo[54] cb_3_1/io_wo[55] cb_3_1/io_wo[56]
+ cb_3_1/io_wo[57] cb_3_1/io_wo[58] cb_3_1/io_wo[59] cb_3_1/io_wo[5] cb_3_1/io_wo[60]
+ cb_3_1/io_wo[61] cb_3_1/io_wo[62] cb_3_1/io_wo[63] cb_3_1/io_wo[6] cb_3_1/io_wo[7]
+ cb_3_1/io_wo[8] cb_3_1/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_7_8 cb_7_9/io_adr_i[0] cb_7_9/io_adr_i[1] cb_7_8/io_cs_i cb_7_9/io_dat_i[0] cb_7_9/io_dat_i[10]
+ cb_7_9/io_dat_i[11] cb_7_9/io_dat_i[12] cb_7_9/io_dat_i[13] cb_7_9/io_dat_i[14]
+ cb_7_9/io_dat_i[15] cb_7_9/io_dat_i[1] cb_7_9/io_dat_i[2] cb_7_9/io_dat_i[3] cb_7_9/io_dat_i[4]
+ cb_7_9/io_dat_i[5] cb_7_9/io_dat_i[6] cb_7_9/io_dat_i[7] cb_7_9/io_dat_i[8] cb_7_9/io_dat_i[9]
+ cb_7_8/io_dat_o[0] cb_7_8/io_dat_o[10] cb_7_8/io_dat_o[11] cb_7_8/io_dat_o[12] cb_7_8/io_dat_o[13]
+ cb_7_8/io_dat_o[14] cb_7_8/io_dat_o[15] cb_7_8/io_dat_o[1] cb_7_8/io_dat_o[2] cb_7_8/io_dat_o[3]
+ cb_7_8/io_dat_o[4] cb_7_8/io_dat_o[5] cb_7_8/io_dat_o[6] cb_7_8/io_dat_o[7] cb_7_8/io_dat_o[8]
+ cb_7_8/io_dat_o[9] cb_7_9/io_wo[0] cb_7_9/io_wo[10] cb_7_9/io_wo[11] cb_7_9/io_wo[12]
+ cb_7_9/io_wo[13] cb_7_9/io_wo[14] cb_7_9/io_wo[15] cb_7_9/io_wo[16] cb_7_9/io_wo[17]
+ cb_7_9/io_wo[18] cb_7_9/io_wo[19] cb_7_9/io_wo[1] cb_7_9/io_wo[20] cb_7_9/io_wo[21]
+ cb_7_9/io_wo[22] cb_7_9/io_wo[23] cb_7_9/io_wo[24] cb_7_9/io_wo[25] cb_7_9/io_wo[26]
+ cb_7_9/io_wo[27] cb_7_9/io_wo[28] cb_7_9/io_wo[29] cb_7_9/io_wo[2] cb_7_9/io_wo[30]
+ cb_7_9/io_wo[31] cb_7_9/io_wo[32] cb_7_9/io_wo[33] cb_7_9/io_wo[34] cb_7_9/io_wo[35]
+ cb_7_9/io_wo[36] cb_7_9/io_wo[37] cb_7_9/io_wo[38] cb_7_9/io_wo[39] cb_7_9/io_wo[3]
+ cb_7_9/io_wo[40] cb_7_9/io_wo[41] cb_7_9/io_wo[42] cb_7_9/io_wo[43] cb_7_9/io_wo[44]
+ cb_7_9/io_wo[45] cb_7_9/io_wo[46] cb_7_9/io_wo[47] cb_7_9/io_wo[48] cb_7_9/io_wo[49]
+ cb_7_9/io_wo[4] cb_7_9/io_wo[50] cb_7_9/io_wo[51] cb_7_9/io_wo[52] cb_7_9/io_wo[53]
+ cb_7_9/io_wo[54] cb_7_9/io_wo[55] cb_7_9/io_wo[56] cb_7_9/io_wo[57] cb_7_9/io_wo[58]
+ cb_7_9/io_wo[59] cb_7_9/io_wo[5] cb_7_9/io_wo[60] cb_7_9/io_wo[61] cb_7_9/io_wo[62]
+ cb_7_9/io_wo[63] cb_7_9/io_wo[6] cb_7_9/io_wo[7] cb_7_9/io_wo[8] cb_7_9/io_wo[9]
+ cb_7_8/io_i_0_ci cb_7_8/io_i_0_in1[0] cb_7_8/io_i_0_in1[1] cb_7_8/io_i_0_in1[2]
+ cb_7_8/io_i_0_in1[3] cb_7_8/io_i_0_in1[4] cb_7_8/io_i_0_in1[5] cb_7_8/io_i_0_in1[6]
+ cb_7_8/io_i_0_in1[7] cb_7_8/io_i_1_ci cb_7_8/io_i_1_in1[0] cb_7_8/io_i_1_in1[1]
+ cb_7_8/io_i_1_in1[2] cb_7_8/io_i_1_in1[3] cb_7_8/io_i_1_in1[4] cb_7_8/io_i_1_in1[5]
+ cb_7_8/io_i_1_in1[6] cb_7_8/io_i_1_in1[7] cb_7_8/io_i_2_ci cb_7_8/io_i_2_in1[0]
+ cb_7_8/io_i_2_in1[1] cb_7_8/io_i_2_in1[2] cb_7_8/io_i_2_in1[3] cb_7_8/io_i_2_in1[4]
+ cb_7_8/io_i_2_in1[5] cb_7_8/io_i_2_in1[6] cb_7_8/io_i_2_in1[7] cb_7_8/io_i_3_ci
+ cb_7_8/io_i_3_in1[0] cb_7_8/io_i_3_in1[1] cb_7_8/io_i_3_in1[2] cb_7_8/io_i_3_in1[3]
+ cb_7_8/io_i_3_in1[4] cb_7_8/io_i_3_in1[5] cb_7_8/io_i_3_in1[6] cb_7_8/io_i_3_in1[7]
+ cb_7_8/io_i_4_ci cb_7_8/io_i_4_in1[0] cb_7_8/io_i_4_in1[1] cb_7_8/io_i_4_in1[2]
+ cb_7_8/io_i_4_in1[3] cb_7_8/io_i_4_in1[4] cb_7_8/io_i_4_in1[5] cb_7_8/io_i_4_in1[6]
+ cb_7_8/io_i_4_in1[7] cb_7_8/io_i_5_ci cb_7_8/io_i_5_in1[0] cb_7_8/io_i_5_in1[1]
+ cb_7_8/io_i_5_in1[2] cb_7_8/io_i_5_in1[3] cb_7_8/io_i_5_in1[4] cb_7_8/io_i_5_in1[5]
+ cb_7_8/io_i_5_in1[6] cb_7_8/io_i_5_in1[7] cb_7_8/io_i_6_ci cb_7_8/io_i_6_in1[0]
+ cb_7_8/io_i_6_in1[1] cb_7_8/io_i_6_in1[2] cb_7_8/io_i_6_in1[3] cb_7_8/io_i_6_in1[4]
+ cb_7_8/io_i_6_in1[5] cb_7_8/io_i_6_in1[6] cb_7_8/io_i_6_in1[7] cb_7_8/io_i_7_ci
+ cb_7_8/io_i_7_in1[0] cb_7_8/io_i_7_in1[1] cb_7_8/io_i_7_in1[2] cb_7_8/io_i_7_in1[3]
+ cb_7_8/io_i_7_in1[4] cb_7_8/io_i_7_in1[5] cb_7_8/io_i_7_in1[6] cb_7_8/io_i_7_in1[7]
+ cb_7_9/io_i_0_ci cb_7_9/io_i_0_in1[0] cb_7_9/io_i_0_in1[1] cb_7_9/io_i_0_in1[2]
+ cb_7_9/io_i_0_in1[3] cb_7_9/io_i_0_in1[4] cb_7_9/io_i_0_in1[5] cb_7_9/io_i_0_in1[6]
+ cb_7_9/io_i_0_in1[7] cb_7_9/io_i_1_ci cb_7_9/io_i_1_in1[0] cb_7_9/io_i_1_in1[1]
+ cb_7_9/io_i_1_in1[2] cb_7_9/io_i_1_in1[3] cb_7_9/io_i_1_in1[4] cb_7_9/io_i_1_in1[5]
+ cb_7_9/io_i_1_in1[6] cb_7_9/io_i_1_in1[7] cb_7_9/io_i_2_ci cb_7_9/io_i_2_in1[0]
+ cb_7_9/io_i_2_in1[1] cb_7_9/io_i_2_in1[2] cb_7_9/io_i_2_in1[3] cb_7_9/io_i_2_in1[4]
+ cb_7_9/io_i_2_in1[5] cb_7_9/io_i_2_in1[6] cb_7_9/io_i_2_in1[7] cb_7_9/io_i_3_ci
+ cb_7_9/io_i_3_in1[0] cb_7_9/io_i_3_in1[1] cb_7_9/io_i_3_in1[2] cb_7_9/io_i_3_in1[3]
+ cb_7_9/io_i_3_in1[4] cb_7_9/io_i_3_in1[5] cb_7_9/io_i_3_in1[6] cb_7_9/io_i_3_in1[7]
+ cb_7_9/io_i_4_ci cb_7_9/io_i_4_in1[0] cb_7_9/io_i_4_in1[1] cb_7_9/io_i_4_in1[2]
+ cb_7_9/io_i_4_in1[3] cb_7_9/io_i_4_in1[4] cb_7_9/io_i_4_in1[5] cb_7_9/io_i_4_in1[6]
+ cb_7_9/io_i_4_in1[7] cb_7_9/io_i_5_ci cb_7_9/io_i_5_in1[0] cb_7_9/io_i_5_in1[1]
+ cb_7_9/io_i_5_in1[2] cb_7_9/io_i_5_in1[3] cb_7_9/io_i_5_in1[4] cb_7_9/io_i_5_in1[5]
+ cb_7_9/io_i_5_in1[6] cb_7_9/io_i_5_in1[7] cb_7_9/io_i_6_ci cb_7_9/io_i_6_in1[0]
+ cb_7_9/io_i_6_in1[1] cb_7_9/io_i_6_in1[2] cb_7_9/io_i_6_in1[3] cb_7_9/io_i_6_in1[4]
+ cb_7_9/io_i_6_in1[5] cb_7_9/io_i_6_in1[6] cb_7_9/io_i_6_in1[7] cb_7_9/io_i_7_ci
+ cb_7_9/io_i_7_in1[0] cb_7_9/io_i_7_in1[1] cb_7_9/io_i_7_in1[2] cb_7_9/io_i_7_in1[3]
+ cb_7_9/io_i_7_in1[4] cb_7_9/io_i_7_in1[5] cb_7_9/io_i_7_in1[6] cb_7_9/io_i_7_in1[7]
+ cb_7_8/io_vci cb_7_9/io_vci cb_7_8/io_vi cb_7_9/io_we_i cb_7_8/io_wo[0] cb_7_8/io_wo[10]
+ cb_7_8/io_wo[11] cb_7_8/io_wo[12] cb_7_8/io_wo[13] cb_7_8/io_wo[14] cb_7_8/io_wo[15]
+ cb_7_8/io_wo[16] cb_7_8/io_wo[17] cb_7_8/io_wo[18] cb_7_8/io_wo[19] cb_7_8/io_wo[1]
+ cb_7_8/io_wo[20] cb_7_8/io_wo[21] cb_7_8/io_wo[22] cb_7_8/io_wo[23] cb_7_8/io_wo[24]
+ cb_7_8/io_wo[25] cb_7_8/io_wo[26] cb_7_8/io_wo[27] cb_7_8/io_wo[28] cb_7_8/io_wo[29]
+ cb_7_8/io_wo[2] cb_7_8/io_wo[30] cb_7_8/io_wo[31] cb_7_8/io_wo[32] cb_7_8/io_wo[33]
+ cb_7_8/io_wo[34] cb_7_8/io_wo[35] cb_7_8/io_wo[36] cb_7_8/io_wo[37] cb_7_8/io_wo[38]
+ cb_7_8/io_wo[39] cb_7_8/io_wo[3] cb_7_8/io_wo[40] cb_7_8/io_wo[41] cb_7_8/io_wo[42]
+ cb_7_8/io_wo[43] cb_7_8/io_wo[44] cb_7_8/io_wo[45] cb_7_8/io_wo[46] cb_7_8/io_wo[47]
+ cb_7_8/io_wo[48] cb_7_8/io_wo[49] cb_7_8/io_wo[4] cb_7_8/io_wo[50] cb_7_8/io_wo[51]
+ cb_7_8/io_wo[52] cb_7_8/io_wo[53] cb_7_8/io_wo[54] cb_7_8/io_wo[55] cb_7_8/io_wo[56]
+ cb_7_8/io_wo[57] cb_7_8/io_wo[58] cb_7_8/io_wo[59] cb_7_8/io_wo[5] cb_7_8/io_wo[60]
+ cb_7_8/io_wo[61] cb_7_8/io_wo[62] cb_7_8/io_wo[63] cb_7_8/io_wo[6] cb_7_8/io_wo[7]
+ cb_7_8/io_wo[8] cb_7_8/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xccon_1 ccon_1/io_ack_o ccon_7/io_adr_i[0] ccon_7/io_adr_i[10] ccon_7/io_adr_i[11]
+ ccon_7/io_adr_i[1] ccon_7/io_adr_i[2] ccon_7/io_adr_i[3] ccon_7/io_adr_i[4] ccon_7/io_adr_i[5]
+ ccon_7/io_adr_i[6] ccon_7/io_adr_i[7] ccon_7/io_adr_i[8] ccon_7/io_adr_i[9] cb_1_9/io_adr_i[0]
+ cb_1_9/io_adr_i[1] cb_1_0/io_cs_i cb_1_1/io_cs_i cb_1_10/io_cs_i cb_1_2/io_cs_i
+ cb_1_3/io_cs_i cb_1_4/io_cs_i cb_1_5/io_cs_i cb_1_6/io_cs_i cb_1_7/io_cs_i cb_1_8/io_cs_i
+ cb_1_9/io_cs_i cb_1_9/io_dat_i[0] cb_1_9/io_dat_i[10] cb_1_9/io_dat_i[11] cb_1_9/io_dat_i[12]
+ cb_1_9/io_dat_i[13] cb_1_9/io_dat_i[14] cb_1_9/io_dat_i[15] cb_1_9/io_dat_i[1] cb_1_9/io_dat_i[2]
+ cb_1_9/io_dat_i[3] cb_1_9/io_dat_i[4] cb_1_9/io_dat_i[5] cb_1_9/io_dat_i[6] cb_1_9/io_dat_i[7]
+ cb_1_9/io_dat_i[8] cb_1_9/io_dat_i[9] cb_1_0/io_dat_o[0] cb_1_0/io_dat_o[10] cb_1_0/io_dat_o[11]
+ cb_1_0/io_dat_o[12] cb_1_0/io_dat_o[13] cb_1_0/io_dat_o[14] cb_1_0/io_dat_o[15]
+ cb_1_0/io_dat_o[1] cb_1_0/io_dat_o[2] cb_1_0/io_dat_o[3] cb_1_0/io_dat_o[4] cb_1_0/io_dat_o[5]
+ cb_1_0/io_dat_o[6] cb_1_0/io_dat_o[7] cb_1_0/io_dat_o[8] cb_1_0/io_dat_o[9] cb_1_10/io_dat_o[0]
+ cb_1_10/io_dat_o[10] cb_1_10/io_dat_o[11] cb_1_10/io_dat_o[12] cb_1_10/io_dat_o[13]
+ cb_1_10/io_dat_o[14] cb_1_10/io_dat_o[15] cb_1_10/io_dat_o[1] cb_1_10/io_dat_o[2]
+ cb_1_10/io_dat_o[3] cb_1_10/io_dat_o[4] cb_1_10/io_dat_o[5] cb_1_10/io_dat_o[6]
+ cb_1_10/io_dat_o[7] cb_1_10/io_dat_o[8] cb_1_10/io_dat_o[9] cb_1_1/io_dat_o[0] cb_1_1/io_dat_o[10]
+ cb_1_1/io_dat_o[11] cb_1_1/io_dat_o[12] cb_1_1/io_dat_o[13] cb_1_1/io_dat_o[14]
+ cb_1_1/io_dat_o[15] cb_1_1/io_dat_o[1] cb_1_1/io_dat_o[2] cb_1_1/io_dat_o[3] cb_1_1/io_dat_o[4]
+ cb_1_1/io_dat_o[5] cb_1_1/io_dat_o[6] cb_1_1/io_dat_o[7] cb_1_1/io_dat_o[8] cb_1_1/io_dat_o[9]
+ cb_1_2/io_dat_o[0] cb_1_2/io_dat_o[10] cb_1_2/io_dat_o[11] cb_1_2/io_dat_o[12] cb_1_2/io_dat_o[13]
+ cb_1_2/io_dat_o[14] cb_1_2/io_dat_o[15] cb_1_2/io_dat_o[1] cb_1_2/io_dat_o[2] cb_1_2/io_dat_o[3]
+ cb_1_2/io_dat_o[4] cb_1_2/io_dat_o[5] cb_1_2/io_dat_o[6] cb_1_2/io_dat_o[7] cb_1_2/io_dat_o[8]
+ cb_1_2/io_dat_o[9] cb_1_3/io_dat_o[0] cb_1_3/io_dat_o[10] cb_1_3/io_dat_o[11] cb_1_3/io_dat_o[12]
+ cb_1_3/io_dat_o[13] cb_1_3/io_dat_o[14] cb_1_3/io_dat_o[15] cb_1_3/io_dat_o[1] cb_1_3/io_dat_o[2]
+ cb_1_3/io_dat_o[3] cb_1_3/io_dat_o[4] cb_1_3/io_dat_o[5] cb_1_3/io_dat_o[6] cb_1_3/io_dat_o[7]
+ cb_1_3/io_dat_o[8] cb_1_3/io_dat_o[9] cb_1_4/io_dat_o[0] cb_1_4/io_dat_o[10] cb_1_4/io_dat_o[11]
+ cb_1_4/io_dat_o[12] cb_1_4/io_dat_o[13] cb_1_4/io_dat_o[14] cb_1_4/io_dat_o[15]
+ cb_1_4/io_dat_o[1] cb_1_4/io_dat_o[2] cb_1_4/io_dat_o[3] cb_1_4/io_dat_o[4] cb_1_4/io_dat_o[5]
+ cb_1_4/io_dat_o[6] cb_1_4/io_dat_o[7] cb_1_4/io_dat_o[8] cb_1_4/io_dat_o[9] cb_1_5/io_dat_o[0]
+ cb_1_5/io_dat_o[10] cb_1_5/io_dat_o[11] cb_1_5/io_dat_o[12] cb_1_5/io_dat_o[13]
+ cb_1_5/io_dat_o[14] cb_1_5/io_dat_o[15] cb_1_5/io_dat_o[1] cb_1_5/io_dat_o[2] cb_1_5/io_dat_o[3]
+ cb_1_5/io_dat_o[4] cb_1_5/io_dat_o[5] cb_1_5/io_dat_o[6] cb_1_5/io_dat_o[7] cb_1_5/io_dat_o[8]
+ cb_1_5/io_dat_o[9] cb_1_6/io_dat_o[0] cb_1_6/io_dat_o[10] cb_1_6/io_dat_o[11] cb_1_6/io_dat_o[12]
+ cb_1_6/io_dat_o[13] cb_1_6/io_dat_o[14] cb_1_6/io_dat_o[15] cb_1_6/io_dat_o[1] cb_1_6/io_dat_o[2]
+ cb_1_6/io_dat_o[3] cb_1_6/io_dat_o[4] cb_1_6/io_dat_o[5] cb_1_6/io_dat_o[6] cb_1_6/io_dat_o[7]
+ cb_1_6/io_dat_o[8] cb_1_6/io_dat_o[9] cb_1_7/io_dat_o[0] cb_1_7/io_dat_o[10] cb_1_7/io_dat_o[11]
+ cb_1_7/io_dat_o[12] cb_1_7/io_dat_o[13] cb_1_7/io_dat_o[14] cb_1_7/io_dat_o[15]
+ cb_1_7/io_dat_o[1] cb_1_7/io_dat_o[2] cb_1_7/io_dat_o[3] cb_1_7/io_dat_o[4] cb_1_7/io_dat_o[5]
+ cb_1_7/io_dat_o[6] cb_1_7/io_dat_o[7] cb_1_7/io_dat_o[8] cb_1_7/io_dat_o[9] cb_1_8/io_dat_o[0]
+ cb_1_8/io_dat_o[10] cb_1_8/io_dat_o[11] cb_1_8/io_dat_o[12] cb_1_8/io_dat_o[13]
+ cb_1_8/io_dat_o[14] cb_1_8/io_dat_o[15] cb_1_8/io_dat_o[1] cb_1_8/io_dat_o[2] cb_1_8/io_dat_o[3]
+ cb_1_8/io_dat_o[4] cb_1_8/io_dat_o[5] cb_1_8/io_dat_o[6] cb_1_8/io_dat_o[7] cb_1_8/io_dat_o[8]
+ cb_1_8/io_dat_o[9] cb_1_9/io_dat_o[0] cb_1_9/io_dat_o[10] cb_1_9/io_dat_o[11] cb_1_9/io_dat_o[12]
+ cb_1_9/io_dat_o[13] cb_1_9/io_dat_o[14] cb_1_9/io_dat_o[15] cb_1_9/io_dat_o[1] cb_1_9/io_dat_o[2]
+ cb_1_9/io_dat_o[3] cb_1_9/io_dat_o[4] cb_1_9/io_dat_o[5] cb_1_9/io_dat_o[6] cb_1_9/io_dat_o[7]
+ cb_1_9/io_dat_o[8] cb_1_9/io_dat_o[9] cb_1_9/io_we_i ccon_1/io_cs_i ccon_7/io_dat_i[0]
+ ccon_7/io_dat_i[10] ccon_7/io_dat_i[11] ccon_7/io_dat_i[12] ccon_7/io_dat_i[13]
+ ccon_7/io_dat_i[14] ccon_7/io_dat_i[15] ccon_7/io_dat_i[16] ccon_7/io_dat_i[17]
+ ccon_7/io_dat_i[18] ccon_7/io_dat_i[19] ccon_7/io_dat_i[1] ccon_7/io_dat_i[20] ccon_7/io_dat_i[21]
+ ccon_7/io_dat_i[22] ccon_7/io_dat_i[23] ccon_7/io_dat_i[24] ccon_7/io_dat_i[25]
+ ccon_7/io_dat_i[26] ccon_7/io_dat_i[27] ccon_7/io_dat_i[28] ccon_7/io_dat_i[29]
+ ccon_7/io_dat_i[2] ccon_7/io_dat_i[30] ccon_7/io_dat_i[31] ccon_7/io_dat_i[3] ccon_7/io_dat_i[4]
+ ccon_7/io_dat_i[5] ccon_7/io_dat_i[6] ccon_7/io_dat_i[7] ccon_7/io_dat_i[8] ccon_7/io_dat_i[9]
+ ccon_1/io_dat_o[0] ccon_1/io_dat_o[10] ccon_1/io_dat_o[11] ccon_1/io_dat_o[12] ccon_1/io_dat_o[13]
+ ccon_1/io_dat_o[14] ccon_1/io_dat_o[15] ccon_1/io_dat_o[16] ccon_1/io_dat_o[17]
+ ccon_1/io_dat_o[18] ccon_1/io_dat_o[19] ccon_1/io_dat_o[1] ccon_1/io_dat_o[20] ccon_1/io_dat_o[21]
+ ccon_1/io_dat_o[22] ccon_1/io_dat_o[23] ccon_1/io_dat_o[24] ccon_1/io_dat_o[25]
+ ccon_1/io_dat_o[26] ccon_1/io_dat_o[27] ccon_1/io_dat_o[28] ccon_1/io_dat_o[29]
+ ccon_1/io_dat_o[2] ccon_1/io_dat_o[30] ccon_1/io_dat_o[31] ccon_1/io_dat_o[3] ccon_1/io_dat_o[4]
+ ccon_1/io_dat_o[5] ccon_1/io_dat_o[6] ccon_1/io_dat_o[7] ccon_1/io_dat_o[8] ccon_1/io_dat_o[9]
+ cb_1_0/io_wo[0] cb_1_0/io_wo[10] cb_1_0/io_wo[11] cb_1_0/io_wo[12] cb_1_0/io_wo[13]
+ cb_1_0/io_wo[14] cb_1_0/io_wo[15] cb_1_0/io_wo[16] cb_1_0/io_wo[17] cb_1_0/io_wo[18]
+ cb_1_0/io_wo[19] cb_1_0/io_wo[1] cb_1_0/io_wo[20] cb_1_0/io_wo[21] cb_1_0/io_wo[22]
+ cb_1_0/io_wo[23] cb_1_0/io_wo[24] cb_1_0/io_wo[25] cb_1_0/io_wo[26] cb_1_0/io_wo[27]
+ cb_1_0/io_wo[28] cb_1_0/io_wo[29] cb_1_0/io_wo[2] cb_1_0/io_wo[30] cb_1_0/io_wo[31]
+ cb_1_0/io_wo[32] cb_1_0/io_wo[33] cb_1_0/io_wo[34] cb_1_0/io_wo[35] cb_1_0/io_wo[36]
+ cb_1_0/io_wo[37] cb_1_0/io_wo[38] cb_1_0/io_wo[39] cb_1_0/io_wo[3] cb_1_0/io_wo[40]
+ cb_1_0/io_wo[41] cb_1_0/io_wo[42] cb_1_0/io_wo[43] cb_1_0/io_wo[44] cb_1_0/io_wo[45]
+ cb_1_0/io_wo[46] cb_1_0/io_wo[47] cb_1_0/io_wo[48] cb_1_0/io_wo[49] cb_1_0/io_wo[4]
+ cb_1_0/io_wo[50] cb_1_0/io_wo[51] cb_1_0/io_wo[52] cb_1_0/io_wo[53] cb_1_0/io_wo[54]
+ cb_1_0/io_wo[55] cb_1_0/io_wo[56] cb_1_0/io_wo[57] cb_1_0/io_wo[58] cb_1_0/io_wo[59]
+ cb_1_0/io_wo[5] cb_1_0/io_wo[60] cb_1_0/io_wo[61] cb_1_0/io_wo[62] cb_1_0/io_wo[63]
+ cb_1_0/io_wo[6] cb_1_0/io_wo[7] cb_1_0/io_wo[8] cb_1_0/io_wo[9] icon/dsi[0] icon/dsi[1]
+ icon/dsi[2] icon/dsi[3] icon/dsi[4] icon/dsi[5] icon/dsi[6] icon/dsi[7] ccon_1/io_dsi_o
+ ccon_1/io_irq cb_1_0/io_vi cb_1_10/io_vi cb_1_1/io_vi cb_1_2/io_vi cb_1_3/io_vi
+ cb_1_4/io_vi cb_1_5/io_vi cb_1_6/io_vi cb_1_7/io_vi cb_1_8/io_vi cb_1_9/io_vi ccon_7/io_we_i
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_con
Xcb_5_5 cb_5_9/io_adr_i[0] cb_5_9/io_adr_i[1] cb_5_5/io_cs_i cb_5_9/io_dat_i[0] cb_5_9/io_dat_i[10]
+ cb_5_9/io_dat_i[11] cb_5_9/io_dat_i[12] cb_5_9/io_dat_i[13] cb_5_9/io_dat_i[14]
+ cb_5_9/io_dat_i[15] cb_5_9/io_dat_i[1] cb_5_9/io_dat_i[2] cb_5_9/io_dat_i[3] cb_5_9/io_dat_i[4]
+ cb_5_9/io_dat_i[5] cb_5_9/io_dat_i[6] cb_5_9/io_dat_i[7] cb_5_9/io_dat_i[8] cb_5_9/io_dat_i[9]
+ cb_5_5/io_dat_o[0] cb_5_5/io_dat_o[10] cb_5_5/io_dat_o[11] cb_5_5/io_dat_o[12] cb_5_5/io_dat_o[13]
+ cb_5_5/io_dat_o[14] cb_5_5/io_dat_o[15] cb_5_5/io_dat_o[1] cb_5_5/io_dat_o[2] cb_5_5/io_dat_o[3]
+ cb_5_5/io_dat_o[4] cb_5_5/io_dat_o[5] cb_5_5/io_dat_o[6] cb_5_5/io_dat_o[7] cb_5_5/io_dat_o[8]
+ cb_5_5/io_dat_o[9] cb_5_6/io_wo[0] cb_5_6/io_wo[10] cb_5_6/io_wo[11] cb_5_6/io_wo[12]
+ cb_5_6/io_wo[13] cb_5_6/io_wo[14] cb_5_6/io_wo[15] cb_5_6/io_wo[16] cb_5_6/io_wo[17]
+ cb_5_6/io_wo[18] cb_5_6/io_wo[19] cb_5_6/io_wo[1] cb_5_6/io_wo[20] cb_5_6/io_wo[21]
+ cb_5_6/io_wo[22] cb_5_6/io_wo[23] cb_5_6/io_wo[24] cb_5_6/io_wo[25] cb_5_6/io_wo[26]
+ cb_5_6/io_wo[27] cb_5_6/io_wo[28] cb_5_6/io_wo[29] cb_5_6/io_wo[2] cb_5_6/io_wo[30]
+ cb_5_6/io_wo[31] cb_5_6/io_wo[32] cb_5_6/io_wo[33] cb_5_6/io_wo[34] cb_5_6/io_wo[35]
+ cb_5_6/io_wo[36] cb_5_6/io_wo[37] cb_5_6/io_wo[38] cb_5_6/io_wo[39] cb_5_6/io_wo[3]
+ cb_5_6/io_wo[40] cb_5_6/io_wo[41] cb_5_6/io_wo[42] cb_5_6/io_wo[43] cb_5_6/io_wo[44]
+ cb_5_6/io_wo[45] cb_5_6/io_wo[46] cb_5_6/io_wo[47] cb_5_6/io_wo[48] cb_5_6/io_wo[49]
+ cb_5_6/io_wo[4] cb_5_6/io_wo[50] cb_5_6/io_wo[51] cb_5_6/io_wo[52] cb_5_6/io_wo[53]
+ cb_5_6/io_wo[54] cb_5_6/io_wo[55] cb_5_6/io_wo[56] cb_5_6/io_wo[57] cb_5_6/io_wo[58]
+ cb_5_6/io_wo[59] cb_5_6/io_wo[5] cb_5_6/io_wo[60] cb_5_6/io_wo[61] cb_5_6/io_wo[62]
+ cb_5_6/io_wo[63] cb_5_6/io_wo[6] cb_5_6/io_wo[7] cb_5_6/io_wo[8] cb_5_6/io_wo[9]
+ cb_5_5/io_i_0_ci cb_5_5/io_i_0_in1[0] cb_5_5/io_i_0_in1[1] cb_5_5/io_i_0_in1[2]
+ cb_5_5/io_i_0_in1[3] cb_5_5/io_i_0_in1[4] cb_5_5/io_i_0_in1[5] cb_5_5/io_i_0_in1[6]
+ cb_5_5/io_i_0_in1[7] cb_5_5/io_i_1_ci cb_5_5/io_i_1_in1[0] cb_5_5/io_i_1_in1[1]
+ cb_5_5/io_i_1_in1[2] cb_5_5/io_i_1_in1[3] cb_5_5/io_i_1_in1[4] cb_5_5/io_i_1_in1[5]
+ cb_5_5/io_i_1_in1[6] cb_5_5/io_i_1_in1[7] cb_5_5/io_i_2_ci cb_5_5/io_i_2_in1[0]
+ cb_5_5/io_i_2_in1[1] cb_5_5/io_i_2_in1[2] cb_5_5/io_i_2_in1[3] cb_5_5/io_i_2_in1[4]
+ cb_5_5/io_i_2_in1[5] cb_5_5/io_i_2_in1[6] cb_5_5/io_i_2_in1[7] cb_5_5/io_i_3_ci
+ cb_5_5/io_i_3_in1[0] cb_5_5/io_i_3_in1[1] cb_5_5/io_i_3_in1[2] cb_5_5/io_i_3_in1[3]
+ cb_5_5/io_i_3_in1[4] cb_5_5/io_i_3_in1[5] cb_5_5/io_i_3_in1[6] cb_5_5/io_i_3_in1[7]
+ cb_5_5/io_i_4_ci cb_5_5/io_i_4_in1[0] cb_5_5/io_i_4_in1[1] cb_5_5/io_i_4_in1[2]
+ cb_5_5/io_i_4_in1[3] cb_5_5/io_i_4_in1[4] cb_5_5/io_i_4_in1[5] cb_5_5/io_i_4_in1[6]
+ cb_5_5/io_i_4_in1[7] cb_5_5/io_i_5_ci cb_5_5/io_i_5_in1[0] cb_5_5/io_i_5_in1[1]
+ cb_5_5/io_i_5_in1[2] cb_5_5/io_i_5_in1[3] cb_5_5/io_i_5_in1[4] cb_5_5/io_i_5_in1[5]
+ cb_5_5/io_i_5_in1[6] cb_5_5/io_i_5_in1[7] cb_5_5/io_i_6_ci cb_5_5/io_i_6_in1[0]
+ cb_5_5/io_i_6_in1[1] cb_5_5/io_i_6_in1[2] cb_5_5/io_i_6_in1[3] cb_5_5/io_i_6_in1[4]
+ cb_5_5/io_i_6_in1[5] cb_5_5/io_i_6_in1[6] cb_5_5/io_i_6_in1[7] cb_5_5/io_i_7_ci
+ cb_5_5/io_i_7_in1[0] cb_5_5/io_i_7_in1[1] cb_5_5/io_i_7_in1[2] cb_5_5/io_i_7_in1[3]
+ cb_5_5/io_i_7_in1[4] cb_5_5/io_i_7_in1[5] cb_5_5/io_i_7_in1[6] cb_5_5/io_i_7_in1[7]
+ cb_5_6/io_i_0_ci cb_5_6/io_i_0_in1[0] cb_5_6/io_i_0_in1[1] cb_5_6/io_i_0_in1[2]
+ cb_5_6/io_i_0_in1[3] cb_5_6/io_i_0_in1[4] cb_5_6/io_i_0_in1[5] cb_5_6/io_i_0_in1[6]
+ cb_5_6/io_i_0_in1[7] cb_5_6/io_i_1_ci cb_5_6/io_i_1_in1[0] cb_5_6/io_i_1_in1[1]
+ cb_5_6/io_i_1_in1[2] cb_5_6/io_i_1_in1[3] cb_5_6/io_i_1_in1[4] cb_5_6/io_i_1_in1[5]
+ cb_5_6/io_i_1_in1[6] cb_5_6/io_i_1_in1[7] cb_5_6/io_i_2_ci cb_5_6/io_i_2_in1[0]
+ cb_5_6/io_i_2_in1[1] cb_5_6/io_i_2_in1[2] cb_5_6/io_i_2_in1[3] cb_5_6/io_i_2_in1[4]
+ cb_5_6/io_i_2_in1[5] cb_5_6/io_i_2_in1[6] cb_5_6/io_i_2_in1[7] cb_5_6/io_i_3_ci
+ cb_5_6/io_i_3_in1[0] cb_5_6/io_i_3_in1[1] cb_5_6/io_i_3_in1[2] cb_5_6/io_i_3_in1[3]
+ cb_5_6/io_i_3_in1[4] cb_5_6/io_i_3_in1[5] cb_5_6/io_i_3_in1[6] cb_5_6/io_i_3_in1[7]
+ cb_5_6/io_i_4_ci cb_5_6/io_i_4_in1[0] cb_5_6/io_i_4_in1[1] cb_5_6/io_i_4_in1[2]
+ cb_5_6/io_i_4_in1[3] cb_5_6/io_i_4_in1[4] cb_5_6/io_i_4_in1[5] cb_5_6/io_i_4_in1[6]
+ cb_5_6/io_i_4_in1[7] cb_5_6/io_i_5_ci cb_5_6/io_i_5_in1[0] cb_5_6/io_i_5_in1[1]
+ cb_5_6/io_i_5_in1[2] cb_5_6/io_i_5_in1[3] cb_5_6/io_i_5_in1[4] cb_5_6/io_i_5_in1[5]
+ cb_5_6/io_i_5_in1[6] cb_5_6/io_i_5_in1[7] cb_5_6/io_i_6_ci cb_5_6/io_i_6_in1[0]
+ cb_5_6/io_i_6_in1[1] cb_5_6/io_i_6_in1[2] cb_5_6/io_i_6_in1[3] cb_5_6/io_i_6_in1[4]
+ cb_5_6/io_i_6_in1[5] cb_5_6/io_i_6_in1[6] cb_5_6/io_i_6_in1[7] cb_5_6/io_i_7_ci
+ cb_5_6/io_i_7_in1[0] cb_5_6/io_i_7_in1[1] cb_5_6/io_i_7_in1[2] cb_5_6/io_i_7_in1[3]
+ cb_5_6/io_i_7_in1[4] cb_5_6/io_i_7_in1[5] cb_5_6/io_i_7_in1[6] cb_5_6/io_i_7_in1[7]
+ cb_5_5/io_vci cb_5_6/io_vci cb_5_5/io_vi cb_5_9/io_we_i cb_5_5/io_wo[0] cb_5_5/io_wo[10]
+ cb_5_5/io_wo[11] cb_5_5/io_wo[12] cb_5_5/io_wo[13] cb_5_5/io_wo[14] cb_5_5/io_wo[15]
+ cb_5_5/io_wo[16] cb_5_5/io_wo[17] cb_5_5/io_wo[18] cb_5_5/io_wo[19] cb_5_5/io_wo[1]
+ cb_5_5/io_wo[20] cb_5_5/io_wo[21] cb_5_5/io_wo[22] cb_5_5/io_wo[23] cb_5_5/io_wo[24]
+ cb_5_5/io_wo[25] cb_5_5/io_wo[26] cb_5_5/io_wo[27] cb_5_5/io_wo[28] cb_5_5/io_wo[29]
+ cb_5_5/io_wo[2] cb_5_5/io_wo[30] cb_5_5/io_wo[31] cb_5_5/io_wo[32] cb_5_5/io_wo[33]
+ cb_5_5/io_wo[34] cb_5_5/io_wo[35] cb_5_5/io_wo[36] cb_5_5/io_wo[37] cb_5_5/io_wo[38]
+ cb_5_5/io_wo[39] cb_5_5/io_wo[3] cb_5_5/io_wo[40] cb_5_5/io_wo[41] cb_5_5/io_wo[42]
+ cb_5_5/io_wo[43] cb_5_5/io_wo[44] cb_5_5/io_wo[45] cb_5_5/io_wo[46] cb_5_5/io_wo[47]
+ cb_5_5/io_wo[48] cb_5_5/io_wo[49] cb_5_5/io_wo[4] cb_5_5/io_wo[50] cb_5_5/io_wo[51]
+ cb_5_5/io_wo[52] cb_5_5/io_wo[53] cb_5_5/io_wo[54] cb_5_5/io_wo[55] cb_5_5/io_wo[56]
+ cb_5_5/io_wo[57] cb_5_5/io_wo[58] cb_5_5/io_wo[59] cb_5_5/io_wo[5] cb_5_5/io_wo[60]
+ cb_5_5/io_wo[61] cb_5_5/io_wo[62] cb_5_5/io_wo[63] cb_5_5/io_wo[6] cb_5_5/io_wo[7]
+ cb_5_5/io_wo[8] cb_5_5/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_3_2 cb_3_9/io_adr_i[0] cb_3_9/io_adr_i[1] cb_3_2/io_cs_i cb_3_9/io_dat_i[0] cb_3_9/io_dat_i[10]
+ cb_3_9/io_dat_i[11] cb_3_9/io_dat_i[12] cb_3_9/io_dat_i[13] cb_3_9/io_dat_i[14]
+ cb_3_9/io_dat_i[15] cb_3_9/io_dat_i[1] cb_3_9/io_dat_i[2] cb_3_9/io_dat_i[3] cb_3_9/io_dat_i[4]
+ cb_3_9/io_dat_i[5] cb_3_9/io_dat_i[6] cb_3_9/io_dat_i[7] cb_3_9/io_dat_i[8] cb_3_9/io_dat_i[9]
+ cb_3_2/io_dat_o[0] cb_3_2/io_dat_o[10] cb_3_2/io_dat_o[11] cb_3_2/io_dat_o[12] cb_3_2/io_dat_o[13]
+ cb_3_2/io_dat_o[14] cb_3_2/io_dat_o[15] cb_3_2/io_dat_o[1] cb_3_2/io_dat_o[2] cb_3_2/io_dat_o[3]
+ cb_3_2/io_dat_o[4] cb_3_2/io_dat_o[5] cb_3_2/io_dat_o[6] cb_3_2/io_dat_o[7] cb_3_2/io_dat_o[8]
+ cb_3_2/io_dat_o[9] cb_3_3/io_wo[0] cb_3_3/io_wo[10] cb_3_3/io_wo[11] cb_3_3/io_wo[12]
+ cb_3_3/io_wo[13] cb_3_3/io_wo[14] cb_3_3/io_wo[15] cb_3_3/io_wo[16] cb_3_3/io_wo[17]
+ cb_3_3/io_wo[18] cb_3_3/io_wo[19] cb_3_3/io_wo[1] cb_3_3/io_wo[20] cb_3_3/io_wo[21]
+ cb_3_3/io_wo[22] cb_3_3/io_wo[23] cb_3_3/io_wo[24] cb_3_3/io_wo[25] cb_3_3/io_wo[26]
+ cb_3_3/io_wo[27] cb_3_3/io_wo[28] cb_3_3/io_wo[29] cb_3_3/io_wo[2] cb_3_3/io_wo[30]
+ cb_3_3/io_wo[31] cb_3_3/io_wo[32] cb_3_3/io_wo[33] cb_3_3/io_wo[34] cb_3_3/io_wo[35]
+ cb_3_3/io_wo[36] cb_3_3/io_wo[37] cb_3_3/io_wo[38] cb_3_3/io_wo[39] cb_3_3/io_wo[3]
+ cb_3_3/io_wo[40] cb_3_3/io_wo[41] cb_3_3/io_wo[42] cb_3_3/io_wo[43] cb_3_3/io_wo[44]
+ cb_3_3/io_wo[45] cb_3_3/io_wo[46] cb_3_3/io_wo[47] cb_3_3/io_wo[48] cb_3_3/io_wo[49]
+ cb_3_3/io_wo[4] cb_3_3/io_wo[50] cb_3_3/io_wo[51] cb_3_3/io_wo[52] cb_3_3/io_wo[53]
+ cb_3_3/io_wo[54] cb_3_3/io_wo[55] cb_3_3/io_wo[56] cb_3_3/io_wo[57] cb_3_3/io_wo[58]
+ cb_3_3/io_wo[59] cb_3_3/io_wo[5] cb_3_3/io_wo[60] cb_3_3/io_wo[61] cb_3_3/io_wo[62]
+ cb_3_3/io_wo[63] cb_3_3/io_wo[6] cb_3_3/io_wo[7] cb_3_3/io_wo[8] cb_3_3/io_wo[9]
+ cb_3_2/io_i_0_ci cb_3_2/io_i_0_in1[0] cb_3_2/io_i_0_in1[1] cb_3_2/io_i_0_in1[2]
+ cb_3_2/io_i_0_in1[3] cb_3_2/io_i_0_in1[4] cb_3_2/io_i_0_in1[5] cb_3_2/io_i_0_in1[6]
+ cb_3_2/io_i_0_in1[7] cb_3_2/io_i_1_ci cb_3_2/io_i_1_in1[0] cb_3_2/io_i_1_in1[1]
+ cb_3_2/io_i_1_in1[2] cb_3_2/io_i_1_in1[3] cb_3_2/io_i_1_in1[4] cb_3_2/io_i_1_in1[5]
+ cb_3_2/io_i_1_in1[6] cb_3_2/io_i_1_in1[7] cb_3_2/io_i_2_ci cb_3_2/io_i_2_in1[0]
+ cb_3_2/io_i_2_in1[1] cb_3_2/io_i_2_in1[2] cb_3_2/io_i_2_in1[3] cb_3_2/io_i_2_in1[4]
+ cb_3_2/io_i_2_in1[5] cb_3_2/io_i_2_in1[6] cb_3_2/io_i_2_in1[7] cb_3_2/io_i_3_ci
+ cb_3_2/io_i_3_in1[0] cb_3_2/io_i_3_in1[1] cb_3_2/io_i_3_in1[2] cb_3_2/io_i_3_in1[3]
+ cb_3_2/io_i_3_in1[4] cb_3_2/io_i_3_in1[5] cb_3_2/io_i_3_in1[6] cb_3_2/io_i_3_in1[7]
+ cb_3_2/io_i_4_ci cb_3_2/io_i_4_in1[0] cb_3_2/io_i_4_in1[1] cb_3_2/io_i_4_in1[2]
+ cb_3_2/io_i_4_in1[3] cb_3_2/io_i_4_in1[4] cb_3_2/io_i_4_in1[5] cb_3_2/io_i_4_in1[6]
+ cb_3_2/io_i_4_in1[7] cb_3_2/io_i_5_ci cb_3_2/io_i_5_in1[0] cb_3_2/io_i_5_in1[1]
+ cb_3_2/io_i_5_in1[2] cb_3_2/io_i_5_in1[3] cb_3_2/io_i_5_in1[4] cb_3_2/io_i_5_in1[5]
+ cb_3_2/io_i_5_in1[6] cb_3_2/io_i_5_in1[7] cb_3_2/io_i_6_ci cb_3_2/io_i_6_in1[0]
+ cb_3_2/io_i_6_in1[1] cb_3_2/io_i_6_in1[2] cb_3_2/io_i_6_in1[3] cb_3_2/io_i_6_in1[4]
+ cb_3_2/io_i_6_in1[5] cb_3_2/io_i_6_in1[6] cb_3_2/io_i_6_in1[7] cb_3_2/io_i_7_ci
+ cb_3_2/io_i_7_in1[0] cb_3_2/io_i_7_in1[1] cb_3_2/io_i_7_in1[2] cb_3_2/io_i_7_in1[3]
+ cb_3_2/io_i_7_in1[4] cb_3_2/io_i_7_in1[5] cb_3_2/io_i_7_in1[6] cb_3_2/io_i_7_in1[7]
+ cb_3_3/io_i_0_ci cb_3_3/io_i_0_in1[0] cb_3_3/io_i_0_in1[1] cb_3_3/io_i_0_in1[2]
+ cb_3_3/io_i_0_in1[3] cb_3_3/io_i_0_in1[4] cb_3_3/io_i_0_in1[5] cb_3_3/io_i_0_in1[6]
+ cb_3_3/io_i_0_in1[7] cb_3_3/io_i_1_ci cb_3_3/io_i_1_in1[0] cb_3_3/io_i_1_in1[1]
+ cb_3_3/io_i_1_in1[2] cb_3_3/io_i_1_in1[3] cb_3_3/io_i_1_in1[4] cb_3_3/io_i_1_in1[5]
+ cb_3_3/io_i_1_in1[6] cb_3_3/io_i_1_in1[7] cb_3_3/io_i_2_ci cb_3_3/io_i_2_in1[0]
+ cb_3_3/io_i_2_in1[1] cb_3_3/io_i_2_in1[2] cb_3_3/io_i_2_in1[3] cb_3_3/io_i_2_in1[4]
+ cb_3_3/io_i_2_in1[5] cb_3_3/io_i_2_in1[6] cb_3_3/io_i_2_in1[7] cb_3_3/io_i_3_ci
+ cb_3_3/io_i_3_in1[0] cb_3_3/io_i_3_in1[1] cb_3_3/io_i_3_in1[2] cb_3_3/io_i_3_in1[3]
+ cb_3_3/io_i_3_in1[4] cb_3_3/io_i_3_in1[5] cb_3_3/io_i_3_in1[6] cb_3_3/io_i_3_in1[7]
+ cb_3_3/io_i_4_ci cb_3_3/io_i_4_in1[0] cb_3_3/io_i_4_in1[1] cb_3_3/io_i_4_in1[2]
+ cb_3_3/io_i_4_in1[3] cb_3_3/io_i_4_in1[4] cb_3_3/io_i_4_in1[5] cb_3_3/io_i_4_in1[6]
+ cb_3_3/io_i_4_in1[7] cb_3_3/io_i_5_ci cb_3_3/io_i_5_in1[0] cb_3_3/io_i_5_in1[1]
+ cb_3_3/io_i_5_in1[2] cb_3_3/io_i_5_in1[3] cb_3_3/io_i_5_in1[4] cb_3_3/io_i_5_in1[5]
+ cb_3_3/io_i_5_in1[6] cb_3_3/io_i_5_in1[7] cb_3_3/io_i_6_ci cb_3_3/io_i_6_in1[0]
+ cb_3_3/io_i_6_in1[1] cb_3_3/io_i_6_in1[2] cb_3_3/io_i_6_in1[3] cb_3_3/io_i_6_in1[4]
+ cb_3_3/io_i_6_in1[5] cb_3_3/io_i_6_in1[6] cb_3_3/io_i_6_in1[7] cb_3_3/io_i_7_ci
+ cb_3_3/io_i_7_in1[0] cb_3_3/io_i_7_in1[1] cb_3_3/io_i_7_in1[2] cb_3_3/io_i_7_in1[3]
+ cb_3_3/io_i_7_in1[4] cb_3_3/io_i_7_in1[5] cb_3_3/io_i_7_in1[6] cb_3_3/io_i_7_in1[7]
+ cb_3_2/io_vci cb_3_3/io_vci cb_3_2/io_vi cb_3_9/io_we_i cb_3_2/io_wo[0] cb_3_2/io_wo[10]
+ cb_3_2/io_wo[11] cb_3_2/io_wo[12] cb_3_2/io_wo[13] cb_3_2/io_wo[14] cb_3_2/io_wo[15]
+ cb_3_2/io_wo[16] cb_3_2/io_wo[17] cb_3_2/io_wo[18] cb_3_2/io_wo[19] cb_3_2/io_wo[1]
+ cb_3_2/io_wo[20] cb_3_2/io_wo[21] cb_3_2/io_wo[22] cb_3_2/io_wo[23] cb_3_2/io_wo[24]
+ cb_3_2/io_wo[25] cb_3_2/io_wo[26] cb_3_2/io_wo[27] cb_3_2/io_wo[28] cb_3_2/io_wo[29]
+ cb_3_2/io_wo[2] cb_3_2/io_wo[30] cb_3_2/io_wo[31] cb_3_2/io_wo[32] cb_3_2/io_wo[33]
+ cb_3_2/io_wo[34] cb_3_2/io_wo[35] cb_3_2/io_wo[36] cb_3_2/io_wo[37] cb_3_2/io_wo[38]
+ cb_3_2/io_wo[39] cb_3_2/io_wo[3] cb_3_2/io_wo[40] cb_3_2/io_wo[41] cb_3_2/io_wo[42]
+ cb_3_2/io_wo[43] cb_3_2/io_wo[44] cb_3_2/io_wo[45] cb_3_2/io_wo[46] cb_3_2/io_wo[47]
+ cb_3_2/io_wo[48] cb_3_2/io_wo[49] cb_3_2/io_wo[4] cb_3_2/io_wo[50] cb_3_2/io_wo[51]
+ cb_3_2/io_wo[52] cb_3_2/io_wo[53] cb_3_2/io_wo[54] cb_3_2/io_wo[55] cb_3_2/io_wo[56]
+ cb_3_2/io_wo[57] cb_3_2/io_wo[58] cb_3_2/io_wo[59] cb_3_2/io_wo[5] cb_3_2/io_wo[60]
+ cb_3_2/io_wo[61] cb_3_2/io_wo[62] cb_3_2/io_wo[63] cb_3_2/io_wo[6] cb_3_2/io_wo[7]
+ cb_3_2/io_wo[8] cb_3_2/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_0_10 cb_0_9/io_adr_i[0] cb_0_9/io_adr_i[1] cb_0_10/io_cs_i cb_0_9/io_dat_i[0]
+ cb_0_9/io_dat_i[10] cb_0_9/io_dat_i[11] cb_0_9/io_dat_i[12] cb_0_9/io_dat_i[13]
+ cb_0_9/io_dat_i[14] cb_0_9/io_dat_i[15] cb_0_9/io_dat_i[1] cb_0_9/io_dat_i[2] cb_0_9/io_dat_i[3]
+ cb_0_9/io_dat_i[4] cb_0_9/io_dat_i[5] cb_0_9/io_dat_i[6] cb_0_9/io_dat_i[7] cb_0_9/io_dat_i[8]
+ cb_0_9/io_dat_i[9] cb_0_10/io_dat_o[0] cb_0_10/io_dat_o[10] cb_0_10/io_dat_o[11]
+ cb_0_10/io_dat_o[12] cb_0_10/io_dat_o[13] cb_0_10/io_dat_o[14] cb_0_10/io_dat_o[15]
+ cb_0_10/io_dat_o[1] cb_0_10/io_dat_o[2] cb_0_10/io_dat_o[3] cb_0_10/io_dat_o[4]
+ cb_0_10/io_dat_o[5] cb_0_10/io_dat_o[6] cb_0_10/io_dat_o[7] cb_0_10/io_dat_o[8]
+ cb_0_10/io_dat_o[9] cb_0_10/io_eo[0] cb_0_10/io_eo[10] cb_0_10/io_eo[11] cb_0_10/io_eo[12]
+ cb_0_10/io_eo[13] cb_0_10/io_eo[14] cb_0_10/io_eo[15] cb_0_10/io_eo[16] cb_0_10/io_eo[17]
+ cb_0_10/io_eo[18] cb_0_10/io_eo[19] cb_0_10/io_eo[1] cb_0_10/io_eo[20] cb_0_10/io_eo[21]
+ cb_0_10/io_eo[22] cb_0_10/io_eo[23] cb_0_10/io_eo[24] cb_0_10/io_eo[25] cb_0_10/io_eo[26]
+ cb_0_10/io_eo[27] cb_0_10/io_eo[28] cb_0_10/io_eo[29] cb_0_10/io_eo[2] cb_0_10/io_eo[30]
+ cb_0_10/io_eo[31] cb_0_10/io_eo[32] cb_0_10/io_eo[33] cb_0_10/io_eo[34] cb_0_10/io_eo[35]
+ cb_0_10/io_eo[36] cb_0_10/io_eo[37] cb_0_10/io_eo[38] cb_0_10/io_eo[39] cb_0_10/io_eo[3]
+ cb_0_10/io_eo[40] cb_0_10/io_eo[41] cb_0_10/io_eo[42] cb_0_10/io_eo[43] cb_0_10/io_eo[44]
+ cb_0_10/io_eo[45] cb_0_10/io_eo[46] cb_0_10/io_eo[47] cb_0_10/io_eo[48] cb_0_10/io_eo[49]
+ cb_0_10/io_eo[4] cb_0_10/io_eo[50] cb_0_10/io_eo[51] cb_0_10/io_eo[52] cb_0_10/io_eo[53]
+ cb_0_10/io_eo[54] cb_0_10/io_eo[55] cb_0_10/io_eo[56] cb_0_10/io_eo[57] cb_0_10/io_eo[58]
+ cb_0_10/io_eo[59] cb_0_10/io_eo[5] cb_0_10/io_eo[60] cb_0_10/io_eo[61] cb_0_10/io_eo[62]
+ cb_0_10/io_eo[63] cb_0_10/io_eo[6] cb_0_10/io_eo[7] cb_0_10/io_eo[8] cb_0_10/io_eo[9]
+ cb_0_9/io_o_0_co cb_0_9/io_o_0_out[0] cb_0_9/io_o_0_out[1] cb_0_9/io_o_0_out[2]
+ cb_0_9/io_o_0_out[3] cb_0_9/io_o_0_out[4] cb_0_9/io_o_0_out[5] cb_0_9/io_o_0_out[6]
+ cb_0_9/io_o_0_out[7] cb_0_9/io_o_1_co cb_0_9/io_o_1_out[0] cb_0_9/io_o_1_out[1]
+ cb_0_9/io_o_1_out[2] cb_0_9/io_o_1_out[3] cb_0_9/io_o_1_out[4] cb_0_9/io_o_1_out[5]
+ cb_0_9/io_o_1_out[6] cb_0_9/io_o_1_out[7] cb_0_9/io_o_2_co cb_0_9/io_o_2_out[0]
+ cb_0_9/io_o_2_out[1] cb_0_9/io_o_2_out[2] cb_0_9/io_o_2_out[3] cb_0_9/io_o_2_out[4]
+ cb_0_9/io_o_2_out[5] cb_0_9/io_o_2_out[6] cb_0_9/io_o_2_out[7] cb_0_9/io_o_3_co
+ cb_0_9/io_o_3_out[0] cb_0_9/io_o_3_out[1] cb_0_9/io_o_3_out[2] cb_0_9/io_o_3_out[3]
+ cb_0_9/io_o_3_out[4] cb_0_9/io_o_3_out[5] cb_0_9/io_o_3_out[6] cb_0_9/io_o_3_out[7]
+ cb_0_9/io_o_4_co cb_0_9/io_o_4_out[0] cb_0_9/io_o_4_out[1] cb_0_9/io_o_4_out[2]
+ cb_0_9/io_o_4_out[3] cb_0_9/io_o_4_out[4] cb_0_9/io_o_4_out[5] cb_0_9/io_o_4_out[6]
+ cb_0_9/io_o_4_out[7] cb_0_9/io_o_5_co cb_0_9/io_o_5_out[0] cb_0_9/io_o_5_out[1]
+ cb_0_9/io_o_5_out[2] cb_0_9/io_o_5_out[3] cb_0_9/io_o_5_out[4] cb_0_9/io_o_5_out[5]
+ cb_0_9/io_o_5_out[6] cb_0_9/io_o_5_out[7] cb_0_9/io_o_6_co cb_0_9/io_o_6_out[0]
+ cb_0_9/io_o_6_out[1] cb_0_9/io_o_6_out[2] cb_0_9/io_o_6_out[3] cb_0_9/io_o_6_out[4]
+ cb_0_9/io_o_6_out[5] cb_0_9/io_o_6_out[6] cb_0_9/io_o_6_out[7] cb_0_9/io_o_7_co
+ cb_0_9/io_o_7_out[0] cb_0_9/io_o_7_out[1] cb_0_9/io_o_7_out[2] cb_0_9/io_o_7_out[3]
+ cb_0_9/io_o_7_out[4] cb_0_9/io_o_7_out[5] cb_0_9/io_o_7_out[6] cb_0_9/io_o_7_out[7]
+ cb_0_10/io_o_0_co cb_0_10/io_eo[0] cb_0_10/io_eo[1] cb_0_10/io_eo[2] cb_0_10/io_eo[3]
+ cb_0_10/io_eo[4] cb_0_10/io_eo[5] cb_0_10/io_eo[6] cb_0_10/io_eo[7] cb_0_10/io_o_1_co
+ cb_0_10/io_eo[8] cb_0_10/io_eo[9] cb_0_10/io_eo[10] cb_0_10/io_eo[11] cb_0_10/io_eo[12]
+ cb_0_10/io_eo[13] cb_0_10/io_eo[14] cb_0_10/io_eo[15] cb_0_10/io_o_2_co cb_0_10/io_eo[16]
+ cb_0_10/io_eo[17] cb_0_10/io_eo[18] cb_0_10/io_eo[19] cb_0_10/io_eo[20] cb_0_10/io_eo[21]
+ cb_0_10/io_eo[22] cb_0_10/io_eo[23] cb_0_10/io_o_3_co cb_0_10/io_eo[24] cb_0_10/io_eo[25]
+ cb_0_10/io_eo[26] cb_0_10/io_eo[27] cb_0_10/io_eo[28] cb_0_10/io_eo[29] cb_0_10/io_eo[30]
+ cb_0_10/io_eo[31] cb_0_10/io_o_4_co cb_0_10/io_eo[32] cb_0_10/io_eo[33] cb_0_10/io_eo[34]
+ cb_0_10/io_eo[35] cb_0_10/io_eo[36] cb_0_10/io_eo[37] cb_0_10/io_eo[38] cb_0_10/io_eo[39]
+ cb_0_10/io_o_5_co cb_0_10/io_eo[40] cb_0_10/io_eo[41] cb_0_10/io_eo[42] cb_0_10/io_eo[43]
+ cb_0_10/io_eo[44] cb_0_10/io_eo[45] cb_0_10/io_eo[46] cb_0_10/io_eo[47] cb_0_10/io_o_6_co
+ cb_0_10/io_eo[48] cb_0_10/io_eo[49] cb_0_10/io_eo[50] cb_0_10/io_eo[51] cb_0_10/io_eo[52]
+ cb_0_10/io_eo[53] cb_0_10/io_eo[54] cb_0_10/io_eo[55] cb_0_10/io_o_7_co cb_0_10/io_eo[56]
+ cb_0_10/io_eo[57] cb_0_10/io_eo[58] cb_0_10/io_eo[59] cb_0_10/io_eo[60] cb_0_10/io_eo[61]
+ cb_0_10/io_eo[62] cb_0_10/io_eo[63] cb_0_9/io_vco cb_0_10/io_vco cb_0_10/io_vi cb_0_9/io_we_i
+ cb_0_9/io_eo[0] cb_0_9/io_eo[10] cb_0_9/io_eo[11] cb_0_9/io_eo[12] cb_0_9/io_eo[13]
+ cb_0_9/io_eo[14] cb_0_9/io_eo[15] cb_0_9/io_eo[16] cb_0_9/io_eo[17] cb_0_9/io_eo[18]
+ cb_0_9/io_eo[19] cb_0_9/io_eo[1] cb_0_9/io_eo[20] cb_0_9/io_eo[21] cb_0_9/io_eo[22]
+ cb_0_9/io_eo[23] cb_0_9/io_eo[24] cb_0_9/io_eo[25] cb_0_9/io_eo[26] cb_0_9/io_eo[27]
+ cb_0_9/io_eo[28] cb_0_9/io_eo[29] cb_0_9/io_eo[2] cb_0_9/io_eo[30] cb_0_9/io_eo[31]
+ cb_0_9/io_eo[32] cb_0_9/io_eo[33] cb_0_9/io_eo[34] cb_0_9/io_eo[35] cb_0_9/io_eo[36]
+ cb_0_9/io_eo[37] cb_0_9/io_eo[38] cb_0_9/io_eo[39] cb_0_9/io_eo[3] cb_0_9/io_eo[40]
+ cb_0_9/io_eo[41] cb_0_9/io_eo[42] cb_0_9/io_eo[43] cb_0_9/io_eo[44] cb_0_9/io_eo[45]
+ cb_0_9/io_eo[46] cb_0_9/io_eo[47] cb_0_9/io_eo[48] cb_0_9/io_eo[49] cb_0_9/io_eo[4]
+ cb_0_9/io_eo[50] cb_0_9/io_eo[51] cb_0_9/io_eo[52] cb_0_9/io_eo[53] cb_0_9/io_eo[54]
+ cb_0_9/io_eo[55] cb_0_9/io_eo[56] cb_0_9/io_eo[57] cb_0_9/io_eo[58] cb_0_9/io_eo[59]
+ cb_0_9/io_eo[5] cb_0_9/io_eo[60] cb_0_9/io_eo[61] cb_0_9/io_eo[62] cb_0_9/io_eo[63]
+ cb_0_9/io_eo[6] cb_0_9/io_eo[7] cb_0_9/io_eo[8] cb_0_9/io_eo[9] mcons_3/clock mcons_3/reset
+ vccd1 vssd1 cic_block
Xcb_7_9 cb_7_9/io_adr_i[0] cb_7_9/io_adr_i[1] cb_7_9/io_cs_i cb_7_9/io_dat_i[0] cb_7_9/io_dat_i[10]
+ cb_7_9/io_dat_i[11] cb_7_9/io_dat_i[12] cb_7_9/io_dat_i[13] cb_7_9/io_dat_i[14]
+ cb_7_9/io_dat_i[15] cb_7_9/io_dat_i[1] cb_7_9/io_dat_i[2] cb_7_9/io_dat_i[3] cb_7_9/io_dat_i[4]
+ cb_7_9/io_dat_i[5] cb_7_9/io_dat_i[6] cb_7_9/io_dat_i[7] cb_7_9/io_dat_i[8] cb_7_9/io_dat_i[9]
+ cb_7_9/io_dat_o[0] cb_7_9/io_dat_o[10] cb_7_9/io_dat_o[11] cb_7_9/io_dat_o[12] cb_7_9/io_dat_o[13]
+ cb_7_9/io_dat_o[14] cb_7_9/io_dat_o[15] cb_7_9/io_dat_o[1] cb_7_9/io_dat_o[2] cb_7_9/io_dat_o[3]
+ cb_7_9/io_dat_o[4] cb_7_9/io_dat_o[5] cb_7_9/io_dat_o[6] cb_7_9/io_dat_o[7] cb_7_9/io_dat_o[8]
+ cb_7_9/io_dat_o[9] cb_7_9/io_eo[0] cb_7_9/io_eo[10] cb_7_9/io_eo[11] cb_7_9/io_eo[12]
+ cb_7_9/io_eo[13] cb_7_9/io_eo[14] cb_7_9/io_eo[15] cb_7_9/io_eo[16] cb_7_9/io_eo[17]
+ cb_7_9/io_eo[18] cb_7_9/io_eo[19] cb_7_9/io_eo[1] cb_7_9/io_eo[20] cb_7_9/io_eo[21]
+ cb_7_9/io_eo[22] cb_7_9/io_eo[23] cb_7_9/io_eo[24] cb_7_9/io_eo[25] cb_7_9/io_eo[26]
+ cb_7_9/io_eo[27] cb_7_9/io_eo[28] cb_7_9/io_eo[29] cb_7_9/io_eo[2] cb_7_9/io_eo[30]
+ cb_7_9/io_eo[31] cb_7_9/io_eo[32] cb_7_9/io_eo[33] cb_7_9/io_eo[34] cb_7_9/io_eo[35]
+ cb_7_9/io_eo[36] cb_7_9/io_eo[37] cb_7_9/io_eo[38] cb_7_9/io_eo[39] cb_7_9/io_eo[3]
+ cb_7_9/io_eo[40] cb_7_9/io_eo[41] cb_7_9/io_eo[42] cb_7_9/io_eo[43] cb_7_9/io_eo[44]
+ cb_7_9/io_eo[45] cb_7_9/io_eo[46] cb_7_9/io_eo[47] cb_7_9/io_eo[48] cb_7_9/io_eo[49]
+ cb_7_9/io_eo[4] cb_7_9/io_eo[50] cb_7_9/io_eo[51] cb_7_9/io_eo[52] cb_7_9/io_eo[53]
+ cb_7_9/io_eo[54] cb_7_9/io_eo[55] cb_7_9/io_eo[56] cb_7_9/io_eo[57] cb_7_9/io_eo[58]
+ cb_7_9/io_eo[59] cb_7_9/io_eo[5] cb_7_9/io_eo[60] cb_7_9/io_eo[61] cb_7_9/io_eo[62]
+ cb_7_9/io_eo[63] cb_7_9/io_eo[6] cb_7_9/io_eo[7] cb_7_9/io_eo[8] cb_7_9/io_eo[9]
+ cb_7_9/io_i_0_ci cb_7_9/io_i_0_in1[0] cb_7_9/io_i_0_in1[1] cb_7_9/io_i_0_in1[2]
+ cb_7_9/io_i_0_in1[3] cb_7_9/io_i_0_in1[4] cb_7_9/io_i_0_in1[5] cb_7_9/io_i_0_in1[6]
+ cb_7_9/io_i_0_in1[7] cb_7_9/io_i_1_ci cb_7_9/io_i_1_in1[0] cb_7_9/io_i_1_in1[1]
+ cb_7_9/io_i_1_in1[2] cb_7_9/io_i_1_in1[3] cb_7_9/io_i_1_in1[4] cb_7_9/io_i_1_in1[5]
+ cb_7_9/io_i_1_in1[6] cb_7_9/io_i_1_in1[7] cb_7_9/io_i_2_ci cb_7_9/io_i_2_in1[0]
+ cb_7_9/io_i_2_in1[1] cb_7_9/io_i_2_in1[2] cb_7_9/io_i_2_in1[3] cb_7_9/io_i_2_in1[4]
+ cb_7_9/io_i_2_in1[5] cb_7_9/io_i_2_in1[6] cb_7_9/io_i_2_in1[7] cb_7_9/io_i_3_ci
+ cb_7_9/io_i_3_in1[0] cb_7_9/io_i_3_in1[1] cb_7_9/io_i_3_in1[2] cb_7_9/io_i_3_in1[3]
+ cb_7_9/io_i_3_in1[4] cb_7_9/io_i_3_in1[5] cb_7_9/io_i_3_in1[6] cb_7_9/io_i_3_in1[7]
+ cb_7_9/io_i_4_ci cb_7_9/io_i_4_in1[0] cb_7_9/io_i_4_in1[1] cb_7_9/io_i_4_in1[2]
+ cb_7_9/io_i_4_in1[3] cb_7_9/io_i_4_in1[4] cb_7_9/io_i_4_in1[5] cb_7_9/io_i_4_in1[6]
+ cb_7_9/io_i_4_in1[7] cb_7_9/io_i_5_ci cb_7_9/io_i_5_in1[0] cb_7_9/io_i_5_in1[1]
+ cb_7_9/io_i_5_in1[2] cb_7_9/io_i_5_in1[3] cb_7_9/io_i_5_in1[4] cb_7_9/io_i_5_in1[5]
+ cb_7_9/io_i_5_in1[6] cb_7_9/io_i_5_in1[7] cb_7_9/io_i_6_ci cb_7_9/io_i_6_in1[0]
+ cb_7_9/io_i_6_in1[1] cb_7_9/io_i_6_in1[2] cb_7_9/io_i_6_in1[3] cb_7_9/io_i_6_in1[4]
+ cb_7_9/io_i_6_in1[5] cb_7_9/io_i_6_in1[6] cb_7_9/io_i_6_in1[7] cb_7_9/io_i_7_ci
+ cb_7_9/io_i_7_in1[0] cb_7_9/io_i_7_in1[1] cb_7_9/io_i_7_in1[2] cb_7_9/io_i_7_in1[3]
+ cb_7_9/io_i_7_in1[4] cb_7_9/io_i_7_in1[5] cb_7_9/io_i_7_in1[6] cb_7_9/io_i_7_in1[7]
+ cb_7_9/io_o_0_co cb_7_9/io_o_0_out[0] cb_7_9/io_o_0_out[1] cb_7_9/io_o_0_out[2]
+ cb_7_9/io_o_0_out[3] cb_7_9/io_o_0_out[4] cb_7_9/io_o_0_out[5] cb_7_9/io_o_0_out[6]
+ cb_7_9/io_o_0_out[7] cb_7_9/io_o_1_co cb_7_9/io_o_1_out[0] cb_7_9/io_o_1_out[1]
+ cb_7_9/io_o_1_out[2] cb_7_9/io_o_1_out[3] cb_7_9/io_o_1_out[4] cb_7_9/io_o_1_out[5]
+ cb_7_9/io_o_1_out[6] cb_7_9/io_o_1_out[7] cb_7_9/io_o_2_co cb_7_9/io_o_2_out[0]
+ cb_7_9/io_o_2_out[1] cb_7_9/io_o_2_out[2] cb_7_9/io_o_2_out[3] cb_7_9/io_o_2_out[4]
+ cb_7_9/io_o_2_out[5] cb_7_9/io_o_2_out[6] cb_7_9/io_o_2_out[7] cb_7_9/io_o_3_co
+ cb_7_9/io_o_3_out[0] cb_7_9/io_o_3_out[1] cb_7_9/io_o_3_out[2] cb_7_9/io_o_3_out[3]
+ cb_7_9/io_o_3_out[4] cb_7_9/io_o_3_out[5] cb_7_9/io_o_3_out[6] cb_7_9/io_o_3_out[7]
+ cb_7_9/io_o_4_co cb_7_9/io_o_4_out[0] cb_7_9/io_o_4_out[1] cb_7_9/io_o_4_out[2]
+ cb_7_9/io_o_4_out[3] cb_7_9/io_o_4_out[4] cb_7_9/io_o_4_out[5] cb_7_9/io_o_4_out[6]
+ cb_7_9/io_o_4_out[7] cb_7_9/io_o_5_co cb_7_9/io_o_5_out[0] cb_7_9/io_o_5_out[1]
+ cb_7_9/io_o_5_out[2] cb_7_9/io_o_5_out[3] cb_7_9/io_o_5_out[4] cb_7_9/io_o_5_out[5]
+ cb_7_9/io_o_5_out[6] cb_7_9/io_o_5_out[7] cb_7_9/io_o_6_co cb_7_9/io_o_6_out[0]
+ cb_7_9/io_o_6_out[1] cb_7_9/io_o_6_out[2] cb_7_9/io_o_6_out[3] cb_7_9/io_o_6_out[4]
+ cb_7_9/io_o_6_out[5] cb_7_9/io_o_6_out[6] cb_7_9/io_o_6_out[7] cb_7_9/io_o_7_co
+ cb_7_9/io_o_7_out[0] cb_7_9/io_o_7_out[1] cb_7_9/io_o_7_out[2] cb_7_9/io_o_7_out[3]
+ cb_7_9/io_o_7_out[4] cb_7_9/io_o_7_out[5] cb_7_9/io_o_7_out[6] cb_7_9/io_o_7_out[7]
+ cb_7_9/io_vci cb_7_9/io_vco cb_7_9/io_vi cb_7_9/io_we_i cb_7_9/io_wo[0] cb_7_9/io_wo[10]
+ cb_7_9/io_wo[11] cb_7_9/io_wo[12] cb_7_9/io_wo[13] cb_7_9/io_wo[14] cb_7_9/io_wo[15]
+ cb_7_9/io_wo[16] cb_7_9/io_wo[17] cb_7_9/io_wo[18] cb_7_9/io_wo[19] cb_7_9/io_wo[1]
+ cb_7_9/io_wo[20] cb_7_9/io_wo[21] cb_7_9/io_wo[22] cb_7_9/io_wo[23] cb_7_9/io_wo[24]
+ cb_7_9/io_wo[25] cb_7_9/io_wo[26] cb_7_9/io_wo[27] cb_7_9/io_wo[28] cb_7_9/io_wo[29]
+ cb_7_9/io_wo[2] cb_7_9/io_wo[30] cb_7_9/io_wo[31] cb_7_9/io_wo[32] cb_7_9/io_wo[33]
+ cb_7_9/io_wo[34] cb_7_9/io_wo[35] cb_7_9/io_wo[36] cb_7_9/io_wo[37] cb_7_9/io_wo[38]
+ cb_7_9/io_wo[39] cb_7_9/io_wo[3] cb_7_9/io_wo[40] cb_7_9/io_wo[41] cb_7_9/io_wo[42]
+ cb_7_9/io_wo[43] cb_7_9/io_wo[44] cb_7_9/io_wo[45] cb_7_9/io_wo[46] cb_7_9/io_wo[47]
+ cb_7_9/io_wo[48] cb_7_9/io_wo[49] cb_7_9/io_wo[4] cb_7_9/io_wo[50] cb_7_9/io_wo[51]
+ cb_7_9/io_wo[52] cb_7_9/io_wo[53] cb_7_9/io_wo[54] cb_7_9/io_wo[55] cb_7_9/io_wo[56]
+ cb_7_9/io_wo[57] cb_7_9/io_wo[58] cb_7_9/io_wo[59] cb_7_9/io_wo[5] cb_7_9/io_wo[60]
+ cb_7_9/io_wo[61] cb_7_9/io_wo[62] cb_7_9/io_wo[63] cb_7_9/io_wo[6] cb_7_9/io_wo[7]
+ cb_7_9/io_wo[8] cb_7_9/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_5_6 cb_5_9/io_adr_i[0] cb_5_9/io_adr_i[1] cb_5_6/io_cs_i cb_5_9/io_dat_i[0] cb_5_9/io_dat_i[10]
+ cb_5_9/io_dat_i[11] cb_5_9/io_dat_i[12] cb_5_9/io_dat_i[13] cb_5_9/io_dat_i[14]
+ cb_5_9/io_dat_i[15] cb_5_9/io_dat_i[1] cb_5_9/io_dat_i[2] cb_5_9/io_dat_i[3] cb_5_9/io_dat_i[4]
+ cb_5_9/io_dat_i[5] cb_5_9/io_dat_i[6] cb_5_9/io_dat_i[7] cb_5_9/io_dat_i[8] cb_5_9/io_dat_i[9]
+ cb_5_6/io_dat_o[0] cb_5_6/io_dat_o[10] cb_5_6/io_dat_o[11] cb_5_6/io_dat_o[12] cb_5_6/io_dat_o[13]
+ cb_5_6/io_dat_o[14] cb_5_6/io_dat_o[15] cb_5_6/io_dat_o[1] cb_5_6/io_dat_o[2] cb_5_6/io_dat_o[3]
+ cb_5_6/io_dat_o[4] cb_5_6/io_dat_o[5] cb_5_6/io_dat_o[6] cb_5_6/io_dat_o[7] cb_5_6/io_dat_o[8]
+ cb_5_6/io_dat_o[9] cb_5_7/io_wo[0] cb_5_7/io_wo[10] cb_5_7/io_wo[11] cb_5_7/io_wo[12]
+ cb_5_7/io_wo[13] cb_5_7/io_wo[14] cb_5_7/io_wo[15] cb_5_7/io_wo[16] cb_5_7/io_wo[17]
+ cb_5_7/io_wo[18] cb_5_7/io_wo[19] cb_5_7/io_wo[1] cb_5_7/io_wo[20] cb_5_7/io_wo[21]
+ cb_5_7/io_wo[22] cb_5_7/io_wo[23] cb_5_7/io_wo[24] cb_5_7/io_wo[25] cb_5_7/io_wo[26]
+ cb_5_7/io_wo[27] cb_5_7/io_wo[28] cb_5_7/io_wo[29] cb_5_7/io_wo[2] cb_5_7/io_wo[30]
+ cb_5_7/io_wo[31] cb_5_7/io_wo[32] cb_5_7/io_wo[33] cb_5_7/io_wo[34] cb_5_7/io_wo[35]
+ cb_5_7/io_wo[36] cb_5_7/io_wo[37] cb_5_7/io_wo[38] cb_5_7/io_wo[39] cb_5_7/io_wo[3]
+ cb_5_7/io_wo[40] cb_5_7/io_wo[41] cb_5_7/io_wo[42] cb_5_7/io_wo[43] cb_5_7/io_wo[44]
+ cb_5_7/io_wo[45] cb_5_7/io_wo[46] cb_5_7/io_wo[47] cb_5_7/io_wo[48] cb_5_7/io_wo[49]
+ cb_5_7/io_wo[4] cb_5_7/io_wo[50] cb_5_7/io_wo[51] cb_5_7/io_wo[52] cb_5_7/io_wo[53]
+ cb_5_7/io_wo[54] cb_5_7/io_wo[55] cb_5_7/io_wo[56] cb_5_7/io_wo[57] cb_5_7/io_wo[58]
+ cb_5_7/io_wo[59] cb_5_7/io_wo[5] cb_5_7/io_wo[60] cb_5_7/io_wo[61] cb_5_7/io_wo[62]
+ cb_5_7/io_wo[63] cb_5_7/io_wo[6] cb_5_7/io_wo[7] cb_5_7/io_wo[8] cb_5_7/io_wo[9]
+ cb_5_6/io_i_0_ci cb_5_6/io_i_0_in1[0] cb_5_6/io_i_0_in1[1] cb_5_6/io_i_0_in1[2]
+ cb_5_6/io_i_0_in1[3] cb_5_6/io_i_0_in1[4] cb_5_6/io_i_0_in1[5] cb_5_6/io_i_0_in1[6]
+ cb_5_6/io_i_0_in1[7] cb_5_6/io_i_1_ci cb_5_6/io_i_1_in1[0] cb_5_6/io_i_1_in1[1]
+ cb_5_6/io_i_1_in1[2] cb_5_6/io_i_1_in1[3] cb_5_6/io_i_1_in1[4] cb_5_6/io_i_1_in1[5]
+ cb_5_6/io_i_1_in1[6] cb_5_6/io_i_1_in1[7] cb_5_6/io_i_2_ci cb_5_6/io_i_2_in1[0]
+ cb_5_6/io_i_2_in1[1] cb_5_6/io_i_2_in1[2] cb_5_6/io_i_2_in1[3] cb_5_6/io_i_2_in1[4]
+ cb_5_6/io_i_2_in1[5] cb_5_6/io_i_2_in1[6] cb_5_6/io_i_2_in1[7] cb_5_6/io_i_3_ci
+ cb_5_6/io_i_3_in1[0] cb_5_6/io_i_3_in1[1] cb_5_6/io_i_3_in1[2] cb_5_6/io_i_3_in1[3]
+ cb_5_6/io_i_3_in1[4] cb_5_6/io_i_3_in1[5] cb_5_6/io_i_3_in1[6] cb_5_6/io_i_3_in1[7]
+ cb_5_6/io_i_4_ci cb_5_6/io_i_4_in1[0] cb_5_6/io_i_4_in1[1] cb_5_6/io_i_4_in1[2]
+ cb_5_6/io_i_4_in1[3] cb_5_6/io_i_4_in1[4] cb_5_6/io_i_4_in1[5] cb_5_6/io_i_4_in1[6]
+ cb_5_6/io_i_4_in1[7] cb_5_6/io_i_5_ci cb_5_6/io_i_5_in1[0] cb_5_6/io_i_5_in1[1]
+ cb_5_6/io_i_5_in1[2] cb_5_6/io_i_5_in1[3] cb_5_6/io_i_5_in1[4] cb_5_6/io_i_5_in1[5]
+ cb_5_6/io_i_5_in1[6] cb_5_6/io_i_5_in1[7] cb_5_6/io_i_6_ci cb_5_6/io_i_6_in1[0]
+ cb_5_6/io_i_6_in1[1] cb_5_6/io_i_6_in1[2] cb_5_6/io_i_6_in1[3] cb_5_6/io_i_6_in1[4]
+ cb_5_6/io_i_6_in1[5] cb_5_6/io_i_6_in1[6] cb_5_6/io_i_6_in1[7] cb_5_6/io_i_7_ci
+ cb_5_6/io_i_7_in1[0] cb_5_6/io_i_7_in1[1] cb_5_6/io_i_7_in1[2] cb_5_6/io_i_7_in1[3]
+ cb_5_6/io_i_7_in1[4] cb_5_6/io_i_7_in1[5] cb_5_6/io_i_7_in1[6] cb_5_6/io_i_7_in1[7]
+ cb_5_7/io_i_0_ci cb_5_7/io_i_0_in1[0] cb_5_7/io_i_0_in1[1] cb_5_7/io_i_0_in1[2]
+ cb_5_7/io_i_0_in1[3] cb_5_7/io_i_0_in1[4] cb_5_7/io_i_0_in1[5] cb_5_7/io_i_0_in1[6]
+ cb_5_7/io_i_0_in1[7] cb_5_7/io_i_1_ci cb_5_7/io_i_1_in1[0] cb_5_7/io_i_1_in1[1]
+ cb_5_7/io_i_1_in1[2] cb_5_7/io_i_1_in1[3] cb_5_7/io_i_1_in1[4] cb_5_7/io_i_1_in1[5]
+ cb_5_7/io_i_1_in1[6] cb_5_7/io_i_1_in1[7] cb_5_7/io_i_2_ci cb_5_7/io_i_2_in1[0]
+ cb_5_7/io_i_2_in1[1] cb_5_7/io_i_2_in1[2] cb_5_7/io_i_2_in1[3] cb_5_7/io_i_2_in1[4]
+ cb_5_7/io_i_2_in1[5] cb_5_7/io_i_2_in1[6] cb_5_7/io_i_2_in1[7] cb_5_7/io_i_3_ci
+ cb_5_7/io_i_3_in1[0] cb_5_7/io_i_3_in1[1] cb_5_7/io_i_3_in1[2] cb_5_7/io_i_3_in1[3]
+ cb_5_7/io_i_3_in1[4] cb_5_7/io_i_3_in1[5] cb_5_7/io_i_3_in1[6] cb_5_7/io_i_3_in1[7]
+ cb_5_7/io_i_4_ci cb_5_7/io_i_4_in1[0] cb_5_7/io_i_4_in1[1] cb_5_7/io_i_4_in1[2]
+ cb_5_7/io_i_4_in1[3] cb_5_7/io_i_4_in1[4] cb_5_7/io_i_4_in1[5] cb_5_7/io_i_4_in1[6]
+ cb_5_7/io_i_4_in1[7] cb_5_7/io_i_5_ci cb_5_7/io_i_5_in1[0] cb_5_7/io_i_5_in1[1]
+ cb_5_7/io_i_5_in1[2] cb_5_7/io_i_5_in1[3] cb_5_7/io_i_5_in1[4] cb_5_7/io_i_5_in1[5]
+ cb_5_7/io_i_5_in1[6] cb_5_7/io_i_5_in1[7] cb_5_7/io_i_6_ci cb_5_7/io_i_6_in1[0]
+ cb_5_7/io_i_6_in1[1] cb_5_7/io_i_6_in1[2] cb_5_7/io_i_6_in1[3] cb_5_7/io_i_6_in1[4]
+ cb_5_7/io_i_6_in1[5] cb_5_7/io_i_6_in1[6] cb_5_7/io_i_6_in1[7] cb_5_7/io_i_7_ci
+ cb_5_7/io_i_7_in1[0] cb_5_7/io_i_7_in1[1] cb_5_7/io_i_7_in1[2] cb_5_7/io_i_7_in1[3]
+ cb_5_7/io_i_7_in1[4] cb_5_7/io_i_7_in1[5] cb_5_7/io_i_7_in1[6] cb_5_7/io_i_7_in1[7]
+ cb_5_6/io_vci cb_5_7/io_vci cb_5_6/io_vi cb_5_9/io_we_i cb_5_6/io_wo[0] cb_5_6/io_wo[10]
+ cb_5_6/io_wo[11] cb_5_6/io_wo[12] cb_5_6/io_wo[13] cb_5_6/io_wo[14] cb_5_6/io_wo[15]
+ cb_5_6/io_wo[16] cb_5_6/io_wo[17] cb_5_6/io_wo[18] cb_5_6/io_wo[19] cb_5_6/io_wo[1]
+ cb_5_6/io_wo[20] cb_5_6/io_wo[21] cb_5_6/io_wo[22] cb_5_6/io_wo[23] cb_5_6/io_wo[24]
+ cb_5_6/io_wo[25] cb_5_6/io_wo[26] cb_5_6/io_wo[27] cb_5_6/io_wo[28] cb_5_6/io_wo[29]
+ cb_5_6/io_wo[2] cb_5_6/io_wo[30] cb_5_6/io_wo[31] cb_5_6/io_wo[32] cb_5_6/io_wo[33]
+ cb_5_6/io_wo[34] cb_5_6/io_wo[35] cb_5_6/io_wo[36] cb_5_6/io_wo[37] cb_5_6/io_wo[38]
+ cb_5_6/io_wo[39] cb_5_6/io_wo[3] cb_5_6/io_wo[40] cb_5_6/io_wo[41] cb_5_6/io_wo[42]
+ cb_5_6/io_wo[43] cb_5_6/io_wo[44] cb_5_6/io_wo[45] cb_5_6/io_wo[46] cb_5_6/io_wo[47]
+ cb_5_6/io_wo[48] cb_5_6/io_wo[49] cb_5_6/io_wo[4] cb_5_6/io_wo[50] cb_5_6/io_wo[51]
+ cb_5_6/io_wo[52] cb_5_6/io_wo[53] cb_5_6/io_wo[54] cb_5_6/io_wo[55] cb_5_6/io_wo[56]
+ cb_5_6/io_wo[57] cb_5_6/io_wo[58] cb_5_6/io_wo[59] cb_5_6/io_wo[5] cb_5_6/io_wo[60]
+ cb_5_6/io_wo[61] cb_5_6/io_wo[62] cb_5_6/io_wo[63] cb_5_6/io_wo[6] cb_5_6/io_wo[7]
+ cb_5_6/io_wo[8] cb_5_6/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xccon_2 ccon_2/io_ack_o ccon_7/io_adr_i[0] ccon_7/io_adr_i[10] ccon_7/io_adr_i[11]
+ ccon_7/io_adr_i[1] ccon_7/io_adr_i[2] ccon_7/io_adr_i[3] ccon_7/io_adr_i[4] ccon_7/io_adr_i[5]
+ ccon_7/io_adr_i[6] ccon_7/io_adr_i[7] ccon_7/io_adr_i[8] ccon_7/io_adr_i[9] cb_2_9/io_adr_i[0]
+ cb_2_9/io_adr_i[1] cb_2_0/io_cs_i cb_2_1/io_cs_i cb_2_10/io_cs_i cb_2_2/io_cs_i
+ cb_2_3/io_cs_i cb_2_4/io_cs_i cb_2_5/io_cs_i cb_2_6/io_cs_i cb_2_7/io_cs_i cb_2_8/io_cs_i
+ cb_2_9/io_cs_i cb_2_9/io_dat_i[0] cb_2_9/io_dat_i[10] cb_2_9/io_dat_i[11] cb_2_9/io_dat_i[12]
+ cb_2_9/io_dat_i[13] cb_2_9/io_dat_i[14] cb_2_9/io_dat_i[15] cb_2_9/io_dat_i[1] cb_2_9/io_dat_i[2]
+ cb_2_9/io_dat_i[3] cb_2_9/io_dat_i[4] cb_2_9/io_dat_i[5] cb_2_9/io_dat_i[6] cb_2_9/io_dat_i[7]
+ cb_2_9/io_dat_i[8] cb_2_9/io_dat_i[9] cb_2_0/io_dat_o[0] cb_2_0/io_dat_o[10] cb_2_0/io_dat_o[11]
+ cb_2_0/io_dat_o[12] cb_2_0/io_dat_o[13] cb_2_0/io_dat_o[14] cb_2_0/io_dat_o[15]
+ cb_2_0/io_dat_o[1] cb_2_0/io_dat_o[2] cb_2_0/io_dat_o[3] cb_2_0/io_dat_o[4] cb_2_0/io_dat_o[5]
+ cb_2_0/io_dat_o[6] cb_2_0/io_dat_o[7] cb_2_0/io_dat_o[8] cb_2_0/io_dat_o[9] cb_2_10/io_dat_o[0]
+ cb_2_10/io_dat_o[10] cb_2_10/io_dat_o[11] cb_2_10/io_dat_o[12] cb_2_10/io_dat_o[13]
+ cb_2_10/io_dat_o[14] cb_2_10/io_dat_o[15] cb_2_10/io_dat_o[1] cb_2_10/io_dat_o[2]
+ cb_2_10/io_dat_o[3] cb_2_10/io_dat_o[4] cb_2_10/io_dat_o[5] cb_2_10/io_dat_o[6]
+ cb_2_10/io_dat_o[7] cb_2_10/io_dat_o[8] cb_2_10/io_dat_o[9] cb_2_1/io_dat_o[0] cb_2_1/io_dat_o[10]
+ cb_2_1/io_dat_o[11] cb_2_1/io_dat_o[12] cb_2_1/io_dat_o[13] cb_2_1/io_dat_o[14]
+ cb_2_1/io_dat_o[15] cb_2_1/io_dat_o[1] cb_2_1/io_dat_o[2] cb_2_1/io_dat_o[3] cb_2_1/io_dat_o[4]
+ cb_2_1/io_dat_o[5] cb_2_1/io_dat_o[6] cb_2_1/io_dat_o[7] cb_2_1/io_dat_o[8] cb_2_1/io_dat_o[9]
+ cb_2_2/io_dat_o[0] cb_2_2/io_dat_o[10] cb_2_2/io_dat_o[11] cb_2_2/io_dat_o[12] cb_2_2/io_dat_o[13]
+ cb_2_2/io_dat_o[14] cb_2_2/io_dat_o[15] cb_2_2/io_dat_o[1] cb_2_2/io_dat_o[2] cb_2_2/io_dat_o[3]
+ cb_2_2/io_dat_o[4] cb_2_2/io_dat_o[5] cb_2_2/io_dat_o[6] cb_2_2/io_dat_o[7] cb_2_2/io_dat_o[8]
+ cb_2_2/io_dat_o[9] cb_2_3/io_dat_o[0] cb_2_3/io_dat_o[10] cb_2_3/io_dat_o[11] cb_2_3/io_dat_o[12]
+ cb_2_3/io_dat_o[13] cb_2_3/io_dat_o[14] cb_2_3/io_dat_o[15] cb_2_3/io_dat_o[1] cb_2_3/io_dat_o[2]
+ cb_2_3/io_dat_o[3] cb_2_3/io_dat_o[4] cb_2_3/io_dat_o[5] cb_2_3/io_dat_o[6] cb_2_3/io_dat_o[7]
+ cb_2_3/io_dat_o[8] cb_2_3/io_dat_o[9] cb_2_4/io_dat_o[0] cb_2_4/io_dat_o[10] cb_2_4/io_dat_o[11]
+ cb_2_4/io_dat_o[12] cb_2_4/io_dat_o[13] cb_2_4/io_dat_o[14] cb_2_4/io_dat_o[15]
+ cb_2_4/io_dat_o[1] cb_2_4/io_dat_o[2] cb_2_4/io_dat_o[3] cb_2_4/io_dat_o[4] cb_2_4/io_dat_o[5]
+ cb_2_4/io_dat_o[6] cb_2_4/io_dat_o[7] cb_2_4/io_dat_o[8] cb_2_4/io_dat_o[9] cb_2_5/io_dat_o[0]
+ cb_2_5/io_dat_o[10] cb_2_5/io_dat_o[11] cb_2_5/io_dat_o[12] cb_2_5/io_dat_o[13]
+ cb_2_5/io_dat_o[14] cb_2_5/io_dat_o[15] cb_2_5/io_dat_o[1] cb_2_5/io_dat_o[2] cb_2_5/io_dat_o[3]
+ cb_2_5/io_dat_o[4] cb_2_5/io_dat_o[5] cb_2_5/io_dat_o[6] cb_2_5/io_dat_o[7] cb_2_5/io_dat_o[8]
+ cb_2_5/io_dat_o[9] cb_2_6/io_dat_o[0] cb_2_6/io_dat_o[10] cb_2_6/io_dat_o[11] cb_2_6/io_dat_o[12]
+ cb_2_6/io_dat_o[13] cb_2_6/io_dat_o[14] cb_2_6/io_dat_o[15] cb_2_6/io_dat_o[1] cb_2_6/io_dat_o[2]
+ cb_2_6/io_dat_o[3] cb_2_6/io_dat_o[4] cb_2_6/io_dat_o[5] cb_2_6/io_dat_o[6] cb_2_6/io_dat_o[7]
+ cb_2_6/io_dat_o[8] cb_2_6/io_dat_o[9] cb_2_7/io_dat_o[0] cb_2_7/io_dat_o[10] cb_2_7/io_dat_o[11]
+ cb_2_7/io_dat_o[12] cb_2_7/io_dat_o[13] cb_2_7/io_dat_o[14] cb_2_7/io_dat_o[15]
+ cb_2_7/io_dat_o[1] cb_2_7/io_dat_o[2] cb_2_7/io_dat_o[3] cb_2_7/io_dat_o[4] cb_2_7/io_dat_o[5]
+ cb_2_7/io_dat_o[6] cb_2_7/io_dat_o[7] cb_2_7/io_dat_o[8] cb_2_7/io_dat_o[9] cb_2_8/io_dat_o[0]
+ cb_2_8/io_dat_o[10] cb_2_8/io_dat_o[11] cb_2_8/io_dat_o[12] cb_2_8/io_dat_o[13]
+ cb_2_8/io_dat_o[14] cb_2_8/io_dat_o[15] cb_2_8/io_dat_o[1] cb_2_8/io_dat_o[2] cb_2_8/io_dat_o[3]
+ cb_2_8/io_dat_o[4] cb_2_8/io_dat_o[5] cb_2_8/io_dat_o[6] cb_2_8/io_dat_o[7] cb_2_8/io_dat_o[8]
+ cb_2_8/io_dat_o[9] cb_2_9/io_dat_o[0] cb_2_9/io_dat_o[10] cb_2_9/io_dat_o[11] cb_2_9/io_dat_o[12]
+ cb_2_9/io_dat_o[13] cb_2_9/io_dat_o[14] cb_2_9/io_dat_o[15] cb_2_9/io_dat_o[1] cb_2_9/io_dat_o[2]
+ cb_2_9/io_dat_o[3] cb_2_9/io_dat_o[4] cb_2_9/io_dat_o[5] cb_2_9/io_dat_o[6] cb_2_9/io_dat_o[7]
+ cb_2_9/io_dat_o[8] cb_2_9/io_dat_o[9] cb_2_9/io_we_i ccon_2/io_cs_i ccon_7/io_dat_i[0]
+ ccon_7/io_dat_i[10] ccon_7/io_dat_i[11] ccon_7/io_dat_i[12] ccon_7/io_dat_i[13]
+ ccon_7/io_dat_i[14] ccon_7/io_dat_i[15] ccon_7/io_dat_i[16] ccon_7/io_dat_i[17]
+ ccon_7/io_dat_i[18] ccon_7/io_dat_i[19] ccon_7/io_dat_i[1] ccon_7/io_dat_i[20] ccon_7/io_dat_i[21]
+ ccon_7/io_dat_i[22] ccon_7/io_dat_i[23] ccon_7/io_dat_i[24] ccon_7/io_dat_i[25]
+ ccon_7/io_dat_i[26] ccon_7/io_dat_i[27] ccon_7/io_dat_i[28] ccon_7/io_dat_i[29]
+ ccon_7/io_dat_i[2] ccon_7/io_dat_i[30] ccon_7/io_dat_i[31] ccon_7/io_dat_i[3] ccon_7/io_dat_i[4]
+ ccon_7/io_dat_i[5] ccon_7/io_dat_i[6] ccon_7/io_dat_i[7] ccon_7/io_dat_i[8] ccon_7/io_dat_i[9]
+ ccon_2/io_dat_o[0] ccon_2/io_dat_o[10] ccon_2/io_dat_o[11] ccon_2/io_dat_o[12] ccon_2/io_dat_o[13]
+ ccon_2/io_dat_o[14] ccon_2/io_dat_o[15] ccon_2/io_dat_o[16] ccon_2/io_dat_o[17]
+ ccon_2/io_dat_o[18] ccon_2/io_dat_o[19] ccon_2/io_dat_o[1] ccon_2/io_dat_o[20] ccon_2/io_dat_o[21]
+ ccon_2/io_dat_o[22] ccon_2/io_dat_o[23] ccon_2/io_dat_o[24] ccon_2/io_dat_o[25]
+ ccon_2/io_dat_o[26] ccon_2/io_dat_o[27] ccon_2/io_dat_o[28] ccon_2/io_dat_o[29]
+ ccon_2/io_dat_o[2] ccon_2/io_dat_o[30] ccon_2/io_dat_o[31] ccon_2/io_dat_o[3] ccon_2/io_dat_o[4]
+ ccon_2/io_dat_o[5] ccon_2/io_dat_o[6] ccon_2/io_dat_o[7] ccon_2/io_dat_o[8] ccon_2/io_dat_o[9]
+ cb_2_0/io_wo[0] cb_2_0/io_wo[10] cb_2_0/io_wo[11] cb_2_0/io_wo[12] cb_2_0/io_wo[13]
+ cb_2_0/io_wo[14] cb_2_0/io_wo[15] cb_2_0/io_wo[16] cb_2_0/io_wo[17] cb_2_0/io_wo[18]
+ cb_2_0/io_wo[19] cb_2_0/io_wo[1] cb_2_0/io_wo[20] cb_2_0/io_wo[21] cb_2_0/io_wo[22]
+ cb_2_0/io_wo[23] cb_2_0/io_wo[24] cb_2_0/io_wo[25] cb_2_0/io_wo[26] cb_2_0/io_wo[27]
+ cb_2_0/io_wo[28] cb_2_0/io_wo[29] cb_2_0/io_wo[2] cb_2_0/io_wo[30] cb_2_0/io_wo[31]
+ cb_2_0/io_wo[32] cb_2_0/io_wo[33] cb_2_0/io_wo[34] cb_2_0/io_wo[35] cb_2_0/io_wo[36]
+ cb_2_0/io_wo[37] cb_2_0/io_wo[38] cb_2_0/io_wo[39] cb_2_0/io_wo[3] cb_2_0/io_wo[40]
+ cb_2_0/io_wo[41] cb_2_0/io_wo[42] cb_2_0/io_wo[43] cb_2_0/io_wo[44] cb_2_0/io_wo[45]
+ cb_2_0/io_wo[46] cb_2_0/io_wo[47] cb_2_0/io_wo[48] cb_2_0/io_wo[49] cb_2_0/io_wo[4]
+ cb_2_0/io_wo[50] cb_2_0/io_wo[51] cb_2_0/io_wo[52] cb_2_0/io_wo[53] cb_2_0/io_wo[54]
+ cb_2_0/io_wo[55] cb_2_0/io_wo[56] cb_2_0/io_wo[57] cb_2_0/io_wo[58] cb_2_0/io_wo[59]
+ cb_2_0/io_wo[5] cb_2_0/io_wo[60] cb_2_0/io_wo[61] cb_2_0/io_wo[62] cb_2_0/io_wo[63]
+ cb_2_0/io_wo[6] cb_2_0/io_wo[7] cb_2_0/io_wo[8] cb_2_0/io_wo[9] icon/dsi[0] icon/dsi[1]
+ icon/dsi[2] icon/dsi[3] icon/dsi[4] icon/dsi[5] icon/dsi[6] icon/dsi[7] ccon_2/io_dsi_o
+ ccon_2/io_irq cb_2_0/io_vi cb_2_10/io_vi cb_2_1/io_vi cb_2_2/io_vi cb_2_3/io_vi
+ cb_2_4/io_vi cb_2_5/io_vi cb_2_6/io_vi cb_2_7/io_vi cb_2_8/io_vi cb_2_9/io_vi ccon_7/io_we_i
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_con
Xcb_3_3 cb_3_9/io_adr_i[0] cb_3_9/io_adr_i[1] cb_3_3/io_cs_i cb_3_9/io_dat_i[0] cb_3_9/io_dat_i[10]
+ cb_3_9/io_dat_i[11] cb_3_9/io_dat_i[12] cb_3_9/io_dat_i[13] cb_3_9/io_dat_i[14]
+ cb_3_9/io_dat_i[15] cb_3_9/io_dat_i[1] cb_3_9/io_dat_i[2] cb_3_9/io_dat_i[3] cb_3_9/io_dat_i[4]
+ cb_3_9/io_dat_i[5] cb_3_9/io_dat_i[6] cb_3_9/io_dat_i[7] cb_3_9/io_dat_i[8] cb_3_9/io_dat_i[9]
+ cb_3_3/io_dat_o[0] cb_3_3/io_dat_o[10] cb_3_3/io_dat_o[11] cb_3_3/io_dat_o[12] cb_3_3/io_dat_o[13]
+ cb_3_3/io_dat_o[14] cb_3_3/io_dat_o[15] cb_3_3/io_dat_o[1] cb_3_3/io_dat_o[2] cb_3_3/io_dat_o[3]
+ cb_3_3/io_dat_o[4] cb_3_3/io_dat_o[5] cb_3_3/io_dat_o[6] cb_3_3/io_dat_o[7] cb_3_3/io_dat_o[8]
+ cb_3_3/io_dat_o[9] cb_3_4/io_wo[0] cb_3_4/io_wo[10] cb_3_4/io_wo[11] cb_3_4/io_wo[12]
+ cb_3_4/io_wo[13] cb_3_4/io_wo[14] cb_3_4/io_wo[15] cb_3_4/io_wo[16] cb_3_4/io_wo[17]
+ cb_3_4/io_wo[18] cb_3_4/io_wo[19] cb_3_4/io_wo[1] cb_3_4/io_wo[20] cb_3_4/io_wo[21]
+ cb_3_4/io_wo[22] cb_3_4/io_wo[23] cb_3_4/io_wo[24] cb_3_4/io_wo[25] cb_3_4/io_wo[26]
+ cb_3_4/io_wo[27] cb_3_4/io_wo[28] cb_3_4/io_wo[29] cb_3_4/io_wo[2] cb_3_4/io_wo[30]
+ cb_3_4/io_wo[31] cb_3_4/io_wo[32] cb_3_4/io_wo[33] cb_3_4/io_wo[34] cb_3_4/io_wo[35]
+ cb_3_4/io_wo[36] cb_3_4/io_wo[37] cb_3_4/io_wo[38] cb_3_4/io_wo[39] cb_3_4/io_wo[3]
+ cb_3_4/io_wo[40] cb_3_4/io_wo[41] cb_3_4/io_wo[42] cb_3_4/io_wo[43] cb_3_4/io_wo[44]
+ cb_3_4/io_wo[45] cb_3_4/io_wo[46] cb_3_4/io_wo[47] cb_3_4/io_wo[48] cb_3_4/io_wo[49]
+ cb_3_4/io_wo[4] cb_3_4/io_wo[50] cb_3_4/io_wo[51] cb_3_4/io_wo[52] cb_3_4/io_wo[53]
+ cb_3_4/io_wo[54] cb_3_4/io_wo[55] cb_3_4/io_wo[56] cb_3_4/io_wo[57] cb_3_4/io_wo[58]
+ cb_3_4/io_wo[59] cb_3_4/io_wo[5] cb_3_4/io_wo[60] cb_3_4/io_wo[61] cb_3_4/io_wo[62]
+ cb_3_4/io_wo[63] cb_3_4/io_wo[6] cb_3_4/io_wo[7] cb_3_4/io_wo[8] cb_3_4/io_wo[9]
+ cb_3_3/io_i_0_ci cb_3_3/io_i_0_in1[0] cb_3_3/io_i_0_in1[1] cb_3_3/io_i_0_in1[2]
+ cb_3_3/io_i_0_in1[3] cb_3_3/io_i_0_in1[4] cb_3_3/io_i_0_in1[5] cb_3_3/io_i_0_in1[6]
+ cb_3_3/io_i_0_in1[7] cb_3_3/io_i_1_ci cb_3_3/io_i_1_in1[0] cb_3_3/io_i_1_in1[1]
+ cb_3_3/io_i_1_in1[2] cb_3_3/io_i_1_in1[3] cb_3_3/io_i_1_in1[4] cb_3_3/io_i_1_in1[5]
+ cb_3_3/io_i_1_in1[6] cb_3_3/io_i_1_in1[7] cb_3_3/io_i_2_ci cb_3_3/io_i_2_in1[0]
+ cb_3_3/io_i_2_in1[1] cb_3_3/io_i_2_in1[2] cb_3_3/io_i_2_in1[3] cb_3_3/io_i_2_in1[4]
+ cb_3_3/io_i_2_in1[5] cb_3_3/io_i_2_in1[6] cb_3_3/io_i_2_in1[7] cb_3_3/io_i_3_ci
+ cb_3_3/io_i_3_in1[0] cb_3_3/io_i_3_in1[1] cb_3_3/io_i_3_in1[2] cb_3_3/io_i_3_in1[3]
+ cb_3_3/io_i_3_in1[4] cb_3_3/io_i_3_in1[5] cb_3_3/io_i_3_in1[6] cb_3_3/io_i_3_in1[7]
+ cb_3_3/io_i_4_ci cb_3_3/io_i_4_in1[0] cb_3_3/io_i_4_in1[1] cb_3_3/io_i_4_in1[2]
+ cb_3_3/io_i_4_in1[3] cb_3_3/io_i_4_in1[4] cb_3_3/io_i_4_in1[5] cb_3_3/io_i_4_in1[6]
+ cb_3_3/io_i_4_in1[7] cb_3_3/io_i_5_ci cb_3_3/io_i_5_in1[0] cb_3_3/io_i_5_in1[1]
+ cb_3_3/io_i_5_in1[2] cb_3_3/io_i_5_in1[3] cb_3_3/io_i_5_in1[4] cb_3_3/io_i_5_in1[5]
+ cb_3_3/io_i_5_in1[6] cb_3_3/io_i_5_in1[7] cb_3_3/io_i_6_ci cb_3_3/io_i_6_in1[0]
+ cb_3_3/io_i_6_in1[1] cb_3_3/io_i_6_in1[2] cb_3_3/io_i_6_in1[3] cb_3_3/io_i_6_in1[4]
+ cb_3_3/io_i_6_in1[5] cb_3_3/io_i_6_in1[6] cb_3_3/io_i_6_in1[7] cb_3_3/io_i_7_ci
+ cb_3_3/io_i_7_in1[0] cb_3_3/io_i_7_in1[1] cb_3_3/io_i_7_in1[2] cb_3_3/io_i_7_in1[3]
+ cb_3_3/io_i_7_in1[4] cb_3_3/io_i_7_in1[5] cb_3_3/io_i_7_in1[6] cb_3_3/io_i_7_in1[7]
+ cb_3_4/io_i_0_ci cb_3_4/io_i_0_in1[0] cb_3_4/io_i_0_in1[1] cb_3_4/io_i_0_in1[2]
+ cb_3_4/io_i_0_in1[3] cb_3_4/io_i_0_in1[4] cb_3_4/io_i_0_in1[5] cb_3_4/io_i_0_in1[6]
+ cb_3_4/io_i_0_in1[7] cb_3_4/io_i_1_ci cb_3_4/io_i_1_in1[0] cb_3_4/io_i_1_in1[1]
+ cb_3_4/io_i_1_in1[2] cb_3_4/io_i_1_in1[3] cb_3_4/io_i_1_in1[4] cb_3_4/io_i_1_in1[5]
+ cb_3_4/io_i_1_in1[6] cb_3_4/io_i_1_in1[7] cb_3_4/io_i_2_ci cb_3_4/io_i_2_in1[0]
+ cb_3_4/io_i_2_in1[1] cb_3_4/io_i_2_in1[2] cb_3_4/io_i_2_in1[3] cb_3_4/io_i_2_in1[4]
+ cb_3_4/io_i_2_in1[5] cb_3_4/io_i_2_in1[6] cb_3_4/io_i_2_in1[7] cb_3_4/io_i_3_ci
+ cb_3_4/io_i_3_in1[0] cb_3_4/io_i_3_in1[1] cb_3_4/io_i_3_in1[2] cb_3_4/io_i_3_in1[3]
+ cb_3_4/io_i_3_in1[4] cb_3_4/io_i_3_in1[5] cb_3_4/io_i_3_in1[6] cb_3_4/io_i_3_in1[7]
+ cb_3_4/io_i_4_ci cb_3_4/io_i_4_in1[0] cb_3_4/io_i_4_in1[1] cb_3_4/io_i_4_in1[2]
+ cb_3_4/io_i_4_in1[3] cb_3_4/io_i_4_in1[4] cb_3_4/io_i_4_in1[5] cb_3_4/io_i_4_in1[6]
+ cb_3_4/io_i_4_in1[7] cb_3_4/io_i_5_ci cb_3_4/io_i_5_in1[0] cb_3_4/io_i_5_in1[1]
+ cb_3_4/io_i_5_in1[2] cb_3_4/io_i_5_in1[3] cb_3_4/io_i_5_in1[4] cb_3_4/io_i_5_in1[5]
+ cb_3_4/io_i_5_in1[6] cb_3_4/io_i_5_in1[7] cb_3_4/io_i_6_ci cb_3_4/io_i_6_in1[0]
+ cb_3_4/io_i_6_in1[1] cb_3_4/io_i_6_in1[2] cb_3_4/io_i_6_in1[3] cb_3_4/io_i_6_in1[4]
+ cb_3_4/io_i_6_in1[5] cb_3_4/io_i_6_in1[6] cb_3_4/io_i_6_in1[7] cb_3_4/io_i_7_ci
+ cb_3_4/io_i_7_in1[0] cb_3_4/io_i_7_in1[1] cb_3_4/io_i_7_in1[2] cb_3_4/io_i_7_in1[3]
+ cb_3_4/io_i_7_in1[4] cb_3_4/io_i_7_in1[5] cb_3_4/io_i_7_in1[6] cb_3_4/io_i_7_in1[7]
+ cb_3_3/io_vci cb_3_4/io_vci cb_3_3/io_vi cb_3_9/io_we_i cb_3_3/io_wo[0] cb_3_3/io_wo[10]
+ cb_3_3/io_wo[11] cb_3_3/io_wo[12] cb_3_3/io_wo[13] cb_3_3/io_wo[14] cb_3_3/io_wo[15]
+ cb_3_3/io_wo[16] cb_3_3/io_wo[17] cb_3_3/io_wo[18] cb_3_3/io_wo[19] cb_3_3/io_wo[1]
+ cb_3_3/io_wo[20] cb_3_3/io_wo[21] cb_3_3/io_wo[22] cb_3_3/io_wo[23] cb_3_3/io_wo[24]
+ cb_3_3/io_wo[25] cb_3_3/io_wo[26] cb_3_3/io_wo[27] cb_3_3/io_wo[28] cb_3_3/io_wo[29]
+ cb_3_3/io_wo[2] cb_3_3/io_wo[30] cb_3_3/io_wo[31] cb_3_3/io_wo[32] cb_3_3/io_wo[33]
+ cb_3_3/io_wo[34] cb_3_3/io_wo[35] cb_3_3/io_wo[36] cb_3_3/io_wo[37] cb_3_3/io_wo[38]
+ cb_3_3/io_wo[39] cb_3_3/io_wo[3] cb_3_3/io_wo[40] cb_3_3/io_wo[41] cb_3_3/io_wo[42]
+ cb_3_3/io_wo[43] cb_3_3/io_wo[44] cb_3_3/io_wo[45] cb_3_3/io_wo[46] cb_3_3/io_wo[47]
+ cb_3_3/io_wo[48] cb_3_3/io_wo[49] cb_3_3/io_wo[4] cb_3_3/io_wo[50] cb_3_3/io_wo[51]
+ cb_3_3/io_wo[52] cb_3_3/io_wo[53] cb_3_3/io_wo[54] cb_3_3/io_wo[55] cb_3_3/io_wo[56]
+ cb_3_3/io_wo[57] cb_3_3/io_wo[58] cb_3_3/io_wo[59] cb_3_3/io_wo[5] cb_3_3/io_wo[60]
+ cb_3_3/io_wo[61] cb_3_3/io_wo[62] cb_3_3/io_wo[63] cb_3_3/io_wo[6] cb_3_3/io_wo[7]
+ cb_3_3/io_wo[8] cb_3_3/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_1_0 cb_1_9/io_adr_i[0] cb_1_9/io_adr_i[1] cb_1_0/io_cs_i cb_1_9/io_dat_i[0] cb_1_9/io_dat_i[10]
+ cb_1_9/io_dat_i[11] cb_1_9/io_dat_i[12] cb_1_9/io_dat_i[13] cb_1_9/io_dat_i[14]
+ cb_1_9/io_dat_i[15] cb_1_9/io_dat_i[1] cb_1_9/io_dat_i[2] cb_1_9/io_dat_i[3] cb_1_9/io_dat_i[4]
+ cb_1_9/io_dat_i[5] cb_1_9/io_dat_i[6] cb_1_9/io_dat_i[7] cb_1_9/io_dat_i[8] cb_1_9/io_dat_i[9]
+ cb_1_0/io_dat_o[0] cb_1_0/io_dat_o[10] cb_1_0/io_dat_o[11] cb_1_0/io_dat_o[12] cb_1_0/io_dat_o[13]
+ cb_1_0/io_dat_o[14] cb_1_0/io_dat_o[15] cb_1_0/io_dat_o[1] cb_1_0/io_dat_o[2] cb_1_0/io_dat_o[3]
+ cb_1_0/io_dat_o[4] cb_1_0/io_dat_o[5] cb_1_0/io_dat_o[6] cb_1_0/io_dat_o[7] cb_1_0/io_dat_o[8]
+ cb_1_0/io_dat_o[9] cb_1_1/io_wo[0] cb_1_1/io_wo[10] cb_1_1/io_wo[11] cb_1_1/io_wo[12]
+ cb_1_1/io_wo[13] cb_1_1/io_wo[14] cb_1_1/io_wo[15] cb_1_1/io_wo[16] cb_1_1/io_wo[17]
+ cb_1_1/io_wo[18] cb_1_1/io_wo[19] cb_1_1/io_wo[1] cb_1_1/io_wo[20] cb_1_1/io_wo[21]
+ cb_1_1/io_wo[22] cb_1_1/io_wo[23] cb_1_1/io_wo[24] cb_1_1/io_wo[25] cb_1_1/io_wo[26]
+ cb_1_1/io_wo[27] cb_1_1/io_wo[28] cb_1_1/io_wo[29] cb_1_1/io_wo[2] cb_1_1/io_wo[30]
+ cb_1_1/io_wo[31] cb_1_1/io_wo[32] cb_1_1/io_wo[33] cb_1_1/io_wo[34] cb_1_1/io_wo[35]
+ cb_1_1/io_wo[36] cb_1_1/io_wo[37] cb_1_1/io_wo[38] cb_1_1/io_wo[39] cb_1_1/io_wo[3]
+ cb_1_1/io_wo[40] cb_1_1/io_wo[41] cb_1_1/io_wo[42] cb_1_1/io_wo[43] cb_1_1/io_wo[44]
+ cb_1_1/io_wo[45] cb_1_1/io_wo[46] cb_1_1/io_wo[47] cb_1_1/io_wo[48] cb_1_1/io_wo[49]
+ cb_1_1/io_wo[4] cb_1_1/io_wo[50] cb_1_1/io_wo[51] cb_1_1/io_wo[52] cb_1_1/io_wo[53]
+ cb_1_1/io_wo[54] cb_1_1/io_wo[55] cb_1_1/io_wo[56] cb_1_1/io_wo[57] cb_1_1/io_wo[58]
+ cb_1_1/io_wo[59] cb_1_1/io_wo[5] cb_1_1/io_wo[60] cb_1_1/io_wo[61] cb_1_1/io_wo[62]
+ cb_1_1/io_wo[63] cb_1_1/io_wo[6] cb_1_1/io_wo[7] cb_1_1/io_wo[8] cb_1_1/io_wo[9]
+ ccon_1/io_dsi_o cb_1_0/io_i_0_in1[0] cb_1_0/io_i_0_in1[1] cb_1_0/io_i_0_in1[2] cb_1_0/io_i_0_in1[3]
+ cb_1_0/io_i_0_in1[4] cb_1_0/io_i_0_in1[5] cb_1_0/io_i_0_in1[6] cb_1_0/io_i_0_in1[7]
+ cb_1_0/io_i_1_ci cb_1_0/io_i_1_in1[0] cb_1_0/io_i_1_in1[1] cb_1_0/io_i_1_in1[2]
+ cb_1_0/io_i_1_in1[3] cb_1_0/io_i_1_in1[4] cb_1_0/io_i_1_in1[5] cb_1_0/io_i_1_in1[6]
+ cb_1_0/io_i_1_in1[7] cb_1_0/io_i_2_ci cb_1_0/io_i_2_in1[0] cb_1_0/io_i_2_in1[1]
+ cb_1_0/io_i_2_in1[2] cb_1_0/io_i_2_in1[3] cb_1_0/io_i_2_in1[4] cb_1_0/io_i_2_in1[5]
+ cb_1_0/io_i_2_in1[6] cb_1_0/io_i_2_in1[7] cb_1_0/io_i_3_ci cb_1_0/io_i_3_in1[0]
+ cb_1_0/io_i_3_in1[1] cb_1_0/io_i_3_in1[2] cb_1_0/io_i_3_in1[3] cb_1_0/io_i_3_in1[4]
+ cb_1_0/io_i_3_in1[5] cb_1_0/io_i_3_in1[6] cb_1_0/io_i_3_in1[7] cb_1_0/io_i_4_ci
+ cb_1_0/io_i_4_in1[0] cb_1_0/io_i_4_in1[1] cb_1_0/io_i_4_in1[2] cb_1_0/io_i_4_in1[3]
+ cb_1_0/io_i_4_in1[4] cb_1_0/io_i_4_in1[5] cb_1_0/io_i_4_in1[6] cb_1_0/io_i_4_in1[7]
+ cb_1_0/io_i_5_ci cb_1_0/io_i_5_in1[0] cb_1_0/io_i_5_in1[1] cb_1_0/io_i_5_in1[2]
+ cb_1_0/io_i_5_in1[3] cb_1_0/io_i_5_in1[4] cb_1_0/io_i_5_in1[5] cb_1_0/io_i_5_in1[6]
+ cb_1_0/io_i_5_in1[7] cb_1_0/io_i_6_ci cb_1_0/io_i_6_in1[0] cb_1_0/io_i_6_in1[1]
+ cb_1_0/io_i_6_in1[2] cb_1_0/io_i_6_in1[3] cb_1_0/io_i_6_in1[4] cb_1_0/io_i_6_in1[5]
+ cb_1_0/io_i_6_in1[6] cb_1_0/io_i_6_in1[7] cb_1_0/io_i_7_ci cb_1_0/io_i_7_in1[0]
+ cb_1_0/io_i_7_in1[1] cb_1_0/io_i_7_in1[2] cb_1_0/io_i_7_in1[3] cb_1_0/io_i_7_in1[4]
+ cb_1_0/io_i_7_in1[5] cb_1_0/io_i_7_in1[6] cb_1_0/io_i_7_in1[7] cb_1_1/io_i_0_ci
+ cb_1_1/io_i_0_in1[0] cb_1_1/io_i_0_in1[1] cb_1_1/io_i_0_in1[2] cb_1_1/io_i_0_in1[3]
+ cb_1_1/io_i_0_in1[4] cb_1_1/io_i_0_in1[5] cb_1_1/io_i_0_in1[6] cb_1_1/io_i_0_in1[7]
+ cb_1_1/io_i_1_ci cb_1_1/io_i_1_in1[0] cb_1_1/io_i_1_in1[1] cb_1_1/io_i_1_in1[2]
+ cb_1_1/io_i_1_in1[3] cb_1_1/io_i_1_in1[4] cb_1_1/io_i_1_in1[5] cb_1_1/io_i_1_in1[6]
+ cb_1_1/io_i_1_in1[7] cb_1_1/io_i_2_ci cb_1_1/io_i_2_in1[0] cb_1_1/io_i_2_in1[1]
+ cb_1_1/io_i_2_in1[2] cb_1_1/io_i_2_in1[3] cb_1_1/io_i_2_in1[4] cb_1_1/io_i_2_in1[5]
+ cb_1_1/io_i_2_in1[6] cb_1_1/io_i_2_in1[7] cb_1_1/io_i_3_ci cb_1_1/io_i_3_in1[0]
+ cb_1_1/io_i_3_in1[1] cb_1_1/io_i_3_in1[2] cb_1_1/io_i_3_in1[3] cb_1_1/io_i_3_in1[4]
+ cb_1_1/io_i_3_in1[5] cb_1_1/io_i_3_in1[6] cb_1_1/io_i_3_in1[7] cb_1_1/io_i_4_ci
+ cb_1_1/io_i_4_in1[0] cb_1_1/io_i_4_in1[1] cb_1_1/io_i_4_in1[2] cb_1_1/io_i_4_in1[3]
+ cb_1_1/io_i_4_in1[4] cb_1_1/io_i_4_in1[5] cb_1_1/io_i_4_in1[6] cb_1_1/io_i_4_in1[7]
+ cb_1_1/io_i_5_ci cb_1_1/io_i_5_in1[0] cb_1_1/io_i_5_in1[1] cb_1_1/io_i_5_in1[2]
+ cb_1_1/io_i_5_in1[3] cb_1_1/io_i_5_in1[4] cb_1_1/io_i_5_in1[5] cb_1_1/io_i_5_in1[6]
+ cb_1_1/io_i_5_in1[7] cb_1_1/io_i_6_ci cb_1_1/io_i_6_in1[0] cb_1_1/io_i_6_in1[1]
+ cb_1_1/io_i_6_in1[2] cb_1_1/io_i_6_in1[3] cb_1_1/io_i_6_in1[4] cb_1_1/io_i_6_in1[5]
+ cb_1_1/io_i_6_in1[6] cb_1_1/io_i_6_in1[7] cb_1_1/io_i_7_ci cb_1_1/io_i_7_in1[0]
+ cb_1_1/io_i_7_in1[1] cb_1_1/io_i_7_in1[2] cb_1_1/io_i_7_in1[3] cb_1_1/io_i_7_in1[4]
+ cb_1_1/io_i_7_in1[5] cb_1_1/io_i_7_in1[6] cb_1_1/io_i_7_in1[7] cb_1_0/io_vci cb_1_1/io_vci
+ cb_1_0/io_vi cb_1_9/io_we_i cb_1_0/io_wo[0] cb_1_0/io_wo[10] cb_1_0/io_wo[11] cb_1_0/io_wo[12]
+ cb_1_0/io_wo[13] cb_1_0/io_wo[14] cb_1_0/io_wo[15] cb_1_0/io_wo[16] cb_1_0/io_wo[17]
+ cb_1_0/io_wo[18] cb_1_0/io_wo[19] cb_1_0/io_wo[1] cb_1_0/io_wo[20] cb_1_0/io_wo[21]
+ cb_1_0/io_wo[22] cb_1_0/io_wo[23] cb_1_0/io_wo[24] cb_1_0/io_wo[25] cb_1_0/io_wo[26]
+ cb_1_0/io_wo[27] cb_1_0/io_wo[28] cb_1_0/io_wo[29] cb_1_0/io_wo[2] cb_1_0/io_wo[30]
+ cb_1_0/io_wo[31] cb_1_0/io_wo[32] cb_1_0/io_wo[33] cb_1_0/io_wo[34] cb_1_0/io_wo[35]
+ cb_1_0/io_wo[36] cb_1_0/io_wo[37] cb_1_0/io_wo[38] cb_1_0/io_wo[39] cb_1_0/io_wo[3]
+ cb_1_0/io_wo[40] cb_1_0/io_wo[41] cb_1_0/io_wo[42] cb_1_0/io_wo[43] cb_1_0/io_wo[44]
+ cb_1_0/io_wo[45] cb_1_0/io_wo[46] cb_1_0/io_wo[47] cb_1_0/io_wo[48] cb_1_0/io_wo[49]
+ cb_1_0/io_wo[4] cb_1_0/io_wo[50] cb_1_0/io_wo[51] cb_1_0/io_wo[52] cb_1_0/io_wo[53]
+ cb_1_0/io_wo[54] cb_1_0/io_wo[55] cb_1_0/io_wo[56] cb_1_0/io_wo[57] cb_1_0/io_wo[58]
+ cb_1_0/io_wo[59] cb_1_0/io_wo[5] cb_1_0/io_wo[60] cb_1_0/io_wo[61] cb_1_0/io_wo[62]
+ cb_1_0/io_wo[63] cb_1_0/io_wo[6] cb_1_0/io_wo[7] cb_1_0/io_wo[8] cb_1_0/io_wo[9]
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xccon_3 ccon_3/io_ack_o ccon_7/io_adr_i[0] ccon_7/io_adr_i[10] ccon_7/io_adr_i[11]
+ ccon_7/io_adr_i[1] ccon_7/io_adr_i[2] ccon_7/io_adr_i[3] ccon_7/io_adr_i[4] ccon_7/io_adr_i[5]
+ ccon_7/io_adr_i[6] ccon_7/io_adr_i[7] ccon_7/io_adr_i[8] ccon_7/io_adr_i[9] cb_3_9/io_adr_i[0]
+ cb_3_9/io_adr_i[1] cb_3_0/io_cs_i cb_3_1/io_cs_i cb_3_10/io_cs_i cb_3_2/io_cs_i
+ cb_3_3/io_cs_i cb_3_4/io_cs_i cb_3_5/io_cs_i cb_3_6/io_cs_i cb_3_7/io_cs_i cb_3_8/io_cs_i
+ cb_3_9/io_cs_i cb_3_9/io_dat_i[0] cb_3_9/io_dat_i[10] cb_3_9/io_dat_i[11] cb_3_9/io_dat_i[12]
+ cb_3_9/io_dat_i[13] cb_3_9/io_dat_i[14] cb_3_9/io_dat_i[15] cb_3_9/io_dat_i[1] cb_3_9/io_dat_i[2]
+ cb_3_9/io_dat_i[3] cb_3_9/io_dat_i[4] cb_3_9/io_dat_i[5] cb_3_9/io_dat_i[6] cb_3_9/io_dat_i[7]
+ cb_3_9/io_dat_i[8] cb_3_9/io_dat_i[9] cb_3_0/io_dat_o[0] cb_3_0/io_dat_o[10] cb_3_0/io_dat_o[11]
+ cb_3_0/io_dat_o[12] cb_3_0/io_dat_o[13] cb_3_0/io_dat_o[14] cb_3_0/io_dat_o[15]
+ cb_3_0/io_dat_o[1] cb_3_0/io_dat_o[2] cb_3_0/io_dat_o[3] cb_3_0/io_dat_o[4] cb_3_0/io_dat_o[5]
+ cb_3_0/io_dat_o[6] cb_3_0/io_dat_o[7] cb_3_0/io_dat_o[8] cb_3_0/io_dat_o[9] cb_3_10/io_dat_o[0]
+ cb_3_10/io_dat_o[10] cb_3_10/io_dat_o[11] cb_3_10/io_dat_o[12] cb_3_10/io_dat_o[13]
+ cb_3_10/io_dat_o[14] cb_3_10/io_dat_o[15] cb_3_10/io_dat_o[1] cb_3_10/io_dat_o[2]
+ cb_3_10/io_dat_o[3] cb_3_10/io_dat_o[4] cb_3_10/io_dat_o[5] cb_3_10/io_dat_o[6]
+ cb_3_10/io_dat_o[7] cb_3_10/io_dat_o[8] cb_3_10/io_dat_o[9] cb_3_1/io_dat_o[0] cb_3_1/io_dat_o[10]
+ cb_3_1/io_dat_o[11] cb_3_1/io_dat_o[12] cb_3_1/io_dat_o[13] cb_3_1/io_dat_o[14]
+ cb_3_1/io_dat_o[15] cb_3_1/io_dat_o[1] cb_3_1/io_dat_o[2] cb_3_1/io_dat_o[3] cb_3_1/io_dat_o[4]
+ cb_3_1/io_dat_o[5] cb_3_1/io_dat_o[6] cb_3_1/io_dat_o[7] cb_3_1/io_dat_o[8] cb_3_1/io_dat_o[9]
+ cb_3_2/io_dat_o[0] cb_3_2/io_dat_o[10] cb_3_2/io_dat_o[11] cb_3_2/io_dat_o[12] cb_3_2/io_dat_o[13]
+ cb_3_2/io_dat_o[14] cb_3_2/io_dat_o[15] cb_3_2/io_dat_o[1] cb_3_2/io_dat_o[2] cb_3_2/io_dat_o[3]
+ cb_3_2/io_dat_o[4] cb_3_2/io_dat_o[5] cb_3_2/io_dat_o[6] cb_3_2/io_dat_o[7] cb_3_2/io_dat_o[8]
+ cb_3_2/io_dat_o[9] cb_3_3/io_dat_o[0] cb_3_3/io_dat_o[10] cb_3_3/io_dat_o[11] cb_3_3/io_dat_o[12]
+ cb_3_3/io_dat_o[13] cb_3_3/io_dat_o[14] cb_3_3/io_dat_o[15] cb_3_3/io_dat_o[1] cb_3_3/io_dat_o[2]
+ cb_3_3/io_dat_o[3] cb_3_3/io_dat_o[4] cb_3_3/io_dat_o[5] cb_3_3/io_dat_o[6] cb_3_3/io_dat_o[7]
+ cb_3_3/io_dat_o[8] cb_3_3/io_dat_o[9] cb_3_4/io_dat_o[0] cb_3_4/io_dat_o[10] cb_3_4/io_dat_o[11]
+ cb_3_4/io_dat_o[12] cb_3_4/io_dat_o[13] cb_3_4/io_dat_o[14] cb_3_4/io_dat_o[15]
+ cb_3_4/io_dat_o[1] cb_3_4/io_dat_o[2] cb_3_4/io_dat_o[3] cb_3_4/io_dat_o[4] cb_3_4/io_dat_o[5]
+ cb_3_4/io_dat_o[6] cb_3_4/io_dat_o[7] cb_3_4/io_dat_o[8] cb_3_4/io_dat_o[9] cb_3_5/io_dat_o[0]
+ cb_3_5/io_dat_o[10] cb_3_5/io_dat_o[11] cb_3_5/io_dat_o[12] cb_3_5/io_dat_o[13]
+ cb_3_5/io_dat_o[14] cb_3_5/io_dat_o[15] cb_3_5/io_dat_o[1] cb_3_5/io_dat_o[2] cb_3_5/io_dat_o[3]
+ cb_3_5/io_dat_o[4] cb_3_5/io_dat_o[5] cb_3_5/io_dat_o[6] cb_3_5/io_dat_o[7] cb_3_5/io_dat_o[8]
+ cb_3_5/io_dat_o[9] cb_3_6/io_dat_o[0] cb_3_6/io_dat_o[10] cb_3_6/io_dat_o[11] cb_3_6/io_dat_o[12]
+ cb_3_6/io_dat_o[13] cb_3_6/io_dat_o[14] cb_3_6/io_dat_o[15] cb_3_6/io_dat_o[1] cb_3_6/io_dat_o[2]
+ cb_3_6/io_dat_o[3] cb_3_6/io_dat_o[4] cb_3_6/io_dat_o[5] cb_3_6/io_dat_o[6] cb_3_6/io_dat_o[7]
+ cb_3_6/io_dat_o[8] cb_3_6/io_dat_o[9] cb_3_7/io_dat_o[0] cb_3_7/io_dat_o[10] cb_3_7/io_dat_o[11]
+ cb_3_7/io_dat_o[12] cb_3_7/io_dat_o[13] cb_3_7/io_dat_o[14] cb_3_7/io_dat_o[15]
+ cb_3_7/io_dat_o[1] cb_3_7/io_dat_o[2] cb_3_7/io_dat_o[3] cb_3_7/io_dat_o[4] cb_3_7/io_dat_o[5]
+ cb_3_7/io_dat_o[6] cb_3_7/io_dat_o[7] cb_3_7/io_dat_o[8] cb_3_7/io_dat_o[9] cb_3_8/io_dat_o[0]
+ cb_3_8/io_dat_o[10] cb_3_8/io_dat_o[11] cb_3_8/io_dat_o[12] cb_3_8/io_dat_o[13]
+ cb_3_8/io_dat_o[14] cb_3_8/io_dat_o[15] cb_3_8/io_dat_o[1] cb_3_8/io_dat_o[2] cb_3_8/io_dat_o[3]
+ cb_3_8/io_dat_o[4] cb_3_8/io_dat_o[5] cb_3_8/io_dat_o[6] cb_3_8/io_dat_o[7] cb_3_8/io_dat_o[8]
+ cb_3_8/io_dat_o[9] cb_3_9/io_dat_o[0] cb_3_9/io_dat_o[10] cb_3_9/io_dat_o[11] cb_3_9/io_dat_o[12]
+ cb_3_9/io_dat_o[13] cb_3_9/io_dat_o[14] cb_3_9/io_dat_o[15] cb_3_9/io_dat_o[1] cb_3_9/io_dat_o[2]
+ cb_3_9/io_dat_o[3] cb_3_9/io_dat_o[4] cb_3_9/io_dat_o[5] cb_3_9/io_dat_o[6] cb_3_9/io_dat_o[7]
+ cb_3_9/io_dat_o[8] cb_3_9/io_dat_o[9] cb_3_9/io_we_i ccon_3/io_cs_i ccon_7/io_dat_i[0]
+ ccon_7/io_dat_i[10] ccon_7/io_dat_i[11] ccon_7/io_dat_i[12] ccon_7/io_dat_i[13]
+ ccon_7/io_dat_i[14] ccon_7/io_dat_i[15] ccon_7/io_dat_i[16] ccon_7/io_dat_i[17]
+ ccon_7/io_dat_i[18] ccon_7/io_dat_i[19] ccon_7/io_dat_i[1] ccon_7/io_dat_i[20] ccon_7/io_dat_i[21]
+ ccon_7/io_dat_i[22] ccon_7/io_dat_i[23] ccon_7/io_dat_i[24] ccon_7/io_dat_i[25]
+ ccon_7/io_dat_i[26] ccon_7/io_dat_i[27] ccon_7/io_dat_i[28] ccon_7/io_dat_i[29]
+ ccon_7/io_dat_i[2] ccon_7/io_dat_i[30] ccon_7/io_dat_i[31] ccon_7/io_dat_i[3] ccon_7/io_dat_i[4]
+ ccon_7/io_dat_i[5] ccon_7/io_dat_i[6] ccon_7/io_dat_i[7] ccon_7/io_dat_i[8] ccon_7/io_dat_i[9]
+ ccon_3/io_dat_o[0] ccon_3/io_dat_o[10] ccon_3/io_dat_o[11] ccon_3/io_dat_o[12] ccon_3/io_dat_o[13]
+ ccon_3/io_dat_o[14] ccon_3/io_dat_o[15] ccon_3/io_dat_o[16] ccon_3/io_dat_o[17]
+ ccon_3/io_dat_o[18] ccon_3/io_dat_o[19] ccon_3/io_dat_o[1] ccon_3/io_dat_o[20] ccon_3/io_dat_o[21]
+ ccon_3/io_dat_o[22] ccon_3/io_dat_o[23] ccon_3/io_dat_o[24] ccon_3/io_dat_o[25]
+ ccon_3/io_dat_o[26] ccon_3/io_dat_o[27] ccon_3/io_dat_o[28] ccon_3/io_dat_o[29]
+ ccon_3/io_dat_o[2] ccon_3/io_dat_o[30] ccon_3/io_dat_o[31] ccon_3/io_dat_o[3] ccon_3/io_dat_o[4]
+ ccon_3/io_dat_o[5] ccon_3/io_dat_o[6] ccon_3/io_dat_o[7] ccon_3/io_dat_o[8] ccon_3/io_dat_o[9]
+ cb_3_0/io_wo[0] cb_3_0/io_wo[10] cb_3_0/io_wo[11] cb_3_0/io_wo[12] cb_3_0/io_wo[13]
+ cb_3_0/io_wo[14] cb_3_0/io_wo[15] cb_3_0/io_wo[16] cb_3_0/io_wo[17] cb_3_0/io_wo[18]
+ cb_3_0/io_wo[19] cb_3_0/io_wo[1] cb_3_0/io_wo[20] cb_3_0/io_wo[21] cb_3_0/io_wo[22]
+ cb_3_0/io_wo[23] cb_3_0/io_wo[24] cb_3_0/io_wo[25] cb_3_0/io_wo[26] cb_3_0/io_wo[27]
+ cb_3_0/io_wo[28] cb_3_0/io_wo[29] cb_3_0/io_wo[2] cb_3_0/io_wo[30] cb_3_0/io_wo[31]
+ cb_3_0/io_wo[32] cb_3_0/io_wo[33] cb_3_0/io_wo[34] cb_3_0/io_wo[35] cb_3_0/io_wo[36]
+ cb_3_0/io_wo[37] cb_3_0/io_wo[38] cb_3_0/io_wo[39] cb_3_0/io_wo[3] cb_3_0/io_wo[40]
+ cb_3_0/io_wo[41] cb_3_0/io_wo[42] cb_3_0/io_wo[43] cb_3_0/io_wo[44] cb_3_0/io_wo[45]
+ cb_3_0/io_wo[46] cb_3_0/io_wo[47] cb_3_0/io_wo[48] cb_3_0/io_wo[49] cb_3_0/io_wo[4]
+ cb_3_0/io_wo[50] cb_3_0/io_wo[51] cb_3_0/io_wo[52] cb_3_0/io_wo[53] cb_3_0/io_wo[54]
+ cb_3_0/io_wo[55] cb_3_0/io_wo[56] cb_3_0/io_wo[57] cb_3_0/io_wo[58] cb_3_0/io_wo[59]
+ cb_3_0/io_wo[5] cb_3_0/io_wo[60] cb_3_0/io_wo[61] cb_3_0/io_wo[62] cb_3_0/io_wo[63]
+ cb_3_0/io_wo[6] cb_3_0/io_wo[7] cb_3_0/io_wo[8] cb_3_0/io_wo[9] icon/dsi[0] icon/dsi[1]
+ icon/dsi[2] icon/dsi[3] icon/dsi[4] icon/dsi[5] icon/dsi[6] icon/dsi[7] ccon_3/io_dsi_o
+ ccon_3/io_irq cb_3_0/io_vi cb_3_10/io_vi cb_3_1/io_vi cb_3_2/io_vi cb_3_3/io_vi
+ cb_3_4/io_vi cb_3_5/io_vi cb_3_6/io_vi cb_3_7/io_vi cb_3_8/io_vi cb_3_9/io_vi ccon_7/io_we_i
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_con
Xcb_3_10 cb_3_9/io_adr_i[0] cb_3_9/io_adr_i[1] cb_3_10/io_cs_i cb_3_9/io_dat_i[0]
+ cb_3_9/io_dat_i[10] cb_3_9/io_dat_i[11] cb_3_9/io_dat_i[12] cb_3_9/io_dat_i[13]
+ cb_3_9/io_dat_i[14] cb_3_9/io_dat_i[15] cb_3_9/io_dat_i[1] cb_3_9/io_dat_i[2] cb_3_9/io_dat_i[3]
+ cb_3_9/io_dat_i[4] cb_3_9/io_dat_i[5] cb_3_9/io_dat_i[6] cb_3_9/io_dat_i[7] cb_3_9/io_dat_i[8]
+ cb_3_9/io_dat_i[9] cb_3_10/io_dat_o[0] cb_3_10/io_dat_o[10] cb_3_10/io_dat_o[11]
+ cb_3_10/io_dat_o[12] cb_3_10/io_dat_o[13] cb_3_10/io_dat_o[14] cb_3_10/io_dat_o[15]
+ cb_3_10/io_dat_o[1] cb_3_10/io_dat_o[2] cb_3_10/io_dat_o[3] cb_3_10/io_dat_o[4]
+ cb_3_10/io_dat_o[5] cb_3_10/io_dat_o[6] cb_3_10/io_dat_o[7] cb_3_10/io_dat_o[8]
+ cb_3_10/io_dat_o[9] cb_3_10/io_eo[0] cb_3_10/io_eo[10] cb_3_10/io_eo[11] cb_3_10/io_eo[12]
+ cb_3_10/io_eo[13] cb_3_10/io_eo[14] cb_3_10/io_eo[15] cb_3_10/io_eo[16] cb_3_10/io_eo[17]
+ cb_3_10/io_eo[18] cb_3_10/io_eo[19] cb_3_10/io_eo[1] cb_3_10/io_eo[20] cb_3_10/io_eo[21]
+ cb_3_10/io_eo[22] cb_3_10/io_eo[23] cb_3_10/io_eo[24] cb_3_10/io_eo[25] cb_3_10/io_eo[26]
+ cb_3_10/io_eo[27] cb_3_10/io_eo[28] cb_3_10/io_eo[29] cb_3_10/io_eo[2] cb_3_10/io_eo[30]
+ cb_3_10/io_eo[31] cb_3_10/io_eo[32] cb_3_10/io_eo[33] cb_3_10/io_eo[34] cb_3_10/io_eo[35]
+ cb_3_10/io_eo[36] cb_3_10/io_eo[37] cb_3_10/io_eo[38] cb_3_10/io_eo[39] cb_3_10/io_eo[3]
+ cb_3_10/io_eo[40] cb_3_10/io_eo[41] cb_3_10/io_eo[42] cb_3_10/io_eo[43] cb_3_10/io_eo[44]
+ cb_3_10/io_eo[45] cb_3_10/io_eo[46] cb_3_10/io_eo[47] cb_3_10/io_eo[48] cb_3_10/io_eo[49]
+ cb_3_10/io_eo[4] cb_3_10/io_eo[50] cb_3_10/io_eo[51] cb_3_10/io_eo[52] cb_3_10/io_eo[53]
+ cb_3_10/io_eo[54] cb_3_10/io_eo[55] cb_3_10/io_eo[56] cb_3_10/io_eo[57] cb_3_10/io_eo[58]
+ cb_3_10/io_eo[59] cb_3_10/io_eo[5] cb_3_10/io_eo[60] cb_3_10/io_eo[61] cb_3_10/io_eo[62]
+ cb_3_10/io_eo[63] cb_3_10/io_eo[6] cb_3_10/io_eo[7] cb_3_10/io_eo[8] cb_3_10/io_eo[9]
+ cb_3_9/io_o_0_co cb_3_9/io_o_0_out[0] cb_3_9/io_o_0_out[1] cb_3_9/io_o_0_out[2]
+ cb_3_9/io_o_0_out[3] cb_3_9/io_o_0_out[4] cb_3_9/io_o_0_out[5] cb_3_9/io_o_0_out[6]
+ cb_3_9/io_o_0_out[7] cb_3_9/io_o_1_co cb_3_9/io_o_1_out[0] cb_3_9/io_o_1_out[1]
+ cb_3_9/io_o_1_out[2] cb_3_9/io_o_1_out[3] cb_3_9/io_o_1_out[4] cb_3_9/io_o_1_out[5]
+ cb_3_9/io_o_1_out[6] cb_3_9/io_o_1_out[7] cb_3_9/io_o_2_co cb_3_9/io_o_2_out[0]
+ cb_3_9/io_o_2_out[1] cb_3_9/io_o_2_out[2] cb_3_9/io_o_2_out[3] cb_3_9/io_o_2_out[4]
+ cb_3_9/io_o_2_out[5] cb_3_9/io_o_2_out[6] cb_3_9/io_o_2_out[7] cb_3_9/io_o_3_co
+ cb_3_9/io_o_3_out[0] cb_3_9/io_o_3_out[1] cb_3_9/io_o_3_out[2] cb_3_9/io_o_3_out[3]
+ cb_3_9/io_o_3_out[4] cb_3_9/io_o_3_out[5] cb_3_9/io_o_3_out[6] cb_3_9/io_o_3_out[7]
+ cb_3_9/io_o_4_co cb_3_9/io_o_4_out[0] cb_3_9/io_o_4_out[1] cb_3_9/io_o_4_out[2]
+ cb_3_9/io_o_4_out[3] cb_3_9/io_o_4_out[4] cb_3_9/io_o_4_out[5] cb_3_9/io_o_4_out[6]
+ cb_3_9/io_o_4_out[7] cb_3_9/io_o_5_co cb_3_9/io_o_5_out[0] cb_3_9/io_o_5_out[1]
+ cb_3_9/io_o_5_out[2] cb_3_9/io_o_5_out[3] cb_3_9/io_o_5_out[4] cb_3_9/io_o_5_out[5]
+ cb_3_9/io_o_5_out[6] cb_3_9/io_o_5_out[7] cb_3_9/io_o_6_co cb_3_9/io_o_6_out[0]
+ cb_3_9/io_o_6_out[1] cb_3_9/io_o_6_out[2] cb_3_9/io_o_6_out[3] cb_3_9/io_o_6_out[4]
+ cb_3_9/io_o_6_out[5] cb_3_9/io_o_6_out[6] cb_3_9/io_o_6_out[7] cb_3_9/io_o_7_co
+ cb_3_9/io_o_7_out[0] cb_3_9/io_o_7_out[1] cb_3_9/io_o_7_out[2] cb_3_9/io_o_7_out[3]
+ cb_3_9/io_o_7_out[4] cb_3_9/io_o_7_out[5] cb_3_9/io_o_7_out[6] cb_3_9/io_o_7_out[7]
+ cb_3_10/io_o_0_co cb_3_10/io_eo[0] cb_3_10/io_eo[1] cb_3_10/io_eo[2] cb_3_10/io_eo[3]
+ cb_3_10/io_eo[4] cb_3_10/io_eo[5] cb_3_10/io_eo[6] cb_3_10/io_eo[7] cb_3_10/io_o_1_co
+ cb_3_10/io_eo[8] cb_3_10/io_eo[9] cb_3_10/io_eo[10] cb_3_10/io_eo[11] cb_3_10/io_eo[12]
+ cb_3_10/io_eo[13] cb_3_10/io_eo[14] cb_3_10/io_eo[15] cb_3_10/io_o_2_co cb_3_10/io_eo[16]
+ cb_3_10/io_eo[17] cb_3_10/io_eo[18] cb_3_10/io_eo[19] cb_3_10/io_eo[20] cb_3_10/io_eo[21]
+ cb_3_10/io_eo[22] cb_3_10/io_eo[23] cb_3_10/io_o_3_co cb_3_10/io_eo[24] cb_3_10/io_eo[25]
+ cb_3_10/io_eo[26] cb_3_10/io_eo[27] cb_3_10/io_eo[28] cb_3_10/io_eo[29] cb_3_10/io_eo[30]
+ cb_3_10/io_eo[31] cb_3_10/io_o_4_co cb_3_10/io_eo[32] cb_3_10/io_eo[33] cb_3_10/io_eo[34]
+ cb_3_10/io_eo[35] cb_3_10/io_eo[36] cb_3_10/io_eo[37] cb_3_10/io_eo[38] cb_3_10/io_eo[39]
+ cb_3_10/io_o_5_co cb_3_10/io_eo[40] cb_3_10/io_eo[41] cb_3_10/io_eo[42] cb_3_10/io_eo[43]
+ cb_3_10/io_eo[44] cb_3_10/io_eo[45] cb_3_10/io_eo[46] cb_3_10/io_eo[47] cb_3_10/io_o_6_co
+ cb_3_10/io_eo[48] cb_3_10/io_eo[49] cb_3_10/io_eo[50] cb_3_10/io_eo[51] cb_3_10/io_eo[52]
+ cb_3_10/io_eo[53] cb_3_10/io_eo[54] cb_3_10/io_eo[55] cb_3_10/io_o_7_co cb_3_10/io_eo[56]
+ cb_3_10/io_eo[57] cb_3_10/io_eo[58] cb_3_10/io_eo[59] cb_3_10/io_eo[60] cb_3_10/io_eo[61]
+ cb_3_10/io_eo[62] cb_3_10/io_eo[63] cb_3_9/io_vco cb_3_10/io_vco cb_3_10/io_vi cb_3_9/io_we_i
+ cb_3_9/io_eo[0] cb_3_9/io_eo[10] cb_3_9/io_eo[11] cb_3_9/io_eo[12] cb_3_9/io_eo[13]
+ cb_3_9/io_eo[14] cb_3_9/io_eo[15] cb_3_9/io_eo[16] cb_3_9/io_eo[17] cb_3_9/io_eo[18]
+ cb_3_9/io_eo[19] cb_3_9/io_eo[1] cb_3_9/io_eo[20] cb_3_9/io_eo[21] cb_3_9/io_eo[22]
+ cb_3_9/io_eo[23] cb_3_9/io_eo[24] cb_3_9/io_eo[25] cb_3_9/io_eo[26] cb_3_9/io_eo[27]
+ cb_3_9/io_eo[28] cb_3_9/io_eo[29] cb_3_9/io_eo[2] cb_3_9/io_eo[30] cb_3_9/io_eo[31]
+ cb_3_9/io_eo[32] cb_3_9/io_eo[33] cb_3_9/io_eo[34] cb_3_9/io_eo[35] cb_3_9/io_eo[36]
+ cb_3_9/io_eo[37] cb_3_9/io_eo[38] cb_3_9/io_eo[39] cb_3_9/io_eo[3] cb_3_9/io_eo[40]
+ cb_3_9/io_eo[41] cb_3_9/io_eo[42] cb_3_9/io_eo[43] cb_3_9/io_eo[44] cb_3_9/io_eo[45]
+ cb_3_9/io_eo[46] cb_3_9/io_eo[47] cb_3_9/io_eo[48] cb_3_9/io_eo[49] cb_3_9/io_eo[4]
+ cb_3_9/io_eo[50] cb_3_9/io_eo[51] cb_3_9/io_eo[52] cb_3_9/io_eo[53] cb_3_9/io_eo[54]
+ cb_3_9/io_eo[55] cb_3_9/io_eo[56] cb_3_9/io_eo[57] cb_3_9/io_eo[58] cb_3_9/io_eo[59]
+ cb_3_9/io_eo[5] cb_3_9/io_eo[60] cb_3_9/io_eo[61] cb_3_9/io_eo[62] cb_3_9/io_eo[63]
+ cb_3_9/io_eo[6] cb_3_9/io_eo[7] cb_3_9/io_eo[8] cb_3_9/io_eo[9] mcons_3/clock mcons_3/reset
+ vccd1 vssd1 cic_block
Xcb_5_7 cb_5_9/io_adr_i[0] cb_5_9/io_adr_i[1] cb_5_7/io_cs_i cb_5_9/io_dat_i[0] cb_5_9/io_dat_i[10]
+ cb_5_9/io_dat_i[11] cb_5_9/io_dat_i[12] cb_5_9/io_dat_i[13] cb_5_9/io_dat_i[14]
+ cb_5_9/io_dat_i[15] cb_5_9/io_dat_i[1] cb_5_9/io_dat_i[2] cb_5_9/io_dat_i[3] cb_5_9/io_dat_i[4]
+ cb_5_9/io_dat_i[5] cb_5_9/io_dat_i[6] cb_5_9/io_dat_i[7] cb_5_9/io_dat_i[8] cb_5_9/io_dat_i[9]
+ cb_5_7/io_dat_o[0] cb_5_7/io_dat_o[10] cb_5_7/io_dat_o[11] cb_5_7/io_dat_o[12] cb_5_7/io_dat_o[13]
+ cb_5_7/io_dat_o[14] cb_5_7/io_dat_o[15] cb_5_7/io_dat_o[1] cb_5_7/io_dat_o[2] cb_5_7/io_dat_o[3]
+ cb_5_7/io_dat_o[4] cb_5_7/io_dat_o[5] cb_5_7/io_dat_o[6] cb_5_7/io_dat_o[7] cb_5_7/io_dat_o[8]
+ cb_5_7/io_dat_o[9] cb_5_8/io_wo[0] cb_5_8/io_wo[10] cb_5_8/io_wo[11] cb_5_8/io_wo[12]
+ cb_5_8/io_wo[13] cb_5_8/io_wo[14] cb_5_8/io_wo[15] cb_5_8/io_wo[16] cb_5_8/io_wo[17]
+ cb_5_8/io_wo[18] cb_5_8/io_wo[19] cb_5_8/io_wo[1] cb_5_8/io_wo[20] cb_5_8/io_wo[21]
+ cb_5_8/io_wo[22] cb_5_8/io_wo[23] cb_5_8/io_wo[24] cb_5_8/io_wo[25] cb_5_8/io_wo[26]
+ cb_5_8/io_wo[27] cb_5_8/io_wo[28] cb_5_8/io_wo[29] cb_5_8/io_wo[2] cb_5_8/io_wo[30]
+ cb_5_8/io_wo[31] cb_5_8/io_wo[32] cb_5_8/io_wo[33] cb_5_8/io_wo[34] cb_5_8/io_wo[35]
+ cb_5_8/io_wo[36] cb_5_8/io_wo[37] cb_5_8/io_wo[38] cb_5_8/io_wo[39] cb_5_8/io_wo[3]
+ cb_5_8/io_wo[40] cb_5_8/io_wo[41] cb_5_8/io_wo[42] cb_5_8/io_wo[43] cb_5_8/io_wo[44]
+ cb_5_8/io_wo[45] cb_5_8/io_wo[46] cb_5_8/io_wo[47] cb_5_8/io_wo[48] cb_5_8/io_wo[49]
+ cb_5_8/io_wo[4] cb_5_8/io_wo[50] cb_5_8/io_wo[51] cb_5_8/io_wo[52] cb_5_8/io_wo[53]
+ cb_5_8/io_wo[54] cb_5_8/io_wo[55] cb_5_8/io_wo[56] cb_5_8/io_wo[57] cb_5_8/io_wo[58]
+ cb_5_8/io_wo[59] cb_5_8/io_wo[5] cb_5_8/io_wo[60] cb_5_8/io_wo[61] cb_5_8/io_wo[62]
+ cb_5_8/io_wo[63] cb_5_8/io_wo[6] cb_5_8/io_wo[7] cb_5_8/io_wo[8] cb_5_8/io_wo[9]
+ cb_5_7/io_i_0_ci cb_5_7/io_i_0_in1[0] cb_5_7/io_i_0_in1[1] cb_5_7/io_i_0_in1[2]
+ cb_5_7/io_i_0_in1[3] cb_5_7/io_i_0_in1[4] cb_5_7/io_i_0_in1[5] cb_5_7/io_i_0_in1[6]
+ cb_5_7/io_i_0_in1[7] cb_5_7/io_i_1_ci cb_5_7/io_i_1_in1[0] cb_5_7/io_i_1_in1[1]
+ cb_5_7/io_i_1_in1[2] cb_5_7/io_i_1_in1[3] cb_5_7/io_i_1_in1[4] cb_5_7/io_i_1_in1[5]
+ cb_5_7/io_i_1_in1[6] cb_5_7/io_i_1_in1[7] cb_5_7/io_i_2_ci cb_5_7/io_i_2_in1[0]
+ cb_5_7/io_i_2_in1[1] cb_5_7/io_i_2_in1[2] cb_5_7/io_i_2_in1[3] cb_5_7/io_i_2_in1[4]
+ cb_5_7/io_i_2_in1[5] cb_5_7/io_i_2_in1[6] cb_5_7/io_i_2_in1[7] cb_5_7/io_i_3_ci
+ cb_5_7/io_i_3_in1[0] cb_5_7/io_i_3_in1[1] cb_5_7/io_i_3_in1[2] cb_5_7/io_i_3_in1[3]
+ cb_5_7/io_i_3_in1[4] cb_5_7/io_i_3_in1[5] cb_5_7/io_i_3_in1[6] cb_5_7/io_i_3_in1[7]
+ cb_5_7/io_i_4_ci cb_5_7/io_i_4_in1[0] cb_5_7/io_i_4_in1[1] cb_5_7/io_i_4_in1[2]
+ cb_5_7/io_i_4_in1[3] cb_5_7/io_i_4_in1[4] cb_5_7/io_i_4_in1[5] cb_5_7/io_i_4_in1[6]
+ cb_5_7/io_i_4_in1[7] cb_5_7/io_i_5_ci cb_5_7/io_i_5_in1[0] cb_5_7/io_i_5_in1[1]
+ cb_5_7/io_i_5_in1[2] cb_5_7/io_i_5_in1[3] cb_5_7/io_i_5_in1[4] cb_5_7/io_i_5_in1[5]
+ cb_5_7/io_i_5_in1[6] cb_5_7/io_i_5_in1[7] cb_5_7/io_i_6_ci cb_5_7/io_i_6_in1[0]
+ cb_5_7/io_i_6_in1[1] cb_5_7/io_i_6_in1[2] cb_5_7/io_i_6_in1[3] cb_5_7/io_i_6_in1[4]
+ cb_5_7/io_i_6_in1[5] cb_5_7/io_i_6_in1[6] cb_5_7/io_i_6_in1[7] cb_5_7/io_i_7_ci
+ cb_5_7/io_i_7_in1[0] cb_5_7/io_i_7_in1[1] cb_5_7/io_i_7_in1[2] cb_5_7/io_i_7_in1[3]
+ cb_5_7/io_i_7_in1[4] cb_5_7/io_i_7_in1[5] cb_5_7/io_i_7_in1[6] cb_5_7/io_i_7_in1[7]
+ cb_5_8/io_i_0_ci cb_5_8/io_i_0_in1[0] cb_5_8/io_i_0_in1[1] cb_5_8/io_i_0_in1[2]
+ cb_5_8/io_i_0_in1[3] cb_5_8/io_i_0_in1[4] cb_5_8/io_i_0_in1[5] cb_5_8/io_i_0_in1[6]
+ cb_5_8/io_i_0_in1[7] cb_5_8/io_i_1_ci cb_5_8/io_i_1_in1[0] cb_5_8/io_i_1_in1[1]
+ cb_5_8/io_i_1_in1[2] cb_5_8/io_i_1_in1[3] cb_5_8/io_i_1_in1[4] cb_5_8/io_i_1_in1[5]
+ cb_5_8/io_i_1_in1[6] cb_5_8/io_i_1_in1[7] cb_5_8/io_i_2_ci cb_5_8/io_i_2_in1[0]
+ cb_5_8/io_i_2_in1[1] cb_5_8/io_i_2_in1[2] cb_5_8/io_i_2_in1[3] cb_5_8/io_i_2_in1[4]
+ cb_5_8/io_i_2_in1[5] cb_5_8/io_i_2_in1[6] cb_5_8/io_i_2_in1[7] cb_5_8/io_i_3_ci
+ cb_5_8/io_i_3_in1[0] cb_5_8/io_i_3_in1[1] cb_5_8/io_i_3_in1[2] cb_5_8/io_i_3_in1[3]
+ cb_5_8/io_i_3_in1[4] cb_5_8/io_i_3_in1[5] cb_5_8/io_i_3_in1[6] cb_5_8/io_i_3_in1[7]
+ cb_5_8/io_i_4_ci cb_5_8/io_i_4_in1[0] cb_5_8/io_i_4_in1[1] cb_5_8/io_i_4_in1[2]
+ cb_5_8/io_i_4_in1[3] cb_5_8/io_i_4_in1[4] cb_5_8/io_i_4_in1[5] cb_5_8/io_i_4_in1[6]
+ cb_5_8/io_i_4_in1[7] cb_5_8/io_i_5_ci cb_5_8/io_i_5_in1[0] cb_5_8/io_i_5_in1[1]
+ cb_5_8/io_i_5_in1[2] cb_5_8/io_i_5_in1[3] cb_5_8/io_i_5_in1[4] cb_5_8/io_i_5_in1[5]
+ cb_5_8/io_i_5_in1[6] cb_5_8/io_i_5_in1[7] cb_5_8/io_i_6_ci cb_5_8/io_i_6_in1[0]
+ cb_5_8/io_i_6_in1[1] cb_5_8/io_i_6_in1[2] cb_5_8/io_i_6_in1[3] cb_5_8/io_i_6_in1[4]
+ cb_5_8/io_i_6_in1[5] cb_5_8/io_i_6_in1[6] cb_5_8/io_i_6_in1[7] cb_5_8/io_i_7_ci
+ cb_5_8/io_i_7_in1[0] cb_5_8/io_i_7_in1[1] cb_5_8/io_i_7_in1[2] cb_5_8/io_i_7_in1[3]
+ cb_5_8/io_i_7_in1[4] cb_5_8/io_i_7_in1[5] cb_5_8/io_i_7_in1[6] cb_5_8/io_i_7_in1[7]
+ cb_5_7/io_vci cb_5_8/io_vci cb_5_7/io_vi cb_5_9/io_we_i cb_5_7/io_wo[0] cb_5_7/io_wo[10]
+ cb_5_7/io_wo[11] cb_5_7/io_wo[12] cb_5_7/io_wo[13] cb_5_7/io_wo[14] cb_5_7/io_wo[15]
+ cb_5_7/io_wo[16] cb_5_7/io_wo[17] cb_5_7/io_wo[18] cb_5_7/io_wo[19] cb_5_7/io_wo[1]
+ cb_5_7/io_wo[20] cb_5_7/io_wo[21] cb_5_7/io_wo[22] cb_5_7/io_wo[23] cb_5_7/io_wo[24]
+ cb_5_7/io_wo[25] cb_5_7/io_wo[26] cb_5_7/io_wo[27] cb_5_7/io_wo[28] cb_5_7/io_wo[29]
+ cb_5_7/io_wo[2] cb_5_7/io_wo[30] cb_5_7/io_wo[31] cb_5_7/io_wo[32] cb_5_7/io_wo[33]
+ cb_5_7/io_wo[34] cb_5_7/io_wo[35] cb_5_7/io_wo[36] cb_5_7/io_wo[37] cb_5_7/io_wo[38]
+ cb_5_7/io_wo[39] cb_5_7/io_wo[3] cb_5_7/io_wo[40] cb_5_7/io_wo[41] cb_5_7/io_wo[42]
+ cb_5_7/io_wo[43] cb_5_7/io_wo[44] cb_5_7/io_wo[45] cb_5_7/io_wo[46] cb_5_7/io_wo[47]
+ cb_5_7/io_wo[48] cb_5_7/io_wo[49] cb_5_7/io_wo[4] cb_5_7/io_wo[50] cb_5_7/io_wo[51]
+ cb_5_7/io_wo[52] cb_5_7/io_wo[53] cb_5_7/io_wo[54] cb_5_7/io_wo[55] cb_5_7/io_wo[56]
+ cb_5_7/io_wo[57] cb_5_7/io_wo[58] cb_5_7/io_wo[59] cb_5_7/io_wo[5] cb_5_7/io_wo[60]
+ cb_5_7/io_wo[61] cb_5_7/io_wo[62] cb_5_7/io_wo[63] cb_5_7/io_wo[6] cb_5_7/io_wo[7]
+ cb_5_7/io_wo[8] cb_5_7/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_6_10 cb_6_9/io_adr_i[0] cb_6_9/io_adr_i[1] cb_6_10/io_cs_i cb_6_9/io_dat_i[0]
+ cb_6_9/io_dat_i[10] cb_6_9/io_dat_i[11] cb_6_9/io_dat_i[12] cb_6_9/io_dat_i[13]
+ cb_6_9/io_dat_i[14] cb_6_9/io_dat_i[15] cb_6_9/io_dat_i[1] cb_6_9/io_dat_i[2] cb_6_9/io_dat_i[3]
+ cb_6_9/io_dat_i[4] cb_6_9/io_dat_i[5] cb_6_9/io_dat_i[6] cb_6_9/io_dat_i[7] cb_6_9/io_dat_i[8]
+ cb_6_9/io_dat_i[9] cb_6_10/io_dat_o[0] cb_6_10/io_dat_o[10] cb_6_10/io_dat_o[11]
+ cb_6_10/io_dat_o[12] cb_6_10/io_dat_o[13] cb_6_10/io_dat_o[14] cb_6_10/io_dat_o[15]
+ cb_6_10/io_dat_o[1] cb_6_10/io_dat_o[2] cb_6_10/io_dat_o[3] cb_6_10/io_dat_o[4]
+ cb_6_10/io_dat_o[5] cb_6_10/io_dat_o[6] cb_6_10/io_dat_o[7] cb_6_10/io_dat_o[8]
+ cb_6_10/io_dat_o[9] cb_6_10/io_eo[0] cb_6_10/io_eo[10] cb_6_10/io_eo[11] cb_6_10/io_eo[12]
+ cb_6_10/io_eo[13] cb_6_10/io_eo[14] cb_6_10/io_eo[15] cb_6_10/io_eo[16] cb_6_10/io_eo[17]
+ cb_6_10/io_eo[18] cb_6_10/io_eo[19] cb_6_10/io_eo[1] cb_6_10/io_eo[20] cb_6_10/io_eo[21]
+ cb_6_10/io_eo[22] cb_6_10/io_eo[23] cb_6_10/io_eo[24] cb_6_10/io_eo[25] cb_6_10/io_eo[26]
+ cb_6_10/io_eo[27] cb_6_10/io_eo[28] cb_6_10/io_eo[29] cb_6_10/io_eo[2] cb_6_10/io_eo[30]
+ cb_6_10/io_eo[31] cb_6_10/io_eo[32] cb_6_10/io_eo[33] cb_6_10/io_eo[34] cb_6_10/io_eo[35]
+ cb_6_10/io_eo[36] cb_6_10/io_eo[37] cb_6_10/io_eo[38] cb_6_10/io_eo[39] cb_6_10/io_eo[3]
+ cb_6_10/io_eo[40] cb_6_10/io_eo[41] cb_6_10/io_eo[42] cb_6_10/io_eo[43] cb_6_10/io_eo[44]
+ cb_6_10/io_eo[45] cb_6_10/io_eo[46] cb_6_10/io_eo[47] cb_6_10/io_eo[48] cb_6_10/io_eo[49]
+ cb_6_10/io_eo[4] cb_6_10/io_eo[50] cb_6_10/io_eo[51] cb_6_10/io_eo[52] cb_6_10/io_eo[53]
+ cb_6_10/io_eo[54] cb_6_10/io_eo[55] cb_6_10/io_eo[56] cb_6_10/io_eo[57] cb_6_10/io_eo[58]
+ cb_6_10/io_eo[59] cb_6_10/io_eo[5] cb_6_10/io_eo[60] cb_6_10/io_eo[61] cb_6_10/io_eo[62]
+ cb_6_10/io_eo[63] cb_6_10/io_eo[6] cb_6_10/io_eo[7] cb_6_10/io_eo[8] cb_6_10/io_eo[9]
+ cb_6_9/io_o_0_co cb_6_9/io_o_0_out[0] cb_6_9/io_o_0_out[1] cb_6_9/io_o_0_out[2]
+ cb_6_9/io_o_0_out[3] cb_6_9/io_o_0_out[4] cb_6_9/io_o_0_out[5] cb_6_9/io_o_0_out[6]
+ cb_6_9/io_o_0_out[7] cb_6_9/io_o_1_co cb_6_9/io_o_1_out[0] cb_6_9/io_o_1_out[1]
+ cb_6_9/io_o_1_out[2] cb_6_9/io_o_1_out[3] cb_6_9/io_o_1_out[4] cb_6_9/io_o_1_out[5]
+ cb_6_9/io_o_1_out[6] cb_6_9/io_o_1_out[7] cb_6_9/io_o_2_co cb_6_9/io_o_2_out[0]
+ cb_6_9/io_o_2_out[1] cb_6_9/io_o_2_out[2] cb_6_9/io_o_2_out[3] cb_6_9/io_o_2_out[4]
+ cb_6_9/io_o_2_out[5] cb_6_9/io_o_2_out[6] cb_6_9/io_o_2_out[7] cb_6_9/io_o_3_co
+ cb_6_9/io_o_3_out[0] cb_6_9/io_o_3_out[1] cb_6_9/io_o_3_out[2] cb_6_9/io_o_3_out[3]
+ cb_6_9/io_o_3_out[4] cb_6_9/io_o_3_out[5] cb_6_9/io_o_3_out[6] cb_6_9/io_o_3_out[7]
+ cb_6_9/io_o_4_co cb_6_9/io_o_4_out[0] cb_6_9/io_o_4_out[1] cb_6_9/io_o_4_out[2]
+ cb_6_9/io_o_4_out[3] cb_6_9/io_o_4_out[4] cb_6_9/io_o_4_out[5] cb_6_9/io_o_4_out[6]
+ cb_6_9/io_o_4_out[7] cb_6_9/io_o_5_co cb_6_9/io_o_5_out[0] cb_6_9/io_o_5_out[1]
+ cb_6_9/io_o_5_out[2] cb_6_9/io_o_5_out[3] cb_6_9/io_o_5_out[4] cb_6_9/io_o_5_out[5]
+ cb_6_9/io_o_5_out[6] cb_6_9/io_o_5_out[7] cb_6_9/io_o_6_co cb_6_9/io_o_6_out[0]
+ cb_6_9/io_o_6_out[1] cb_6_9/io_o_6_out[2] cb_6_9/io_o_6_out[3] cb_6_9/io_o_6_out[4]
+ cb_6_9/io_o_6_out[5] cb_6_9/io_o_6_out[6] cb_6_9/io_o_6_out[7] cb_6_9/io_o_7_co
+ cb_6_9/io_o_7_out[0] cb_6_9/io_o_7_out[1] cb_6_9/io_o_7_out[2] cb_6_9/io_o_7_out[3]
+ cb_6_9/io_o_7_out[4] cb_6_9/io_o_7_out[5] cb_6_9/io_o_7_out[6] cb_6_9/io_o_7_out[7]
+ cb_6_10/io_o_0_co cb_6_10/io_eo[0] cb_6_10/io_eo[1] cb_6_10/io_eo[2] cb_6_10/io_eo[3]
+ cb_6_10/io_eo[4] cb_6_10/io_eo[5] cb_6_10/io_eo[6] cb_6_10/io_eo[7] cb_6_10/io_o_1_co
+ cb_6_10/io_eo[8] cb_6_10/io_eo[9] cb_6_10/io_eo[10] cb_6_10/io_eo[11] cb_6_10/io_eo[12]
+ cb_6_10/io_eo[13] cb_6_10/io_eo[14] cb_6_10/io_eo[15] cb_6_10/io_o_2_co cb_6_10/io_eo[16]
+ cb_6_10/io_eo[17] cb_6_10/io_eo[18] cb_6_10/io_eo[19] cb_6_10/io_eo[20] cb_6_10/io_eo[21]
+ cb_6_10/io_eo[22] cb_6_10/io_eo[23] cb_6_10/io_o_3_co cb_6_10/io_eo[24] cb_6_10/io_eo[25]
+ cb_6_10/io_eo[26] cb_6_10/io_eo[27] cb_6_10/io_eo[28] cb_6_10/io_eo[29] cb_6_10/io_eo[30]
+ cb_6_10/io_eo[31] cb_6_10/io_o_4_co cb_6_10/io_eo[32] cb_6_10/io_eo[33] cb_6_10/io_eo[34]
+ cb_6_10/io_eo[35] cb_6_10/io_eo[36] cb_6_10/io_eo[37] cb_6_10/io_eo[38] cb_6_10/io_eo[39]
+ cb_6_10/io_o_5_co cb_6_10/io_eo[40] cb_6_10/io_eo[41] cb_6_10/io_eo[42] cb_6_10/io_eo[43]
+ cb_6_10/io_eo[44] cb_6_10/io_eo[45] cb_6_10/io_eo[46] cb_6_10/io_eo[47] cb_6_10/io_o_6_co
+ cb_6_10/io_eo[48] cb_6_10/io_eo[49] cb_6_10/io_eo[50] cb_6_10/io_eo[51] cb_6_10/io_eo[52]
+ cb_6_10/io_eo[53] cb_6_10/io_eo[54] cb_6_10/io_eo[55] cb_6_10/io_o_7_co cb_6_10/io_eo[56]
+ cb_6_10/io_eo[57] cb_6_10/io_eo[58] cb_6_10/io_eo[59] cb_6_10/io_eo[60] cb_6_10/io_eo[61]
+ cb_6_10/io_eo[62] cb_6_10/io_eo[63] cb_6_9/io_vco cb_6_10/io_vco cb_6_10/io_vi cb_6_9/io_we_i
+ cb_6_9/io_eo[0] cb_6_9/io_eo[10] cb_6_9/io_eo[11] cb_6_9/io_eo[12] cb_6_9/io_eo[13]
+ cb_6_9/io_eo[14] cb_6_9/io_eo[15] cb_6_9/io_eo[16] cb_6_9/io_eo[17] cb_6_9/io_eo[18]
+ cb_6_9/io_eo[19] cb_6_9/io_eo[1] cb_6_9/io_eo[20] cb_6_9/io_eo[21] cb_6_9/io_eo[22]
+ cb_6_9/io_eo[23] cb_6_9/io_eo[24] cb_6_9/io_eo[25] cb_6_9/io_eo[26] cb_6_9/io_eo[27]
+ cb_6_9/io_eo[28] cb_6_9/io_eo[29] cb_6_9/io_eo[2] cb_6_9/io_eo[30] cb_6_9/io_eo[31]
+ cb_6_9/io_eo[32] cb_6_9/io_eo[33] cb_6_9/io_eo[34] cb_6_9/io_eo[35] cb_6_9/io_eo[36]
+ cb_6_9/io_eo[37] cb_6_9/io_eo[38] cb_6_9/io_eo[39] cb_6_9/io_eo[3] cb_6_9/io_eo[40]
+ cb_6_9/io_eo[41] cb_6_9/io_eo[42] cb_6_9/io_eo[43] cb_6_9/io_eo[44] cb_6_9/io_eo[45]
+ cb_6_9/io_eo[46] cb_6_9/io_eo[47] cb_6_9/io_eo[48] cb_6_9/io_eo[49] cb_6_9/io_eo[4]
+ cb_6_9/io_eo[50] cb_6_9/io_eo[51] cb_6_9/io_eo[52] cb_6_9/io_eo[53] cb_6_9/io_eo[54]
+ cb_6_9/io_eo[55] cb_6_9/io_eo[56] cb_6_9/io_eo[57] cb_6_9/io_eo[58] cb_6_9/io_eo[59]
+ cb_6_9/io_eo[5] cb_6_9/io_eo[60] cb_6_9/io_eo[61] cb_6_9/io_eo[62] cb_6_9/io_eo[63]
+ cb_6_9/io_eo[6] cb_6_9/io_eo[7] cb_6_9/io_eo[8] cb_6_9/io_eo[9] mcons_3/clock mcons_3/reset
+ vccd1 vssd1 cic_block
Xcb_3_4 cb_3_9/io_adr_i[0] cb_3_9/io_adr_i[1] cb_3_4/io_cs_i cb_3_9/io_dat_i[0] cb_3_9/io_dat_i[10]
+ cb_3_9/io_dat_i[11] cb_3_9/io_dat_i[12] cb_3_9/io_dat_i[13] cb_3_9/io_dat_i[14]
+ cb_3_9/io_dat_i[15] cb_3_9/io_dat_i[1] cb_3_9/io_dat_i[2] cb_3_9/io_dat_i[3] cb_3_9/io_dat_i[4]
+ cb_3_9/io_dat_i[5] cb_3_9/io_dat_i[6] cb_3_9/io_dat_i[7] cb_3_9/io_dat_i[8] cb_3_9/io_dat_i[9]
+ cb_3_4/io_dat_o[0] cb_3_4/io_dat_o[10] cb_3_4/io_dat_o[11] cb_3_4/io_dat_o[12] cb_3_4/io_dat_o[13]
+ cb_3_4/io_dat_o[14] cb_3_4/io_dat_o[15] cb_3_4/io_dat_o[1] cb_3_4/io_dat_o[2] cb_3_4/io_dat_o[3]
+ cb_3_4/io_dat_o[4] cb_3_4/io_dat_o[5] cb_3_4/io_dat_o[6] cb_3_4/io_dat_o[7] cb_3_4/io_dat_o[8]
+ cb_3_4/io_dat_o[9] cb_3_5/io_wo[0] cb_3_5/io_wo[10] cb_3_5/io_wo[11] cb_3_5/io_wo[12]
+ cb_3_5/io_wo[13] cb_3_5/io_wo[14] cb_3_5/io_wo[15] cb_3_5/io_wo[16] cb_3_5/io_wo[17]
+ cb_3_5/io_wo[18] cb_3_5/io_wo[19] cb_3_5/io_wo[1] cb_3_5/io_wo[20] cb_3_5/io_wo[21]
+ cb_3_5/io_wo[22] cb_3_5/io_wo[23] cb_3_5/io_wo[24] cb_3_5/io_wo[25] cb_3_5/io_wo[26]
+ cb_3_5/io_wo[27] cb_3_5/io_wo[28] cb_3_5/io_wo[29] cb_3_5/io_wo[2] cb_3_5/io_wo[30]
+ cb_3_5/io_wo[31] cb_3_5/io_wo[32] cb_3_5/io_wo[33] cb_3_5/io_wo[34] cb_3_5/io_wo[35]
+ cb_3_5/io_wo[36] cb_3_5/io_wo[37] cb_3_5/io_wo[38] cb_3_5/io_wo[39] cb_3_5/io_wo[3]
+ cb_3_5/io_wo[40] cb_3_5/io_wo[41] cb_3_5/io_wo[42] cb_3_5/io_wo[43] cb_3_5/io_wo[44]
+ cb_3_5/io_wo[45] cb_3_5/io_wo[46] cb_3_5/io_wo[47] cb_3_5/io_wo[48] cb_3_5/io_wo[49]
+ cb_3_5/io_wo[4] cb_3_5/io_wo[50] cb_3_5/io_wo[51] cb_3_5/io_wo[52] cb_3_5/io_wo[53]
+ cb_3_5/io_wo[54] cb_3_5/io_wo[55] cb_3_5/io_wo[56] cb_3_5/io_wo[57] cb_3_5/io_wo[58]
+ cb_3_5/io_wo[59] cb_3_5/io_wo[5] cb_3_5/io_wo[60] cb_3_5/io_wo[61] cb_3_5/io_wo[62]
+ cb_3_5/io_wo[63] cb_3_5/io_wo[6] cb_3_5/io_wo[7] cb_3_5/io_wo[8] cb_3_5/io_wo[9]
+ cb_3_4/io_i_0_ci cb_3_4/io_i_0_in1[0] cb_3_4/io_i_0_in1[1] cb_3_4/io_i_0_in1[2]
+ cb_3_4/io_i_0_in1[3] cb_3_4/io_i_0_in1[4] cb_3_4/io_i_0_in1[5] cb_3_4/io_i_0_in1[6]
+ cb_3_4/io_i_0_in1[7] cb_3_4/io_i_1_ci cb_3_4/io_i_1_in1[0] cb_3_4/io_i_1_in1[1]
+ cb_3_4/io_i_1_in1[2] cb_3_4/io_i_1_in1[3] cb_3_4/io_i_1_in1[4] cb_3_4/io_i_1_in1[5]
+ cb_3_4/io_i_1_in1[6] cb_3_4/io_i_1_in1[7] cb_3_4/io_i_2_ci cb_3_4/io_i_2_in1[0]
+ cb_3_4/io_i_2_in1[1] cb_3_4/io_i_2_in1[2] cb_3_4/io_i_2_in1[3] cb_3_4/io_i_2_in1[4]
+ cb_3_4/io_i_2_in1[5] cb_3_4/io_i_2_in1[6] cb_3_4/io_i_2_in1[7] cb_3_4/io_i_3_ci
+ cb_3_4/io_i_3_in1[0] cb_3_4/io_i_3_in1[1] cb_3_4/io_i_3_in1[2] cb_3_4/io_i_3_in1[3]
+ cb_3_4/io_i_3_in1[4] cb_3_4/io_i_3_in1[5] cb_3_4/io_i_3_in1[6] cb_3_4/io_i_3_in1[7]
+ cb_3_4/io_i_4_ci cb_3_4/io_i_4_in1[0] cb_3_4/io_i_4_in1[1] cb_3_4/io_i_4_in1[2]
+ cb_3_4/io_i_4_in1[3] cb_3_4/io_i_4_in1[4] cb_3_4/io_i_4_in1[5] cb_3_4/io_i_4_in1[6]
+ cb_3_4/io_i_4_in1[7] cb_3_4/io_i_5_ci cb_3_4/io_i_5_in1[0] cb_3_4/io_i_5_in1[1]
+ cb_3_4/io_i_5_in1[2] cb_3_4/io_i_5_in1[3] cb_3_4/io_i_5_in1[4] cb_3_4/io_i_5_in1[5]
+ cb_3_4/io_i_5_in1[6] cb_3_4/io_i_5_in1[7] cb_3_4/io_i_6_ci cb_3_4/io_i_6_in1[0]
+ cb_3_4/io_i_6_in1[1] cb_3_4/io_i_6_in1[2] cb_3_4/io_i_6_in1[3] cb_3_4/io_i_6_in1[4]
+ cb_3_4/io_i_6_in1[5] cb_3_4/io_i_6_in1[6] cb_3_4/io_i_6_in1[7] cb_3_4/io_i_7_ci
+ cb_3_4/io_i_7_in1[0] cb_3_4/io_i_7_in1[1] cb_3_4/io_i_7_in1[2] cb_3_4/io_i_7_in1[3]
+ cb_3_4/io_i_7_in1[4] cb_3_4/io_i_7_in1[5] cb_3_4/io_i_7_in1[6] cb_3_4/io_i_7_in1[7]
+ cb_3_5/io_i_0_ci cb_3_5/io_i_0_in1[0] cb_3_5/io_i_0_in1[1] cb_3_5/io_i_0_in1[2]
+ cb_3_5/io_i_0_in1[3] cb_3_5/io_i_0_in1[4] cb_3_5/io_i_0_in1[5] cb_3_5/io_i_0_in1[6]
+ cb_3_5/io_i_0_in1[7] cb_3_5/io_i_1_ci cb_3_5/io_i_1_in1[0] cb_3_5/io_i_1_in1[1]
+ cb_3_5/io_i_1_in1[2] cb_3_5/io_i_1_in1[3] cb_3_5/io_i_1_in1[4] cb_3_5/io_i_1_in1[5]
+ cb_3_5/io_i_1_in1[6] cb_3_5/io_i_1_in1[7] cb_3_5/io_i_2_ci cb_3_5/io_i_2_in1[0]
+ cb_3_5/io_i_2_in1[1] cb_3_5/io_i_2_in1[2] cb_3_5/io_i_2_in1[3] cb_3_5/io_i_2_in1[4]
+ cb_3_5/io_i_2_in1[5] cb_3_5/io_i_2_in1[6] cb_3_5/io_i_2_in1[7] cb_3_5/io_i_3_ci
+ cb_3_5/io_i_3_in1[0] cb_3_5/io_i_3_in1[1] cb_3_5/io_i_3_in1[2] cb_3_5/io_i_3_in1[3]
+ cb_3_5/io_i_3_in1[4] cb_3_5/io_i_3_in1[5] cb_3_5/io_i_3_in1[6] cb_3_5/io_i_3_in1[7]
+ cb_3_5/io_i_4_ci cb_3_5/io_i_4_in1[0] cb_3_5/io_i_4_in1[1] cb_3_5/io_i_4_in1[2]
+ cb_3_5/io_i_4_in1[3] cb_3_5/io_i_4_in1[4] cb_3_5/io_i_4_in1[5] cb_3_5/io_i_4_in1[6]
+ cb_3_5/io_i_4_in1[7] cb_3_5/io_i_5_ci cb_3_5/io_i_5_in1[0] cb_3_5/io_i_5_in1[1]
+ cb_3_5/io_i_5_in1[2] cb_3_5/io_i_5_in1[3] cb_3_5/io_i_5_in1[4] cb_3_5/io_i_5_in1[5]
+ cb_3_5/io_i_5_in1[6] cb_3_5/io_i_5_in1[7] cb_3_5/io_i_6_ci cb_3_5/io_i_6_in1[0]
+ cb_3_5/io_i_6_in1[1] cb_3_5/io_i_6_in1[2] cb_3_5/io_i_6_in1[3] cb_3_5/io_i_6_in1[4]
+ cb_3_5/io_i_6_in1[5] cb_3_5/io_i_6_in1[6] cb_3_5/io_i_6_in1[7] cb_3_5/io_i_7_ci
+ cb_3_5/io_i_7_in1[0] cb_3_5/io_i_7_in1[1] cb_3_5/io_i_7_in1[2] cb_3_5/io_i_7_in1[3]
+ cb_3_5/io_i_7_in1[4] cb_3_5/io_i_7_in1[5] cb_3_5/io_i_7_in1[6] cb_3_5/io_i_7_in1[7]
+ cb_3_4/io_vci cb_3_5/io_vci cb_3_4/io_vi cb_3_9/io_we_i cb_3_4/io_wo[0] cb_3_4/io_wo[10]
+ cb_3_4/io_wo[11] cb_3_4/io_wo[12] cb_3_4/io_wo[13] cb_3_4/io_wo[14] cb_3_4/io_wo[15]
+ cb_3_4/io_wo[16] cb_3_4/io_wo[17] cb_3_4/io_wo[18] cb_3_4/io_wo[19] cb_3_4/io_wo[1]
+ cb_3_4/io_wo[20] cb_3_4/io_wo[21] cb_3_4/io_wo[22] cb_3_4/io_wo[23] cb_3_4/io_wo[24]
+ cb_3_4/io_wo[25] cb_3_4/io_wo[26] cb_3_4/io_wo[27] cb_3_4/io_wo[28] cb_3_4/io_wo[29]
+ cb_3_4/io_wo[2] cb_3_4/io_wo[30] cb_3_4/io_wo[31] cb_3_4/io_wo[32] cb_3_4/io_wo[33]
+ cb_3_4/io_wo[34] cb_3_4/io_wo[35] cb_3_4/io_wo[36] cb_3_4/io_wo[37] cb_3_4/io_wo[38]
+ cb_3_4/io_wo[39] cb_3_4/io_wo[3] cb_3_4/io_wo[40] cb_3_4/io_wo[41] cb_3_4/io_wo[42]
+ cb_3_4/io_wo[43] cb_3_4/io_wo[44] cb_3_4/io_wo[45] cb_3_4/io_wo[46] cb_3_4/io_wo[47]
+ cb_3_4/io_wo[48] cb_3_4/io_wo[49] cb_3_4/io_wo[4] cb_3_4/io_wo[50] cb_3_4/io_wo[51]
+ cb_3_4/io_wo[52] cb_3_4/io_wo[53] cb_3_4/io_wo[54] cb_3_4/io_wo[55] cb_3_4/io_wo[56]
+ cb_3_4/io_wo[57] cb_3_4/io_wo[58] cb_3_4/io_wo[59] cb_3_4/io_wo[5] cb_3_4/io_wo[60]
+ cb_3_4/io_wo[61] cb_3_4/io_wo[62] cb_3_4/io_wo[63] cb_3_4/io_wo[6] cb_3_4/io_wo[7]
+ cb_3_4/io_wo[8] cb_3_4/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_1_1 cb_1_9/io_adr_i[0] cb_1_9/io_adr_i[1] cb_1_1/io_cs_i cb_1_9/io_dat_i[0] cb_1_9/io_dat_i[10]
+ cb_1_9/io_dat_i[11] cb_1_9/io_dat_i[12] cb_1_9/io_dat_i[13] cb_1_9/io_dat_i[14]
+ cb_1_9/io_dat_i[15] cb_1_9/io_dat_i[1] cb_1_9/io_dat_i[2] cb_1_9/io_dat_i[3] cb_1_9/io_dat_i[4]
+ cb_1_9/io_dat_i[5] cb_1_9/io_dat_i[6] cb_1_9/io_dat_i[7] cb_1_9/io_dat_i[8] cb_1_9/io_dat_i[9]
+ cb_1_1/io_dat_o[0] cb_1_1/io_dat_o[10] cb_1_1/io_dat_o[11] cb_1_1/io_dat_o[12] cb_1_1/io_dat_o[13]
+ cb_1_1/io_dat_o[14] cb_1_1/io_dat_o[15] cb_1_1/io_dat_o[1] cb_1_1/io_dat_o[2] cb_1_1/io_dat_o[3]
+ cb_1_1/io_dat_o[4] cb_1_1/io_dat_o[5] cb_1_1/io_dat_o[6] cb_1_1/io_dat_o[7] cb_1_1/io_dat_o[8]
+ cb_1_1/io_dat_o[9] cb_1_2/io_wo[0] cb_1_2/io_wo[10] cb_1_2/io_wo[11] cb_1_2/io_wo[12]
+ cb_1_2/io_wo[13] cb_1_2/io_wo[14] cb_1_2/io_wo[15] cb_1_2/io_wo[16] cb_1_2/io_wo[17]
+ cb_1_2/io_wo[18] cb_1_2/io_wo[19] cb_1_2/io_wo[1] cb_1_2/io_wo[20] cb_1_2/io_wo[21]
+ cb_1_2/io_wo[22] cb_1_2/io_wo[23] cb_1_2/io_wo[24] cb_1_2/io_wo[25] cb_1_2/io_wo[26]
+ cb_1_2/io_wo[27] cb_1_2/io_wo[28] cb_1_2/io_wo[29] cb_1_2/io_wo[2] cb_1_2/io_wo[30]
+ cb_1_2/io_wo[31] cb_1_2/io_wo[32] cb_1_2/io_wo[33] cb_1_2/io_wo[34] cb_1_2/io_wo[35]
+ cb_1_2/io_wo[36] cb_1_2/io_wo[37] cb_1_2/io_wo[38] cb_1_2/io_wo[39] cb_1_2/io_wo[3]
+ cb_1_2/io_wo[40] cb_1_2/io_wo[41] cb_1_2/io_wo[42] cb_1_2/io_wo[43] cb_1_2/io_wo[44]
+ cb_1_2/io_wo[45] cb_1_2/io_wo[46] cb_1_2/io_wo[47] cb_1_2/io_wo[48] cb_1_2/io_wo[49]
+ cb_1_2/io_wo[4] cb_1_2/io_wo[50] cb_1_2/io_wo[51] cb_1_2/io_wo[52] cb_1_2/io_wo[53]
+ cb_1_2/io_wo[54] cb_1_2/io_wo[55] cb_1_2/io_wo[56] cb_1_2/io_wo[57] cb_1_2/io_wo[58]
+ cb_1_2/io_wo[59] cb_1_2/io_wo[5] cb_1_2/io_wo[60] cb_1_2/io_wo[61] cb_1_2/io_wo[62]
+ cb_1_2/io_wo[63] cb_1_2/io_wo[6] cb_1_2/io_wo[7] cb_1_2/io_wo[8] cb_1_2/io_wo[9]
+ cb_1_1/io_i_0_ci cb_1_1/io_i_0_in1[0] cb_1_1/io_i_0_in1[1] cb_1_1/io_i_0_in1[2]
+ cb_1_1/io_i_0_in1[3] cb_1_1/io_i_0_in1[4] cb_1_1/io_i_0_in1[5] cb_1_1/io_i_0_in1[6]
+ cb_1_1/io_i_0_in1[7] cb_1_1/io_i_1_ci cb_1_1/io_i_1_in1[0] cb_1_1/io_i_1_in1[1]
+ cb_1_1/io_i_1_in1[2] cb_1_1/io_i_1_in1[3] cb_1_1/io_i_1_in1[4] cb_1_1/io_i_1_in1[5]
+ cb_1_1/io_i_1_in1[6] cb_1_1/io_i_1_in1[7] cb_1_1/io_i_2_ci cb_1_1/io_i_2_in1[0]
+ cb_1_1/io_i_2_in1[1] cb_1_1/io_i_2_in1[2] cb_1_1/io_i_2_in1[3] cb_1_1/io_i_2_in1[4]
+ cb_1_1/io_i_2_in1[5] cb_1_1/io_i_2_in1[6] cb_1_1/io_i_2_in1[7] cb_1_1/io_i_3_ci
+ cb_1_1/io_i_3_in1[0] cb_1_1/io_i_3_in1[1] cb_1_1/io_i_3_in1[2] cb_1_1/io_i_3_in1[3]
+ cb_1_1/io_i_3_in1[4] cb_1_1/io_i_3_in1[5] cb_1_1/io_i_3_in1[6] cb_1_1/io_i_3_in1[7]
+ cb_1_1/io_i_4_ci cb_1_1/io_i_4_in1[0] cb_1_1/io_i_4_in1[1] cb_1_1/io_i_4_in1[2]
+ cb_1_1/io_i_4_in1[3] cb_1_1/io_i_4_in1[4] cb_1_1/io_i_4_in1[5] cb_1_1/io_i_4_in1[6]
+ cb_1_1/io_i_4_in1[7] cb_1_1/io_i_5_ci cb_1_1/io_i_5_in1[0] cb_1_1/io_i_5_in1[1]
+ cb_1_1/io_i_5_in1[2] cb_1_1/io_i_5_in1[3] cb_1_1/io_i_5_in1[4] cb_1_1/io_i_5_in1[5]
+ cb_1_1/io_i_5_in1[6] cb_1_1/io_i_5_in1[7] cb_1_1/io_i_6_ci cb_1_1/io_i_6_in1[0]
+ cb_1_1/io_i_6_in1[1] cb_1_1/io_i_6_in1[2] cb_1_1/io_i_6_in1[3] cb_1_1/io_i_6_in1[4]
+ cb_1_1/io_i_6_in1[5] cb_1_1/io_i_6_in1[6] cb_1_1/io_i_6_in1[7] cb_1_1/io_i_7_ci
+ cb_1_1/io_i_7_in1[0] cb_1_1/io_i_7_in1[1] cb_1_1/io_i_7_in1[2] cb_1_1/io_i_7_in1[3]
+ cb_1_1/io_i_7_in1[4] cb_1_1/io_i_7_in1[5] cb_1_1/io_i_7_in1[6] cb_1_1/io_i_7_in1[7]
+ cb_1_2/io_i_0_ci cb_1_2/io_i_0_in1[0] cb_1_2/io_i_0_in1[1] cb_1_2/io_i_0_in1[2]
+ cb_1_2/io_i_0_in1[3] cb_1_2/io_i_0_in1[4] cb_1_2/io_i_0_in1[5] cb_1_2/io_i_0_in1[6]
+ cb_1_2/io_i_0_in1[7] cb_1_2/io_i_1_ci cb_1_2/io_i_1_in1[0] cb_1_2/io_i_1_in1[1]
+ cb_1_2/io_i_1_in1[2] cb_1_2/io_i_1_in1[3] cb_1_2/io_i_1_in1[4] cb_1_2/io_i_1_in1[5]
+ cb_1_2/io_i_1_in1[6] cb_1_2/io_i_1_in1[7] cb_1_2/io_i_2_ci cb_1_2/io_i_2_in1[0]
+ cb_1_2/io_i_2_in1[1] cb_1_2/io_i_2_in1[2] cb_1_2/io_i_2_in1[3] cb_1_2/io_i_2_in1[4]
+ cb_1_2/io_i_2_in1[5] cb_1_2/io_i_2_in1[6] cb_1_2/io_i_2_in1[7] cb_1_2/io_i_3_ci
+ cb_1_2/io_i_3_in1[0] cb_1_2/io_i_3_in1[1] cb_1_2/io_i_3_in1[2] cb_1_2/io_i_3_in1[3]
+ cb_1_2/io_i_3_in1[4] cb_1_2/io_i_3_in1[5] cb_1_2/io_i_3_in1[6] cb_1_2/io_i_3_in1[7]
+ cb_1_2/io_i_4_ci cb_1_2/io_i_4_in1[0] cb_1_2/io_i_4_in1[1] cb_1_2/io_i_4_in1[2]
+ cb_1_2/io_i_4_in1[3] cb_1_2/io_i_4_in1[4] cb_1_2/io_i_4_in1[5] cb_1_2/io_i_4_in1[6]
+ cb_1_2/io_i_4_in1[7] cb_1_2/io_i_5_ci cb_1_2/io_i_5_in1[0] cb_1_2/io_i_5_in1[1]
+ cb_1_2/io_i_5_in1[2] cb_1_2/io_i_5_in1[3] cb_1_2/io_i_5_in1[4] cb_1_2/io_i_5_in1[5]
+ cb_1_2/io_i_5_in1[6] cb_1_2/io_i_5_in1[7] cb_1_2/io_i_6_ci cb_1_2/io_i_6_in1[0]
+ cb_1_2/io_i_6_in1[1] cb_1_2/io_i_6_in1[2] cb_1_2/io_i_6_in1[3] cb_1_2/io_i_6_in1[4]
+ cb_1_2/io_i_6_in1[5] cb_1_2/io_i_6_in1[6] cb_1_2/io_i_6_in1[7] cb_1_2/io_i_7_ci
+ cb_1_2/io_i_7_in1[0] cb_1_2/io_i_7_in1[1] cb_1_2/io_i_7_in1[2] cb_1_2/io_i_7_in1[3]
+ cb_1_2/io_i_7_in1[4] cb_1_2/io_i_7_in1[5] cb_1_2/io_i_7_in1[6] cb_1_2/io_i_7_in1[7]
+ cb_1_1/io_vci cb_1_2/io_vci cb_1_1/io_vi cb_1_9/io_we_i cb_1_1/io_wo[0] cb_1_1/io_wo[10]
+ cb_1_1/io_wo[11] cb_1_1/io_wo[12] cb_1_1/io_wo[13] cb_1_1/io_wo[14] cb_1_1/io_wo[15]
+ cb_1_1/io_wo[16] cb_1_1/io_wo[17] cb_1_1/io_wo[18] cb_1_1/io_wo[19] cb_1_1/io_wo[1]
+ cb_1_1/io_wo[20] cb_1_1/io_wo[21] cb_1_1/io_wo[22] cb_1_1/io_wo[23] cb_1_1/io_wo[24]
+ cb_1_1/io_wo[25] cb_1_1/io_wo[26] cb_1_1/io_wo[27] cb_1_1/io_wo[28] cb_1_1/io_wo[29]
+ cb_1_1/io_wo[2] cb_1_1/io_wo[30] cb_1_1/io_wo[31] cb_1_1/io_wo[32] cb_1_1/io_wo[33]
+ cb_1_1/io_wo[34] cb_1_1/io_wo[35] cb_1_1/io_wo[36] cb_1_1/io_wo[37] cb_1_1/io_wo[38]
+ cb_1_1/io_wo[39] cb_1_1/io_wo[3] cb_1_1/io_wo[40] cb_1_1/io_wo[41] cb_1_1/io_wo[42]
+ cb_1_1/io_wo[43] cb_1_1/io_wo[44] cb_1_1/io_wo[45] cb_1_1/io_wo[46] cb_1_1/io_wo[47]
+ cb_1_1/io_wo[48] cb_1_1/io_wo[49] cb_1_1/io_wo[4] cb_1_1/io_wo[50] cb_1_1/io_wo[51]
+ cb_1_1/io_wo[52] cb_1_1/io_wo[53] cb_1_1/io_wo[54] cb_1_1/io_wo[55] cb_1_1/io_wo[56]
+ cb_1_1/io_wo[57] cb_1_1/io_wo[58] cb_1_1/io_wo[59] cb_1_1/io_wo[5] cb_1_1/io_wo[60]
+ cb_1_1/io_wo[61] cb_1_1/io_wo[62] cb_1_1/io_wo[63] cb_1_1/io_wo[6] cb_1_1/io_wo[7]
+ cb_1_1/io_wo[8] cb_1_1/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xccon_4 ccon_4/io_ack_o ccon_7/io_adr_i[0] ccon_7/io_adr_i[10] ccon_7/io_adr_i[11]
+ ccon_7/io_adr_i[1] ccon_7/io_adr_i[2] ccon_7/io_adr_i[3] ccon_7/io_adr_i[4] ccon_7/io_adr_i[5]
+ ccon_7/io_adr_i[6] ccon_7/io_adr_i[7] ccon_7/io_adr_i[8] ccon_7/io_adr_i[9] cb_4_9/io_adr_i[0]
+ cb_4_9/io_adr_i[1] cb_4_0/io_cs_i cb_4_1/io_cs_i cb_4_10/io_cs_i cb_4_2/io_cs_i
+ cb_4_3/io_cs_i cb_4_4/io_cs_i cb_4_5/io_cs_i cb_4_6/io_cs_i cb_4_7/io_cs_i cb_4_8/io_cs_i
+ cb_4_9/io_cs_i cb_4_9/io_dat_i[0] cb_4_9/io_dat_i[10] cb_4_9/io_dat_i[11] cb_4_9/io_dat_i[12]
+ cb_4_9/io_dat_i[13] cb_4_9/io_dat_i[14] cb_4_9/io_dat_i[15] cb_4_9/io_dat_i[1] cb_4_9/io_dat_i[2]
+ cb_4_9/io_dat_i[3] cb_4_9/io_dat_i[4] cb_4_9/io_dat_i[5] cb_4_9/io_dat_i[6] cb_4_9/io_dat_i[7]
+ cb_4_9/io_dat_i[8] cb_4_9/io_dat_i[9] cb_4_0/io_dat_o[0] cb_4_0/io_dat_o[10] cb_4_0/io_dat_o[11]
+ cb_4_0/io_dat_o[12] cb_4_0/io_dat_o[13] cb_4_0/io_dat_o[14] cb_4_0/io_dat_o[15]
+ cb_4_0/io_dat_o[1] cb_4_0/io_dat_o[2] cb_4_0/io_dat_o[3] cb_4_0/io_dat_o[4] cb_4_0/io_dat_o[5]
+ cb_4_0/io_dat_o[6] cb_4_0/io_dat_o[7] cb_4_0/io_dat_o[8] cb_4_0/io_dat_o[9] cb_4_10/io_dat_o[0]
+ cb_4_10/io_dat_o[10] cb_4_10/io_dat_o[11] cb_4_10/io_dat_o[12] cb_4_10/io_dat_o[13]
+ cb_4_10/io_dat_o[14] cb_4_10/io_dat_o[15] cb_4_10/io_dat_o[1] cb_4_10/io_dat_o[2]
+ cb_4_10/io_dat_o[3] cb_4_10/io_dat_o[4] cb_4_10/io_dat_o[5] cb_4_10/io_dat_o[6]
+ cb_4_10/io_dat_o[7] cb_4_10/io_dat_o[8] cb_4_10/io_dat_o[9] cb_4_1/io_dat_o[0] cb_4_1/io_dat_o[10]
+ cb_4_1/io_dat_o[11] cb_4_1/io_dat_o[12] cb_4_1/io_dat_o[13] cb_4_1/io_dat_o[14]
+ cb_4_1/io_dat_o[15] cb_4_1/io_dat_o[1] cb_4_1/io_dat_o[2] cb_4_1/io_dat_o[3] cb_4_1/io_dat_o[4]
+ cb_4_1/io_dat_o[5] cb_4_1/io_dat_o[6] cb_4_1/io_dat_o[7] cb_4_1/io_dat_o[8] cb_4_1/io_dat_o[9]
+ cb_4_2/io_dat_o[0] cb_4_2/io_dat_o[10] cb_4_2/io_dat_o[11] cb_4_2/io_dat_o[12] cb_4_2/io_dat_o[13]
+ cb_4_2/io_dat_o[14] cb_4_2/io_dat_o[15] cb_4_2/io_dat_o[1] cb_4_2/io_dat_o[2] cb_4_2/io_dat_o[3]
+ cb_4_2/io_dat_o[4] cb_4_2/io_dat_o[5] cb_4_2/io_dat_o[6] cb_4_2/io_dat_o[7] cb_4_2/io_dat_o[8]
+ cb_4_2/io_dat_o[9] cb_4_3/io_dat_o[0] cb_4_3/io_dat_o[10] cb_4_3/io_dat_o[11] cb_4_3/io_dat_o[12]
+ cb_4_3/io_dat_o[13] cb_4_3/io_dat_o[14] cb_4_3/io_dat_o[15] cb_4_3/io_dat_o[1] cb_4_3/io_dat_o[2]
+ cb_4_3/io_dat_o[3] cb_4_3/io_dat_o[4] cb_4_3/io_dat_o[5] cb_4_3/io_dat_o[6] cb_4_3/io_dat_o[7]
+ cb_4_3/io_dat_o[8] cb_4_3/io_dat_o[9] cb_4_4/io_dat_o[0] cb_4_4/io_dat_o[10] cb_4_4/io_dat_o[11]
+ cb_4_4/io_dat_o[12] cb_4_4/io_dat_o[13] cb_4_4/io_dat_o[14] cb_4_4/io_dat_o[15]
+ cb_4_4/io_dat_o[1] cb_4_4/io_dat_o[2] cb_4_4/io_dat_o[3] cb_4_4/io_dat_o[4] cb_4_4/io_dat_o[5]
+ cb_4_4/io_dat_o[6] cb_4_4/io_dat_o[7] cb_4_4/io_dat_o[8] cb_4_4/io_dat_o[9] cb_4_5/io_dat_o[0]
+ cb_4_5/io_dat_o[10] cb_4_5/io_dat_o[11] cb_4_5/io_dat_o[12] cb_4_5/io_dat_o[13]
+ cb_4_5/io_dat_o[14] cb_4_5/io_dat_o[15] cb_4_5/io_dat_o[1] cb_4_5/io_dat_o[2] cb_4_5/io_dat_o[3]
+ cb_4_5/io_dat_o[4] cb_4_5/io_dat_o[5] cb_4_5/io_dat_o[6] cb_4_5/io_dat_o[7] cb_4_5/io_dat_o[8]
+ cb_4_5/io_dat_o[9] cb_4_6/io_dat_o[0] cb_4_6/io_dat_o[10] cb_4_6/io_dat_o[11] cb_4_6/io_dat_o[12]
+ cb_4_6/io_dat_o[13] cb_4_6/io_dat_o[14] cb_4_6/io_dat_o[15] cb_4_6/io_dat_o[1] cb_4_6/io_dat_o[2]
+ cb_4_6/io_dat_o[3] cb_4_6/io_dat_o[4] cb_4_6/io_dat_o[5] cb_4_6/io_dat_o[6] cb_4_6/io_dat_o[7]
+ cb_4_6/io_dat_o[8] cb_4_6/io_dat_o[9] cb_4_7/io_dat_o[0] cb_4_7/io_dat_o[10] cb_4_7/io_dat_o[11]
+ cb_4_7/io_dat_o[12] cb_4_7/io_dat_o[13] cb_4_7/io_dat_o[14] cb_4_7/io_dat_o[15]
+ cb_4_7/io_dat_o[1] cb_4_7/io_dat_o[2] cb_4_7/io_dat_o[3] cb_4_7/io_dat_o[4] cb_4_7/io_dat_o[5]
+ cb_4_7/io_dat_o[6] cb_4_7/io_dat_o[7] cb_4_7/io_dat_o[8] cb_4_7/io_dat_o[9] cb_4_8/io_dat_o[0]
+ cb_4_8/io_dat_o[10] cb_4_8/io_dat_o[11] cb_4_8/io_dat_o[12] cb_4_8/io_dat_o[13]
+ cb_4_8/io_dat_o[14] cb_4_8/io_dat_o[15] cb_4_8/io_dat_o[1] cb_4_8/io_dat_o[2] cb_4_8/io_dat_o[3]
+ cb_4_8/io_dat_o[4] cb_4_8/io_dat_o[5] cb_4_8/io_dat_o[6] cb_4_8/io_dat_o[7] cb_4_8/io_dat_o[8]
+ cb_4_8/io_dat_o[9] cb_4_9/io_dat_o[0] cb_4_9/io_dat_o[10] cb_4_9/io_dat_o[11] cb_4_9/io_dat_o[12]
+ cb_4_9/io_dat_o[13] cb_4_9/io_dat_o[14] cb_4_9/io_dat_o[15] cb_4_9/io_dat_o[1] cb_4_9/io_dat_o[2]
+ cb_4_9/io_dat_o[3] cb_4_9/io_dat_o[4] cb_4_9/io_dat_o[5] cb_4_9/io_dat_o[6] cb_4_9/io_dat_o[7]
+ cb_4_9/io_dat_o[8] cb_4_9/io_dat_o[9] cb_4_9/io_we_i ccon_4/io_cs_i ccon_7/io_dat_i[0]
+ ccon_7/io_dat_i[10] ccon_7/io_dat_i[11] ccon_7/io_dat_i[12] ccon_7/io_dat_i[13]
+ ccon_7/io_dat_i[14] ccon_7/io_dat_i[15] ccon_7/io_dat_i[16] ccon_7/io_dat_i[17]
+ ccon_7/io_dat_i[18] ccon_7/io_dat_i[19] ccon_7/io_dat_i[1] ccon_7/io_dat_i[20] ccon_7/io_dat_i[21]
+ ccon_7/io_dat_i[22] ccon_7/io_dat_i[23] ccon_7/io_dat_i[24] ccon_7/io_dat_i[25]
+ ccon_7/io_dat_i[26] ccon_7/io_dat_i[27] ccon_7/io_dat_i[28] ccon_7/io_dat_i[29]
+ ccon_7/io_dat_i[2] ccon_7/io_dat_i[30] ccon_7/io_dat_i[31] ccon_7/io_dat_i[3] ccon_7/io_dat_i[4]
+ ccon_7/io_dat_i[5] ccon_7/io_dat_i[6] ccon_7/io_dat_i[7] ccon_7/io_dat_i[8] ccon_7/io_dat_i[9]
+ ccon_4/io_dat_o[0] ccon_4/io_dat_o[10] ccon_4/io_dat_o[11] ccon_4/io_dat_o[12] ccon_4/io_dat_o[13]
+ ccon_4/io_dat_o[14] ccon_4/io_dat_o[15] ccon_4/io_dat_o[16] ccon_4/io_dat_o[17]
+ ccon_4/io_dat_o[18] ccon_4/io_dat_o[19] ccon_4/io_dat_o[1] ccon_4/io_dat_o[20] ccon_4/io_dat_o[21]
+ ccon_4/io_dat_o[22] ccon_4/io_dat_o[23] ccon_4/io_dat_o[24] ccon_4/io_dat_o[25]
+ ccon_4/io_dat_o[26] ccon_4/io_dat_o[27] ccon_4/io_dat_o[28] ccon_4/io_dat_o[29]
+ ccon_4/io_dat_o[2] ccon_4/io_dat_o[30] ccon_4/io_dat_o[31] ccon_4/io_dat_o[3] ccon_4/io_dat_o[4]
+ ccon_4/io_dat_o[5] ccon_4/io_dat_o[6] ccon_4/io_dat_o[7] ccon_4/io_dat_o[8] ccon_4/io_dat_o[9]
+ cb_4_0/io_wo[0] cb_4_0/io_wo[10] cb_4_0/io_wo[11] cb_4_0/io_wo[12] cb_4_0/io_wo[13]
+ cb_4_0/io_wo[14] cb_4_0/io_wo[15] cb_4_0/io_wo[16] cb_4_0/io_wo[17] cb_4_0/io_wo[18]
+ cb_4_0/io_wo[19] cb_4_0/io_wo[1] cb_4_0/io_wo[20] cb_4_0/io_wo[21] cb_4_0/io_wo[22]
+ cb_4_0/io_wo[23] cb_4_0/io_wo[24] cb_4_0/io_wo[25] cb_4_0/io_wo[26] cb_4_0/io_wo[27]
+ cb_4_0/io_wo[28] cb_4_0/io_wo[29] cb_4_0/io_wo[2] cb_4_0/io_wo[30] cb_4_0/io_wo[31]
+ cb_4_0/io_wo[32] cb_4_0/io_wo[33] cb_4_0/io_wo[34] cb_4_0/io_wo[35] cb_4_0/io_wo[36]
+ cb_4_0/io_wo[37] cb_4_0/io_wo[38] cb_4_0/io_wo[39] cb_4_0/io_wo[3] cb_4_0/io_wo[40]
+ cb_4_0/io_wo[41] cb_4_0/io_wo[42] cb_4_0/io_wo[43] cb_4_0/io_wo[44] cb_4_0/io_wo[45]
+ cb_4_0/io_wo[46] cb_4_0/io_wo[47] cb_4_0/io_wo[48] cb_4_0/io_wo[49] cb_4_0/io_wo[4]
+ cb_4_0/io_wo[50] cb_4_0/io_wo[51] cb_4_0/io_wo[52] cb_4_0/io_wo[53] cb_4_0/io_wo[54]
+ cb_4_0/io_wo[55] cb_4_0/io_wo[56] cb_4_0/io_wo[57] cb_4_0/io_wo[58] cb_4_0/io_wo[59]
+ cb_4_0/io_wo[5] cb_4_0/io_wo[60] cb_4_0/io_wo[61] cb_4_0/io_wo[62] cb_4_0/io_wo[63]
+ cb_4_0/io_wo[6] cb_4_0/io_wo[7] cb_4_0/io_wo[8] cb_4_0/io_wo[9] icon/dsi[0] icon/dsi[1]
+ icon/dsi[2] icon/dsi[3] icon/dsi[4] icon/dsi[5] icon/dsi[6] icon/dsi[7] ccon_4/io_dsi_o
+ ccon_4/io_irq cb_4_0/io_vi cb_4_10/io_vi cb_4_1/io_vi cb_4_2/io_vi cb_4_3/io_vi
+ cb_4_4/io_vi cb_4_5/io_vi cb_4_6/io_vi cb_4_7/io_vi cb_4_8/io_vi cb_4_9/io_vi ccon_7/io_we_i
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_con
Xcb_5_8 cb_5_9/io_adr_i[0] cb_5_9/io_adr_i[1] cb_5_8/io_cs_i cb_5_9/io_dat_i[0] cb_5_9/io_dat_i[10]
+ cb_5_9/io_dat_i[11] cb_5_9/io_dat_i[12] cb_5_9/io_dat_i[13] cb_5_9/io_dat_i[14]
+ cb_5_9/io_dat_i[15] cb_5_9/io_dat_i[1] cb_5_9/io_dat_i[2] cb_5_9/io_dat_i[3] cb_5_9/io_dat_i[4]
+ cb_5_9/io_dat_i[5] cb_5_9/io_dat_i[6] cb_5_9/io_dat_i[7] cb_5_9/io_dat_i[8] cb_5_9/io_dat_i[9]
+ cb_5_8/io_dat_o[0] cb_5_8/io_dat_o[10] cb_5_8/io_dat_o[11] cb_5_8/io_dat_o[12] cb_5_8/io_dat_o[13]
+ cb_5_8/io_dat_o[14] cb_5_8/io_dat_o[15] cb_5_8/io_dat_o[1] cb_5_8/io_dat_o[2] cb_5_8/io_dat_o[3]
+ cb_5_8/io_dat_o[4] cb_5_8/io_dat_o[5] cb_5_8/io_dat_o[6] cb_5_8/io_dat_o[7] cb_5_8/io_dat_o[8]
+ cb_5_8/io_dat_o[9] cb_5_9/io_wo[0] cb_5_9/io_wo[10] cb_5_9/io_wo[11] cb_5_9/io_wo[12]
+ cb_5_9/io_wo[13] cb_5_9/io_wo[14] cb_5_9/io_wo[15] cb_5_9/io_wo[16] cb_5_9/io_wo[17]
+ cb_5_9/io_wo[18] cb_5_9/io_wo[19] cb_5_9/io_wo[1] cb_5_9/io_wo[20] cb_5_9/io_wo[21]
+ cb_5_9/io_wo[22] cb_5_9/io_wo[23] cb_5_9/io_wo[24] cb_5_9/io_wo[25] cb_5_9/io_wo[26]
+ cb_5_9/io_wo[27] cb_5_9/io_wo[28] cb_5_9/io_wo[29] cb_5_9/io_wo[2] cb_5_9/io_wo[30]
+ cb_5_9/io_wo[31] cb_5_9/io_wo[32] cb_5_9/io_wo[33] cb_5_9/io_wo[34] cb_5_9/io_wo[35]
+ cb_5_9/io_wo[36] cb_5_9/io_wo[37] cb_5_9/io_wo[38] cb_5_9/io_wo[39] cb_5_9/io_wo[3]
+ cb_5_9/io_wo[40] cb_5_9/io_wo[41] cb_5_9/io_wo[42] cb_5_9/io_wo[43] cb_5_9/io_wo[44]
+ cb_5_9/io_wo[45] cb_5_9/io_wo[46] cb_5_9/io_wo[47] cb_5_9/io_wo[48] cb_5_9/io_wo[49]
+ cb_5_9/io_wo[4] cb_5_9/io_wo[50] cb_5_9/io_wo[51] cb_5_9/io_wo[52] cb_5_9/io_wo[53]
+ cb_5_9/io_wo[54] cb_5_9/io_wo[55] cb_5_9/io_wo[56] cb_5_9/io_wo[57] cb_5_9/io_wo[58]
+ cb_5_9/io_wo[59] cb_5_9/io_wo[5] cb_5_9/io_wo[60] cb_5_9/io_wo[61] cb_5_9/io_wo[62]
+ cb_5_9/io_wo[63] cb_5_9/io_wo[6] cb_5_9/io_wo[7] cb_5_9/io_wo[8] cb_5_9/io_wo[9]
+ cb_5_8/io_i_0_ci cb_5_8/io_i_0_in1[0] cb_5_8/io_i_0_in1[1] cb_5_8/io_i_0_in1[2]
+ cb_5_8/io_i_0_in1[3] cb_5_8/io_i_0_in1[4] cb_5_8/io_i_0_in1[5] cb_5_8/io_i_0_in1[6]
+ cb_5_8/io_i_0_in1[7] cb_5_8/io_i_1_ci cb_5_8/io_i_1_in1[0] cb_5_8/io_i_1_in1[1]
+ cb_5_8/io_i_1_in1[2] cb_5_8/io_i_1_in1[3] cb_5_8/io_i_1_in1[4] cb_5_8/io_i_1_in1[5]
+ cb_5_8/io_i_1_in1[6] cb_5_8/io_i_1_in1[7] cb_5_8/io_i_2_ci cb_5_8/io_i_2_in1[0]
+ cb_5_8/io_i_2_in1[1] cb_5_8/io_i_2_in1[2] cb_5_8/io_i_2_in1[3] cb_5_8/io_i_2_in1[4]
+ cb_5_8/io_i_2_in1[5] cb_5_8/io_i_2_in1[6] cb_5_8/io_i_2_in1[7] cb_5_8/io_i_3_ci
+ cb_5_8/io_i_3_in1[0] cb_5_8/io_i_3_in1[1] cb_5_8/io_i_3_in1[2] cb_5_8/io_i_3_in1[3]
+ cb_5_8/io_i_3_in1[4] cb_5_8/io_i_3_in1[5] cb_5_8/io_i_3_in1[6] cb_5_8/io_i_3_in1[7]
+ cb_5_8/io_i_4_ci cb_5_8/io_i_4_in1[0] cb_5_8/io_i_4_in1[1] cb_5_8/io_i_4_in1[2]
+ cb_5_8/io_i_4_in1[3] cb_5_8/io_i_4_in1[4] cb_5_8/io_i_4_in1[5] cb_5_8/io_i_4_in1[6]
+ cb_5_8/io_i_4_in1[7] cb_5_8/io_i_5_ci cb_5_8/io_i_5_in1[0] cb_5_8/io_i_5_in1[1]
+ cb_5_8/io_i_5_in1[2] cb_5_8/io_i_5_in1[3] cb_5_8/io_i_5_in1[4] cb_5_8/io_i_5_in1[5]
+ cb_5_8/io_i_5_in1[6] cb_5_8/io_i_5_in1[7] cb_5_8/io_i_6_ci cb_5_8/io_i_6_in1[0]
+ cb_5_8/io_i_6_in1[1] cb_5_8/io_i_6_in1[2] cb_5_8/io_i_6_in1[3] cb_5_8/io_i_6_in1[4]
+ cb_5_8/io_i_6_in1[5] cb_5_8/io_i_6_in1[6] cb_5_8/io_i_6_in1[7] cb_5_8/io_i_7_ci
+ cb_5_8/io_i_7_in1[0] cb_5_8/io_i_7_in1[1] cb_5_8/io_i_7_in1[2] cb_5_8/io_i_7_in1[3]
+ cb_5_8/io_i_7_in1[4] cb_5_8/io_i_7_in1[5] cb_5_8/io_i_7_in1[6] cb_5_8/io_i_7_in1[7]
+ cb_5_9/io_i_0_ci cb_5_9/io_i_0_in1[0] cb_5_9/io_i_0_in1[1] cb_5_9/io_i_0_in1[2]
+ cb_5_9/io_i_0_in1[3] cb_5_9/io_i_0_in1[4] cb_5_9/io_i_0_in1[5] cb_5_9/io_i_0_in1[6]
+ cb_5_9/io_i_0_in1[7] cb_5_9/io_i_1_ci cb_5_9/io_i_1_in1[0] cb_5_9/io_i_1_in1[1]
+ cb_5_9/io_i_1_in1[2] cb_5_9/io_i_1_in1[3] cb_5_9/io_i_1_in1[4] cb_5_9/io_i_1_in1[5]
+ cb_5_9/io_i_1_in1[6] cb_5_9/io_i_1_in1[7] cb_5_9/io_i_2_ci cb_5_9/io_i_2_in1[0]
+ cb_5_9/io_i_2_in1[1] cb_5_9/io_i_2_in1[2] cb_5_9/io_i_2_in1[3] cb_5_9/io_i_2_in1[4]
+ cb_5_9/io_i_2_in1[5] cb_5_9/io_i_2_in1[6] cb_5_9/io_i_2_in1[7] cb_5_9/io_i_3_ci
+ cb_5_9/io_i_3_in1[0] cb_5_9/io_i_3_in1[1] cb_5_9/io_i_3_in1[2] cb_5_9/io_i_3_in1[3]
+ cb_5_9/io_i_3_in1[4] cb_5_9/io_i_3_in1[5] cb_5_9/io_i_3_in1[6] cb_5_9/io_i_3_in1[7]
+ cb_5_9/io_i_4_ci cb_5_9/io_i_4_in1[0] cb_5_9/io_i_4_in1[1] cb_5_9/io_i_4_in1[2]
+ cb_5_9/io_i_4_in1[3] cb_5_9/io_i_4_in1[4] cb_5_9/io_i_4_in1[5] cb_5_9/io_i_4_in1[6]
+ cb_5_9/io_i_4_in1[7] cb_5_9/io_i_5_ci cb_5_9/io_i_5_in1[0] cb_5_9/io_i_5_in1[1]
+ cb_5_9/io_i_5_in1[2] cb_5_9/io_i_5_in1[3] cb_5_9/io_i_5_in1[4] cb_5_9/io_i_5_in1[5]
+ cb_5_9/io_i_5_in1[6] cb_5_9/io_i_5_in1[7] cb_5_9/io_i_6_ci cb_5_9/io_i_6_in1[0]
+ cb_5_9/io_i_6_in1[1] cb_5_9/io_i_6_in1[2] cb_5_9/io_i_6_in1[3] cb_5_9/io_i_6_in1[4]
+ cb_5_9/io_i_6_in1[5] cb_5_9/io_i_6_in1[6] cb_5_9/io_i_6_in1[7] cb_5_9/io_i_7_ci
+ cb_5_9/io_i_7_in1[0] cb_5_9/io_i_7_in1[1] cb_5_9/io_i_7_in1[2] cb_5_9/io_i_7_in1[3]
+ cb_5_9/io_i_7_in1[4] cb_5_9/io_i_7_in1[5] cb_5_9/io_i_7_in1[6] cb_5_9/io_i_7_in1[7]
+ cb_5_8/io_vci cb_5_9/io_vci cb_5_8/io_vi cb_5_9/io_we_i cb_5_8/io_wo[0] cb_5_8/io_wo[10]
+ cb_5_8/io_wo[11] cb_5_8/io_wo[12] cb_5_8/io_wo[13] cb_5_8/io_wo[14] cb_5_8/io_wo[15]
+ cb_5_8/io_wo[16] cb_5_8/io_wo[17] cb_5_8/io_wo[18] cb_5_8/io_wo[19] cb_5_8/io_wo[1]
+ cb_5_8/io_wo[20] cb_5_8/io_wo[21] cb_5_8/io_wo[22] cb_5_8/io_wo[23] cb_5_8/io_wo[24]
+ cb_5_8/io_wo[25] cb_5_8/io_wo[26] cb_5_8/io_wo[27] cb_5_8/io_wo[28] cb_5_8/io_wo[29]
+ cb_5_8/io_wo[2] cb_5_8/io_wo[30] cb_5_8/io_wo[31] cb_5_8/io_wo[32] cb_5_8/io_wo[33]
+ cb_5_8/io_wo[34] cb_5_8/io_wo[35] cb_5_8/io_wo[36] cb_5_8/io_wo[37] cb_5_8/io_wo[38]
+ cb_5_8/io_wo[39] cb_5_8/io_wo[3] cb_5_8/io_wo[40] cb_5_8/io_wo[41] cb_5_8/io_wo[42]
+ cb_5_8/io_wo[43] cb_5_8/io_wo[44] cb_5_8/io_wo[45] cb_5_8/io_wo[46] cb_5_8/io_wo[47]
+ cb_5_8/io_wo[48] cb_5_8/io_wo[49] cb_5_8/io_wo[4] cb_5_8/io_wo[50] cb_5_8/io_wo[51]
+ cb_5_8/io_wo[52] cb_5_8/io_wo[53] cb_5_8/io_wo[54] cb_5_8/io_wo[55] cb_5_8/io_wo[56]
+ cb_5_8/io_wo[57] cb_5_8/io_wo[58] cb_5_8/io_wo[59] cb_5_8/io_wo[5] cb_5_8/io_wo[60]
+ cb_5_8/io_wo[61] cb_5_8/io_wo[62] cb_5_8/io_wo[63] cb_5_8/io_wo[6] cb_5_8/io_wo[7]
+ cb_5_8/io_wo[8] cb_5_8/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_3_5 cb_3_9/io_adr_i[0] cb_3_9/io_adr_i[1] cb_3_5/io_cs_i cb_3_9/io_dat_i[0] cb_3_9/io_dat_i[10]
+ cb_3_9/io_dat_i[11] cb_3_9/io_dat_i[12] cb_3_9/io_dat_i[13] cb_3_9/io_dat_i[14]
+ cb_3_9/io_dat_i[15] cb_3_9/io_dat_i[1] cb_3_9/io_dat_i[2] cb_3_9/io_dat_i[3] cb_3_9/io_dat_i[4]
+ cb_3_9/io_dat_i[5] cb_3_9/io_dat_i[6] cb_3_9/io_dat_i[7] cb_3_9/io_dat_i[8] cb_3_9/io_dat_i[9]
+ cb_3_5/io_dat_o[0] cb_3_5/io_dat_o[10] cb_3_5/io_dat_o[11] cb_3_5/io_dat_o[12] cb_3_5/io_dat_o[13]
+ cb_3_5/io_dat_o[14] cb_3_5/io_dat_o[15] cb_3_5/io_dat_o[1] cb_3_5/io_dat_o[2] cb_3_5/io_dat_o[3]
+ cb_3_5/io_dat_o[4] cb_3_5/io_dat_o[5] cb_3_5/io_dat_o[6] cb_3_5/io_dat_o[7] cb_3_5/io_dat_o[8]
+ cb_3_5/io_dat_o[9] cb_3_6/io_wo[0] cb_3_6/io_wo[10] cb_3_6/io_wo[11] cb_3_6/io_wo[12]
+ cb_3_6/io_wo[13] cb_3_6/io_wo[14] cb_3_6/io_wo[15] cb_3_6/io_wo[16] cb_3_6/io_wo[17]
+ cb_3_6/io_wo[18] cb_3_6/io_wo[19] cb_3_6/io_wo[1] cb_3_6/io_wo[20] cb_3_6/io_wo[21]
+ cb_3_6/io_wo[22] cb_3_6/io_wo[23] cb_3_6/io_wo[24] cb_3_6/io_wo[25] cb_3_6/io_wo[26]
+ cb_3_6/io_wo[27] cb_3_6/io_wo[28] cb_3_6/io_wo[29] cb_3_6/io_wo[2] cb_3_6/io_wo[30]
+ cb_3_6/io_wo[31] cb_3_6/io_wo[32] cb_3_6/io_wo[33] cb_3_6/io_wo[34] cb_3_6/io_wo[35]
+ cb_3_6/io_wo[36] cb_3_6/io_wo[37] cb_3_6/io_wo[38] cb_3_6/io_wo[39] cb_3_6/io_wo[3]
+ cb_3_6/io_wo[40] cb_3_6/io_wo[41] cb_3_6/io_wo[42] cb_3_6/io_wo[43] cb_3_6/io_wo[44]
+ cb_3_6/io_wo[45] cb_3_6/io_wo[46] cb_3_6/io_wo[47] cb_3_6/io_wo[48] cb_3_6/io_wo[49]
+ cb_3_6/io_wo[4] cb_3_6/io_wo[50] cb_3_6/io_wo[51] cb_3_6/io_wo[52] cb_3_6/io_wo[53]
+ cb_3_6/io_wo[54] cb_3_6/io_wo[55] cb_3_6/io_wo[56] cb_3_6/io_wo[57] cb_3_6/io_wo[58]
+ cb_3_6/io_wo[59] cb_3_6/io_wo[5] cb_3_6/io_wo[60] cb_3_6/io_wo[61] cb_3_6/io_wo[62]
+ cb_3_6/io_wo[63] cb_3_6/io_wo[6] cb_3_6/io_wo[7] cb_3_6/io_wo[8] cb_3_6/io_wo[9]
+ cb_3_5/io_i_0_ci cb_3_5/io_i_0_in1[0] cb_3_5/io_i_0_in1[1] cb_3_5/io_i_0_in1[2]
+ cb_3_5/io_i_0_in1[3] cb_3_5/io_i_0_in1[4] cb_3_5/io_i_0_in1[5] cb_3_5/io_i_0_in1[6]
+ cb_3_5/io_i_0_in1[7] cb_3_5/io_i_1_ci cb_3_5/io_i_1_in1[0] cb_3_5/io_i_1_in1[1]
+ cb_3_5/io_i_1_in1[2] cb_3_5/io_i_1_in1[3] cb_3_5/io_i_1_in1[4] cb_3_5/io_i_1_in1[5]
+ cb_3_5/io_i_1_in1[6] cb_3_5/io_i_1_in1[7] cb_3_5/io_i_2_ci cb_3_5/io_i_2_in1[0]
+ cb_3_5/io_i_2_in1[1] cb_3_5/io_i_2_in1[2] cb_3_5/io_i_2_in1[3] cb_3_5/io_i_2_in1[4]
+ cb_3_5/io_i_2_in1[5] cb_3_5/io_i_2_in1[6] cb_3_5/io_i_2_in1[7] cb_3_5/io_i_3_ci
+ cb_3_5/io_i_3_in1[0] cb_3_5/io_i_3_in1[1] cb_3_5/io_i_3_in1[2] cb_3_5/io_i_3_in1[3]
+ cb_3_5/io_i_3_in1[4] cb_3_5/io_i_3_in1[5] cb_3_5/io_i_3_in1[6] cb_3_5/io_i_3_in1[7]
+ cb_3_5/io_i_4_ci cb_3_5/io_i_4_in1[0] cb_3_5/io_i_4_in1[1] cb_3_5/io_i_4_in1[2]
+ cb_3_5/io_i_4_in1[3] cb_3_5/io_i_4_in1[4] cb_3_5/io_i_4_in1[5] cb_3_5/io_i_4_in1[6]
+ cb_3_5/io_i_4_in1[7] cb_3_5/io_i_5_ci cb_3_5/io_i_5_in1[0] cb_3_5/io_i_5_in1[1]
+ cb_3_5/io_i_5_in1[2] cb_3_5/io_i_5_in1[3] cb_3_5/io_i_5_in1[4] cb_3_5/io_i_5_in1[5]
+ cb_3_5/io_i_5_in1[6] cb_3_5/io_i_5_in1[7] cb_3_5/io_i_6_ci cb_3_5/io_i_6_in1[0]
+ cb_3_5/io_i_6_in1[1] cb_3_5/io_i_6_in1[2] cb_3_5/io_i_6_in1[3] cb_3_5/io_i_6_in1[4]
+ cb_3_5/io_i_6_in1[5] cb_3_5/io_i_6_in1[6] cb_3_5/io_i_6_in1[7] cb_3_5/io_i_7_ci
+ cb_3_5/io_i_7_in1[0] cb_3_5/io_i_7_in1[1] cb_3_5/io_i_7_in1[2] cb_3_5/io_i_7_in1[3]
+ cb_3_5/io_i_7_in1[4] cb_3_5/io_i_7_in1[5] cb_3_5/io_i_7_in1[6] cb_3_5/io_i_7_in1[7]
+ cb_3_6/io_i_0_ci cb_3_6/io_i_0_in1[0] cb_3_6/io_i_0_in1[1] cb_3_6/io_i_0_in1[2]
+ cb_3_6/io_i_0_in1[3] cb_3_6/io_i_0_in1[4] cb_3_6/io_i_0_in1[5] cb_3_6/io_i_0_in1[6]
+ cb_3_6/io_i_0_in1[7] cb_3_6/io_i_1_ci cb_3_6/io_i_1_in1[0] cb_3_6/io_i_1_in1[1]
+ cb_3_6/io_i_1_in1[2] cb_3_6/io_i_1_in1[3] cb_3_6/io_i_1_in1[4] cb_3_6/io_i_1_in1[5]
+ cb_3_6/io_i_1_in1[6] cb_3_6/io_i_1_in1[7] cb_3_6/io_i_2_ci cb_3_6/io_i_2_in1[0]
+ cb_3_6/io_i_2_in1[1] cb_3_6/io_i_2_in1[2] cb_3_6/io_i_2_in1[3] cb_3_6/io_i_2_in1[4]
+ cb_3_6/io_i_2_in1[5] cb_3_6/io_i_2_in1[6] cb_3_6/io_i_2_in1[7] cb_3_6/io_i_3_ci
+ cb_3_6/io_i_3_in1[0] cb_3_6/io_i_3_in1[1] cb_3_6/io_i_3_in1[2] cb_3_6/io_i_3_in1[3]
+ cb_3_6/io_i_3_in1[4] cb_3_6/io_i_3_in1[5] cb_3_6/io_i_3_in1[6] cb_3_6/io_i_3_in1[7]
+ cb_3_6/io_i_4_ci cb_3_6/io_i_4_in1[0] cb_3_6/io_i_4_in1[1] cb_3_6/io_i_4_in1[2]
+ cb_3_6/io_i_4_in1[3] cb_3_6/io_i_4_in1[4] cb_3_6/io_i_4_in1[5] cb_3_6/io_i_4_in1[6]
+ cb_3_6/io_i_4_in1[7] cb_3_6/io_i_5_ci cb_3_6/io_i_5_in1[0] cb_3_6/io_i_5_in1[1]
+ cb_3_6/io_i_5_in1[2] cb_3_6/io_i_5_in1[3] cb_3_6/io_i_5_in1[4] cb_3_6/io_i_5_in1[5]
+ cb_3_6/io_i_5_in1[6] cb_3_6/io_i_5_in1[7] cb_3_6/io_i_6_ci cb_3_6/io_i_6_in1[0]
+ cb_3_6/io_i_6_in1[1] cb_3_6/io_i_6_in1[2] cb_3_6/io_i_6_in1[3] cb_3_6/io_i_6_in1[4]
+ cb_3_6/io_i_6_in1[5] cb_3_6/io_i_6_in1[6] cb_3_6/io_i_6_in1[7] cb_3_6/io_i_7_ci
+ cb_3_6/io_i_7_in1[0] cb_3_6/io_i_7_in1[1] cb_3_6/io_i_7_in1[2] cb_3_6/io_i_7_in1[3]
+ cb_3_6/io_i_7_in1[4] cb_3_6/io_i_7_in1[5] cb_3_6/io_i_7_in1[6] cb_3_6/io_i_7_in1[7]
+ cb_3_5/io_vci cb_3_6/io_vci cb_3_5/io_vi cb_3_9/io_we_i cb_3_5/io_wo[0] cb_3_5/io_wo[10]
+ cb_3_5/io_wo[11] cb_3_5/io_wo[12] cb_3_5/io_wo[13] cb_3_5/io_wo[14] cb_3_5/io_wo[15]
+ cb_3_5/io_wo[16] cb_3_5/io_wo[17] cb_3_5/io_wo[18] cb_3_5/io_wo[19] cb_3_5/io_wo[1]
+ cb_3_5/io_wo[20] cb_3_5/io_wo[21] cb_3_5/io_wo[22] cb_3_5/io_wo[23] cb_3_5/io_wo[24]
+ cb_3_5/io_wo[25] cb_3_5/io_wo[26] cb_3_5/io_wo[27] cb_3_5/io_wo[28] cb_3_5/io_wo[29]
+ cb_3_5/io_wo[2] cb_3_5/io_wo[30] cb_3_5/io_wo[31] cb_3_5/io_wo[32] cb_3_5/io_wo[33]
+ cb_3_5/io_wo[34] cb_3_5/io_wo[35] cb_3_5/io_wo[36] cb_3_5/io_wo[37] cb_3_5/io_wo[38]
+ cb_3_5/io_wo[39] cb_3_5/io_wo[3] cb_3_5/io_wo[40] cb_3_5/io_wo[41] cb_3_5/io_wo[42]
+ cb_3_5/io_wo[43] cb_3_5/io_wo[44] cb_3_5/io_wo[45] cb_3_5/io_wo[46] cb_3_5/io_wo[47]
+ cb_3_5/io_wo[48] cb_3_5/io_wo[49] cb_3_5/io_wo[4] cb_3_5/io_wo[50] cb_3_5/io_wo[51]
+ cb_3_5/io_wo[52] cb_3_5/io_wo[53] cb_3_5/io_wo[54] cb_3_5/io_wo[55] cb_3_5/io_wo[56]
+ cb_3_5/io_wo[57] cb_3_5/io_wo[58] cb_3_5/io_wo[59] cb_3_5/io_wo[5] cb_3_5/io_wo[60]
+ cb_3_5/io_wo[61] cb_3_5/io_wo[62] cb_3_5/io_wo[63] cb_3_5/io_wo[6] cb_3_5/io_wo[7]
+ cb_3_5/io_wo[8] cb_3_5/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_1_2 cb_1_9/io_adr_i[0] cb_1_9/io_adr_i[1] cb_1_2/io_cs_i cb_1_9/io_dat_i[0] cb_1_9/io_dat_i[10]
+ cb_1_9/io_dat_i[11] cb_1_9/io_dat_i[12] cb_1_9/io_dat_i[13] cb_1_9/io_dat_i[14]
+ cb_1_9/io_dat_i[15] cb_1_9/io_dat_i[1] cb_1_9/io_dat_i[2] cb_1_9/io_dat_i[3] cb_1_9/io_dat_i[4]
+ cb_1_9/io_dat_i[5] cb_1_9/io_dat_i[6] cb_1_9/io_dat_i[7] cb_1_9/io_dat_i[8] cb_1_9/io_dat_i[9]
+ cb_1_2/io_dat_o[0] cb_1_2/io_dat_o[10] cb_1_2/io_dat_o[11] cb_1_2/io_dat_o[12] cb_1_2/io_dat_o[13]
+ cb_1_2/io_dat_o[14] cb_1_2/io_dat_o[15] cb_1_2/io_dat_o[1] cb_1_2/io_dat_o[2] cb_1_2/io_dat_o[3]
+ cb_1_2/io_dat_o[4] cb_1_2/io_dat_o[5] cb_1_2/io_dat_o[6] cb_1_2/io_dat_o[7] cb_1_2/io_dat_o[8]
+ cb_1_2/io_dat_o[9] cb_1_3/io_wo[0] cb_1_3/io_wo[10] cb_1_3/io_wo[11] cb_1_3/io_wo[12]
+ cb_1_3/io_wo[13] cb_1_3/io_wo[14] cb_1_3/io_wo[15] cb_1_3/io_wo[16] cb_1_3/io_wo[17]
+ cb_1_3/io_wo[18] cb_1_3/io_wo[19] cb_1_3/io_wo[1] cb_1_3/io_wo[20] cb_1_3/io_wo[21]
+ cb_1_3/io_wo[22] cb_1_3/io_wo[23] cb_1_3/io_wo[24] cb_1_3/io_wo[25] cb_1_3/io_wo[26]
+ cb_1_3/io_wo[27] cb_1_3/io_wo[28] cb_1_3/io_wo[29] cb_1_3/io_wo[2] cb_1_3/io_wo[30]
+ cb_1_3/io_wo[31] cb_1_3/io_wo[32] cb_1_3/io_wo[33] cb_1_3/io_wo[34] cb_1_3/io_wo[35]
+ cb_1_3/io_wo[36] cb_1_3/io_wo[37] cb_1_3/io_wo[38] cb_1_3/io_wo[39] cb_1_3/io_wo[3]
+ cb_1_3/io_wo[40] cb_1_3/io_wo[41] cb_1_3/io_wo[42] cb_1_3/io_wo[43] cb_1_3/io_wo[44]
+ cb_1_3/io_wo[45] cb_1_3/io_wo[46] cb_1_3/io_wo[47] cb_1_3/io_wo[48] cb_1_3/io_wo[49]
+ cb_1_3/io_wo[4] cb_1_3/io_wo[50] cb_1_3/io_wo[51] cb_1_3/io_wo[52] cb_1_3/io_wo[53]
+ cb_1_3/io_wo[54] cb_1_3/io_wo[55] cb_1_3/io_wo[56] cb_1_3/io_wo[57] cb_1_3/io_wo[58]
+ cb_1_3/io_wo[59] cb_1_3/io_wo[5] cb_1_3/io_wo[60] cb_1_3/io_wo[61] cb_1_3/io_wo[62]
+ cb_1_3/io_wo[63] cb_1_3/io_wo[6] cb_1_3/io_wo[7] cb_1_3/io_wo[8] cb_1_3/io_wo[9]
+ cb_1_2/io_i_0_ci cb_1_2/io_i_0_in1[0] cb_1_2/io_i_0_in1[1] cb_1_2/io_i_0_in1[2]
+ cb_1_2/io_i_0_in1[3] cb_1_2/io_i_0_in1[4] cb_1_2/io_i_0_in1[5] cb_1_2/io_i_0_in1[6]
+ cb_1_2/io_i_0_in1[7] cb_1_2/io_i_1_ci cb_1_2/io_i_1_in1[0] cb_1_2/io_i_1_in1[1]
+ cb_1_2/io_i_1_in1[2] cb_1_2/io_i_1_in1[3] cb_1_2/io_i_1_in1[4] cb_1_2/io_i_1_in1[5]
+ cb_1_2/io_i_1_in1[6] cb_1_2/io_i_1_in1[7] cb_1_2/io_i_2_ci cb_1_2/io_i_2_in1[0]
+ cb_1_2/io_i_2_in1[1] cb_1_2/io_i_2_in1[2] cb_1_2/io_i_2_in1[3] cb_1_2/io_i_2_in1[4]
+ cb_1_2/io_i_2_in1[5] cb_1_2/io_i_2_in1[6] cb_1_2/io_i_2_in1[7] cb_1_2/io_i_3_ci
+ cb_1_2/io_i_3_in1[0] cb_1_2/io_i_3_in1[1] cb_1_2/io_i_3_in1[2] cb_1_2/io_i_3_in1[3]
+ cb_1_2/io_i_3_in1[4] cb_1_2/io_i_3_in1[5] cb_1_2/io_i_3_in1[6] cb_1_2/io_i_3_in1[7]
+ cb_1_2/io_i_4_ci cb_1_2/io_i_4_in1[0] cb_1_2/io_i_4_in1[1] cb_1_2/io_i_4_in1[2]
+ cb_1_2/io_i_4_in1[3] cb_1_2/io_i_4_in1[4] cb_1_2/io_i_4_in1[5] cb_1_2/io_i_4_in1[6]
+ cb_1_2/io_i_4_in1[7] cb_1_2/io_i_5_ci cb_1_2/io_i_5_in1[0] cb_1_2/io_i_5_in1[1]
+ cb_1_2/io_i_5_in1[2] cb_1_2/io_i_5_in1[3] cb_1_2/io_i_5_in1[4] cb_1_2/io_i_5_in1[5]
+ cb_1_2/io_i_5_in1[6] cb_1_2/io_i_5_in1[7] cb_1_2/io_i_6_ci cb_1_2/io_i_6_in1[0]
+ cb_1_2/io_i_6_in1[1] cb_1_2/io_i_6_in1[2] cb_1_2/io_i_6_in1[3] cb_1_2/io_i_6_in1[4]
+ cb_1_2/io_i_6_in1[5] cb_1_2/io_i_6_in1[6] cb_1_2/io_i_6_in1[7] cb_1_2/io_i_7_ci
+ cb_1_2/io_i_7_in1[0] cb_1_2/io_i_7_in1[1] cb_1_2/io_i_7_in1[2] cb_1_2/io_i_7_in1[3]
+ cb_1_2/io_i_7_in1[4] cb_1_2/io_i_7_in1[5] cb_1_2/io_i_7_in1[6] cb_1_2/io_i_7_in1[7]
+ cb_1_3/io_i_0_ci cb_1_3/io_i_0_in1[0] cb_1_3/io_i_0_in1[1] cb_1_3/io_i_0_in1[2]
+ cb_1_3/io_i_0_in1[3] cb_1_3/io_i_0_in1[4] cb_1_3/io_i_0_in1[5] cb_1_3/io_i_0_in1[6]
+ cb_1_3/io_i_0_in1[7] cb_1_3/io_i_1_ci cb_1_3/io_i_1_in1[0] cb_1_3/io_i_1_in1[1]
+ cb_1_3/io_i_1_in1[2] cb_1_3/io_i_1_in1[3] cb_1_3/io_i_1_in1[4] cb_1_3/io_i_1_in1[5]
+ cb_1_3/io_i_1_in1[6] cb_1_3/io_i_1_in1[7] cb_1_3/io_i_2_ci cb_1_3/io_i_2_in1[0]
+ cb_1_3/io_i_2_in1[1] cb_1_3/io_i_2_in1[2] cb_1_3/io_i_2_in1[3] cb_1_3/io_i_2_in1[4]
+ cb_1_3/io_i_2_in1[5] cb_1_3/io_i_2_in1[6] cb_1_3/io_i_2_in1[7] cb_1_3/io_i_3_ci
+ cb_1_3/io_i_3_in1[0] cb_1_3/io_i_3_in1[1] cb_1_3/io_i_3_in1[2] cb_1_3/io_i_3_in1[3]
+ cb_1_3/io_i_3_in1[4] cb_1_3/io_i_3_in1[5] cb_1_3/io_i_3_in1[6] cb_1_3/io_i_3_in1[7]
+ cb_1_3/io_i_4_ci cb_1_3/io_i_4_in1[0] cb_1_3/io_i_4_in1[1] cb_1_3/io_i_4_in1[2]
+ cb_1_3/io_i_4_in1[3] cb_1_3/io_i_4_in1[4] cb_1_3/io_i_4_in1[5] cb_1_3/io_i_4_in1[6]
+ cb_1_3/io_i_4_in1[7] cb_1_3/io_i_5_ci cb_1_3/io_i_5_in1[0] cb_1_3/io_i_5_in1[1]
+ cb_1_3/io_i_5_in1[2] cb_1_3/io_i_5_in1[3] cb_1_3/io_i_5_in1[4] cb_1_3/io_i_5_in1[5]
+ cb_1_3/io_i_5_in1[6] cb_1_3/io_i_5_in1[7] cb_1_3/io_i_6_ci cb_1_3/io_i_6_in1[0]
+ cb_1_3/io_i_6_in1[1] cb_1_3/io_i_6_in1[2] cb_1_3/io_i_6_in1[3] cb_1_3/io_i_6_in1[4]
+ cb_1_3/io_i_6_in1[5] cb_1_3/io_i_6_in1[6] cb_1_3/io_i_6_in1[7] cb_1_3/io_i_7_ci
+ cb_1_3/io_i_7_in1[0] cb_1_3/io_i_7_in1[1] cb_1_3/io_i_7_in1[2] cb_1_3/io_i_7_in1[3]
+ cb_1_3/io_i_7_in1[4] cb_1_3/io_i_7_in1[5] cb_1_3/io_i_7_in1[6] cb_1_3/io_i_7_in1[7]
+ cb_1_2/io_vci cb_1_3/io_vci cb_1_2/io_vi cb_1_9/io_we_i cb_1_2/io_wo[0] cb_1_2/io_wo[10]
+ cb_1_2/io_wo[11] cb_1_2/io_wo[12] cb_1_2/io_wo[13] cb_1_2/io_wo[14] cb_1_2/io_wo[15]
+ cb_1_2/io_wo[16] cb_1_2/io_wo[17] cb_1_2/io_wo[18] cb_1_2/io_wo[19] cb_1_2/io_wo[1]
+ cb_1_2/io_wo[20] cb_1_2/io_wo[21] cb_1_2/io_wo[22] cb_1_2/io_wo[23] cb_1_2/io_wo[24]
+ cb_1_2/io_wo[25] cb_1_2/io_wo[26] cb_1_2/io_wo[27] cb_1_2/io_wo[28] cb_1_2/io_wo[29]
+ cb_1_2/io_wo[2] cb_1_2/io_wo[30] cb_1_2/io_wo[31] cb_1_2/io_wo[32] cb_1_2/io_wo[33]
+ cb_1_2/io_wo[34] cb_1_2/io_wo[35] cb_1_2/io_wo[36] cb_1_2/io_wo[37] cb_1_2/io_wo[38]
+ cb_1_2/io_wo[39] cb_1_2/io_wo[3] cb_1_2/io_wo[40] cb_1_2/io_wo[41] cb_1_2/io_wo[42]
+ cb_1_2/io_wo[43] cb_1_2/io_wo[44] cb_1_2/io_wo[45] cb_1_2/io_wo[46] cb_1_2/io_wo[47]
+ cb_1_2/io_wo[48] cb_1_2/io_wo[49] cb_1_2/io_wo[4] cb_1_2/io_wo[50] cb_1_2/io_wo[51]
+ cb_1_2/io_wo[52] cb_1_2/io_wo[53] cb_1_2/io_wo[54] cb_1_2/io_wo[55] cb_1_2/io_wo[56]
+ cb_1_2/io_wo[57] cb_1_2/io_wo[58] cb_1_2/io_wo[59] cb_1_2/io_wo[5] cb_1_2/io_wo[60]
+ cb_1_2/io_wo[61] cb_1_2/io_wo[62] cb_1_2/io_wo[63] cb_1_2/io_wo[6] cb_1_2/io_wo[7]
+ cb_1_2/io_wo[8] cb_1_2/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xccon_5 ccon_5/io_ack_o ccon_7/io_adr_i[0] ccon_7/io_adr_i[10] ccon_7/io_adr_i[11]
+ ccon_7/io_adr_i[1] ccon_7/io_adr_i[2] ccon_7/io_adr_i[3] ccon_7/io_adr_i[4] ccon_7/io_adr_i[5]
+ ccon_7/io_adr_i[6] ccon_7/io_adr_i[7] ccon_7/io_adr_i[8] ccon_7/io_adr_i[9] cb_5_9/io_adr_i[0]
+ cb_5_9/io_adr_i[1] cb_5_0/io_cs_i cb_5_1/io_cs_i cb_5_10/io_cs_i cb_5_2/io_cs_i
+ cb_5_3/io_cs_i cb_5_4/io_cs_i cb_5_5/io_cs_i cb_5_6/io_cs_i cb_5_7/io_cs_i cb_5_8/io_cs_i
+ cb_5_9/io_cs_i cb_5_9/io_dat_i[0] cb_5_9/io_dat_i[10] cb_5_9/io_dat_i[11] cb_5_9/io_dat_i[12]
+ cb_5_9/io_dat_i[13] cb_5_9/io_dat_i[14] cb_5_9/io_dat_i[15] cb_5_9/io_dat_i[1] cb_5_9/io_dat_i[2]
+ cb_5_9/io_dat_i[3] cb_5_9/io_dat_i[4] cb_5_9/io_dat_i[5] cb_5_9/io_dat_i[6] cb_5_9/io_dat_i[7]
+ cb_5_9/io_dat_i[8] cb_5_9/io_dat_i[9] cb_5_0/io_dat_o[0] cb_5_0/io_dat_o[10] cb_5_0/io_dat_o[11]
+ cb_5_0/io_dat_o[12] cb_5_0/io_dat_o[13] cb_5_0/io_dat_o[14] cb_5_0/io_dat_o[15]
+ cb_5_0/io_dat_o[1] cb_5_0/io_dat_o[2] cb_5_0/io_dat_o[3] cb_5_0/io_dat_o[4] cb_5_0/io_dat_o[5]
+ cb_5_0/io_dat_o[6] cb_5_0/io_dat_o[7] cb_5_0/io_dat_o[8] cb_5_0/io_dat_o[9] cb_5_10/io_dat_o[0]
+ cb_5_10/io_dat_o[10] cb_5_10/io_dat_o[11] cb_5_10/io_dat_o[12] cb_5_10/io_dat_o[13]
+ cb_5_10/io_dat_o[14] cb_5_10/io_dat_o[15] cb_5_10/io_dat_o[1] cb_5_10/io_dat_o[2]
+ cb_5_10/io_dat_o[3] cb_5_10/io_dat_o[4] cb_5_10/io_dat_o[5] cb_5_10/io_dat_o[6]
+ cb_5_10/io_dat_o[7] cb_5_10/io_dat_o[8] cb_5_10/io_dat_o[9] cb_5_1/io_dat_o[0] cb_5_1/io_dat_o[10]
+ cb_5_1/io_dat_o[11] cb_5_1/io_dat_o[12] cb_5_1/io_dat_o[13] cb_5_1/io_dat_o[14]
+ cb_5_1/io_dat_o[15] cb_5_1/io_dat_o[1] cb_5_1/io_dat_o[2] cb_5_1/io_dat_o[3] cb_5_1/io_dat_o[4]
+ cb_5_1/io_dat_o[5] cb_5_1/io_dat_o[6] cb_5_1/io_dat_o[7] cb_5_1/io_dat_o[8] cb_5_1/io_dat_o[9]
+ cb_5_2/io_dat_o[0] cb_5_2/io_dat_o[10] cb_5_2/io_dat_o[11] cb_5_2/io_dat_o[12] cb_5_2/io_dat_o[13]
+ cb_5_2/io_dat_o[14] cb_5_2/io_dat_o[15] cb_5_2/io_dat_o[1] cb_5_2/io_dat_o[2] cb_5_2/io_dat_o[3]
+ cb_5_2/io_dat_o[4] cb_5_2/io_dat_o[5] cb_5_2/io_dat_o[6] cb_5_2/io_dat_o[7] cb_5_2/io_dat_o[8]
+ cb_5_2/io_dat_o[9] cb_5_3/io_dat_o[0] cb_5_3/io_dat_o[10] cb_5_3/io_dat_o[11] cb_5_3/io_dat_o[12]
+ cb_5_3/io_dat_o[13] cb_5_3/io_dat_o[14] cb_5_3/io_dat_o[15] cb_5_3/io_dat_o[1] cb_5_3/io_dat_o[2]
+ cb_5_3/io_dat_o[3] cb_5_3/io_dat_o[4] cb_5_3/io_dat_o[5] cb_5_3/io_dat_o[6] cb_5_3/io_dat_o[7]
+ cb_5_3/io_dat_o[8] cb_5_3/io_dat_o[9] cb_5_4/io_dat_o[0] cb_5_4/io_dat_o[10] cb_5_4/io_dat_o[11]
+ cb_5_4/io_dat_o[12] cb_5_4/io_dat_o[13] cb_5_4/io_dat_o[14] cb_5_4/io_dat_o[15]
+ cb_5_4/io_dat_o[1] cb_5_4/io_dat_o[2] cb_5_4/io_dat_o[3] cb_5_4/io_dat_o[4] cb_5_4/io_dat_o[5]
+ cb_5_4/io_dat_o[6] cb_5_4/io_dat_o[7] cb_5_4/io_dat_o[8] cb_5_4/io_dat_o[9] cb_5_5/io_dat_o[0]
+ cb_5_5/io_dat_o[10] cb_5_5/io_dat_o[11] cb_5_5/io_dat_o[12] cb_5_5/io_dat_o[13]
+ cb_5_5/io_dat_o[14] cb_5_5/io_dat_o[15] cb_5_5/io_dat_o[1] cb_5_5/io_dat_o[2] cb_5_5/io_dat_o[3]
+ cb_5_5/io_dat_o[4] cb_5_5/io_dat_o[5] cb_5_5/io_dat_o[6] cb_5_5/io_dat_o[7] cb_5_5/io_dat_o[8]
+ cb_5_5/io_dat_o[9] cb_5_6/io_dat_o[0] cb_5_6/io_dat_o[10] cb_5_6/io_dat_o[11] cb_5_6/io_dat_o[12]
+ cb_5_6/io_dat_o[13] cb_5_6/io_dat_o[14] cb_5_6/io_dat_o[15] cb_5_6/io_dat_o[1] cb_5_6/io_dat_o[2]
+ cb_5_6/io_dat_o[3] cb_5_6/io_dat_o[4] cb_5_6/io_dat_o[5] cb_5_6/io_dat_o[6] cb_5_6/io_dat_o[7]
+ cb_5_6/io_dat_o[8] cb_5_6/io_dat_o[9] cb_5_7/io_dat_o[0] cb_5_7/io_dat_o[10] cb_5_7/io_dat_o[11]
+ cb_5_7/io_dat_o[12] cb_5_7/io_dat_o[13] cb_5_7/io_dat_o[14] cb_5_7/io_dat_o[15]
+ cb_5_7/io_dat_o[1] cb_5_7/io_dat_o[2] cb_5_7/io_dat_o[3] cb_5_7/io_dat_o[4] cb_5_7/io_dat_o[5]
+ cb_5_7/io_dat_o[6] cb_5_7/io_dat_o[7] cb_5_7/io_dat_o[8] cb_5_7/io_dat_o[9] cb_5_8/io_dat_o[0]
+ cb_5_8/io_dat_o[10] cb_5_8/io_dat_o[11] cb_5_8/io_dat_o[12] cb_5_8/io_dat_o[13]
+ cb_5_8/io_dat_o[14] cb_5_8/io_dat_o[15] cb_5_8/io_dat_o[1] cb_5_8/io_dat_o[2] cb_5_8/io_dat_o[3]
+ cb_5_8/io_dat_o[4] cb_5_8/io_dat_o[5] cb_5_8/io_dat_o[6] cb_5_8/io_dat_o[7] cb_5_8/io_dat_o[8]
+ cb_5_8/io_dat_o[9] cb_5_9/io_dat_o[0] cb_5_9/io_dat_o[10] cb_5_9/io_dat_o[11] cb_5_9/io_dat_o[12]
+ cb_5_9/io_dat_o[13] cb_5_9/io_dat_o[14] cb_5_9/io_dat_o[15] cb_5_9/io_dat_o[1] cb_5_9/io_dat_o[2]
+ cb_5_9/io_dat_o[3] cb_5_9/io_dat_o[4] cb_5_9/io_dat_o[5] cb_5_9/io_dat_o[6] cb_5_9/io_dat_o[7]
+ cb_5_9/io_dat_o[8] cb_5_9/io_dat_o[9] cb_5_9/io_we_i ccon_5/io_cs_i ccon_7/io_dat_i[0]
+ ccon_7/io_dat_i[10] ccon_7/io_dat_i[11] ccon_7/io_dat_i[12] ccon_7/io_dat_i[13]
+ ccon_7/io_dat_i[14] ccon_7/io_dat_i[15] ccon_7/io_dat_i[16] ccon_7/io_dat_i[17]
+ ccon_7/io_dat_i[18] ccon_7/io_dat_i[19] ccon_7/io_dat_i[1] ccon_7/io_dat_i[20] ccon_7/io_dat_i[21]
+ ccon_7/io_dat_i[22] ccon_7/io_dat_i[23] ccon_7/io_dat_i[24] ccon_7/io_dat_i[25]
+ ccon_7/io_dat_i[26] ccon_7/io_dat_i[27] ccon_7/io_dat_i[28] ccon_7/io_dat_i[29]
+ ccon_7/io_dat_i[2] ccon_7/io_dat_i[30] ccon_7/io_dat_i[31] ccon_7/io_dat_i[3] ccon_7/io_dat_i[4]
+ ccon_7/io_dat_i[5] ccon_7/io_dat_i[6] ccon_7/io_dat_i[7] ccon_7/io_dat_i[8] ccon_7/io_dat_i[9]
+ ccon_5/io_dat_o[0] ccon_5/io_dat_o[10] ccon_5/io_dat_o[11] ccon_5/io_dat_o[12] ccon_5/io_dat_o[13]
+ ccon_5/io_dat_o[14] ccon_5/io_dat_o[15] ccon_5/io_dat_o[16] ccon_5/io_dat_o[17]
+ ccon_5/io_dat_o[18] ccon_5/io_dat_o[19] ccon_5/io_dat_o[1] ccon_5/io_dat_o[20] ccon_5/io_dat_o[21]
+ ccon_5/io_dat_o[22] ccon_5/io_dat_o[23] ccon_5/io_dat_o[24] ccon_5/io_dat_o[25]
+ ccon_5/io_dat_o[26] ccon_5/io_dat_o[27] ccon_5/io_dat_o[28] ccon_5/io_dat_o[29]
+ ccon_5/io_dat_o[2] ccon_5/io_dat_o[30] ccon_5/io_dat_o[31] ccon_5/io_dat_o[3] ccon_5/io_dat_o[4]
+ ccon_5/io_dat_o[5] ccon_5/io_dat_o[6] ccon_5/io_dat_o[7] ccon_5/io_dat_o[8] ccon_5/io_dat_o[9]
+ cb_5_0/io_wo[0] cb_5_0/io_wo[10] cb_5_0/io_wo[11] cb_5_0/io_wo[12] cb_5_0/io_wo[13]
+ cb_5_0/io_wo[14] cb_5_0/io_wo[15] cb_5_0/io_wo[16] cb_5_0/io_wo[17] cb_5_0/io_wo[18]
+ cb_5_0/io_wo[19] cb_5_0/io_wo[1] cb_5_0/io_wo[20] cb_5_0/io_wo[21] cb_5_0/io_wo[22]
+ cb_5_0/io_wo[23] cb_5_0/io_wo[24] cb_5_0/io_wo[25] cb_5_0/io_wo[26] cb_5_0/io_wo[27]
+ cb_5_0/io_wo[28] cb_5_0/io_wo[29] cb_5_0/io_wo[2] cb_5_0/io_wo[30] cb_5_0/io_wo[31]
+ cb_5_0/io_wo[32] cb_5_0/io_wo[33] cb_5_0/io_wo[34] cb_5_0/io_wo[35] cb_5_0/io_wo[36]
+ cb_5_0/io_wo[37] cb_5_0/io_wo[38] cb_5_0/io_wo[39] cb_5_0/io_wo[3] cb_5_0/io_wo[40]
+ cb_5_0/io_wo[41] cb_5_0/io_wo[42] cb_5_0/io_wo[43] cb_5_0/io_wo[44] cb_5_0/io_wo[45]
+ cb_5_0/io_wo[46] cb_5_0/io_wo[47] cb_5_0/io_wo[48] cb_5_0/io_wo[49] cb_5_0/io_wo[4]
+ cb_5_0/io_wo[50] cb_5_0/io_wo[51] cb_5_0/io_wo[52] cb_5_0/io_wo[53] cb_5_0/io_wo[54]
+ cb_5_0/io_wo[55] cb_5_0/io_wo[56] cb_5_0/io_wo[57] cb_5_0/io_wo[58] cb_5_0/io_wo[59]
+ cb_5_0/io_wo[5] cb_5_0/io_wo[60] cb_5_0/io_wo[61] cb_5_0/io_wo[62] cb_5_0/io_wo[63]
+ cb_5_0/io_wo[6] cb_5_0/io_wo[7] cb_5_0/io_wo[8] cb_5_0/io_wo[9] icon/dsi[0] icon/dsi[1]
+ icon/dsi[2] icon/dsi[3] icon/dsi[4] icon/dsi[5] icon/dsi[6] icon/dsi[7] ccon_5/io_dsi_o
+ ccon_5/io_irq cb_5_0/io_vi cb_5_10/io_vi cb_5_1/io_vi cb_5_2/io_vi cb_5_3/io_vi
+ cb_5_4/io_vi cb_5_5/io_vi cb_5_6/io_vi cb_5_7/io_vi cb_5_8/io_vi cb_5_9/io_vi ccon_7/io_we_i
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_con
Xcb_5_9 cb_5_9/io_adr_i[0] cb_5_9/io_adr_i[1] cb_5_9/io_cs_i cb_5_9/io_dat_i[0] cb_5_9/io_dat_i[10]
+ cb_5_9/io_dat_i[11] cb_5_9/io_dat_i[12] cb_5_9/io_dat_i[13] cb_5_9/io_dat_i[14]
+ cb_5_9/io_dat_i[15] cb_5_9/io_dat_i[1] cb_5_9/io_dat_i[2] cb_5_9/io_dat_i[3] cb_5_9/io_dat_i[4]
+ cb_5_9/io_dat_i[5] cb_5_9/io_dat_i[6] cb_5_9/io_dat_i[7] cb_5_9/io_dat_i[8] cb_5_9/io_dat_i[9]
+ cb_5_9/io_dat_o[0] cb_5_9/io_dat_o[10] cb_5_9/io_dat_o[11] cb_5_9/io_dat_o[12] cb_5_9/io_dat_o[13]
+ cb_5_9/io_dat_o[14] cb_5_9/io_dat_o[15] cb_5_9/io_dat_o[1] cb_5_9/io_dat_o[2] cb_5_9/io_dat_o[3]
+ cb_5_9/io_dat_o[4] cb_5_9/io_dat_o[5] cb_5_9/io_dat_o[6] cb_5_9/io_dat_o[7] cb_5_9/io_dat_o[8]
+ cb_5_9/io_dat_o[9] cb_5_9/io_eo[0] cb_5_9/io_eo[10] cb_5_9/io_eo[11] cb_5_9/io_eo[12]
+ cb_5_9/io_eo[13] cb_5_9/io_eo[14] cb_5_9/io_eo[15] cb_5_9/io_eo[16] cb_5_9/io_eo[17]
+ cb_5_9/io_eo[18] cb_5_9/io_eo[19] cb_5_9/io_eo[1] cb_5_9/io_eo[20] cb_5_9/io_eo[21]
+ cb_5_9/io_eo[22] cb_5_9/io_eo[23] cb_5_9/io_eo[24] cb_5_9/io_eo[25] cb_5_9/io_eo[26]
+ cb_5_9/io_eo[27] cb_5_9/io_eo[28] cb_5_9/io_eo[29] cb_5_9/io_eo[2] cb_5_9/io_eo[30]
+ cb_5_9/io_eo[31] cb_5_9/io_eo[32] cb_5_9/io_eo[33] cb_5_9/io_eo[34] cb_5_9/io_eo[35]
+ cb_5_9/io_eo[36] cb_5_9/io_eo[37] cb_5_9/io_eo[38] cb_5_9/io_eo[39] cb_5_9/io_eo[3]
+ cb_5_9/io_eo[40] cb_5_9/io_eo[41] cb_5_9/io_eo[42] cb_5_9/io_eo[43] cb_5_9/io_eo[44]
+ cb_5_9/io_eo[45] cb_5_9/io_eo[46] cb_5_9/io_eo[47] cb_5_9/io_eo[48] cb_5_9/io_eo[49]
+ cb_5_9/io_eo[4] cb_5_9/io_eo[50] cb_5_9/io_eo[51] cb_5_9/io_eo[52] cb_5_9/io_eo[53]
+ cb_5_9/io_eo[54] cb_5_9/io_eo[55] cb_5_9/io_eo[56] cb_5_9/io_eo[57] cb_5_9/io_eo[58]
+ cb_5_9/io_eo[59] cb_5_9/io_eo[5] cb_5_9/io_eo[60] cb_5_9/io_eo[61] cb_5_9/io_eo[62]
+ cb_5_9/io_eo[63] cb_5_9/io_eo[6] cb_5_9/io_eo[7] cb_5_9/io_eo[8] cb_5_9/io_eo[9]
+ cb_5_9/io_i_0_ci cb_5_9/io_i_0_in1[0] cb_5_9/io_i_0_in1[1] cb_5_9/io_i_0_in1[2]
+ cb_5_9/io_i_0_in1[3] cb_5_9/io_i_0_in1[4] cb_5_9/io_i_0_in1[5] cb_5_9/io_i_0_in1[6]
+ cb_5_9/io_i_0_in1[7] cb_5_9/io_i_1_ci cb_5_9/io_i_1_in1[0] cb_5_9/io_i_1_in1[1]
+ cb_5_9/io_i_1_in1[2] cb_5_9/io_i_1_in1[3] cb_5_9/io_i_1_in1[4] cb_5_9/io_i_1_in1[5]
+ cb_5_9/io_i_1_in1[6] cb_5_9/io_i_1_in1[7] cb_5_9/io_i_2_ci cb_5_9/io_i_2_in1[0]
+ cb_5_9/io_i_2_in1[1] cb_5_9/io_i_2_in1[2] cb_5_9/io_i_2_in1[3] cb_5_9/io_i_2_in1[4]
+ cb_5_9/io_i_2_in1[5] cb_5_9/io_i_2_in1[6] cb_5_9/io_i_2_in1[7] cb_5_9/io_i_3_ci
+ cb_5_9/io_i_3_in1[0] cb_5_9/io_i_3_in1[1] cb_5_9/io_i_3_in1[2] cb_5_9/io_i_3_in1[3]
+ cb_5_9/io_i_3_in1[4] cb_5_9/io_i_3_in1[5] cb_5_9/io_i_3_in1[6] cb_5_9/io_i_3_in1[7]
+ cb_5_9/io_i_4_ci cb_5_9/io_i_4_in1[0] cb_5_9/io_i_4_in1[1] cb_5_9/io_i_4_in1[2]
+ cb_5_9/io_i_4_in1[3] cb_5_9/io_i_4_in1[4] cb_5_9/io_i_4_in1[5] cb_5_9/io_i_4_in1[6]
+ cb_5_9/io_i_4_in1[7] cb_5_9/io_i_5_ci cb_5_9/io_i_5_in1[0] cb_5_9/io_i_5_in1[1]
+ cb_5_9/io_i_5_in1[2] cb_5_9/io_i_5_in1[3] cb_5_9/io_i_5_in1[4] cb_5_9/io_i_5_in1[5]
+ cb_5_9/io_i_5_in1[6] cb_5_9/io_i_5_in1[7] cb_5_9/io_i_6_ci cb_5_9/io_i_6_in1[0]
+ cb_5_9/io_i_6_in1[1] cb_5_9/io_i_6_in1[2] cb_5_9/io_i_6_in1[3] cb_5_9/io_i_6_in1[4]
+ cb_5_9/io_i_6_in1[5] cb_5_9/io_i_6_in1[6] cb_5_9/io_i_6_in1[7] cb_5_9/io_i_7_ci
+ cb_5_9/io_i_7_in1[0] cb_5_9/io_i_7_in1[1] cb_5_9/io_i_7_in1[2] cb_5_9/io_i_7_in1[3]
+ cb_5_9/io_i_7_in1[4] cb_5_9/io_i_7_in1[5] cb_5_9/io_i_7_in1[6] cb_5_9/io_i_7_in1[7]
+ cb_5_9/io_o_0_co cb_5_9/io_o_0_out[0] cb_5_9/io_o_0_out[1] cb_5_9/io_o_0_out[2]
+ cb_5_9/io_o_0_out[3] cb_5_9/io_o_0_out[4] cb_5_9/io_o_0_out[5] cb_5_9/io_o_0_out[6]
+ cb_5_9/io_o_0_out[7] cb_5_9/io_o_1_co cb_5_9/io_o_1_out[0] cb_5_9/io_o_1_out[1]
+ cb_5_9/io_o_1_out[2] cb_5_9/io_o_1_out[3] cb_5_9/io_o_1_out[4] cb_5_9/io_o_1_out[5]
+ cb_5_9/io_o_1_out[6] cb_5_9/io_o_1_out[7] cb_5_9/io_o_2_co cb_5_9/io_o_2_out[0]
+ cb_5_9/io_o_2_out[1] cb_5_9/io_o_2_out[2] cb_5_9/io_o_2_out[3] cb_5_9/io_o_2_out[4]
+ cb_5_9/io_o_2_out[5] cb_5_9/io_o_2_out[6] cb_5_9/io_o_2_out[7] cb_5_9/io_o_3_co
+ cb_5_9/io_o_3_out[0] cb_5_9/io_o_3_out[1] cb_5_9/io_o_3_out[2] cb_5_9/io_o_3_out[3]
+ cb_5_9/io_o_3_out[4] cb_5_9/io_o_3_out[5] cb_5_9/io_o_3_out[6] cb_5_9/io_o_3_out[7]
+ cb_5_9/io_o_4_co cb_5_9/io_o_4_out[0] cb_5_9/io_o_4_out[1] cb_5_9/io_o_4_out[2]
+ cb_5_9/io_o_4_out[3] cb_5_9/io_o_4_out[4] cb_5_9/io_o_4_out[5] cb_5_9/io_o_4_out[6]
+ cb_5_9/io_o_4_out[7] cb_5_9/io_o_5_co cb_5_9/io_o_5_out[0] cb_5_9/io_o_5_out[1]
+ cb_5_9/io_o_5_out[2] cb_5_9/io_o_5_out[3] cb_5_9/io_o_5_out[4] cb_5_9/io_o_5_out[5]
+ cb_5_9/io_o_5_out[6] cb_5_9/io_o_5_out[7] cb_5_9/io_o_6_co cb_5_9/io_o_6_out[0]
+ cb_5_9/io_o_6_out[1] cb_5_9/io_o_6_out[2] cb_5_9/io_o_6_out[3] cb_5_9/io_o_6_out[4]
+ cb_5_9/io_o_6_out[5] cb_5_9/io_o_6_out[6] cb_5_9/io_o_6_out[7] cb_5_9/io_o_7_co
+ cb_5_9/io_o_7_out[0] cb_5_9/io_o_7_out[1] cb_5_9/io_o_7_out[2] cb_5_9/io_o_7_out[3]
+ cb_5_9/io_o_7_out[4] cb_5_9/io_o_7_out[5] cb_5_9/io_o_7_out[6] cb_5_9/io_o_7_out[7]
+ cb_5_9/io_vci cb_5_9/io_vco cb_5_9/io_vi cb_5_9/io_we_i cb_5_9/io_wo[0] cb_5_9/io_wo[10]
+ cb_5_9/io_wo[11] cb_5_9/io_wo[12] cb_5_9/io_wo[13] cb_5_9/io_wo[14] cb_5_9/io_wo[15]
+ cb_5_9/io_wo[16] cb_5_9/io_wo[17] cb_5_9/io_wo[18] cb_5_9/io_wo[19] cb_5_9/io_wo[1]
+ cb_5_9/io_wo[20] cb_5_9/io_wo[21] cb_5_9/io_wo[22] cb_5_9/io_wo[23] cb_5_9/io_wo[24]
+ cb_5_9/io_wo[25] cb_5_9/io_wo[26] cb_5_9/io_wo[27] cb_5_9/io_wo[28] cb_5_9/io_wo[29]
+ cb_5_9/io_wo[2] cb_5_9/io_wo[30] cb_5_9/io_wo[31] cb_5_9/io_wo[32] cb_5_9/io_wo[33]
+ cb_5_9/io_wo[34] cb_5_9/io_wo[35] cb_5_9/io_wo[36] cb_5_9/io_wo[37] cb_5_9/io_wo[38]
+ cb_5_9/io_wo[39] cb_5_9/io_wo[3] cb_5_9/io_wo[40] cb_5_9/io_wo[41] cb_5_9/io_wo[42]
+ cb_5_9/io_wo[43] cb_5_9/io_wo[44] cb_5_9/io_wo[45] cb_5_9/io_wo[46] cb_5_9/io_wo[47]
+ cb_5_9/io_wo[48] cb_5_9/io_wo[49] cb_5_9/io_wo[4] cb_5_9/io_wo[50] cb_5_9/io_wo[51]
+ cb_5_9/io_wo[52] cb_5_9/io_wo[53] cb_5_9/io_wo[54] cb_5_9/io_wo[55] cb_5_9/io_wo[56]
+ cb_5_9/io_wo[57] cb_5_9/io_wo[58] cb_5_9/io_wo[59] cb_5_9/io_wo[5] cb_5_9/io_wo[60]
+ cb_5_9/io_wo[61] cb_5_9/io_wo[62] cb_5_9/io_wo[63] cb_5_9/io_wo[6] cb_5_9/io_wo[7]
+ cb_5_9/io_wo[8] cb_5_9/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xicon icon/dsi[0] icon/dsi[1] icon/dsi[2] icon/dsi[3] icon/dsi[4] icon/dsi[5] icon/dsi[6]
+ icon/dsi[7] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] user_irq[0]
+ user_irq[1] user_irq[2] mcons_0/io_irq ccon_6/io_irq ccon_7/io_irq mcons_1/io_irq
+ mcons_2/io_irq mcons_3/io_irq ccon_0/io_irq ccon_1/io_irq ccon_2/io_irq ccon_3/io_irq
+ ccon_4/io_irq ccon_5/io_irq mcons_3/clock mcons_3/reset mcons_0/io_wb_ack_o ccon_6/io_ack_o
+ ccon_7/io_ack_o mcons_1/io_wb_ack_o mcons_2/io_wb_ack_o mcons_3/io_wb_ack_o ccon_0/io_ack_o
+ ccon_1/io_ack_o ccon_2/io_ack_o ccon_3/io_ack_o ccon_4/io_ack_o ccon_5/io_ack_o
+ ccon_7/io_adr_i[0] ccon_7/io_adr_i[10] ccon_7/io_adr_i[11] ccon_7/io_adr_i[1] ccon_7/io_adr_i[2]
+ ccon_7/io_adr_i[3] ccon_7/io_adr_i[4] ccon_7/io_adr_i[5] ccon_7/io_adr_i[6] ccon_7/io_adr_i[7]
+ ccon_7/io_adr_i[8] ccon_7/io_adr_i[9] mcons_0/io_wb_cs_i ccon_6/io_cs_i ccon_7/io_cs_i
+ mcons_1/io_wb_cs_i mcons_2/io_wb_cs_i mcons_3/io_wb_cs_i ccon_0/io_cs_i ccon_1/io_cs_i
+ ccon_2/io_cs_i ccon_3/io_cs_i ccon_4/io_cs_i ccon_5/io_cs_i ccon_7/io_dat_i[0] ccon_7/io_dat_i[10]
+ ccon_7/io_dat_i[11] ccon_7/io_dat_i[12] ccon_7/io_dat_i[13] ccon_7/io_dat_i[14]
+ ccon_7/io_dat_i[15] ccon_7/io_dat_i[16] ccon_7/io_dat_i[17] ccon_7/io_dat_i[18]
+ ccon_7/io_dat_i[19] ccon_7/io_dat_i[1] ccon_7/io_dat_i[20] ccon_7/io_dat_i[21] ccon_7/io_dat_i[22]
+ ccon_7/io_dat_i[23] ccon_7/io_dat_i[24] ccon_7/io_dat_i[25] ccon_7/io_dat_i[26]
+ ccon_7/io_dat_i[27] ccon_7/io_dat_i[28] ccon_7/io_dat_i[29] ccon_7/io_dat_i[2] ccon_7/io_dat_i[30]
+ ccon_7/io_dat_i[31] ccon_7/io_dat_i[3] ccon_7/io_dat_i[4] ccon_7/io_dat_i[5] ccon_7/io_dat_i[6]
+ ccon_7/io_dat_i[7] ccon_7/io_dat_i[8] ccon_7/io_dat_i[9] icon/m_wbs_dat_o_0[0] icon/m_wbs_dat_o_0[10]
+ icon/m_wbs_dat_o_0[11] icon/m_wbs_dat_o_0[12] icon/m_wbs_dat_o_0[13] icon/m_wbs_dat_o_0[14]
+ icon/m_wbs_dat_o_0[15] icon/m_wbs_dat_o_0[16] icon/m_wbs_dat_o_0[17] icon/m_wbs_dat_o_0[18]
+ icon/m_wbs_dat_o_0[19] icon/m_wbs_dat_o_0[1] icon/m_wbs_dat_o_0[20] icon/m_wbs_dat_o_0[21]
+ icon/m_wbs_dat_o_0[22] icon/m_wbs_dat_o_0[23] icon/m_wbs_dat_o_0[24] icon/m_wbs_dat_o_0[25]
+ icon/m_wbs_dat_o_0[26] icon/m_wbs_dat_o_0[27] icon/m_wbs_dat_o_0[28] icon/m_wbs_dat_o_0[29]
+ icon/m_wbs_dat_o_0[2] icon/m_wbs_dat_o_0[30] icon/m_wbs_dat_o_0[31] icon/m_wbs_dat_o_0[3]
+ icon/m_wbs_dat_o_0[4] icon/m_wbs_dat_o_0[5] icon/m_wbs_dat_o_0[6] icon/m_wbs_dat_o_0[7]
+ icon/m_wbs_dat_o_0[8] icon/m_wbs_dat_o_0[9] ccon_6/io_dat_o[0] ccon_6/io_dat_o[10]
+ ccon_6/io_dat_o[11] ccon_6/io_dat_o[12] ccon_6/io_dat_o[13] ccon_6/io_dat_o[14]
+ ccon_6/io_dat_o[15] ccon_6/io_dat_o[16] ccon_6/io_dat_o[17] ccon_6/io_dat_o[18]
+ ccon_6/io_dat_o[19] ccon_6/io_dat_o[1] ccon_6/io_dat_o[20] ccon_6/io_dat_o[21] ccon_6/io_dat_o[22]
+ ccon_6/io_dat_o[23] ccon_6/io_dat_o[24] ccon_6/io_dat_o[25] ccon_6/io_dat_o[26]
+ ccon_6/io_dat_o[27] ccon_6/io_dat_o[28] ccon_6/io_dat_o[29] ccon_6/io_dat_o[2] ccon_6/io_dat_o[30]
+ ccon_6/io_dat_o[31] ccon_6/io_dat_o[3] ccon_6/io_dat_o[4] ccon_6/io_dat_o[5] ccon_6/io_dat_o[6]
+ ccon_6/io_dat_o[7] ccon_6/io_dat_o[8] ccon_6/io_dat_o[9] ccon_7/io_dat_o[0] ccon_7/io_dat_o[10]
+ ccon_7/io_dat_o[11] ccon_7/io_dat_o[12] ccon_7/io_dat_o[13] ccon_7/io_dat_o[14]
+ ccon_7/io_dat_o[15] ccon_7/io_dat_o[16] ccon_7/io_dat_o[17] ccon_7/io_dat_o[18]
+ ccon_7/io_dat_o[19] ccon_7/io_dat_o[1] ccon_7/io_dat_o[20] ccon_7/io_dat_o[21] ccon_7/io_dat_o[22]
+ ccon_7/io_dat_o[23] ccon_7/io_dat_o[24] ccon_7/io_dat_o[25] ccon_7/io_dat_o[26]
+ ccon_7/io_dat_o[27] ccon_7/io_dat_o[28] ccon_7/io_dat_o[29] ccon_7/io_dat_o[2] ccon_7/io_dat_o[30]
+ ccon_7/io_dat_o[31] ccon_7/io_dat_o[3] ccon_7/io_dat_o[4] ccon_7/io_dat_o[5] ccon_7/io_dat_o[6]
+ ccon_7/io_dat_o[7] ccon_7/io_dat_o[8] ccon_7/io_dat_o[9] icon/m_wbs_dat_o_1[0] icon/m_wbs_dat_o_1[10]
+ icon/m_wbs_dat_o_1[11] icon/m_wbs_dat_o_1[12] icon/m_wbs_dat_o_1[13] icon/m_wbs_dat_o_1[14]
+ icon/m_wbs_dat_o_1[15] icon/m_wbs_dat_o_1[16] icon/m_wbs_dat_o_1[17] icon/m_wbs_dat_o_1[18]
+ icon/m_wbs_dat_o_1[19] icon/m_wbs_dat_o_1[1] icon/m_wbs_dat_o_1[20] icon/m_wbs_dat_o_1[21]
+ icon/m_wbs_dat_o_1[22] icon/m_wbs_dat_o_1[23] icon/m_wbs_dat_o_1[24] icon/m_wbs_dat_o_1[25]
+ icon/m_wbs_dat_o_1[26] icon/m_wbs_dat_o_1[27] icon/m_wbs_dat_o_1[28] icon/m_wbs_dat_o_1[29]
+ icon/m_wbs_dat_o_1[2] icon/m_wbs_dat_o_1[30] icon/m_wbs_dat_o_1[31] icon/m_wbs_dat_o_1[3]
+ icon/m_wbs_dat_o_1[4] icon/m_wbs_dat_o_1[5] icon/m_wbs_dat_o_1[6] icon/m_wbs_dat_o_1[7]
+ icon/m_wbs_dat_o_1[8] icon/m_wbs_dat_o_1[9] icon/m_wbs_dat_o_2[0] icon/m_wbs_dat_o_2[10]
+ icon/m_wbs_dat_o_2[11] icon/m_wbs_dat_o_2[12] icon/m_wbs_dat_o_2[13] icon/m_wbs_dat_o_2[14]
+ icon/m_wbs_dat_o_2[15] icon/m_wbs_dat_o_2[16] icon/m_wbs_dat_o_2[17] icon/m_wbs_dat_o_2[18]
+ icon/m_wbs_dat_o_2[19] icon/m_wbs_dat_o_2[1] icon/m_wbs_dat_o_2[20] icon/m_wbs_dat_o_2[21]
+ icon/m_wbs_dat_o_2[22] icon/m_wbs_dat_o_2[23] icon/m_wbs_dat_o_2[24] icon/m_wbs_dat_o_2[25]
+ icon/m_wbs_dat_o_2[26] icon/m_wbs_dat_o_2[27] icon/m_wbs_dat_o_2[28] icon/m_wbs_dat_o_2[29]
+ icon/m_wbs_dat_o_2[2] icon/m_wbs_dat_o_2[30] icon/m_wbs_dat_o_2[31] icon/m_wbs_dat_o_2[3]
+ icon/m_wbs_dat_o_2[4] icon/m_wbs_dat_o_2[5] icon/m_wbs_dat_o_2[6] icon/m_wbs_dat_o_2[7]
+ icon/m_wbs_dat_o_2[8] icon/m_wbs_dat_o_2[9] icon/m_wbs_dat_o_3[0] icon/m_wbs_dat_o_3[10]
+ icon/m_wbs_dat_o_3[11] icon/m_wbs_dat_o_3[12] icon/m_wbs_dat_o_3[13] icon/m_wbs_dat_o_3[14]
+ icon/m_wbs_dat_o_3[15] icon/m_wbs_dat_o_3[16] icon/m_wbs_dat_o_3[17] icon/m_wbs_dat_o_3[18]
+ icon/m_wbs_dat_o_3[19] icon/m_wbs_dat_o_3[1] icon/m_wbs_dat_o_3[20] icon/m_wbs_dat_o_3[21]
+ icon/m_wbs_dat_o_3[22] icon/m_wbs_dat_o_3[23] icon/m_wbs_dat_o_3[24] icon/m_wbs_dat_o_3[25]
+ icon/m_wbs_dat_o_3[26] icon/m_wbs_dat_o_3[27] icon/m_wbs_dat_o_3[28] icon/m_wbs_dat_o_3[29]
+ icon/m_wbs_dat_o_3[2] icon/m_wbs_dat_o_3[30] icon/m_wbs_dat_o_3[31] icon/m_wbs_dat_o_3[3]
+ icon/m_wbs_dat_o_3[4] icon/m_wbs_dat_o_3[5] icon/m_wbs_dat_o_3[6] icon/m_wbs_dat_o_3[7]
+ icon/m_wbs_dat_o_3[8] icon/m_wbs_dat_o_3[9] ccon_0/io_dat_o[0] ccon_0/io_dat_o[10]
+ ccon_0/io_dat_o[11] ccon_0/io_dat_o[12] ccon_0/io_dat_o[13] ccon_0/io_dat_o[14]
+ ccon_0/io_dat_o[15] ccon_0/io_dat_o[16] ccon_0/io_dat_o[17] ccon_0/io_dat_o[18]
+ ccon_0/io_dat_o[19] ccon_0/io_dat_o[1] ccon_0/io_dat_o[20] ccon_0/io_dat_o[21] ccon_0/io_dat_o[22]
+ ccon_0/io_dat_o[23] ccon_0/io_dat_o[24] ccon_0/io_dat_o[25] ccon_0/io_dat_o[26]
+ ccon_0/io_dat_o[27] ccon_0/io_dat_o[28] ccon_0/io_dat_o[29] ccon_0/io_dat_o[2] ccon_0/io_dat_o[30]
+ ccon_0/io_dat_o[31] ccon_0/io_dat_o[3] ccon_0/io_dat_o[4] ccon_0/io_dat_o[5] ccon_0/io_dat_o[6]
+ ccon_0/io_dat_o[7] ccon_0/io_dat_o[8] ccon_0/io_dat_o[9] ccon_1/io_dat_o[0] ccon_1/io_dat_o[10]
+ ccon_1/io_dat_o[11] ccon_1/io_dat_o[12] ccon_1/io_dat_o[13] ccon_1/io_dat_o[14]
+ ccon_1/io_dat_o[15] ccon_1/io_dat_o[16] ccon_1/io_dat_o[17] ccon_1/io_dat_o[18]
+ ccon_1/io_dat_o[19] ccon_1/io_dat_o[1] ccon_1/io_dat_o[20] ccon_1/io_dat_o[21] ccon_1/io_dat_o[22]
+ ccon_1/io_dat_o[23] ccon_1/io_dat_o[24] ccon_1/io_dat_o[25] ccon_1/io_dat_o[26]
+ ccon_1/io_dat_o[27] ccon_1/io_dat_o[28] ccon_1/io_dat_o[29] ccon_1/io_dat_o[2] ccon_1/io_dat_o[30]
+ ccon_1/io_dat_o[31] ccon_1/io_dat_o[3] ccon_1/io_dat_o[4] ccon_1/io_dat_o[5] ccon_1/io_dat_o[6]
+ ccon_1/io_dat_o[7] ccon_1/io_dat_o[8] ccon_1/io_dat_o[9] ccon_2/io_dat_o[0] ccon_2/io_dat_o[10]
+ ccon_2/io_dat_o[11] ccon_2/io_dat_o[12] ccon_2/io_dat_o[13] ccon_2/io_dat_o[14]
+ ccon_2/io_dat_o[15] ccon_2/io_dat_o[16] ccon_2/io_dat_o[17] ccon_2/io_dat_o[18]
+ ccon_2/io_dat_o[19] ccon_2/io_dat_o[1] ccon_2/io_dat_o[20] ccon_2/io_dat_o[21] ccon_2/io_dat_o[22]
+ ccon_2/io_dat_o[23] ccon_2/io_dat_o[24] ccon_2/io_dat_o[25] ccon_2/io_dat_o[26]
+ ccon_2/io_dat_o[27] ccon_2/io_dat_o[28] ccon_2/io_dat_o[29] ccon_2/io_dat_o[2] ccon_2/io_dat_o[30]
+ ccon_2/io_dat_o[31] ccon_2/io_dat_o[3] ccon_2/io_dat_o[4] ccon_2/io_dat_o[5] ccon_2/io_dat_o[6]
+ ccon_2/io_dat_o[7] ccon_2/io_dat_o[8] ccon_2/io_dat_o[9] ccon_3/io_dat_o[0] ccon_3/io_dat_o[10]
+ ccon_3/io_dat_o[11] ccon_3/io_dat_o[12] ccon_3/io_dat_o[13] ccon_3/io_dat_o[14]
+ ccon_3/io_dat_o[15] ccon_3/io_dat_o[16] ccon_3/io_dat_o[17] ccon_3/io_dat_o[18]
+ ccon_3/io_dat_o[19] ccon_3/io_dat_o[1] ccon_3/io_dat_o[20] ccon_3/io_dat_o[21] ccon_3/io_dat_o[22]
+ ccon_3/io_dat_o[23] ccon_3/io_dat_o[24] ccon_3/io_dat_o[25] ccon_3/io_dat_o[26]
+ ccon_3/io_dat_o[27] ccon_3/io_dat_o[28] ccon_3/io_dat_o[29] ccon_3/io_dat_o[2] ccon_3/io_dat_o[30]
+ ccon_3/io_dat_o[31] ccon_3/io_dat_o[3] ccon_3/io_dat_o[4] ccon_3/io_dat_o[5] ccon_3/io_dat_o[6]
+ ccon_3/io_dat_o[7] ccon_3/io_dat_o[8] ccon_3/io_dat_o[9] ccon_4/io_dat_o[0] ccon_4/io_dat_o[10]
+ ccon_4/io_dat_o[11] ccon_4/io_dat_o[12] ccon_4/io_dat_o[13] ccon_4/io_dat_o[14]
+ ccon_4/io_dat_o[15] ccon_4/io_dat_o[16] ccon_4/io_dat_o[17] ccon_4/io_dat_o[18]
+ ccon_4/io_dat_o[19] ccon_4/io_dat_o[1] ccon_4/io_dat_o[20] ccon_4/io_dat_o[21] ccon_4/io_dat_o[22]
+ ccon_4/io_dat_o[23] ccon_4/io_dat_o[24] ccon_4/io_dat_o[25] ccon_4/io_dat_o[26]
+ ccon_4/io_dat_o[27] ccon_4/io_dat_o[28] ccon_4/io_dat_o[29] ccon_4/io_dat_o[2] ccon_4/io_dat_o[30]
+ ccon_4/io_dat_o[31] ccon_4/io_dat_o[3] ccon_4/io_dat_o[4] ccon_4/io_dat_o[5] ccon_4/io_dat_o[6]
+ ccon_4/io_dat_o[7] ccon_4/io_dat_o[8] ccon_4/io_dat_o[9] ccon_5/io_dat_o[0] ccon_5/io_dat_o[10]
+ ccon_5/io_dat_o[11] ccon_5/io_dat_o[12] ccon_5/io_dat_o[13] ccon_5/io_dat_o[14]
+ ccon_5/io_dat_o[15] ccon_5/io_dat_o[16] ccon_5/io_dat_o[17] ccon_5/io_dat_o[18]
+ ccon_5/io_dat_o[19] ccon_5/io_dat_o[1] ccon_5/io_dat_o[20] ccon_5/io_dat_o[21] ccon_5/io_dat_o[22]
+ ccon_5/io_dat_o[23] ccon_5/io_dat_o[24] ccon_5/io_dat_o[25] ccon_5/io_dat_o[26]
+ ccon_5/io_dat_o[27] ccon_5/io_dat_o[28] ccon_5/io_dat_o[29] ccon_5/io_dat_o[2] ccon_5/io_dat_o[30]
+ ccon_5/io_dat_o[31] ccon_5/io_dat_o[3] ccon_5/io_dat_o[4] ccon_5/io_dat_o[5] ccon_5/io_dat_o[6]
+ ccon_5/io_dat_o[7] ccon_5/io_dat_o[8] ccon_5/io_dat_o[9] ccon_7/io_we_i icon/mt_QEI_ChA_0
+ icon/mt_QEI_ChA_1 icon/mt_QEI_ChA_2 icon/mt_QEI_ChA_3 icon/mt_QEI_ChB_0 icon/mt_QEI_ChB_1
+ icon/mt_QEI_ChB_2 icon/mt_QEI_ChB_3 icon/mt_pwm_h_0 icon/mt_pwm_h_1 icon/mt_pwm_h_2
+ icon/mt_pwm_h_3 icon/mt_pwm_l_0 icon/mt_pwm_l_1 icon/mt_pwm_l_2 icon/mt_pwm_l_3
+ wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i vccd1 vssd1
+ wb_local
Xcb_3_6 cb_3_9/io_adr_i[0] cb_3_9/io_adr_i[1] cb_3_6/io_cs_i cb_3_9/io_dat_i[0] cb_3_9/io_dat_i[10]
+ cb_3_9/io_dat_i[11] cb_3_9/io_dat_i[12] cb_3_9/io_dat_i[13] cb_3_9/io_dat_i[14]
+ cb_3_9/io_dat_i[15] cb_3_9/io_dat_i[1] cb_3_9/io_dat_i[2] cb_3_9/io_dat_i[3] cb_3_9/io_dat_i[4]
+ cb_3_9/io_dat_i[5] cb_3_9/io_dat_i[6] cb_3_9/io_dat_i[7] cb_3_9/io_dat_i[8] cb_3_9/io_dat_i[9]
+ cb_3_6/io_dat_o[0] cb_3_6/io_dat_o[10] cb_3_6/io_dat_o[11] cb_3_6/io_dat_o[12] cb_3_6/io_dat_o[13]
+ cb_3_6/io_dat_o[14] cb_3_6/io_dat_o[15] cb_3_6/io_dat_o[1] cb_3_6/io_dat_o[2] cb_3_6/io_dat_o[3]
+ cb_3_6/io_dat_o[4] cb_3_6/io_dat_o[5] cb_3_6/io_dat_o[6] cb_3_6/io_dat_o[7] cb_3_6/io_dat_o[8]
+ cb_3_6/io_dat_o[9] cb_3_7/io_wo[0] cb_3_7/io_wo[10] cb_3_7/io_wo[11] cb_3_7/io_wo[12]
+ cb_3_7/io_wo[13] cb_3_7/io_wo[14] cb_3_7/io_wo[15] cb_3_7/io_wo[16] cb_3_7/io_wo[17]
+ cb_3_7/io_wo[18] cb_3_7/io_wo[19] cb_3_7/io_wo[1] cb_3_7/io_wo[20] cb_3_7/io_wo[21]
+ cb_3_7/io_wo[22] cb_3_7/io_wo[23] cb_3_7/io_wo[24] cb_3_7/io_wo[25] cb_3_7/io_wo[26]
+ cb_3_7/io_wo[27] cb_3_7/io_wo[28] cb_3_7/io_wo[29] cb_3_7/io_wo[2] cb_3_7/io_wo[30]
+ cb_3_7/io_wo[31] cb_3_7/io_wo[32] cb_3_7/io_wo[33] cb_3_7/io_wo[34] cb_3_7/io_wo[35]
+ cb_3_7/io_wo[36] cb_3_7/io_wo[37] cb_3_7/io_wo[38] cb_3_7/io_wo[39] cb_3_7/io_wo[3]
+ cb_3_7/io_wo[40] cb_3_7/io_wo[41] cb_3_7/io_wo[42] cb_3_7/io_wo[43] cb_3_7/io_wo[44]
+ cb_3_7/io_wo[45] cb_3_7/io_wo[46] cb_3_7/io_wo[47] cb_3_7/io_wo[48] cb_3_7/io_wo[49]
+ cb_3_7/io_wo[4] cb_3_7/io_wo[50] cb_3_7/io_wo[51] cb_3_7/io_wo[52] cb_3_7/io_wo[53]
+ cb_3_7/io_wo[54] cb_3_7/io_wo[55] cb_3_7/io_wo[56] cb_3_7/io_wo[57] cb_3_7/io_wo[58]
+ cb_3_7/io_wo[59] cb_3_7/io_wo[5] cb_3_7/io_wo[60] cb_3_7/io_wo[61] cb_3_7/io_wo[62]
+ cb_3_7/io_wo[63] cb_3_7/io_wo[6] cb_3_7/io_wo[7] cb_3_7/io_wo[8] cb_3_7/io_wo[9]
+ cb_3_6/io_i_0_ci cb_3_6/io_i_0_in1[0] cb_3_6/io_i_0_in1[1] cb_3_6/io_i_0_in1[2]
+ cb_3_6/io_i_0_in1[3] cb_3_6/io_i_0_in1[4] cb_3_6/io_i_0_in1[5] cb_3_6/io_i_0_in1[6]
+ cb_3_6/io_i_0_in1[7] cb_3_6/io_i_1_ci cb_3_6/io_i_1_in1[0] cb_3_6/io_i_1_in1[1]
+ cb_3_6/io_i_1_in1[2] cb_3_6/io_i_1_in1[3] cb_3_6/io_i_1_in1[4] cb_3_6/io_i_1_in1[5]
+ cb_3_6/io_i_1_in1[6] cb_3_6/io_i_1_in1[7] cb_3_6/io_i_2_ci cb_3_6/io_i_2_in1[0]
+ cb_3_6/io_i_2_in1[1] cb_3_6/io_i_2_in1[2] cb_3_6/io_i_2_in1[3] cb_3_6/io_i_2_in1[4]
+ cb_3_6/io_i_2_in1[5] cb_3_6/io_i_2_in1[6] cb_3_6/io_i_2_in1[7] cb_3_6/io_i_3_ci
+ cb_3_6/io_i_3_in1[0] cb_3_6/io_i_3_in1[1] cb_3_6/io_i_3_in1[2] cb_3_6/io_i_3_in1[3]
+ cb_3_6/io_i_3_in1[4] cb_3_6/io_i_3_in1[5] cb_3_6/io_i_3_in1[6] cb_3_6/io_i_3_in1[7]
+ cb_3_6/io_i_4_ci cb_3_6/io_i_4_in1[0] cb_3_6/io_i_4_in1[1] cb_3_6/io_i_4_in1[2]
+ cb_3_6/io_i_4_in1[3] cb_3_6/io_i_4_in1[4] cb_3_6/io_i_4_in1[5] cb_3_6/io_i_4_in1[6]
+ cb_3_6/io_i_4_in1[7] cb_3_6/io_i_5_ci cb_3_6/io_i_5_in1[0] cb_3_6/io_i_5_in1[1]
+ cb_3_6/io_i_5_in1[2] cb_3_6/io_i_5_in1[3] cb_3_6/io_i_5_in1[4] cb_3_6/io_i_5_in1[5]
+ cb_3_6/io_i_5_in1[6] cb_3_6/io_i_5_in1[7] cb_3_6/io_i_6_ci cb_3_6/io_i_6_in1[0]
+ cb_3_6/io_i_6_in1[1] cb_3_6/io_i_6_in1[2] cb_3_6/io_i_6_in1[3] cb_3_6/io_i_6_in1[4]
+ cb_3_6/io_i_6_in1[5] cb_3_6/io_i_6_in1[6] cb_3_6/io_i_6_in1[7] cb_3_6/io_i_7_ci
+ cb_3_6/io_i_7_in1[0] cb_3_6/io_i_7_in1[1] cb_3_6/io_i_7_in1[2] cb_3_6/io_i_7_in1[3]
+ cb_3_6/io_i_7_in1[4] cb_3_6/io_i_7_in1[5] cb_3_6/io_i_7_in1[6] cb_3_6/io_i_7_in1[7]
+ cb_3_7/io_i_0_ci cb_3_7/io_i_0_in1[0] cb_3_7/io_i_0_in1[1] cb_3_7/io_i_0_in1[2]
+ cb_3_7/io_i_0_in1[3] cb_3_7/io_i_0_in1[4] cb_3_7/io_i_0_in1[5] cb_3_7/io_i_0_in1[6]
+ cb_3_7/io_i_0_in1[7] cb_3_7/io_i_1_ci cb_3_7/io_i_1_in1[0] cb_3_7/io_i_1_in1[1]
+ cb_3_7/io_i_1_in1[2] cb_3_7/io_i_1_in1[3] cb_3_7/io_i_1_in1[4] cb_3_7/io_i_1_in1[5]
+ cb_3_7/io_i_1_in1[6] cb_3_7/io_i_1_in1[7] cb_3_7/io_i_2_ci cb_3_7/io_i_2_in1[0]
+ cb_3_7/io_i_2_in1[1] cb_3_7/io_i_2_in1[2] cb_3_7/io_i_2_in1[3] cb_3_7/io_i_2_in1[4]
+ cb_3_7/io_i_2_in1[5] cb_3_7/io_i_2_in1[6] cb_3_7/io_i_2_in1[7] cb_3_7/io_i_3_ci
+ cb_3_7/io_i_3_in1[0] cb_3_7/io_i_3_in1[1] cb_3_7/io_i_3_in1[2] cb_3_7/io_i_3_in1[3]
+ cb_3_7/io_i_3_in1[4] cb_3_7/io_i_3_in1[5] cb_3_7/io_i_3_in1[6] cb_3_7/io_i_3_in1[7]
+ cb_3_7/io_i_4_ci cb_3_7/io_i_4_in1[0] cb_3_7/io_i_4_in1[1] cb_3_7/io_i_4_in1[2]
+ cb_3_7/io_i_4_in1[3] cb_3_7/io_i_4_in1[4] cb_3_7/io_i_4_in1[5] cb_3_7/io_i_4_in1[6]
+ cb_3_7/io_i_4_in1[7] cb_3_7/io_i_5_ci cb_3_7/io_i_5_in1[0] cb_3_7/io_i_5_in1[1]
+ cb_3_7/io_i_5_in1[2] cb_3_7/io_i_5_in1[3] cb_3_7/io_i_5_in1[4] cb_3_7/io_i_5_in1[5]
+ cb_3_7/io_i_5_in1[6] cb_3_7/io_i_5_in1[7] cb_3_7/io_i_6_ci cb_3_7/io_i_6_in1[0]
+ cb_3_7/io_i_6_in1[1] cb_3_7/io_i_6_in1[2] cb_3_7/io_i_6_in1[3] cb_3_7/io_i_6_in1[4]
+ cb_3_7/io_i_6_in1[5] cb_3_7/io_i_6_in1[6] cb_3_7/io_i_6_in1[7] cb_3_7/io_i_7_ci
+ cb_3_7/io_i_7_in1[0] cb_3_7/io_i_7_in1[1] cb_3_7/io_i_7_in1[2] cb_3_7/io_i_7_in1[3]
+ cb_3_7/io_i_7_in1[4] cb_3_7/io_i_7_in1[5] cb_3_7/io_i_7_in1[6] cb_3_7/io_i_7_in1[7]
+ cb_3_6/io_vci cb_3_7/io_vci cb_3_6/io_vi cb_3_9/io_we_i cb_3_6/io_wo[0] cb_3_6/io_wo[10]
+ cb_3_6/io_wo[11] cb_3_6/io_wo[12] cb_3_6/io_wo[13] cb_3_6/io_wo[14] cb_3_6/io_wo[15]
+ cb_3_6/io_wo[16] cb_3_6/io_wo[17] cb_3_6/io_wo[18] cb_3_6/io_wo[19] cb_3_6/io_wo[1]
+ cb_3_6/io_wo[20] cb_3_6/io_wo[21] cb_3_6/io_wo[22] cb_3_6/io_wo[23] cb_3_6/io_wo[24]
+ cb_3_6/io_wo[25] cb_3_6/io_wo[26] cb_3_6/io_wo[27] cb_3_6/io_wo[28] cb_3_6/io_wo[29]
+ cb_3_6/io_wo[2] cb_3_6/io_wo[30] cb_3_6/io_wo[31] cb_3_6/io_wo[32] cb_3_6/io_wo[33]
+ cb_3_6/io_wo[34] cb_3_6/io_wo[35] cb_3_6/io_wo[36] cb_3_6/io_wo[37] cb_3_6/io_wo[38]
+ cb_3_6/io_wo[39] cb_3_6/io_wo[3] cb_3_6/io_wo[40] cb_3_6/io_wo[41] cb_3_6/io_wo[42]
+ cb_3_6/io_wo[43] cb_3_6/io_wo[44] cb_3_6/io_wo[45] cb_3_6/io_wo[46] cb_3_6/io_wo[47]
+ cb_3_6/io_wo[48] cb_3_6/io_wo[49] cb_3_6/io_wo[4] cb_3_6/io_wo[50] cb_3_6/io_wo[51]
+ cb_3_6/io_wo[52] cb_3_6/io_wo[53] cb_3_6/io_wo[54] cb_3_6/io_wo[55] cb_3_6/io_wo[56]
+ cb_3_6/io_wo[57] cb_3_6/io_wo[58] cb_3_6/io_wo[59] cb_3_6/io_wo[5] cb_3_6/io_wo[60]
+ cb_3_6/io_wo[61] cb_3_6/io_wo[62] cb_3_6/io_wo[63] cb_3_6/io_wo[6] cb_3_6/io_wo[7]
+ cb_3_6/io_wo[8] cb_3_6/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_1_3 cb_1_9/io_adr_i[0] cb_1_9/io_adr_i[1] cb_1_3/io_cs_i cb_1_9/io_dat_i[0] cb_1_9/io_dat_i[10]
+ cb_1_9/io_dat_i[11] cb_1_9/io_dat_i[12] cb_1_9/io_dat_i[13] cb_1_9/io_dat_i[14]
+ cb_1_9/io_dat_i[15] cb_1_9/io_dat_i[1] cb_1_9/io_dat_i[2] cb_1_9/io_dat_i[3] cb_1_9/io_dat_i[4]
+ cb_1_9/io_dat_i[5] cb_1_9/io_dat_i[6] cb_1_9/io_dat_i[7] cb_1_9/io_dat_i[8] cb_1_9/io_dat_i[9]
+ cb_1_3/io_dat_o[0] cb_1_3/io_dat_o[10] cb_1_3/io_dat_o[11] cb_1_3/io_dat_o[12] cb_1_3/io_dat_o[13]
+ cb_1_3/io_dat_o[14] cb_1_3/io_dat_o[15] cb_1_3/io_dat_o[1] cb_1_3/io_dat_o[2] cb_1_3/io_dat_o[3]
+ cb_1_3/io_dat_o[4] cb_1_3/io_dat_o[5] cb_1_3/io_dat_o[6] cb_1_3/io_dat_o[7] cb_1_3/io_dat_o[8]
+ cb_1_3/io_dat_o[9] cb_1_4/io_wo[0] cb_1_4/io_wo[10] cb_1_4/io_wo[11] cb_1_4/io_wo[12]
+ cb_1_4/io_wo[13] cb_1_4/io_wo[14] cb_1_4/io_wo[15] cb_1_4/io_wo[16] cb_1_4/io_wo[17]
+ cb_1_4/io_wo[18] cb_1_4/io_wo[19] cb_1_4/io_wo[1] cb_1_4/io_wo[20] cb_1_4/io_wo[21]
+ cb_1_4/io_wo[22] cb_1_4/io_wo[23] cb_1_4/io_wo[24] cb_1_4/io_wo[25] cb_1_4/io_wo[26]
+ cb_1_4/io_wo[27] cb_1_4/io_wo[28] cb_1_4/io_wo[29] cb_1_4/io_wo[2] cb_1_4/io_wo[30]
+ cb_1_4/io_wo[31] cb_1_4/io_wo[32] cb_1_4/io_wo[33] cb_1_4/io_wo[34] cb_1_4/io_wo[35]
+ cb_1_4/io_wo[36] cb_1_4/io_wo[37] cb_1_4/io_wo[38] cb_1_4/io_wo[39] cb_1_4/io_wo[3]
+ cb_1_4/io_wo[40] cb_1_4/io_wo[41] cb_1_4/io_wo[42] cb_1_4/io_wo[43] cb_1_4/io_wo[44]
+ cb_1_4/io_wo[45] cb_1_4/io_wo[46] cb_1_4/io_wo[47] cb_1_4/io_wo[48] cb_1_4/io_wo[49]
+ cb_1_4/io_wo[4] cb_1_4/io_wo[50] cb_1_4/io_wo[51] cb_1_4/io_wo[52] cb_1_4/io_wo[53]
+ cb_1_4/io_wo[54] cb_1_4/io_wo[55] cb_1_4/io_wo[56] cb_1_4/io_wo[57] cb_1_4/io_wo[58]
+ cb_1_4/io_wo[59] cb_1_4/io_wo[5] cb_1_4/io_wo[60] cb_1_4/io_wo[61] cb_1_4/io_wo[62]
+ cb_1_4/io_wo[63] cb_1_4/io_wo[6] cb_1_4/io_wo[7] cb_1_4/io_wo[8] cb_1_4/io_wo[9]
+ cb_1_3/io_i_0_ci cb_1_3/io_i_0_in1[0] cb_1_3/io_i_0_in1[1] cb_1_3/io_i_0_in1[2]
+ cb_1_3/io_i_0_in1[3] cb_1_3/io_i_0_in1[4] cb_1_3/io_i_0_in1[5] cb_1_3/io_i_0_in1[6]
+ cb_1_3/io_i_0_in1[7] cb_1_3/io_i_1_ci cb_1_3/io_i_1_in1[0] cb_1_3/io_i_1_in1[1]
+ cb_1_3/io_i_1_in1[2] cb_1_3/io_i_1_in1[3] cb_1_3/io_i_1_in1[4] cb_1_3/io_i_1_in1[5]
+ cb_1_3/io_i_1_in1[6] cb_1_3/io_i_1_in1[7] cb_1_3/io_i_2_ci cb_1_3/io_i_2_in1[0]
+ cb_1_3/io_i_2_in1[1] cb_1_3/io_i_2_in1[2] cb_1_3/io_i_2_in1[3] cb_1_3/io_i_2_in1[4]
+ cb_1_3/io_i_2_in1[5] cb_1_3/io_i_2_in1[6] cb_1_3/io_i_2_in1[7] cb_1_3/io_i_3_ci
+ cb_1_3/io_i_3_in1[0] cb_1_3/io_i_3_in1[1] cb_1_3/io_i_3_in1[2] cb_1_3/io_i_3_in1[3]
+ cb_1_3/io_i_3_in1[4] cb_1_3/io_i_3_in1[5] cb_1_3/io_i_3_in1[6] cb_1_3/io_i_3_in1[7]
+ cb_1_3/io_i_4_ci cb_1_3/io_i_4_in1[0] cb_1_3/io_i_4_in1[1] cb_1_3/io_i_4_in1[2]
+ cb_1_3/io_i_4_in1[3] cb_1_3/io_i_4_in1[4] cb_1_3/io_i_4_in1[5] cb_1_3/io_i_4_in1[6]
+ cb_1_3/io_i_4_in1[7] cb_1_3/io_i_5_ci cb_1_3/io_i_5_in1[0] cb_1_3/io_i_5_in1[1]
+ cb_1_3/io_i_5_in1[2] cb_1_3/io_i_5_in1[3] cb_1_3/io_i_5_in1[4] cb_1_3/io_i_5_in1[5]
+ cb_1_3/io_i_5_in1[6] cb_1_3/io_i_5_in1[7] cb_1_3/io_i_6_ci cb_1_3/io_i_6_in1[0]
+ cb_1_3/io_i_6_in1[1] cb_1_3/io_i_6_in1[2] cb_1_3/io_i_6_in1[3] cb_1_3/io_i_6_in1[4]
+ cb_1_3/io_i_6_in1[5] cb_1_3/io_i_6_in1[6] cb_1_3/io_i_6_in1[7] cb_1_3/io_i_7_ci
+ cb_1_3/io_i_7_in1[0] cb_1_3/io_i_7_in1[1] cb_1_3/io_i_7_in1[2] cb_1_3/io_i_7_in1[3]
+ cb_1_3/io_i_7_in1[4] cb_1_3/io_i_7_in1[5] cb_1_3/io_i_7_in1[6] cb_1_3/io_i_7_in1[7]
+ cb_1_4/io_i_0_ci cb_1_4/io_i_0_in1[0] cb_1_4/io_i_0_in1[1] cb_1_4/io_i_0_in1[2]
+ cb_1_4/io_i_0_in1[3] cb_1_4/io_i_0_in1[4] cb_1_4/io_i_0_in1[5] cb_1_4/io_i_0_in1[6]
+ cb_1_4/io_i_0_in1[7] cb_1_4/io_i_1_ci cb_1_4/io_i_1_in1[0] cb_1_4/io_i_1_in1[1]
+ cb_1_4/io_i_1_in1[2] cb_1_4/io_i_1_in1[3] cb_1_4/io_i_1_in1[4] cb_1_4/io_i_1_in1[5]
+ cb_1_4/io_i_1_in1[6] cb_1_4/io_i_1_in1[7] cb_1_4/io_i_2_ci cb_1_4/io_i_2_in1[0]
+ cb_1_4/io_i_2_in1[1] cb_1_4/io_i_2_in1[2] cb_1_4/io_i_2_in1[3] cb_1_4/io_i_2_in1[4]
+ cb_1_4/io_i_2_in1[5] cb_1_4/io_i_2_in1[6] cb_1_4/io_i_2_in1[7] cb_1_4/io_i_3_ci
+ cb_1_4/io_i_3_in1[0] cb_1_4/io_i_3_in1[1] cb_1_4/io_i_3_in1[2] cb_1_4/io_i_3_in1[3]
+ cb_1_4/io_i_3_in1[4] cb_1_4/io_i_3_in1[5] cb_1_4/io_i_3_in1[6] cb_1_4/io_i_3_in1[7]
+ cb_1_4/io_i_4_ci cb_1_4/io_i_4_in1[0] cb_1_4/io_i_4_in1[1] cb_1_4/io_i_4_in1[2]
+ cb_1_4/io_i_4_in1[3] cb_1_4/io_i_4_in1[4] cb_1_4/io_i_4_in1[5] cb_1_4/io_i_4_in1[6]
+ cb_1_4/io_i_4_in1[7] cb_1_4/io_i_5_ci cb_1_4/io_i_5_in1[0] cb_1_4/io_i_5_in1[1]
+ cb_1_4/io_i_5_in1[2] cb_1_4/io_i_5_in1[3] cb_1_4/io_i_5_in1[4] cb_1_4/io_i_5_in1[5]
+ cb_1_4/io_i_5_in1[6] cb_1_4/io_i_5_in1[7] cb_1_4/io_i_6_ci cb_1_4/io_i_6_in1[0]
+ cb_1_4/io_i_6_in1[1] cb_1_4/io_i_6_in1[2] cb_1_4/io_i_6_in1[3] cb_1_4/io_i_6_in1[4]
+ cb_1_4/io_i_6_in1[5] cb_1_4/io_i_6_in1[6] cb_1_4/io_i_6_in1[7] cb_1_4/io_i_7_ci
+ cb_1_4/io_i_7_in1[0] cb_1_4/io_i_7_in1[1] cb_1_4/io_i_7_in1[2] cb_1_4/io_i_7_in1[3]
+ cb_1_4/io_i_7_in1[4] cb_1_4/io_i_7_in1[5] cb_1_4/io_i_7_in1[6] cb_1_4/io_i_7_in1[7]
+ cb_1_3/io_vci cb_1_4/io_vci cb_1_3/io_vi cb_1_9/io_we_i cb_1_3/io_wo[0] cb_1_3/io_wo[10]
+ cb_1_3/io_wo[11] cb_1_3/io_wo[12] cb_1_3/io_wo[13] cb_1_3/io_wo[14] cb_1_3/io_wo[15]
+ cb_1_3/io_wo[16] cb_1_3/io_wo[17] cb_1_3/io_wo[18] cb_1_3/io_wo[19] cb_1_3/io_wo[1]
+ cb_1_3/io_wo[20] cb_1_3/io_wo[21] cb_1_3/io_wo[22] cb_1_3/io_wo[23] cb_1_3/io_wo[24]
+ cb_1_3/io_wo[25] cb_1_3/io_wo[26] cb_1_3/io_wo[27] cb_1_3/io_wo[28] cb_1_3/io_wo[29]
+ cb_1_3/io_wo[2] cb_1_3/io_wo[30] cb_1_3/io_wo[31] cb_1_3/io_wo[32] cb_1_3/io_wo[33]
+ cb_1_3/io_wo[34] cb_1_3/io_wo[35] cb_1_3/io_wo[36] cb_1_3/io_wo[37] cb_1_3/io_wo[38]
+ cb_1_3/io_wo[39] cb_1_3/io_wo[3] cb_1_3/io_wo[40] cb_1_3/io_wo[41] cb_1_3/io_wo[42]
+ cb_1_3/io_wo[43] cb_1_3/io_wo[44] cb_1_3/io_wo[45] cb_1_3/io_wo[46] cb_1_3/io_wo[47]
+ cb_1_3/io_wo[48] cb_1_3/io_wo[49] cb_1_3/io_wo[4] cb_1_3/io_wo[50] cb_1_3/io_wo[51]
+ cb_1_3/io_wo[52] cb_1_3/io_wo[53] cb_1_3/io_wo[54] cb_1_3/io_wo[55] cb_1_3/io_wo[56]
+ cb_1_3/io_wo[57] cb_1_3/io_wo[58] cb_1_3/io_wo[59] cb_1_3/io_wo[5] cb_1_3/io_wo[60]
+ cb_1_3/io_wo[61] cb_1_3/io_wo[62] cb_1_3/io_wo[63] cb_1_3/io_wo[6] cb_1_3/io_wo[7]
+ cb_1_3/io_wo[8] cb_1_3/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xccon_6 ccon_6/io_ack_o ccon_7/io_adr_i[0] ccon_7/io_adr_i[10] ccon_7/io_adr_i[11]
+ ccon_7/io_adr_i[1] ccon_7/io_adr_i[2] ccon_7/io_adr_i[3] ccon_7/io_adr_i[4] ccon_7/io_adr_i[5]
+ ccon_7/io_adr_i[6] ccon_7/io_adr_i[7] ccon_7/io_adr_i[8] ccon_7/io_adr_i[9] cb_6_9/io_adr_i[0]
+ cb_6_9/io_adr_i[1] cb_6_0/io_cs_i cb_6_1/io_cs_i cb_6_10/io_cs_i cb_6_2/io_cs_i
+ cb_6_3/io_cs_i cb_6_4/io_cs_i cb_6_5/io_cs_i cb_6_6/io_cs_i cb_6_7/io_cs_i cb_6_8/io_cs_i
+ cb_6_9/io_cs_i cb_6_9/io_dat_i[0] cb_6_9/io_dat_i[10] cb_6_9/io_dat_i[11] cb_6_9/io_dat_i[12]
+ cb_6_9/io_dat_i[13] cb_6_9/io_dat_i[14] cb_6_9/io_dat_i[15] cb_6_9/io_dat_i[1] cb_6_9/io_dat_i[2]
+ cb_6_9/io_dat_i[3] cb_6_9/io_dat_i[4] cb_6_9/io_dat_i[5] cb_6_9/io_dat_i[6] cb_6_9/io_dat_i[7]
+ cb_6_9/io_dat_i[8] cb_6_9/io_dat_i[9] cb_6_0/io_dat_o[0] cb_6_0/io_dat_o[10] cb_6_0/io_dat_o[11]
+ cb_6_0/io_dat_o[12] cb_6_0/io_dat_o[13] cb_6_0/io_dat_o[14] cb_6_0/io_dat_o[15]
+ cb_6_0/io_dat_o[1] cb_6_0/io_dat_o[2] cb_6_0/io_dat_o[3] cb_6_0/io_dat_o[4] cb_6_0/io_dat_o[5]
+ cb_6_0/io_dat_o[6] cb_6_0/io_dat_o[7] cb_6_0/io_dat_o[8] cb_6_0/io_dat_o[9] cb_6_10/io_dat_o[0]
+ cb_6_10/io_dat_o[10] cb_6_10/io_dat_o[11] cb_6_10/io_dat_o[12] cb_6_10/io_dat_o[13]
+ cb_6_10/io_dat_o[14] cb_6_10/io_dat_o[15] cb_6_10/io_dat_o[1] cb_6_10/io_dat_o[2]
+ cb_6_10/io_dat_o[3] cb_6_10/io_dat_o[4] cb_6_10/io_dat_o[5] cb_6_10/io_dat_o[6]
+ cb_6_10/io_dat_o[7] cb_6_10/io_dat_o[8] cb_6_10/io_dat_o[9] cb_6_1/io_dat_o[0] cb_6_1/io_dat_o[10]
+ cb_6_1/io_dat_o[11] cb_6_1/io_dat_o[12] cb_6_1/io_dat_o[13] cb_6_1/io_dat_o[14]
+ cb_6_1/io_dat_o[15] cb_6_1/io_dat_o[1] cb_6_1/io_dat_o[2] cb_6_1/io_dat_o[3] cb_6_1/io_dat_o[4]
+ cb_6_1/io_dat_o[5] cb_6_1/io_dat_o[6] cb_6_1/io_dat_o[7] cb_6_1/io_dat_o[8] cb_6_1/io_dat_o[9]
+ cb_6_2/io_dat_o[0] cb_6_2/io_dat_o[10] cb_6_2/io_dat_o[11] cb_6_2/io_dat_o[12] cb_6_2/io_dat_o[13]
+ cb_6_2/io_dat_o[14] cb_6_2/io_dat_o[15] cb_6_2/io_dat_o[1] cb_6_2/io_dat_o[2] cb_6_2/io_dat_o[3]
+ cb_6_2/io_dat_o[4] cb_6_2/io_dat_o[5] cb_6_2/io_dat_o[6] cb_6_2/io_dat_o[7] cb_6_2/io_dat_o[8]
+ cb_6_2/io_dat_o[9] cb_6_3/io_dat_o[0] cb_6_3/io_dat_o[10] cb_6_3/io_dat_o[11] cb_6_3/io_dat_o[12]
+ cb_6_3/io_dat_o[13] cb_6_3/io_dat_o[14] cb_6_3/io_dat_o[15] cb_6_3/io_dat_o[1] cb_6_3/io_dat_o[2]
+ cb_6_3/io_dat_o[3] cb_6_3/io_dat_o[4] cb_6_3/io_dat_o[5] cb_6_3/io_dat_o[6] cb_6_3/io_dat_o[7]
+ cb_6_3/io_dat_o[8] cb_6_3/io_dat_o[9] cb_6_4/io_dat_o[0] cb_6_4/io_dat_o[10] cb_6_4/io_dat_o[11]
+ cb_6_4/io_dat_o[12] cb_6_4/io_dat_o[13] cb_6_4/io_dat_o[14] cb_6_4/io_dat_o[15]
+ cb_6_4/io_dat_o[1] cb_6_4/io_dat_o[2] cb_6_4/io_dat_o[3] cb_6_4/io_dat_o[4] cb_6_4/io_dat_o[5]
+ cb_6_4/io_dat_o[6] cb_6_4/io_dat_o[7] cb_6_4/io_dat_o[8] cb_6_4/io_dat_o[9] cb_6_5/io_dat_o[0]
+ cb_6_5/io_dat_o[10] cb_6_5/io_dat_o[11] cb_6_5/io_dat_o[12] cb_6_5/io_dat_o[13]
+ cb_6_5/io_dat_o[14] cb_6_5/io_dat_o[15] cb_6_5/io_dat_o[1] cb_6_5/io_dat_o[2] cb_6_5/io_dat_o[3]
+ cb_6_5/io_dat_o[4] cb_6_5/io_dat_o[5] cb_6_5/io_dat_o[6] cb_6_5/io_dat_o[7] cb_6_5/io_dat_o[8]
+ cb_6_5/io_dat_o[9] cb_6_6/io_dat_o[0] cb_6_6/io_dat_o[10] cb_6_6/io_dat_o[11] cb_6_6/io_dat_o[12]
+ cb_6_6/io_dat_o[13] cb_6_6/io_dat_o[14] cb_6_6/io_dat_o[15] cb_6_6/io_dat_o[1] cb_6_6/io_dat_o[2]
+ cb_6_6/io_dat_o[3] cb_6_6/io_dat_o[4] cb_6_6/io_dat_o[5] cb_6_6/io_dat_o[6] cb_6_6/io_dat_o[7]
+ cb_6_6/io_dat_o[8] cb_6_6/io_dat_o[9] cb_6_7/io_dat_o[0] cb_6_7/io_dat_o[10] cb_6_7/io_dat_o[11]
+ cb_6_7/io_dat_o[12] cb_6_7/io_dat_o[13] cb_6_7/io_dat_o[14] cb_6_7/io_dat_o[15]
+ cb_6_7/io_dat_o[1] cb_6_7/io_dat_o[2] cb_6_7/io_dat_o[3] cb_6_7/io_dat_o[4] cb_6_7/io_dat_o[5]
+ cb_6_7/io_dat_o[6] cb_6_7/io_dat_o[7] cb_6_7/io_dat_o[8] cb_6_7/io_dat_o[9] cb_6_8/io_dat_o[0]
+ cb_6_8/io_dat_o[10] cb_6_8/io_dat_o[11] cb_6_8/io_dat_o[12] cb_6_8/io_dat_o[13]
+ cb_6_8/io_dat_o[14] cb_6_8/io_dat_o[15] cb_6_8/io_dat_o[1] cb_6_8/io_dat_o[2] cb_6_8/io_dat_o[3]
+ cb_6_8/io_dat_o[4] cb_6_8/io_dat_o[5] cb_6_8/io_dat_o[6] cb_6_8/io_dat_o[7] cb_6_8/io_dat_o[8]
+ cb_6_8/io_dat_o[9] cb_6_9/io_dat_o[0] cb_6_9/io_dat_o[10] cb_6_9/io_dat_o[11] cb_6_9/io_dat_o[12]
+ cb_6_9/io_dat_o[13] cb_6_9/io_dat_o[14] cb_6_9/io_dat_o[15] cb_6_9/io_dat_o[1] cb_6_9/io_dat_o[2]
+ cb_6_9/io_dat_o[3] cb_6_9/io_dat_o[4] cb_6_9/io_dat_o[5] cb_6_9/io_dat_o[6] cb_6_9/io_dat_o[7]
+ cb_6_9/io_dat_o[8] cb_6_9/io_dat_o[9] cb_6_9/io_we_i ccon_6/io_cs_i ccon_7/io_dat_i[0]
+ ccon_7/io_dat_i[10] ccon_7/io_dat_i[11] ccon_7/io_dat_i[12] ccon_7/io_dat_i[13]
+ ccon_7/io_dat_i[14] ccon_7/io_dat_i[15] ccon_7/io_dat_i[16] ccon_7/io_dat_i[17]
+ ccon_7/io_dat_i[18] ccon_7/io_dat_i[19] ccon_7/io_dat_i[1] ccon_7/io_dat_i[20] ccon_7/io_dat_i[21]
+ ccon_7/io_dat_i[22] ccon_7/io_dat_i[23] ccon_7/io_dat_i[24] ccon_7/io_dat_i[25]
+ ccon_7/io_dat_i[26] ccon_7/io_dat_i[27] ccon_7/io_dat_i[28] ccon_7/io_dat_i[29]
+ ccon_7/io_dat_i[2] ccon_7/io_dat_i[30] ccon_7/io_dat_i[31] ccon_7/io_dat_i[3] ccon_7/io_dat_i[4]
+ ccon_7/io_dat_i[5] ccon_7/io_dat_i[6] ccon_7/io_dat_i[7] ccon_7/io_dat_i[8] ccon_7/io_dat_i[9]
+ ccon_6/io_dat_o[0] ccon_6/io_dat_o[10] ccon_6/io_dat_o[11] ccon_6/io_dat_o[12] ccon_6/io_dat_o[13]
+ ccon_6/io_dat_o[14] ccon_6/io_dat_o[15] ccon_6/io_dat_o[16] ccon_6/io_dat_o[17]
+ ccon_6/io_dat_o[18] ccon_6/io_dat_o[19] ccon_6/io_dat_o[1] ccon_6/io_dat_o[20] ccon_6/io_dat_o[21]
+ ccon_6/io_dat_o[22] ccon_6/io_dat_o[23] ccon_6/io_dat_o[24] ccon_6/io_dat_o[25]
+ ccon_6/io_dat_o[26] ccon_6/io_dat_o[27] ccon_6/io_dat_o[28] ccon_6/io_dat_o[29]
+ ccon_6/io_dat_o[2] ccon_6/io_dat_o[30] ccon_6/io_dat_o[31] ccon_6/io_dat_o[3] ccon_6/io_dat_o[4]
+ ccon_6/io_dat_o[5] ccon_6/io_dat_o[6] ccon_6/io_dat_o[7] ccon_6/io_dat_o[8] ccon_6/io_dat_o[9]
+ cb_6_0/io_wo[0] cb_6_0/io_wo[10] cb_6_0/io_wo[11] cb_6_0/io_wo[12] cb_6_0/io_wo[13]
+ cb_6_0/io_wo[14] cb_6_0/io_wo[15] cb_6_0/io_wo[16] cb_6_0/io_wo[17] cb_6_0/io_wo[18]
+ cb_6_0/io_wo[19] cb_6_0/io_wo[1] cb_6_0/io_wo[20] cb_6_0/io_wo[21] cb_6_0/io_wo[22]
+ cb_6_0/io_wo[23] cb_6_0/io_wo[24] cb_6_0/io_wo[25] cb_6_0/io_wo[26] cb_6_0/io_wo[27]
+ cb_6_0/io_wo[28] cb_6_0/io_wo[29] cb_6_0/io_wo[2] cb_6_0/io_wo[30] cb_6_0/io_wo[31]
+ cb_6_0/io_wo[32] cb_6_0/io_wo[33] cb_6_0/io_wo[34] cb_6_0/io_wo[35] cb_6_0/io_wo[36]
+ cb_6_0/io_wo[37] cb_6_0/io_wo[38] cb_6_0/io_wo[39] cb_6_0/io_wo[3] cb_6_0/io_wo[40]
+ cb_6_0/io_wo[41] cb_6_0/io_wo[42] cb_6_0/io_wo[43] cb_6_0/io_wo[44] cb_6_0/io_wo[45]
+ cb_6_0/io_wo[46] cb_6_0/io_wo[47] cb_6_0/io_wo[48] cb_6_0/io_wo[49] cb_6_0/io_wo[4]
+ cb_6_0/io_wo[50] cb_6_0/io_wo[51] cb_6_0/io_wo[52] cb_6_0/io_wo[53] cb_6_0/io_wo[54]
+ cb_6_0/io_wo[55] cb_6_0/io_wo[56] cb_6_0/io_wo[57] cb_6_0/io_wo[58] cb_6_0/io_wo[59]
+ cb_6_0/io_wo[5] cb_6_0/io_wo[60] cb_6_0/io_wo[61] cb_6_0/io_wo[62] cb_6_0/io_wo[63]
+ cb_6_0/io_wo[6] cb_6_0/io_wo[7] cb_6_0/io_wo[8] cb_6_0/io_wo[9] icon/dsi[0] icon/dsi[1]
+ icon/dsi[2] icon/dsi[3] icon/dsi[4] icon/dsi[5] icon/dsi[6] icon/dsi[7] ccon_6/io_dsi_o
+ ccon_6/io_irq cb_6_0/io_vi cb_6_10/io_vi cb_6_1/io_vi cb_6_2/io_vi cb_6_3/io_vi
+ cb_6_4/io_vi cb_6_5/io_vi cb_6_6/io_vi cb_6_7/io_vi cb_6_8/io_vi cb_6_9/io_vi ccon_7/io_we_i
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_con
Xcb_3_7 cb_3_9/io_adr_i[0] cb_3_9/io_adr_i[1] cb_3_7/io_cs_i cb_3_9/io_dat_i[0] cb_3_9/io_dat_i[10]
+ cb_3_9/io_dat_i[11] cb_3_9/io_dat_i[12] cb_3_9/io_dat_i[13] cb_3_9/io_dat_i[14]
+ cb_3_9/io_dat_i[15] cb_3_9/io_dat_i[1] cb_3_9/io_dat_i[2] cb_3_9/io_dat_i[3] cb_3_9/io_dat_i[4]
+ cb_3_9/io_dat_i[5] cb_3_9/io_dat_i[6] cb_3_9/io_dat_i[7] cb_3_9/io_dat_i[8] cb_3_9/io_dat_i[9]
+ cb_3_7/io_dat_o[0] cb_3_7/io_dat_o[10] cb_3_7/io_dat_o[11] cb_3_7/io_dat_o[12] cb_3_7/io_dat_o[13]
+ cb_3_7/io_dat_o[14] cb_3_7/io_dat_o[15] cb_3_7/io_dat_o[1] cb_3_7/io_dat_o[2] cb_3_7/io_dat_o[3]
+ cb_3_7/io_dat_o[4] cb_3_7/io_dat_o[5] cb_3_7/io_dat_o[6] cb_3_7/io_dat_o[7] cb_3_7/io_dat_o[8]
+ cb_3_7/io_dat_o[9] cb_3_8/io_wo[0] cb_3_8/io_wo[10] cb_3_8/io_wo[11] cb_3_8/io_wo[12]
+ cb_3_8/io_wo[13] cb_3_8/io_wo[14] cb_3_8/io_wo[15] cb_3_8/io_wo[16] cb_3_8/io_wo[17]
+ cb_3_8/io_wo[18] cb_3_8/io_wo[19] cb_3_8/io_wo[1] cb_3_8/io_wo[20] cb_3_8/io_wo[21]
+ cb_3_8/io_wo[22] cb_3_8/io_wo[23] cb_3_8/io_wo[24] cb_3_8/io_wo[25] cb_3_8/io_wo[26]
+ cb_3_8/io_wo[27] cb_3_8/io_wo[28] cb_3_8/io_wo[29] cb_3_8/io_wo[2] cb_3_8/io_wo[30]
+ cb_3_8/io_wo[31] cb_3_8/io_wo[32] cb_3_8/io_wo[33] cb_3_8/io_wo[34] cb_3_8/io_wo[35]
+ cb_3_8/io_wo[36] cb_3_8/io_wo[37] cb_3_8/io_wo[38] cb_3_8/io_wo[39] cb_3_8/io_wo[3]
+ cb_3_8/io_wo[40] cb_3_8/io_wo[41] cb_3_8/io_wo[42] cb_3_8/io_wo[43] cb_3_8/io_wo[44]
+ cb_3_8/io_wo[45] cb_3_8/io_wo[46] cb_3_8/io_wo[47] cb_3_8/io_wo[48] cb_3_8/io_wo[49]
+ cb_3_8/io_wo[4] cb_3_8/io_wo[50] cb_3_8/io_wo[51] cb_3_8/io_wo[52] cb_3_8/io_wo[53]
+ cb_3_8/io_wo[54] cb_3_8/io_wo[55] cb_3_8/io_wo[56] cb_3_8/io_wo[57] cb_3_8/io_wo[58]
+ cb_3_8/io_wo[59] cb_3_8/io_wo[5] cb_3_8/io_wo[60] cb_3_8/io_wo[61] cb_3_8/io_wo[62]
+ cb_3_8/io_wo[63] cb_3_8/io_wo[6] cb_3_8/io_wo[7] cb_3_8/io_wo[8] cb_3_8/io_wo[9]
+ cb_3_7/io_i_0_ci cb_3_7/io_i_0_in1[0] cb_3_7/io_i_0_in1[1] cb_3_7/io_i_0_in1[2]
+ cb_3_7/io_i_0_in1[3] cb_3_7/io_i_0_in1[4] cb_3_7/io_i_0_in1[5] cb_3_7/io_i_0_in1[6]
+ cb_3_7/io_i_0_in1[7] cb_3_7/io_i_1_ci cb_3_7/io_i_1_in1[0] cb_3_7/io_i_1_in1[1]
+ cb_3_7/io_i_1_in1[2] cb_3_7/io_i_1_in1[3] cb_3_7/io_i_1_in1[4] cb_3_7/io_i_1_in1[5]
+ cb_3_7/io_i_1_in1[6] cb_3_7/io_i_1_in1[7] cb_3_7/io_i_2_ci cb_3_7/io_i_2_in1[0]
+ cb_3_7/io_i_2_in1[1] cb_3_7/io_i_2_in1[2] cb_3_7/io_i_2_in1[3] cb_3_7/io_i_2_in1[4]
+ cb_3_7/io_i_2_in1[5] cb_3_7/io_i_2_in1[6] cb_3_7/io_i_2_in1[7] cb_3_7/io_i_3_ci
+ cb_3_7/io_i_3_in1[0] cb_3_7/io_i_3_in1[1] cb_3_7/io_i_3_in1[2] cb_3_7/io_i_3_in1[3]
+ cb_3_7/io_i_3_in1[4] cb_3_7/io_i_3_in1[5] cb_3_7/io_i_3_in1[6] cb_3_7/io_i_3_in1[7]
+ cb_3_7/io_i_4_ci cb_3_7/io_i_4_in1[0] cb_3_7/io_i_4_in1[1] cb_3_7/io_i_4_in1[2]
+ cb_3_7/io_i_4_in1[3] cb_3_7/io_i_4_in1[4] cb_3_7/io_i_4_in1[5] cb_3_7/io_i_4_in1[6]
+ cb_3_7/io_i_4_in1[7] cb_3_7/io_i_5_ci cb_3_7/io_i_5_in1[0] cb_3_7/io_i_5_in1[1]
+ cb_3_7/io_i_5_in1[2] cb_3_7/io_i_5_in1[3] cb_3_7/io_i_5_in1[4] cb_3_7/io_i_5_in1[5]
+ cb_3_7/io_i_5_in1[6] cb_3_7/io_i_5_in1[7] cb_3_7/io_i_6_ci cb_3_7/io_i_6_in1[0]
+ cb_3_7/io_i_6_in1[1] cb_3_7/io_i_6_in1[2] cb_3_7/io_i_6_in1[3] cb_3_7/io_i_6_in1[4]
+ cb_3_7/io_i_6_in1[5] cb_3_7/io_i_6_in1[6] cb_3_7/io_i_6_in1[7] cb_3_7/io_i_7_ci
+ cb_3_7/io_i_7_in1[0] cb_3_7/io_i_7_in1[1] cb_3_7/io_i_7_in1[2] cb_3_7/io_i_7_in1[3]
+ cb_3_7/io_i_7_in1[4] cb_3_7/io_i_7_in1[5] cb_3_7/io_i_7_in1[6] cb_3_7/io_i_7_in1[7]
+ cb_3_8/io_i_0_ci cb_3_8/io_i_0_in1[0] cb_3_8/io_i_0_in1[1] cb_3_8/io_i_0_in1[2]
+ cb_3_8/io_i_0_in1[3] cb_3_8/io_i_0_in1[4] cb_3_8/io_i_0_in1[5] cb_3_8/io_i_0_in1[6]
+ cb_3_8/io_i_0_in1[7] cb_3_8/io_i_1_ci cb_3_8/io_i_1_in1[0] cb_3_8/io_i_1_in1[1]
+ cb_3_8/io_i_1_in1[2] cb_3_8/io_i_1_in1[3] cb_3_8/io_i_1_in1[4] cb_3_8/io_i_1_in1[5]
+ cb_3_8/io_i_1_in1[6] cb_3_8/io_i_1_in1[7] cb_3_8/io_i_2_ci cb_3_8/io_i_2_in1[0]
+ cb_3_8/io_i_2_in1[1] cb_3_8/io_i_2_in1[2] cb_3_8/io_i_2_in1[3] cb_3_8/io_i_2_in1[4]
+ cb_3_8/io_i_2_in1[5] cb_3_8/io_i_2_in1[6] cb_3_8/io_i_2_in1[7] cb_3_8/io_i_3_ci
+ cb_3_8/io_i_3_in1[0] cb_3_8/io_i_3_in1[1] cb_3_8/io_i_3_in1[2] cb_3_8/io_i_3_in1[3]
+ cb_3_8/io_i_3_in1[4] cb_3_8/io_i_3_in1[5] cb_3_8/io_i_3_in1[6] cb_3_8/io_i_3_in1[7]
+ cb_3_8/io_i_4_ci cb_3_8/io_i_4_in1[0] cb_3_8/io_i_4_in1[1] cb_3_8/io_i_4_in1[2]
+ cb_3_8/io_i_4_in1[3] cb_3_8/io_i_4_in1[4] cb_3_8/io_i_4_in1[5] cb_3_8/io_i_4_in1[6]
+ cb_3_8/io_i_4_in1[7] cb_3_8/io_i_5_ci cb_3_8/io_i_5_in1[0] cb_3_8/io_i_5_in1[1]
+ cb_3_8/io_i_5_in1[2] cb_3_8/io_i_5_in1[3] cb_3_8/io_i_5_in1[4] cb_3_8/io_i_5_in1[5]
+ cb_3_8/io_i_5_in1[6] cb_3_8/io_i_5_in1[7] cb_3_8/io_i_6_ci cb_3_8/io_i_6_in1[0]
+ cb_3_8/io_i_6_in1[1] cb_3_8/io_i_6_in1[2] cb_3_8/io_i_6_in1[3] cb_3_8/io_i_6_in1[4]
+ cb_3_8/io_i_6_in1[5] cb_3_8/io_i_6_in1[6] cb_3_8/io_i_6_in1[7] cb_3_8/io_i_7_ci
+ cb_3_8/io_i_7_in1[0] cb_3_8/io_i_7_in1[1] cb_3_8/io_i_7_in1[2] cb_3_8/io_i_7_in1[3]
+ cb_3_8/io_i_7_in1[4] cb_3_8/io_i_7_in1[5] cb_3_8/io_i_7_in1[6] cb_3_8/io_i_7_in1[7]
+ cb_3_7/io_vci cb_3_8/io_vci cb_3_7/io_vi cb_3_9/io_we_i cb_3_7/io_wo[0] cb_3_7/io_wo[10]
+ cb_3_7/io_wo[11] cb_3_7/io_wo[12] cb_3_7/io_wo[13] cb_3_7/io_wo[14] cb_3_7/io_wo[15]
+ cb_3_7/io_wo[16] cb_3_7/io_wo[17] cb_3_7/io_wo[18] cb_3_7/io_wo[19] cb_3_7/io_wo[1]
+ cb_3_7/io_wo[20] cb_3_7/io_wo[21] cb_3_7/io_wo[22] cb_3_7/io_wo[23] cb_3_7/io_wo[24]
+ cb_3_7/io_wo[25] cb_3_7/io_wo[26] cb_3_7/io_wo[27] cb_3_7/io_wo[28] cb_3_7/io_wo[29]
+ cb_3_7/io_wo[2] cb_3_7/io_wo[30] cb_3_7/io_wo[31] cb_3_7/io_wo[32] cb_3_7/io_wo[33]
+ cb_3_7/io_wo[34] cb_3_7/io_wo[35] cb_3_7/io_wo[36] cb_3_7/io_wo[37] cb_3_7/io_wo[38]
+ cb_3_7/io_wo[39] cb_3_7/io_wo[3] cb_3_7/io_wo[40] cb_3_7/io_wo[41] cb_3_7/io_wo[42]
+ cb_3_7/io_wo[43] cb_3_7/io_wo[44] cb_3_7/io_wo[45] cb_3_7/io_wo[46] cb_3_7/io_wo[47]
+ cb_3_7/io_wo[48] cb_3_7/io_wo[49] cb_3_7/io_wo[4] cb_3_7/io_wo[50] cb_3_7/io_wo[51]
+ cb_3_7/io_wo[52] cb_3_7/io_wo[53] cb_3_7/io_wo[54] cb_3_7/io_wo[55] cb_3_7/io_wo[56]
+ cb_3_7/io_wo[57] cb_3_7/io_wo[58] cb_3_7/io_wo[59] cb_3_7/io_wo[5] cb_3_7/io_wo[60]
+ cb_3_7/io_wo[61] cb_3_7/io_wo[62] cb_3_7/io_wo[63] cb_3_7/io_wo[6] cb_3_7/io_wo[7]
+ cb_3_7/io_wo[8] cb_3_7/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_1_4 cb_1_9/io_adr_i[0] cb_1_9/io_adr_i[1] cb_1_4/io_cs_i cb_1_9/io_dat_i[0] cb_1_9/io_dat_i[10]
+ cb_1_9/io_dat_i[11] cb_1_9/io_dat_i[12] cb_1_9/io_dat_i[13] cb_1_9/io_dat_i[14]
+ cb_1_9/io_dat_i[15] cb_1_9/io_dat_i[1] cb_1_9/io_dat_i[2] cb_1_9/io_dat_i[3] cb_1_9/io_dat_i[4]
+ cb_1_9/io_dat_i[5] cb_1_9/io_dat_i[6] cb_1_9/io_dat_i[7] cb_1_9/io_dat_i[8] cb_1_9/io_dat_i[9]
+ cb_1_4/io_dat_o[0] cb_1_4/io_dat_o[10] cb_1_4/io_dat_o[11] cb_1_4/io_dat_o[12] cb_1_4/io_dat_o[13]
+ cb_1_4/io_dat_o[14] cb_1_4/io_dat_o[15] cb_1_4/io_dat_o[1] cb_1_4/io_dat_o[2] cb_1_4/io_dat_o[3]
+ cb_1_4/io_dat_o[4] cb_1_4/io_dat_o[5] cb_1_4/io_dat_o[6] cb_1_4/io_dat_o[7] cb_1_4/io_dat_o[8]
+ cb_1_4/io_dat_o[9] cb_1_5/io_wo[0] cb_1_5/io_wo[10] cb_1_5/io_wo[11] cb_1_5/io_wo[12]
+ cb_1_5/io_wo[13] cb_1_5/io_wo[14] cb_1_5/io_wo[15] cb_1_5/io_wo[16] cb_1_5/io_wo[17]
+ cb_1_5/io_wo[18] cb_1_5/io_wo[19] cb_1_5/io_wo[1] cb_1_5/io_wo[20] cb_1_5/io_wo[21]
+ cb_1_5/io_wo[22] cb_1_5/io_wo[23] cb_1_5/io_wo[24] cb_1_5/io_wo[25] cb_1_5/io_wo[26]
+ cb_1_5/io_wo[27] cb_1_5/io_wo[28] cb_1_5/io_wo[29] cb_1_5/io_wo[2] cb_1_5/io_wo[30]
+ cb_1_5/io_wo[31] cb_1_5/io_wo[32] cb_1_5/io_wo[33] cb_1_5/io_wo[34] cb_1_5/io_wo[35]
+ cb_1_5/io_wo[36] cb_1_5/io_wo[37] cb_1_5/io_wo[38] cb_1_5/io_wo[39] cb_1_5/io_wo[3]
+ cb_1_5/io_wo[40] cb_1_5/io_wo[41] cb_1_5/io_wo[42] cb_1_5/io_wo[43] cb_1_5/io_wo[44]
+ cb_1_5/io_wo[45] cb_1_5/io_wo[46] cb_1_5/io_wo[47] cb_1_5/io_wo[48] cb_1_5/io_wo[49]
+ cb_1_5/io_wo[4] cb_1_5/io_wo[50] cb_1_5/io_wo[51] cb_1_5/io_wo[52] cb_1_5/io_wo[53]
+ cb_1_5/io_wo[54] cb_1_5/io_wo[55] cb_1_5/io_wo[56] cb_1_5/io_wo[57] cb_1_5/io_wo[58]
+ cb_1_5/io_wo[59] cb_1_5/io_wo[5] cb_1_5/io_wo[60] cb_1_5/io_wo[61] cb_1_5/io_wo[62]
+ cb_1_5/io_wo[63] cb_1_5/io_wo[6] cb_1_5/io_wo[7] cb_1_5/io_wo[8] cb_1_5/io_wo[9]
+ cb_1_4/io_i_0_ci cb_1_4/io_i_0_in1[0] cb_1_4/io_i_0_in1[1] cb_1_4/io_i_0_in1[2]
+ cb_1_4/io_i_0_in1[3] cb_1_4/io_i_0_in1[4] cb_1_4/io_i_0_in1[5] cb_1_4/io_i_0_in1[6]
+ cb_1_4/io_i_0_in1[7] cb_1_4/io_i_1_ci cb_1_4/io_i_1_in1[0] cb_1_4/io_i_1_in1[1]
+ cb_1_4/io_i_1_in1[2] cb_1_4/io_i_1_in1[3] cb_1_4/io_i_1_in1[4] cb_1_4/io_i_1_in1[5]
+ cb_1_4/io_i_1_in1[6] cb_1_4/io_i_1_in1[7] cb_1_4/io_i_2_ci cb_1_4/io_i_2_in1[0]
+ cb_1_4/io_i_2_in1[1] cb_1_4/io_i_2_in1[2] cb_1_4/io_i_2_in1[3] cb_1_4/io_i_2_in1[4]
+ cb_1_4/io_i_2_in1[5] cb_1_4/io_i_2_in1[6] cb_1_4/io_i_2_in1[7] cb_1_4/io_i_3_ci
+ cb_1_4/io_i_3_in1[0] cb_1_4/io_i_3_in1[1] cb_1_4/io_i_3_in1[2] cb_1_4/io_i_3_in1[3]
+ cb_1_4/io_i_3_in1[4] cb_1_4/io_i_3_in1[5] cb_1_4/io_i_3_in1[6] cb_1_4/io_i_3_in1[7]
+ cb_1_4/io_i_4_ci cb_1_4/io_i_4_in1[0] cb_1_4/io_i_4_in1[1] cb_1_4/io_i_4_in1[2]
+ cb_1_4/io_i_4_in1[3] cb_1_4/io_i_4_in1[4] cb_1_4/io_i_4_in1[5] cb_1_4/io_i_4_in1[6]
+ cb_1_4/io_i_4_in1[7] cb_1_4/io_i_5_ci cb_1_4/io_i_5_in1[0] cb_1_4/io_i_5_in1[1]
+ cb_1_4/io_i_5_in1[2] cb_1_4/io_i_5_in1[3] cb_1_4/io_i_5_in1[4] cb_1_4/io_i_5_in1[5]
+ cb_1_4/io_i_5_in1[6] cb_1_4/io_i_5_in1[7] cb_1_4/io_i_6_ci cb_1_4/io_i_6_in1[0]
+ cb_1_4/io_i_6_in1[1] cb_1_4/io_i_6_in1[2] cb_1_4/io_i_6_in1[3] cb_1_4/io_i_6_in1[4]
+ cb_1_4/io_i_6_in1[5] cb_1_4/io_i_6_in1[6] cb_1_4/io_i_6_in1[7] cb_1_4/io_i_7_ci
+ cb_1_4/io_i_7_in1[0] cb_1_4/io_i_7_in1[1] cb_1_4/io_i_7_in1[2] cb_1_4/io_i_7_in1[3]
+ cb_1_4/io_i_7_in1[4] cb_1_4/io_i_7_in1[5] cb_1_4/io_i_7_in1[6] cb_1_4/io_i_7_in1[7]
+ cb_1_5/io_i_0_ci cb_1_5/io_i_0_in1[0] cb_1_5/io_i_0_in1[1] cb_1_5/io_i_0_in1[2]
+ cb_1_5/io_i_0_in1[3] cb_1_5/io_i_0_in1[4] cb_1_5/io_i_0_in1[5] cb_1_5/io_i_0_in1[6]
+ cb_1_5/io_i_0_in1[7] cb_1_5/io_i_1_ci cb_1_5/io_i_1_in1[0] cb_1_5/io_i_1_in1[1]
+ cb_1_5/io_i_1_in1[2] cb_1_5/io_i_1_in1[3] cb_1_5/io_i_1_in1[4] cb_1_5/io_i_1_in1[5]
+ cb_1_5/io_i_1_in1[6] cb_1_5/io_i_1_in1[7] cb_1_5/io_i_2_ci cb_1_5/io_i_2_in1[0]
+ cb_1_5/io_i_2_in1[1] cb_1_5/io_i_2_in1[2] cb_1_5/io_i_2_in1[3] cb_1_5/io_i_2_in1[4]
+ cb_1_5/io_i_2_in1[5] cb_1_5/io_i_2_in1[6] cb_1_5/io_i_2_in1[7] cb_1_5/io_i_3_ci
+ cb_1_5/io_i_3_in1[0] cb_1_5/io_i_3_in1[1] cb_1_5/io_i_3_in1[2] cb_1_5/io_i_3_in1[3]
+ cb_1_5/io_i_3_in1[4] cb_1_5/io_i_3_in1[5] cb_1_5/io_i_3_in1[6] cb_1_5/io_i_3_in1[7]
+ cb_1_5/io_i_4_ci cb_1_5/io_i_4_in1[0] cb_1_5/io_i_4_in1[1] cb_1_5/io_i_4_in1[2]
+ cb_1_5/io_i_4_in1[3] cb_1_5/io_i_4_in1[4] cb_1_5/io_i_4_in1[5] cb_1_5/io_i_4_in1[6]
+ cb_1_5/io_i_4_in1[7] cb_1_5/io_i_5_ci cb_1_5/io_i_5_in1[0] cb_1_5/io_i_5_in1[1]
+ cb_1_5/io_i_5_in1[2] cb_1_5/io_i_5_in1[3] cb_1_5/io_i_5_in1[4] cb_1_5/io_i_5_in1[5]
+ cb_1_5/io_i_5_in1[6] cb_1_5/io_i_5_in1[7] cb_1_5/io_i_6_ci cb_1_5/io_i_6_in1[0]
+ cb_1_5/io_i_6_in1[1] cb_1_5/io_i_6_in1[2] cb_1_5/io_i_6_in1[3] cb_1_5/io_i_6_in1[4]
+ cb_1_5/io_i_6_in1[5] cb_1_5/io_i_6_in1[6] cb_1_5/io_i_6_in1[7] cb_1_5/io_i_7_ci
+ cb_1_5/io_i_7_in1[0] cb_1_5/io_i_7_in1[1] cb_1_5/io_i_7_in1[2] cb_1_5/io_i_7_in1[3]
+ cb_1_5/io_i_7_in1[4] cb_1_5/io_i_7_in1[5] cb_1_5/io_i_7_in1[6] cb_1_5/io_i_7_in1[7]
+ cb_1_4/io_vci cb_1_5/io_vci cb_1_4/io_vi cb_1_9/io_we_i cb_1_4/io_wo[0] cb_1_4/io_wo[10]
+ cb_1_4/io_wo[11] cb_1_4/io_wo[12] cb_1_4/io_wo[13] cb_1_4/io_wo[14] cb_1_4/io_wo[15]
+ cb_1_4/io_wo[16] cb_1_4/io_wo[17] cb_1_4/io_wo[18] cb_1_4/io_wo[19] cb_1_4/io_wo[1]
+ cb_1_4/io_wo[20] cb_1_4/io_wo[21] cb_1_4/io_wo[22] cb_1_4/io_wo[23] cb_1_4/io_wo[24]
+ cb_1_4/io_wo[25] cb_1_4/io_wo[26] cb_1_4/io_wo[27] cb_1_4/io_wo[28] cb_1_4/io_wo[29]
+ cb_1_4/io_wo[2] cb_1_4/io_wo[30] cb_1_4/io_wo[31] cb_1_4/io_wo[32] cb_1_4/io_wo[33]
+ cb_1_4/io_wo[34] cb_1_4/io_wo[35] cb_1_4/io_wo[36] cb_1_4/io_wo[37] cb_1_4/io_wo[38]
+ cb_1_4/io_wo[39] cb_1_4/io_wo[3] cb_1_4/io_wo[40] cb_1_4/io_wo[41] cb_1_4/io_wo[42]
+ cb_1_4/io_wo[43] cb_1_4/io_wo[44] cb_1_4/io_wo[45] cb_1_4/io_wo[46] cb_1_4/io_wo[47]
+ cb_1_4/io_wo[48] cb_1_4/io_wo[49] cb_1_4/io_wo[4] cb_1_4/io_wo[50] cb_1_4/io_wo[51]
+ cb_1_4/io_wo[52] cb_1_4/io_wo[53] cb_1_4/io_wo[54] cb_1_4/io_wo[55] cb_1_4/io_wo[56]
+ cb_1_4/io_wo[57] cb_1_4/io_wo[58] cb_1_4/io_wo[59] cb_1_4/io_wo[5] cb_1_4/io_wo[60]
+ cb_1_4/io_wo[61] cb_1_4/io_wo[62] cb_1_4/io_wo[63] cb_1_4/io_wo[6] cb_1_4/io_wo[7]
+ cb_1_4/io_wo[8] cb_1_4/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xccon_7 ccon_7/io_ack_o ccon_7/io_adr_i[0] ccon_7/io_adr_i[10] ccon_7/io_adr_i[11]
+ ccon_7/io_adr_i[1] ccon_7/io_adr_i[2] ccon_7/io_adr_i[3] ccon_7/io_adr_i[4] ccon_7/io_adr_i[5]
+ ccon_7/io_adr_i[6] ccon_7/io_adr_i[7] ccon_7/io_adr_i[8] ccon_7/io_adr_i[9] cb_7_9/io_adr_i[0]
+ cb_7_9/io_adr_i[1] cb_7_0/io_cs_i cb_7_1/io_cs_i cb_7_10/io_cs_i cb_7_2/io_cs_i
+ cb_7_3/io_cs_i cb_7_4/io_cs_i cb_7_5/io_cs_i cb_7_6/io_cs_i cb_7_7/io_cs_i cb_7_8/io_cs_i
+ cb_7_9/io_cs_i cb_7_9/io_dat_i[0] cb_7_9/io_dat_i[10] cb_7_9/io_dat_i[11] cb_7_9/io_dat_i[12]
+ cb_7_9/io_dat_i[13] cb_7_9/io_dat_i[14] cb_7_9/io_dat_i[15] cb_7_9/io_dat_i[1] cb_7_9/io_dat_i[2]
+ cb_7_9/io_dat_i[3] cb_7_9/io_dat_i[4] cb_7_9/io_dat_i[5] cb_7_9/io_dat_i[6] cb_7_9/io_dat_i[7]
+ cb_7_9/io_dat_i[8] cb_7_9/io_dat_i[9] cb_7_0/io_dat_o[0] cb_7_0/io_dat_o[10] cb_7_0/io_dat_o[11]
+ cb_7_0/io_dat_o[12] cb_7_0/io_dat_o[13] cb_7_0/io_dat_o[14] cb_7_0/io_dat_o[15]
+ cb_7_0/io_dat_o[1] cb_7_0/io_dat_o[2] cb_7_0/io_dat_o[3] cb_7_0/io_dat_o[4] cb_7_0/io_dat_o[5]
+ cb_7_0/io_dat_o[6] cb_7_0/io_dat_o[7] cb_7_0/io_dat_o[8] cb_7_0/io_dat_o[9] cb_7_10/io_dat_o[0]
+ cb_7_10/io_dat_o[10] cb_7_10/io_dat_o[11] cb_7_10/io_dat_o[12] cb_7_10/io_dat_o[13]
+ cb_7_10/io_dat_o[14] cb_7_10/io_dat_o[15] cb_7_10/io_dat_o[1] cb_7_10/io_dat_o[2]
+ cb_7_10/io_dat_o[3] cb_7_10/io_dat_o[4] cb_7_10/io_dat_o[5] cb_7_10/io_dat_o[6]
+ cb_7_10/io_dat_o[7] cb_7_10/io_dat_o[8] cb_7_10/io_dat_o[9] cb_7_1/io_dat_o[0] cb_7_1/io_dat_o[10]
+ cb_7_1/io_dat_o[11] cb_7_1/io_dat_o[12] cb_7_1/io_dat_o[13] cb_7_1/io_dat_o[14]
+ cb_7_1/io_dat_o[15] cb_7_1/io_dat_o[1] cb_7_1/io_dat_o[2] cb_7_1/io_dat_o[3] cb_7_1/io_dat_o[4]
+ cb_7_1/io_dat_o[5] cb_7_1/io_dat_o[6] cb_7_1/io_dat_o[7] cb_7_1/io_dat_o[8] cb_7_1/io_dat_o[9]
+ cb_7_2/io_dat_o[0] cb_7_2/io_dat_o[10] cb_7_2/io_dat_o[11] cb_7_2/io_dat_o[12] cb_7_2/io_dat_o[13]
+ cb_7_2/io_dat_o[14] cb_7_2/io_dat_o[15] cb_7_2/io_dat_o[1] cb_7_2/io_dat_o[2] cb_7_2/io_dat_o[3]
+ cb_7_2/io_dat_o[4] cb_7_2/io_dat_o[5] cb_7_2/io_dat_o[6] cb_7_2/io_dat_o[7] cb_7_2/io_dat_o[8]
+ cb_7_2/io_dat_o[9] cb_7_3/io_dat_o[0] cb_7_3/io_dat_o[10] cb_7_3/io_dat_o[11] cb_7_3/io_dat_o[12]
+ cb_7_3/io_dat_o[13] cb_7_3/io_dat_o[14] cb_7_3/io_dat_o[15] cb_7_3/io_dat_o[1] cb_7_3/io_dat_o[2]
+ cb_7_3/io_dat_o[3] cb_7_3/io_dat_o[4] cb_7_3/io_dat_o[5] cb_7_3/io_dat_o[6] cb_7_3/io_dat_o[7]
+ cb_7_3/io_dat_o[8] cb_7_3/io_dat_o[9] cb_7_4/io_dat_o[0] cb_7_4/io_dat_o[10] cb_7_4/io_dat_o[11]
+ cb_7_4/io_dat_o[12] cb_7_4/io_dat_o[13] cb_7_4/io_dat_o[14] cb_7_4/io_dat_o[15]
+ cb_7_4/io_dat_o[1] cb_7_4/io_dat_o[2] cb_7_4/io_dat_o[3] cb_7_4/io_dat_o[4] cb_7_4/io_dat_o[5]
+ cb_7_4/io_dat_o[6] cb_7_4/io_dat_o[7] cb_7_4/io_dat_o[8] cb_7_4/io_dat_o[9] cb_7_5/io_dat_o[0]
+ cb_7_5/io_dat_o[10] cb_7_5/io_dat_o[11] cb_7_5/io_dat_o[12] cb_7_5/io_dat_o[13]
+ cb_7_5/io_dat_o[14] cb_7_5/io_dat_o[15] cb_7_5/io_dat_o[1] cb_7_5/io_dat_o[2] cb_7_5/io_dat_o[3]
+ cb_7_5/io_dat_o[4] cb_7_5/io_dat_o[5] cb_7_5/io_dat_o[6] cb_7_5/io_dat_o[7] cb_7_5/io_dat_o[8]
+ cb_7_5/io_dat_o[9] cb_7_6/io_dat_o[0] cb_7_6/io_dat_o[10] cb_7_6/io_dat_o[11] cb_7_6/io_dat_o[12]
+ cb_7_6/io_dat_o[13] cb_7_6/io_dat_o[14] cb_7_6/io_dat_o[15] cb_7_6/io_dat_o[1] cb_7_6/io_dat_o[2]
+ cb_7_6/io_dat_o[3] cb_7_6/io_dat_o[4] cb_7_6/io_dat_o[5] cb_7_6/io_dat_o[6] cb_7_6/io_dat_o[7]
+ cb_7_6/io_dat_o[8] cb_7_6/io_dat_o[9] cb_7_7/io_dat_o[0] cb_7_7/io_dat_o[10] cb_7_7/io_dat_o[11]
+ cb_7_7/io_dat_o[12] cb_7_7/io_dat_o[13] cb_7_7/io_dat_o[14] cb_7_7/io_dat_o[15]
+ cb_7_7/io_dat_o[1] cb_7_7/io_dat_o[2] cb_7_7/io_dat_o[3] cb_7_7/io_dat_o[4] cb_7_7/io_dat_o[5]
+ cb_7_7/io_dat_o[6] cb_7_7/io_dat_o[7] cb_7_7/io_dat_o[8] cb_7_7/io_dat_o[9] cb_7_8/io_dat_o[0]
+ cb_7_8/io_dat_o[10] cb_7_8/io_dat_o[11] cb_7_8/io_dat_o[12] cb_7_8/io_dat_o[13]
+ cb_7_8/io_dat_o[14] cb_7_8/io_dat_o[15] cb_7_8/io_dat_o[1] cb_7_8/io_dat_o[2] cb_7_8/io_dat_o[3]
+ cb_7_8/io_dat_o[4] cb_7_8/io_dat_o[5] cb_7_8/io_dat_o[6] cb_7_8/io_dat_o[7] cb_7_8/io_dat_o[8]
+ cb_7_8/io_dat_o[9] cb_7_9/io_dat_o[0] cb_7_9/io_dat_o[10] cb_7_9/io_dat_o[11] cb_7_9/io_dat_o[12]
+ cb_7_9/io_dat_o[13] cb_7_9/io_dat_o[14] cb_7_9/io_dat_o[15] cb_7_9/io_dat_o[1] cb_7_9/io_dat_o[2]
+ cb_7_9/io_dat_o[3] cb_7_9/io_dat_o[4] cb_7_9/io_dat_o[5] cb_7_9/io_dat_o[6] cb_7_9/io_dat_o[7]
+ cb_7_9/io_dat_o[8] cb_7_9/io_dat_o[9] cb_7_9/io_we_i ccon_7/io_cs_i ccon_7/io_dat_i[0]
+ ccon_7/io_dat_i[10] ccon_7/io_dat_i[11] ccon_7/io_dat_i[12] ccon_7/io_dat_i[13]
+ ccon_7/io_dat_i[14] ccon_7/io_dat_i[15] ccon_7/io_dat_i[16] ccon_7/io_dat_i[17]
+ ccon_7/io_dat_i[18] ccon_7/io_dat_i[19] ccon_7/io_dat_i[1] ccon_7/io_dat_i[20] ccon_7/io_dat_i[21]
+ ccon_7/io_dat_i[22] ccon_7/io_dat_i[23] ccon_7/io_dat_i[24] ccon_7/io_dat_i[25]
+ ccon_7/io_dat_i[26] ccon_7/io_dat_i[27] ccon_7/io_dat_i[28] ccon_7/io_dat_i[29]
+ ccon_7/io_dat_i[2] ccon_7/io_dat_i[30] ccon_7/io_dat_i[31] ccon_7/io_dat_i[3] ccon_7/io_dat_i[4]
+ ccon_7/io_dat_i[5] ccon_7/io_dat_i[6] ccon_7/io_dat_i[7] ccon_7/io_dat_i[8] ccon_7/io_dat_i[9]
+ ccon_7/io_dat_o[0] ccon_7/io_dat_o[10] ccon_7/io_dat_o[11] ccon_7/io_dat_o[12] ccon_7/io_dat_o[13]
+ ccon_7/io_dat_o[14] ccon_7/io_dat_o[15] ccon_7/io_dat_o[16] ccon_7/io_dat_o[17]
+ ccon_7/io_dat_o[18] ccon_7/io_dat_o[19] ccon_7/io_dat_o[1] ccon_7/io_dat_o[20] ccon_7/io_dat_o[21]
+ ccon_7/io_dat_o[22] ccon_7/io_dat_o[23] ccon_7/io_dat_o[24] ccon_7/io_dat_o[25]
+ ccon_7/io_dat_o[26] ccon_7/io_dat_o[27] ccon_7/io_dat_o[28] ccon_7/io_dat_o[29]
+ ccon_7/io_dat_o[2] ccon_7/io_dat_o[30] ccon_7/io_dat_o[31] ccon_7/io_dat_o[3] ccon_7/io_dat_o[4]
+ ccon_7/io_dat_o[5] ccon_7/io_dat_o[6] ccon_7/io_dat_o[7] ccon_7/io_dat_o[8] ccon_7/io_dat_o[9]
+ cb_7_0/io_wo[0] cb_7_0/io_wo[10] cb_7_0/io_wo[11] cb_7_0/io_wo[12] cb_7_0/io_wo[13]
+ cb_7_0/io_wo[14] cb_7_0/io_wo[15] cb_7_0/io_wo[16] cb_7_0/io_wo[17] cb_7_0/io_wo[18]
+ cb_7_0/io_wo[19] cb_7_0/io_wo[1] cb_7_0/io_wo[20] cb_7_0/io_wo[21] cb_7_0/io_wo[22]
+ cb_7_0/io_wo[23] cb_7_0/io_wo[24] cb_7_0/io_wo[25] cb_7_0/io_wo[26] cb_7_0/io_wo[27]
+ cb_7_0/io_wo[28] cb_7_0/io_wo[29] cb_7_0/io_wo[2] cb_7_0/io_wo[30] cb_7_0/io_wo[31]
+ cb_7_0/io_wo[32] cb_7_0/io_wo[33] cb_7_0/io_wo[34] cb_7_0/io_wo[35] cb_7_0/io_wo[36]
+ cb_7_0/io_wo[37] cb_7_0/io_wo[38] cb_7_0/io_wo[39] cb_7_0/io_wo[3] cb_7_0/io_wo[40]
+ cb_7_0/io_wo[41] cb_7_0/io_wo[42] cb_7_0/io_wo[43] cb_7_0/io_wo[44] cb_7_0/io_wo[45]
+ cb_7_0/io_wo[46] cb_7_0/io_wo[47] cb_7_0/io_wo[48] cb_7_0/io_wo[49] cb_7_0/io_wo[4]
+ cb_7_0/io_wo[50] cb_7_0/io_wo[51] cb_7_0/io_wo[52] cb_7_0/io_wo[53] cb_7_0/io_wo[54]
+ cb_7_0/io_wo[55] cb_7_0/io_wo[56] cb_7_0/io_wo[57] cb_7_0/io_wo[58] cb_7_0/io_wo[59]
+ cb_7_0/io_wo[5] cb_7_0/io_wo[60] cb_7_0/io_wo[61] cb_7_0/io_wo[62] cb_7_0/io_wo[63]
+ cb_7_0/io_wo[6] cb_7_0/io_wo[7] cb_7_0/io_wo[8] cb_7_0/io_wo[9] icon/dsi[0] icon/dsi[1]
+ icon/dsi[2] icon/dsi[3] icon/dsi[4] icon/dsi[5] icon/dsi[6] icon/dsi[7] ccon_7/io_dsi_o
+ ccon_7/io_irq cb_7_0/io_vi cb_7_10/io_vi cb_7_1/io_vi cb_7_2/io_vi cb_7_3/io_vi
+ cb_7_4/io_vi cb_7_5/io_vi cb_7_6/io_vi cb_7_7/io_vi cb_7_8/io_vi cb_7_9/io_vi ccon_7/io_we_i
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_con
Xcb_3_8 cb_3_9/io_adr_i[0] cb_3_9/io_adr_i[1] cb_3_8/io_cs_i cb_3_9/io_dat_i[0] cb_3_9/io_dat_i[10]
+ cb_3_9/io_dat_i[11] cb_3_9/io_dat_i[12] cb_3_9/io_dat_i[13] cb_3_9/io_dat_i[14]
+ cb_3_9/io_dat_i[15] cb_3_9/io_dat_i[1] cb_3_9/io_dat_i[2] cb_3_9/io_dat_i[3] cb_3_9/io_dat_i[4]
+ cb_3_9/io_dat_i[5] cb_3_9/io_dat_i[6] cb_3_9/io_dat_i[7] cb_3_9/io_dat_i[8] cb_3_9/io_dat_i[9]
+ cb_3_8/io_dat_o[0] cb_3_8/io_dat_o[10] cb_3_8/io_dat_o[11] cb_3_8/io_dat_o[12] cb_3_8/io_dat_o[13]
+ cb_3_8/io_dat_o[14] cb_3_8/io_dat_o[15] cb_3_8/io_dat_o[1] cb_3_8/io_dat_o[2] cb_3_8/io_dat_o[3]
+ cb_3_8/io_dat_o[4] cb_3_8/io_dat_o[5] cb_3_8/io_dat_o[6] cb_3_8/io_dat_o[7] cb_3_8/io_dat_o[8]
+ cb_3_8/io_dat_o[9] cb_3_9/io_wo[0] cb_3_9/io_wo[10] cb_3_9/io_wo[11] cb_3_9/io_wo[12]
+ cb_3_9/io_wo[13] cb_3_9/io_wo[14] cb_3_9/io_wo[15] cb_3_9/io_wo[16] cb_3_9/io_wo[17]
+ cb_3_9/io_wo[18] cb_3_9/io_wo[19] cb_3_9/io_wo[1] cb_3_9/io_wo[20] cb_3_9/io_wo[21]
+ cb_3_9/io_wo[22] cb_3_9/io_wo[23] cb_3_9/io_wo[24] cb_3_9/io_wo[25] cb_3_9/io_wo[26]
+ cb_3_9/io_wo[27] cb_3_9/io_wo[28] cb_3_9/io_wo[29] cb_3_9/io_wo[2] cb_3_9/io_wo[30]
+ cb_3_9/io_wo[31] cb_3_9/io_wo[32] cb_3_9/io_wo[33] cb_3_9/io_wo[34] cb_3_9/io_wo[35]
+ cb_3_9/io_wo[36] cb_3_9/io_wo[37] cb_3_9/io_wo[38] cb_3_9/io_wo[39] cb_3_9/io_wo[3]
+ cb_3_9/io_wo[40] cb_3_9/io_wo[41] cb_3_9/io_wo[42] cb_3_9/io_wo[43] cb_3_9/io_wo[44]
+ cb_3_9/io_wo[45] cb_3_9/io_wo[46] cb_3_9/io_wo[47] cb_3_9/io_wo[48] cb_3_9/io_wo[49]
+ cb_3_9/io_wo[4] cb_3_9/io_wo[50] cb_3_9/io_wo[51] cb_3_9/io_wo[52] cb_3_9/io_wo[53]
+ cb_3_9/io_wo[54] cb_3_9/io_wo[55] cb_3_9/io_wo[56] cb_3_9/io_wo[57] cb_3_9/io_wo[58]
+ cb_3_9/io_wo[59] cb_3_9/io_wo[5] cb_3_9/io_wo[60] cb_3_9/io_wo[61] cb_3_9/io_wo[62]
+ cb_3_9/io_wo[63] cb_3_9/io_wo[6] cb_3_9/io_wo[7] cb_3_9/io_wo[8] cb_3_9/io_wo[9]
+ cb_3_8/io_i_0_ci cb_3_8/io_i_0_in1[0] cb_3_8/io_i_0_in1[1] cb_3_8/io_i_0_in1[2]
+ cb_3_8/io_i_0_in1[3] cb_3_8/io_i_0_in1[4] cb_3_8/io_i_0_in1[5] cb_3_8/io_i_0_in1[6]
+ cb_3_8/io_i_0_in1[7] cb_3_8/io_i_1_ci cb_3_8/io_i_1_in1[0] cb_3_8/io_i_1_in1[1]
+ cb_3_8/io_i_1_in1[2] cb_3_8/io_i_1_in1[3] cb_3_8/io_i_1_in1[4] cb_3_8/io_i_1_in1[5]
+ cb_3_8/io_i_1_in1[6] cb_3_8/io_i_1_in1[7] cb_3_8/io_i_2_ci cb_3_8/io_i_2_in1[0]
+ cb_3_8/io_i_2_in1[1] cb_3_8/io_i_2_in1[2] cb_3_8/io_i_2_in1[3] cb_3_8/io_i_2_in1[4]
+ cb_3_8/io_i_2_in1[5] cb_3_8/io_i_2_in1[6] cb_3_8/io_i_2_in1[7] cb_3_8/io_i_3_ci
+ cb_3_8/io_i_3_in1[0] cb_3_8/io_i_3_in1[1] cb_3_8/io_i_3_in1[2] cb_3_8/io_i_3_in1[3]
+ cb_3_8/io_i_3_in1[4] cb_3_8/io_i_3_in1[5] cb_3_8/io_i_3_in1[6] cb_3_8/io_i_3_in1[7]
+ cb_3_8/io_i_4_ci cb_3_8/io_i_4_in1[0] cb_3_8/io_i_4_in1[1] cb_3_8/io_i_4_in1[2]
+ cb_3_8/io_i_4_in1[3] cb_3_8/io_i_4_in1[4] cb_3_8/io_i_4_in1[5] cb_3_8/io_i_4_in1[6]
+ cb_3_8/io_i_4_in1[7] cb_3_8/io_i_5_ci cb_3_8/io_i_5_in1[0] cb_3_8/io_i_5_in1[1]
+ cb_3_8/io_i_5_in1[2] cb_3_8/io_i_5_in1[3] cb_3_8/io_i_5_in1[4] cb_3_8/io_i_5_in1[5]
+ cb_3_8/io_i_5_in1[6] cb_3_8/io_i_5_in1[7] cb_3_8/io_i_6_ci cb_3_8/io_i_6_in1[0]
+ cb_3_8/io_i_6_in1[1] cb_3_8/io_i_6_in1[2] cb_3_8/io_i_6_in1[3] cb_3_8/io_i_6_in1[4]
+ cb_3_8/io_i_6_in1[5] cb_3_8/io_i_6_in1[6] cb_3_8/io_i_6_in1[7] cb_3_8/io_i_7_ci
+ cb_3_8/io_i_7_in1[0] cb_3_8/io_i_7_in1[1] cb_3_8/io_i_7_in1[2] cb_3_8/io_i_7_in1[3]
+ cb_3_8/io_i_7_in1[4] cb_3_8/io_i_7_in1[5] cb_3_8/io_i_7_in1[6] cb_3_8/io_i_7_in1[7]
+ cb_3_9/io_i_0_ci cb_3_9/io_i_0_in1[0] cb_3_9/io_i_0_in1[1] cb_3_9/io_i_0_in1[2]
+ cb_3_9/io_i_0_in1[3] cb_3_9/io_i_0_in1[4] cb_3_9/io_i_0_in1[5] cb_3_9/io_i_0_in1[6]
+ cb_3_9/io_i_0_in1[7] cb_3_9/io_i_1_ci cb_3_9/io_i_1_in1[0] cb_3_9/io_i_1_in1[1]
+ cb_3_9/io_i_1_in1[2] cb_3_9/io_i_1_in1[3] cb_3_9/io_i_1_in1[4] cb_3_9/io_i_1_in1[5]
+ cb_3_9/io_i_1_in1[6] cb_3_9/io_i_1_in1[7] cb_3_9/io_i_2_ci cb_3_9/io_i_2_in1[0]
+ cb_3_9/io_i_2_in1[1] cb_3_9/io_i_2_in1[2] cb_3_9/io_i_2_in1[3] cb_3_9/io_i_2_in1[4]
+ cb_3_9/io_i_2_in1[5] cb_3_9/io_i_2_in1[6] cb_3_9/io_i_2_in1[7] cb_3_9/io_i_3_ci
+ cb_3_9/io_i_3_in1[0] cb_3_9/io_i_3_in1[1] cb_3_9/io_i_3_in1[2] cb_3_9/io_i_3_in1[3]
+ cb_3_9/io_i_3_in1[4] cb_3_9/io_i_3_in1[5] cb_3_9/io_i_3_in1[6] cb_3_9/io_i_3_in1[7]
+ cb_3_9/io_i_4_ci cb_3_9/io_i_4_in1[0] cb_3_9/io_i_4_in1[1] cb_3_9/io_i_4_in1[2]
+ cb_3_9/io_i_4_in1[3] cb_3_9/io_i_4_in1[4] cb_3_9/io_i_4_in1[5] cb_3_9/io_i_4_in1[6]
+ cb_3_9/io_i_4_in1[7] cb_3_9/io_i_5_ci cb_3_9/io_i_5_in1[0] cb_3_9/io_i_5_in1[1]
+ cb_3_9/io_i_5_in1[2] cb_3_9/io_i_5_in1[3] cb_3_9/io_i_5_in1[4] cb_3_9/io_i_5_in1[5]
+ cb_3_9/io_i_5_in1[6] cb_3_9/io_i_5_in1[7] cb_3_9/io_i_6_ci cb_3_9/io_i_6_in1[0]
+ cb_3_9/io_i_6_in1[1] cb_3_9/io_i_6_in1[2] cb_3_9/io_i_6_in1[3] cb_3_9/io_i_6_in1[4]
+ cb_3_9/io_i_6_in1[5] cb_3_9/io_i_6_in1[6] cb_3_9/io_i_6_in1[7] cb_3_9/io_i_7_ci
+ cb_3_9/io_i_7_in1[0] cb_3_9/io_i_7_in1[1] cb_3_9/io_i_7_in1[2] cb_3_9/io_i_7_in1[3]
+ cb_3_9/io_i_7_in1[4] cb_3_9/io_i_7_in1[5] cb_3_9/io_i_7_in1[6] cb_3_9/io_i_7_in1[7]
+ cb_3_8/io_vci cb_3_9/io_vci cb_3_8/io_vi cb_3_9/io_we_i cb_3_8/io_wo[0] cb_3_8/io_wo[10]
+ cb_3_8/io_wo[11] cb_3_8/io_wo[12] cb_3_8/io_wo[13] cb_3_8/io_wo[14] cb_3_8/io_wo[15]
+ cb_3_8/io_wo[16] cb_3_8/io_wo[17] cb_3_8/io_wo[18] cb_3_8/io_wo[19] cb_3_8/io_wo[1]
+ cb_3_8/io_wo[20] cb_3_8/io_wo[21] cb_3_8/io_wo[22] cb_3_8/io_wo[23] cb_3_8/io_wo[24]
+ cb_3_8/io_wo[25] cb_3_8/io_wo[26] cb_3_8/io_wo[27] cb_3_8/io_wo[28] cb_3_8/io_wo[29]
+ cb_3_8/io_wo[2] cb_3_8/io_wo[30] cb_3_8/io_wo[31] cb_3_8/io_wo[32] cb_3_8/io_wo[33]
+ cb_3_8/io_wo[34] cb_3_8/io_wo[35] cb_3_8/io_wo[36] cb_3_8/io_wo[37] cb_3_8/io_wo[38]
+ cb_3_8/io_wo[39] cb_3_8/io_wo[3] cb_3_8/io_wo[40] cb_3_8/io_wo[41] cb_3_8/io_wo[42]
+ cb_3_8/io_wo[43] cb_3_8/io_wo[44] cb_3_8/io_wo[45] cb_3_8/io_wo[46] cb_3_8/io_wo[47]
+ cb_3_8/io_wo[48] cb_3_8/io_wo[49] cb_3_8/io_wo[4] cb_3_8/io_wo[50] cb_3_8/io_wo[51]
+ cb_3_8/io_wo[52] cb_3_8/io_wo[53] cb_3_8/io_wo[54] cb_3_8/io_wo[55] cb_3_8/io_wo[56]
+ cb_3_8/io_wo[57] cb_3_8/io_wo[58] cb_3_8/io_wo[59] cb_3_8/io_wo[5] cb_3_8/io_wo[60]
+ cb_3_8/io_wo[61] cb_3_8/io_wo[62] cb_3_8/io_wo[63] cb_3_8/io_wo[6] cb_3_8/io_wo[7]
+ cb_3_8/io_wo[8] cb_3_8/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_1_5 cb_1_9/io_adr_i[0] cb_1_9/io_adr_i[1] cb_1_5/io_cs_i cb_1_9/io_dat_i[0] cb_1_9/io_dat_i[10]
+ cb_1_9/io_dat_i[11] cb_1_9/io_dat_i[12] cb_1_9/io_dat_i[13] cb_1_9/io_dat_i[14]
+ cb_1_9/io_dat_i[15] cb_1_9/io_dat_i[1] cb_1_9/io_dat_i[2] cb_1_9/io_dat_i[3] cb_1_9/io_dat_i[4]
+ cb_1_9/io_dat_i[5] cb_1_9/io_dat_i[6] cb_1_9/io_dat_i[7] cb_1_9/io_dat_i[8] cb_1_9/io_dat_i[9]
+ cb_1_5/io_dat_o[0] cb_1_5/io_dat_o[10] cb_1_5/io_dat_o[11] cb_1_5/io_dat_o[12] cb_1_5/io_dat_o[13]
+ cb_1_5/io_dat_o[14] cb_1_5/io_dat_o[15] cb_1_5/io_dat_o[1] cb_1_5/io_dat_o[2] cb_1_5/io_dat_o[3]
+ cb_1_5/io_dat_o[4] cb_1_5/io_dat_o[5] cb_1_5/io_dat_o[6] cb_1_5/io_dat_o[7] cb_1_5/io_dat_o[8]
+ cb_1_5/io_dat_o[9] cb_1_6/io_wo[0] cb_1_6/io_wo[10] cb_1_6/io_wo[11] cb_1_6/io_wo[12]
+ cb_1_6/io_wo[13] cb_1_6/io_wo[14] cb_1_6/io_wo[15] cb_1_6/io_wo[16] cb_1_6/io_wo[17]
+ cb_1_6/io_wo[18] cb_1_6/io_wo[19] cb_1_6/io_wo[1] cb_1_6/io_wo[20] cb_1_6/io_wo[21]
+ cb_1_6/io_wo[22] cb_1_6/io_wo[23] cb_1_6/io_wo[24] cb_1_6/io_wo[25] cb_1_6/io_wo[26]
+ cb_1_6/io_wo[27] cb_1_6/io_wo[28] cb_1_6/io_wo[29] cb_1_6/io_wo[2] cb_1_6/io_wo[30]
+ cb_1_6/io_wo[31] cb_1_6/io_wo[32] cb_1_6/io_wo[33] cb_1_6/io_wo[34] cb_1_6/io_wo[35]
+ cb_1_6/io_wo[36] cb_1_6/io_wo[37] cb_1_6/io_wo[38] cb_1_6/io_wo[39] cb_1_6/io_wo[3]
+ cb_1_6/io_wo[40] cb_1_6/io_wo[41] cb_1_6/io_wo[42] cb_1_6/io_wo[43] cb_1_6/io_wo[44]
+ cb_1_6/io_wo[45] cb_1_6/io_wo[46] cb_1_6/io_wo[47] cb_1_6/io_wo[48] cb_1_6/io_wo[49]
+ cb_1_6/io_wo[4] cb_1_6/io_wo[50] cb_1_6/io_wo[51] cb_1_6/io_wo[52] cb_1_6/io_wo[53]
+ cb_1_6/io_wo[54] cb_1_6/io_wo[55] cb_1_6/io_wo[56] cb_1_6/io_wo[57] cb_1_6/io_wo[58]
+ cb_1_6/io_wo[59] cb_1_6/io_wo[5] cb_1_6/io_wo[60] cb_1_6/io_wo[61] cb_1_6/io_wo[62]
+ cb_1_6/io_wo[63] cb_1_6/io_wo[6] cb_1_6/io_wo[7] cb_1_6/io_wo[8] cb_1_6/io_wo[9]
+ cb_1_5/io_i_0_ci cb_1_5/io_i_0_in1[0] cb_1_5/io_i_0_in1[1] cb_1_5/io_i_0_in1[2]
+ cb_1_5/io_i_0_in1[3] cb_1_5/io_i_0_in1[4] cb_1_5/io_i_0_in1[5] cb_1_5/io_i_0_in1[6]
+ cb_1_5/io_i_0_in1[7] cb_1_5/io_i_1_ci cb_1_5/io_i_1_in1[0] cb_1_5/io_i_1_in1[1]
+ cb_1_5/io_i_1_in1[2] cb_1_5/io_i_1_in1[3] cb_1_5/io_i_1_in1[4] cb_1_5/io_i_1_in1[5]
+ cb_1_5/io_i_1_in1[6] cb_1_5/io_i_1_in1[7] cb_1_5/io_i_2_ci cb_1_5/io_i_2_in1[0]
+ cb_1_5/io_i_2_in1[1] cb_1_5/io_i_2_in1[2] cb_1_5/io_i_2_in1[3] cb_1_5/io_i_2_in1[4]
+ cb_1_5/io_i_2_in1[5] cb_1_5/io_i_2_in1[6] cb_1_5/io_i_2_in1[7] cb_1_5/io_i_3_ci
+ cb_1_5/io_i_3_in1[0] cb_1_5/io_i_3_in1[1] cb_1_5/io_i_3_in1[2] cb_1_5/io_i_3_in1[3]
+ cb_1_5/io_i_3_in1[4] cb_1_5/io_i_3_in1[5] cb_1_5/io_i_3_in1[6] cb_1_5/io_i_3_in1[7]
+ cb_1_5/io_i_4_ci cb_1_5/io_i_4_in1[0] cb_1_5/io_i_4_in1[1] cb_1_5/io_i_4_in1[2]
+ cb_1_5/io_i_4_in1[3] cb_1_5/io_i_4_in1[4] cb_1_5/io_i_4_in1[5] cb_1_5/io_i_4_in1[6]
+ cb_1_5/io_i_4_in1[7] cb_1_5/io_i_5_ci cb_1_5/io_i_5_in1[0] cb_1_5/io_i_5_in1[1]
+ cb_1_5/io_i_5_in1[2] cb_1_5/io_i_5_in1[3] cb_1_5/io_i_5_in1[4] cb_1_5/io_i_5_in1[5]
+ cb_1_5/io_i_5_in1[6] cb_1_5/io_i_5_in1[7] cb_1_5/io_i_6_ci cb_1_5/io_i_6_in1[0]
+ cb_1_5/io_i_6_in1[1] cb_1_5/io_i_6_in1[2] cb_1_5/io_i_6_in1[3] cb_1_5/io_i_6_in1[4]
+ cb_1_5/io_i_6_in1[5] cb_1_5/io_i_6_in1[6] cb_1_5/io_i_6_in1[7] cb_1_5/io_i_7_ci
+ cb_1_5/io_i_7_in1[0] cb_1_5/io_i_7_in1[1] cb_1_5/io_i_7_in1[2] cb_1_5/io_i_7_in1[3]
+ cb_1_5/io_i_7_in1[4] cb_1_5/io_i_7_in1[5] cb_1_5/io_i_7_in1[6] cb_1_5/io_i_7_in1[7]
+ cb_1_6/io_i_0_ci cb_1_6/io_i_0_in1[0] cb_1_6/io_i_0_in1[1] cb_1_6/io_i_0_in1[2]
+ cb_1_6/io_i_0_in1[3] cb_1_6/io_i_0_in1[4] cb_1_6/io_i_0_in1[5] cb_1_6/io_i_0_in1[6]
+ cb_1_6/io_i_0_in1[7] cb_1_6/io_i_1_ci cb_1_6/io_i_1_in1[0] cb_1_6/io_i_1_in1[1]
+ cb_1_6/io_i_1_in1[2] cb_1_6/io_i_1_in1[3] cb_1_6/io_i_1_in1[4] cb_1_6/io_i_1_in1[5]
+ cb_1_6/io_i_1_in1[6] cb_1_6/io_i_1_in1[7] cb_1_6/io_i_2_ci cb_1_6/io_i_2_in1[0]
+ cb_1_6/io_i_2_in1[1] cb_1_6/io_i_2_in1[2] cb_1_6/io_i_2_in1[3] cb_1_6/io_i_2_in1[4]
+ cb_1_6/io_i_2_in1[5] cb_1_6/io_i_2_in1[6] cb_1_6/io_i_2_in1[7] cb_1_6/io_i_3_ci
+ cb_1_6/io_i_3_in1[0] cb_1_6/io_i_3_in1[1] cb_1_6/io_i_3_in1[2] cb_1_6/io_i_3_in1[3]
+ cb_1_6/io_i_3_in1[4] cb_1_6/io_i_3_in1[5] cb_1_6/io_i_3_in1[6] cb_1_6/io_i_3_in1[7]
+ cb_1_6/io_i_4_ci cb_1_6/io_i_4_in1[0] cb_1_6/io_i_4_in1[1] cb_1_6/io_i_4_in1[2]
+ cb_1_6/io_i_4_in1[3] cb_1_6/io_i_4_in1[4] cb_1_6/io_i_4_in1[5] cb_1_6/io_i_4_in1[6]
+ cb_1_6/io_i_4_in1[7] cb_1_6/io_i_5_ci cb_1_6/io_i_5_in1[0] cb_1_6/io_i_5_in1[1]
+ cb_1_6/io_i_5_in1[2] cb_1_6/io_i_5_in1[3] cb_1_6/io_i_5_in1[4] cb_1_6/io_i_5_in1[5]
+ cb_1_6/io_i_5_in1[6] cb_1_6/io_i_5_in1[7] cb_1_6/io_i_6_ci cb_1_6/io_i_6_in1[0]
+ cb_1_6/io_i_6_in1[1] cb_1_6/io_i_6_in1[2] cb_1_6/io_i_6_in1[3] cb_1_6/io_i_6_in1[4]
+ cb_1_6/io_i_6_in1[5] cb_1_6/io_i_6_in1[6] cb_1_6/io_i_6_in1[7] cb_1_6/io_i_7_ci
+ cb_1_6/io_i_7_in1[0] cb_1_6/io_i_7_in1[1] cb_1_6/io_i_7_in1[2] cb_1_6/io_i_7_in1[3]
+ cb_1_6/io_i_7_in1[4] cb_1_6/io_i_7_in1[5] cb_1_6/io_i_7_in1[6] cb_1_6/io_i_7_in1[7]
+ cb_1_5/io_vci cb_1_6/io_vci cb_1_5/io_vi cb_1_9/io_we_i cb_1_5/io_wo[0] cb_1_5/io_wo[10]
+ cb_1_5/io_wo[11] cb_1_5/io_wo[12] cb_1_5/io_wo[13] cb_1_5/io_wo[14] cb_1_5/io_wo[15]
+ cb_1_5/io_wo[16] cb_1_5/io_wo[17] cb_1_5/io_wo[18] cb_1_5/io_wo[19] cb_1_5/io_wo[1]
+ cb_1_5/io_wo[20] cb_1_5/io_wo[21] cb_1_5/io_wo[22] cb_1_5/io_wo[23] cb_1_5/io_wo[24]
+ cb_1_5/io_wo[25] cb_1_5/io_wo[26] cb_1_5/io_wo[27] cb_1_5/io_wo[28] cb_1_5/io_wo[29]
+ cb_1_5/io_wo[2] cb_1_5/io_wo[30] cb_1_5/io_wo[31] cb_1_5/io_wo[32] cb_1_5/io_wo[33]
+ cb_1_5/io_wo[34] cb_1_5/io_wo[35] cb_1_5/io_wo[36] cb_1_5/io_wo[37] cb_1_5/io_wo[38]
+ cb_1_5/io_wo[39] cb_1_5/io_wo[3] cb_1_5/io_wo[40] cb_1_5/io_wo[41] cb_1_5/io_wo[42]
+ cb_1_5/io_wo[43] cb_1_5/io_wo[44] cb_1_5/io_wo[45] cb_1_5/io_wo[46] cb_1_5/io_wo[47]
+ cb_1_5/io_wo[48] cb_1_5/io_wo[49] cb_1_5/io_wo[4] cb_1_5/io_wo[50] cb_1_5/io_wo[51]
+ cb_1_5/io_wo[52] cb_1_5/io_wo[53] cb_1_5/io_wo[54] cb_1_5/io_wo[55] cb_1_5/io_wo[56]
+ cb_1_5/io_wo[57] cb_1_5/io_wo[58] cb_1_5/io_wo[59] cb_1_5/io_wo[5] cb_1_5/io_wo[60]
+ cb_1_5/io_wo[61] cb_1_5/io_wo[62] cb_1_5/io_wo[63] cb_1_5/io_wo[6] cb_1_5/io_wo[7]
+ cb_1_5/io_wo[8] cb_1_5/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_3_9 cb_3_9/io_adr_i[0] cb_3_9/io_adr_i[1] cb_3_9/io_cs_i cb_3_9/io_dat_i[0] cb_3_9/io_dat_i[10]
+ cb_3_9/io_dat_i[11] cb_3_9/io_dat_i[12] cb_3_9/io_dat_i[13] cb_3_9/io_dat_i[14]
+ cb_3_9/io_dat_i[15] cb_3_9/io_dat_i[1] cb_3_9/io_dat_i[2] cb_3_9/io_dat_i[3] cb_3_9/io_dat_i[4]
+ cb_3_9/io_dat_i[5] cb_3_9/io_dat_i[6] cb_3_9/io_dat_i[7] cb_3_9/io_dat_i[8] cb_3_9/io_dat_i[9]
+ cb_3_9/io_dat_o[0] cb_3_9/io_dat_o[10] cb_3_9/io_dat_o[11] cb_3_9/io_dat_o[12] cb_3_9/io_dat_o[13]
+ cb_3_9/io_dat_o[14] cb_3_9/io_dat_o[15] cb_3_9/io_dat_o[1] cb_3_9/io_dat_o[2] cb_3_9/io_dat_o[3]
+ cb_3_9/io_dat_o[4] cb_3_9/io_dat_o[5] cb_3_9/io_dat_o[6] cb_3_9/io_dat_o[7] cb_3_9/io_dat_o[8]
+ cb_3_9/io_dat_o[9] cb_3_9/io_eo[0] cb_3_9/io_eo[10] cb_3_9/io_eo[11] cb_3_9/io_eo[12]
+ cb_3_9/io_eo[13] cb_3_9/io_eo[14] cb_3_9/io_eo[15] cb_3_9/io_eo[16] cb_3_9/io_eo[17]
+ cb_3_9/io_eo[18] cb_3_9/io_eo[19] cb_3_9/io_eo[1] cb_3_9/io_eo[20] cb_3_9/io_eo[21]
+ cb_3_9/io_eo[22] cb_3_9/io_eo[23] cb_3_9/io_eo[24] cb_3_9/io_eo[25] cb_3_9/io_eo[26]
+ cb_3_9/io_eo[27] cb_3_9/io_eo[28] cb_3_9/io_eo[29] cb_3_9/io_eo[2] cb_3_9/io_eo[30]
+ cb_3_9/io_eo[31] cb_3_9/io_eo[32] cb_3_9/io_eo[33] cb_3_9/io_eo[34] cb_3_9/io_eo[35]
+ cb_3_9/io_eo[36] cb_3_9/io_eo[37] cb_3_9/io_eo[38] cb_3_9/io_eo[39] cb_3_9/io_eo[3]
+ cb_3_9/io_eo[40] cb_3_9/io_eo[41] cb_3_9/io_eo[42] cb_3_9/io_eo[43] cb_3_9/io_eo[44]
+ cb_3_9/io_eo[45] cb_3_9/io_eo[46] cb_3_9/io_eo[47] cb_3_9/io_eo[48] cb_3_9/io_eo[49]
+ cb_3_9/io_eo[4] cb_3_9/io_eo[50] cb_3_9/io_eo[51] cb_3_9/io_eo[52] cb_3_9/io_eo[53]
+ cb_3_9/io_eo[54] cb_3_9/io_eo[55] cb_3_9/io_eo[56] cb_3_9/io_eo[57] cb_3_9/io_eo[58]
+ cb_3_9/io_eo[59] cb_3_9/io_eo[5] cb_3_9/io_eo[60] cb_3_9/io_eo[61] cb_3_9/io_eo[62]
+ cb_3_9/io_eo[63] cb_3_9/io_eo[6] cb_3_9/io_eo[7] cb_3_9/io_eo[8] cb_3_9/io_eo[9]
+ cb_3_9/io_i_0_ci cb_3_9/io_i_0_in1[0] cb_3_9/io_i_0_in1[1] cb_3_9/io_i_0_in1[2]
+ cb_3_9/io_i_0_in1[3] cb_3_9/io_i_0_in1[4] cb_3_9/io_i_0_in1[5] cb_3_9/io_i_0_in1[6]
+ cb_3_9/io_i_0_in1[7] cb_3_9/io_i_1_ci cb_3_9/io_i_1_in1[0] cb_3_9/io_i_1_in1[1]
+ cb_3_9/io_i_1_in1[2] cb_3_9/io_i_1_in1[3] cb_3_9/io_i_1_in1[4] cb_3_9/io_i_1_in1[5]
+ cb_3_9/io_i_1_in1[6] cb_3_9/io_i_1_in1[7] cb_3_9/io_i_2_ci cb_3_9/io_i_2_in1[0]
+ cb_3_9/io_i_2_in1[1] cb_3_9/io_i_2_in1[2] cb_3_9/io_i_2_in1[3] cb_3_9/io_i_2_in1[4]
+ cb_3_9/io_i_2_in1[5] cb_3_9/io_i_2_in1[6] cb_3_9/io_i_2_in1[7] cb_3_9/io_i_3_ci
+ cb_3_9/io_i_3_in1[0] cb_3_9/io_i_3_in1[1] cb_3_9/io_i_3_in1[2] cb_3_9/io_i_3_in1[3]
+ cb_3_9/io_i_3_in1[4] cb_3_9/io_i_3_in1[5] cb_3_9/io_i_3_in1[6] cb_3_9/io_i_3_in1[7]
+ cb_3_9/io_i_4_ci cb_3_9/io_i_4_in1[0] cb_3_9/io_i_4_in1[1] cb_3_9/io_i_4_in1[2]
+ cb_3_9/io_i_4_in1[3] cb_3_9/io_i_4_in1[4] cb_3_9/io_i_4_in1[5] cb_3_9/io_i_4_in1[6]
+ cb_3_9/io_i_4_in1[7] cb_3_9/io_i_5_ci cb_3_9/io_i_5_in1[0] cb_3_9/io_i_5_in1[1]
+ cb_3_9/io_i_5_in1[2] cb_3_9/io_i_5_in1[3] cb_3_9/io_i_5_in1[4] cb_3_9/io_i_5_in1[5]
+ cb_3_9/io_i_5_in1[6] cb_3_9/io_i_5_in1[7] cb_3_9/io_i_6_ci cb_3_9/io_i_6_in1[0]
+ cb_3_9/io_i_6_in1[1] cb_3_9/io_i_6_in1[2] cb_3_9/io_i_6_in1[3] cb_3_9/io_i_6_in1[4]
+ cb_3_9/io_i_6_in1[5] cb_3_9/io_i_6_in1[6] cb_3_9/io_i_6_in1[7] cb_3_9/io_i_7_ci
+ cb_3_9/io_i_7_in1[0] cb_3_9/io_i_7_in1[1] cb_3_9/io_i_7_in1[2] cb_3_9/io_i_7_in1[3]
+ cb_3_9/io_i_7_in1[4] cb_3_9/io_i_7_in1[5] cb_3_9/io_i_7_in1[6] cb_3_9/io_i_7_in1[7]
+ cb_3_9/io_o_0_co cb_3_9/io_o_0_out[0] cb_3_9/io_o_0_out[1] cb_3_9/io_o_0_out[2]
+ cb_3_9/io_o_0_out[3] cb_3_9/io_o_0_out[4] cb_3_9/io_o_0_out[5] cb_3_9/io_o_0_out[6]
+ cb_3_9/io_o_0_out[7] cb_3_9/io_o_1_co cb_3_9/io_o_1_out[0] cb_3_9/io_o_1_out[1]
+ cb_3_9/io_o_1_out[2] cb_3_9/io_o_1_out[3] cb_3_9/io_o_1_out[4] cb_3_9/io_o_1_out[5]
+ cb_3_9/io_o_1_out[6] cb_3_9/io_o_1_out[7] cb_3_9/io_o_2_co cb_3_9/io_o_2_out[0]
+ cb_3_9/io_o_2_out[1] cb_3_9/io_o_2_out[2] cb_3_9/io_o_2_out[3] cb_3_9/io_o_2_out[4]
+ cb_3_9/io_o_2_out[5] cb_3_9/io_o_2_out[6] cb_3_9/io_o_2_out[7] cb_3_9/io_o_3_co
+ cb_3_9/io_o_3_out[0] cb_3_9/io_o_3_out[1] cb_3_9/io_o_3_out[2] cb_3_9/io_o_3_out[3]
+ cb_3_9/io_o_3_out[4] cb_3_9/io_o_3_out[5] cb_3_9/io_o_3_out[6] cb_3_9/io_o_3_out[7]
+ cb_3_9/io_o_4_co cb_3_9/io_o_4_out[0] cb_3_9/io_o_4_out[1] cb_3_9/io_o_4_out[2]
+ cb_3_9/io_o_4_out[3] cb_3_9/io_o_4_out[4] cb_3_9/io_o_4_out[5] cb_3_9/io_o_4_out[6]
+ cb_3_9/io_o_4_out[7] cb_3_9/io_o_5_co cb_3_9/io_o_5_out[0] cb_3_9/io_o_5_out[1]
+ cb_3_9/io_o_5_out[2] cb_3_9/io_o_5_out[3] cb_3_9/io_o_5_out[4] cb_3_9/io_o_5_out[5]
+ cb_3_9/io_o_5_out[6] cb_3_9/io_o_5_out[7] cb_3_9/io_o_6_co cb_3_9/io_o_6_out[0]
+ cb_3_9/io_o_6_out[1] cb_3_9/io_o_6_out[2] cb_3_9/io_o_6_out[3] cb_3_9/io_o_6_out[4]
+ cb_3_9/io_o_6_out[5] cb_3_9/io_o_6_out[6] cb_3_9/io_o_6_out[7] cb_3_9/io_o_7_co
+ cb_3_9/io_o_7_out[0] cb_3_9/io_o_7_out[1] cb_3_9/io_o_7_out[2] cb_3_9/io_o_7_out[3]
+ cb_3_9/io_o_7_out[4] cb_3_9/io_o_7_out[5] cb_3_9/io_o_7_out[6] cb_3_9/io_o_7_out[7]
+ cb_3_9/io_vci cb_3_9/io_vco cb_3_9/io_vi cb_3_9/io_we_i cb_3_9/io_wo[0] cb_3_9/io_wo[10]
+ cb_3_9/io_wo[11] cb_3_9/io_wo[12] cb_3_9/io_wo[13] cb_3_9/io_wo[14] cb_3_9/io_wo[15]
+ cb_3_9/io_wo[16] cb_3_9/io_wo[17] cb_3_9/io_wo[18] cb_3_9/io_wo[19] cb_3_9/io_wo[1]
+ cb_3_9/io_wo[20] cb_3_9/io_wo[21] cb_3_9/io_wo[22] cb_3_9/io_wo[23] cb_3_9/io_wo[24]
+ cb_3_9/io_wo[25] cb_3_9/io_wo[26] cb_3_9/io_wo[27] cb_3_9/io_wo[28] cb_3_9/io_wo[29]
+ cb_3_9/io_wo[2] cb_3_9/io_wo[30] cb_3_9/io_wo[31] cb_3_9/io_wo[32] cb_3_9/io_wo[33]
+ cb_3_9/io_wo[34] cb_3_9/io_wo[35] cb_3_9/io_wo[36] cb_3_9/io_wo[37] cb_3_9/io_wo[38]
+ cb_3_9/io_wo[39] cb_3_9/io_wo[3] cb_3_9/io_wo[40] cb_3_9/io_wo[41] cb_3_9/io_wo[42]
+ cb_3_9/io_wo[43] cb_3_9/io_wo[44] cb_3_9/io_wo[45] cb_3_9/io_wo[46] cb_3_9/io_wo[47]
+ cb_3_9/io_wo[48] cb_3_9/io_wo[49] cb_3_9/io_wo[4] cb_3_9/io_wo[50] cb_3_9/io_wo[51]
+ cb_3_9/io_wo[52] cb_3_9/io_wo[53] cb_3_9/io_wo[54] cb_3_9/io_wo[55] cb_3_9/io_wo[56]
+ cb_3_9/io_wo[57] cb_3_9/io_wo[58] cb_3_9/io_wo[59] cb_3_9/io_wo[5] cb_3_9/io_wo[60]
+ cb_3_9/io_wo[61] cb_3_9/io_wo[62] cb_3_9/io_wo[63] cb_3_9/io_wo[6] cb_3_9/io_wo[7]
+ cb_3_9/io_wo[8] cb_3_9/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_1_6 cb_1_9/io_adr_i[0] cb_1_9/io_adr_i[1] cb_1_6/io_cs_i cb_1_9/io_dat_i[0] cb_1_9/io_dat_i[10]
+ cb_1_9/io_dat_i[11] cb_1_9/io_dat_i[12] cb_1_9/io_dat_i[13] cb_1_9/io_dat_i[14]
+ cb_1_9/io_dat_i[15] cb_1_9/io_dat_i[1] cb_1_9/io_dat_i[2] cb_1_9/io_dat_i[3] cb_1_9/io_dat_i[4]
+ cb_1_9/io_dat_i[5] cb_1_9/io_dat_i[6] cb_1_9/io_dat_i[7] cb_1_9/io_dat_i[8] cb_1_9/io_dat_i[9]
+ cb_1_6/io_dat_o[0] cb_1_6/io_dat_o[10] cb_1_6/io_dat_o[11] cb_1_6/io_dat_o[12] cb_1_6/io_dat_o[13]
+ cb_1_6/io_dat_o[14] cb_1_6/io_dat_o[15] cb_1_6/io_dat_o[1] cb_1_6/io_dat_o[2] cb_1_6/io_dat_o[3]
+ cb_1_6/io_dat_o[4] cb_1_6/io_dat_o[5] cb_1_6/io_dat_o[6] cb_1_6/io_dat_o[7] cb_1_6/io_dat_o[8]
+ cb_1_6/io_dat_o[9] cb_1_7/io_wo[0] cb_1_7/io_wo[10] cb_1_7/io_wo[11] cb_1_7/io_wo[12]
+ cb_1_7/io_wo[13] cb_1_7/io_wo[14] cb_1_7/io_wo[15] cb_1_7/io_wo[16] cb_1_7/io_wo[17]
+ cb_1_7/io_wo[18] cb_1_7/io_wo[19] cb_1_7/io_wo[1] cb_1_7/io_wo[20] cb_1_7/io_wo[21]
+ cb_1_7/io_wo[22] cb_1_7/io_wo[23] cb_1_7/io_wo[24] cb_1_7/io_wo[25] cb_1_7/io_wo[26]
+ cb_1_7/io_wo[27] cb_1_7/io_wo[28] cb_1_7/io_wo[29] cb_1_7/io_wo[2] cb_1_7/io_wo[30]
+ cb_1_7/io_wo[31] cb_1_7/io_wo[32] cb_1_7/io_wo[33] cb_1_7/io_wo[34] cb_1_7/io_wo[35]
+ cb_1_7/io_wo[36] cb_1_7/io_wo[37] cb_1_7/io_wo[38] cb_1_7/io_wo[39] cb_1_7/io_wo[3]
+ cb_1_7/io_wo[40] cb_1_7/io_wo[41] cb_1_7/io_wo[42] cb_1_7/io_wo[43] cb_1_7/io_wo[44]
+ cb_1_7/io_wo[45] cb_1_7/io_wo[46] cb_1_7/io_wo[47] cb_1_7/io_wo[48] cb_1_7/io_wo[49]
+ cb_1_7/io_wo[4] cb_1_7/io_wo[50] cb_1_7/io_wo[51] cb_1_7/io_wo[52] cb_1_7/io_wo[53]
+ cb_1_7/io_wo[54] cb_1_7/io_wo[55] cb_1_7/io_wo[56] cb_1_7/io_wo[57] cb_1_7/io_wo[58]
+ cb_1_7/io_wo[59] cb_1_7/io_wo[5] cb_1_7/io_wo[60] cb_1_7/io_wo[61] cb_1_7/io_wo[62]
+ cb_1_7/io_wo[63] cb_1_7/io_wo[6] cb_1_7/io_wo[7] cb_1_7/io_wo[8] cb_1_7/io_wo[9]
+ cb_1_6/io_i_0_ci cb_1_6/io_i_0_in1[0] cb_1_6/io_i_0_in1[1] cb_1_6/io_i_0_in1[2]
+ cb_1_6/io_i_0_in1[3] cb_1_6/io_i_0_in1[4] cb_1_6/io_i_0_in1[5] cb_1_6/io_i_0_in1[6]
+ cb_1_6/io_i_0_in1[7] cb_1_6/io_i_1_ci cb_1_6/io_i_1_in1[0] cb_1_6/io_i_1_in1[1]
+ cb_1_6/io_i_1_in1[2] cb_1_6/io_i_1_in1[3] cb_1_6/io_i_1_in1[4] cb_1_6/io_i_1_in1[5]
+ cb_1_6/io_i_1_in1[6] cb_1_6/io_i_1_in1[7] cb_1_6/io_i_2_ci cb_1_6/io_i_2_in1[0]
+ cb_1_6/io_i_2_in1[1] cb_1_6/io_i_2_in1[2] cb_1_6/io_i_2_in1[3] cb_1_6/io_i_2_in1[4]
+ cb_1_6/io_i_2_in1[5] cb_1_6/io_i_2_in1[6] cb_1_6/io_i_2_in1[7] cb_1_6/io_i_3_ci
+ cb_1_6/io_i_3_in1[0] cb_1_6/io_i_3_in1[1] cb_1_6/io_i_3_in1[2] cb_1_6/io_i_3_in1[3]
+ cb_1_6/io_i_3_in1[4] cb_1_6/io_i_3_in1[5] cb_1_6/io_i_3_in1[6] cb_1_6/io_i_3_in1[7]
+ cb_1_6/io_i_4_ci cb_1_6/io_i_4_in1[0] cb_1_6/io_i_4_in1[1] cb_1_6/io_i_4_in1[2]
+ cb_1_6/io_i_4_in1[3] cb_1_6/io_i_4_in1[4] cb_1_6/io_i_4_in1[5] cb_1_6/io_i_4_in1[6]
+ cb_1_6/io_i_4_in1[7] cb_1_6/io_i_5_ci cb_1_6/io_i_5_in1[0] cb_1_6/io_i_5_in1[1]
+ cb_1_6/io_i_5_in1[2] cb_1_6/io_i_5_in1[3] cb_1_6/io_i_5_in1[4] cb_1_6/io_i_5_in1[5]
+ cb_1_6/io_i_5_in1[6] cb_1_6/io_i_5_in1[7] cb_1_6/io_i_6_ci cb_1_6/io_i_6_in1[0]
+ cb_1_6/io_i_6_in1[1] cb_1_6/io_i_6_in1[2] cb_1_6/io_i_6_in1[3] cb_1_6/io_i_6_in1[4]
+ cb_1_6/io_i_6_in1[5] cb_1_6/io_i_6_in1[6] cb_1_6/io_i_6_in1[7] cb_1_6/io_i_7_ci
+ cb_1_6/io_i_7_in1[0] cb_1_6/io_i_7_in1[1] cb_1_6/io_i_7_in1[2] cb_1_6/io_i_7_in1[3]
+ cb_1_6/io_i_7_in1[4] cb_1_6/io_i_7_in1[5] cb_1_6/io_i_7_in1[6] cb_1_6/io_i_7_in1[7]
+ cb_1_7/io_i_0_ci cb_1_7/io_i_0_in1[0] cb_1_7/io_i_0_in1[1] cb_1_7/io_i_0_in1[2]
+ cb_1_7/io_i_0_in1[3] cb_1_7/io_i_0_in1[4] cb_1_7/io_i_0_in1[5] cb_1_7/io_i_0_in1[6]
+ cb_1_7/io_i_0_in1[7] cb_1_7/io_i_1_ci cb_1_7/io_i_1_in1[0] cb_1_7/io_i_1_in1[1]
+ cb_1_7/io_i_1_in1[2] cb_1_7/io_i_1_in1[3] cb_1_7/io_i_1_in1[4] cb_1_7/io_i_1_in1[5]
+ cb_1_7/io_i_1_in1[6] cb_1_7/io_i_1_in1[7] cb_1_7/io_i_2_ci cb_1_7/io_i_2_in1[0]
+ cb_1_7/io_i_2_in1[1] cb_1_7/io_i_2_in1[2] cb_1_7/io_i_2_in1[3] cb_1_7/io_i_2_in1[4]
+ cb_1_7/io_i_2_in1[5] cb_1_7/io_i_2_in1[6] cb_1_7/io_i_2_in1[7] cb_1_7/io_i_3_ci
+ cb_1_7/io_i_3_in1[0] cb_1_7/io_i_3_in1[1] cb_1_7/io_i_3_in1[2] cb_1_7/io_i_3_in1[3]
+ cb_1_7/io_i_3_in1[4] cb_1_7/io_i_3_in1[5] cb_1_7/io_i_3_in1[6] cb_1_7/io_i_3_in1[7]
+ cb_1_7/io_i_4_ci cb_1_7/io_i_4_in1[0] cb_1_7/io_i_4_in1[1] cb_1_7/io_i_4_in1[2]
+ cb_1_7/io_i_4_in1[3] cb_1_7/io_i_4_in1[4] cb_1_7/io_i_4_in1[5] cb_1_7/io_i_4_in1[6]
+ cb_1_7/io_i_4_in1[7] cb_1_7/io_i_5_ci cb_1_7/io_i_5_in1[0] cb_1_7/io_i_5_in1[1]
+ cb_1_7/io_i_5_in1[2] cb_1_7/io_i_5_in1[3] cb_1_7/io_i_5_in1[4] cb_1_7/io_i_5_in1[5]
+ cb_1_7/io_i_5_in1[6] cb_1_7/io_i_5_in1[7] cb_1_7/io_i_6_ci cb_1_7/io_i_6_in1[0]
+ cb_1_7/io_i_6_in1[1] cb_1_7/io_i_6_in1[2] cb_1_7/io_i_6_in1[3] cb_1_7/io_i_6_in1[4]
+ cb_1_7/io_i_6_in1[5] cb_1_7/io_i_6_in1[6] cb_1_7/io_i_6_in1[7] cb_1_7/io_i_7_ci
+ cb_1_7/io_i_7_in1[0] cb_1_7/io_i_7_in1[1] cb_1_7/io_i_7_in1[2] cb_1_7/io_i_7_in1[3]
+ cb_1_7/io_i_7_in1[4] cb_1_7/io_i_7_in1[5] cb_1_7/io_i_7_in1[6] cb_1_7/io_i_7_in1[7]
+ cb_1_6/io_vci cb_1_7/io_vci cb_1_6/io_vi cb_1_9/io_we_i cb_1_6/io_wo[0] cb_1_6/io_wo[10]
+ cb_1_6/io_wo[11] cb_1_6/io_wo[12] cb_1_6/io_wo[13] cb_1_6/io_wo[14] cb_1_6/io_wo[15]
+ cb_1_6/io_wo[16] cb_1_6/io_wo[17] cb_1_6/io_wo[18] cb_1_6/io_wo[19] cb_1_6/io_wo[1]
+ cb_1_6/io_wo[20] cb_1_6/io_wo[21] cb_1_6/io_wo[22] cb_1_6/io_wo[23] cb_1_6/io_wo[24]
+ cb_1_6/io_wo[25] cb_1_6/io_wo[26] cb_1_6/io_wo[27] cb_1_6/io_wo[28] cb_1_6/io_wo[29]
+ cb_1_6/io_wo[2] cb_1_6/io_wo[30] cb_1_6/io_wo[31] cb_1_6/io_wo[32] cb_1_6/io_wo[33]
+ cb_1_6/io_wo[34] cb_1_6/io_wo[35] cb_1_6/io_wo[36] cb_1_6/io_wo[37] cb_1_6/io_wo[38]
+ cb_1_6/io_wo[39] cb_1_6/io_wo[3] cb_1_6/io_wo[40] cb_1_6/io_wo[41] cb_1_6/io_wo[42]
+ cb_1_6/io_wo[43] cb_1_6/io_wo[44] cb_1_6/io_wo[45] cb_1_6/io_wo[46] cb_1_6/io_wo[47]
+ cb_1_6/io_wo[48] cb_1_6/io_wo[49] cb_1_6/io_wo[4] cb_1_6/io_wo[50] cb_1_6/io_wo[51]
+ cb_1_6/io_wo[52] cb_1_6/io_wo[53] cb_1_6/io_wo[54] cb_1_6/io_wo[55] cb_1_6/io_wo[56]
+ cb_1_6/io_wo[57] cb_1_6/io_wo[58] cb_1_6/io_wo[59] cb_1_6/io_wo[5] cb_1_6/io_wo[60]
+ cb_1_6/io_wo[61] cb_1_6/io_wo[62] cb_1_6/io_wo[63] cb_1_6/io_wo[6] cb_1_6/io_wo[7]
+ cb_1_6/io_wo[8] cb_1_6/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_1_7 cb_1_9/io_adr_i[0] cb_1_9/io_adr_i[1] cb_1_7/io_cs_i cb_1_9/io_dat_i[0] cb_1_9/io_dat_i[10]
+ cb_1_9/io_dat_i[11] cb_1_9/io_dat_i[12] cb_1_9/io_dat_i[13] cb_1_9/io_dat_i[14]
+ cb_1_9/io_dat_i[15] cb_1_9/io_dat_i[1] cb_1_9/io_dat_i[2] cb_1_9/io_dat_i[3] cb_1_9/io_dat_i[4]
+ cb_1_9/io_dat_i[5] cb_1_9/io_dat_i[6] cb_1_9/io_dat_i[7] cb_1_9/io_dat_i[8] cb_1_9/io_dat_i[9]
+ cb_1_7/io_dat_o[0] cb_1_7/io_dat_o[10] cb_1_7/io_dat_o[11] cb_1_7/io_dat_o[12] cb_1_7/io_dat_o[13]
+ cb_1_7/io_dat_o[14] cb_1_7/io_dat_o[15] cb_1_7/io_dat_o[1] cb_1_7/io_dat_o[2] cb_1_7/io_dat_o[3]
+ cb_1_7/io_dat_o[4] cb_1_7/io_dat_o[5] cb_1_7/io_dat_o[6] cb_1_7/io_dat_o[7] cb_1_7/io_dat_o[8]
+ cb_1_7/io_dat_o[9] cb_1_8/io_wo[0] cb_1_8/io_wo[10] cb_1_8/io_wo[11] cb_1_8/io_wo[12]
+ cb_1_8/io_wo[13] cb_1_8/io_wo[14] cb_1_8/io_wo[15] cb_1_8/io_wo[16] cb_1_8/io_wo[17]
+ cb_1_8/io_wo[18] cb_1_8/io_wo[19] cb_1_8/io_wo[1] cb_1_8/io_wo[20] cb_1_8/io_wo[21]
+ cb_1_8/io_wo[22] cb_1_8/io_wo[23] cb_1_8/io_wo[24] cb_1_8/io_wo[25] cb_1_8/io_wo[26]
+ cb_1_8/io_wo[27] cb_1_8/io_wo[28] cb_1_8/io_wo[29] cb_1_8/io_wo[2] cb_1_8/io_wo[30]
+ cb_1_8/io_wo[31] cb_1_8/io_wo[32] cb_1_8/io_wo[33] cb_1_8/io_wo[34] cb_1_8/io_wo[35]
+ cb_1_8/io_wo[36] cb_1_8/io_wo[37] cb_1_8/io_wo[38] cb_1_8/io_wo[39] cb_1_8/io_wo[3]
+ cb_1_8/io_wo[40] cb_1_8/io_wo[41] cb_1_8/io_wo[42] cb_1_8/io_wo[43] cb_1_8/io_wo[44]
+ cb_1_8/io_wo[45] cb_1_8/io_wo[46] cb_1_8/io_wo[47] cb_1_8/io_wo[48] cb_1_8/io_wo[49]
+ cb_1_8/io_wo[4] cb_1_8/io_wo[50] cb_1_8/io_wo[51] cb_1_8/io_wo[52] cb_1_8/io_wo[53]
+ cb_1_8/io_wo[54] cb_1_8/io_wo[55] cb_1_8/io_wo[56] cb_1_8/io_wo[57] cb_1_8/io_wo[58]
+ cb_1_8/io_wo[59] cb_1_8/io_wo[5] cb_1_8/io_wo[60] cb_1_8/io_wo[61] cb_1_8/io_wo[62]
+ cb_1_8/io_wo[63] cb_1_8/io_wo[6] cb_1_8/io_wo[7] cb_1_8/io_wo[8] cb_1_8/io_wo[9]
+ cb_1_7/io_i_0_ci cb_1_7/io_i_0_in1[0] cb_1_7/io_i_0_in1[1] cb_1_7/io_i_0_in1[2]
+ cb_1_7/io_i_0_in1[3] cb_1_7/io_i_0_in1[4] cb_1_7/io_i_0_in1[5] cb_1_7/io_i_0_in1[6]
+ cb_1_7/io_i_0_in1[7] cb_1_7/io_i_1_ci cb_1_7/io_i_1_in1[0] cb_1_7/io_i_1_in1[1]
+ cb_1_7/io_i_1_in1[2] cb_1_7/io_i_1_in1[3] cb_1_7/io_i_1_in1[4] cb_1_7/io_i_1_in1[5]
+ cb_1_7/io_i_1_in1[6] cb_1_7/io_i_1_in1[7] cb_1_7/io_i_2_ci cb_1_7/io_i_2_in1[0]
+ cb_1_7/io_i_2_in1[1] cb_1_7/io_i_2_in1[2] cb_1_7/io_i_2_in1[3] cb_1_7/io_i_2_in1[4]
+ cb_1_7/io_i_2_in1[5] cb_1_7/io_i_2_in1[6] cb_1_7/io_i_2_in1[7] cb_1_7/io_i_3_ci
+ cb_1_7/io_i_3_in1[0] cb_1_7/io_i_3_in1[1] cb_1_7/io_i_3_in1[2] cb_1_7/io_i_3_in1[3]
+ cb_1_7/io_i_3_in1[4] cb_1_7/io_i_3_in1[5] cb_1_7/io_i_3_in1[6] cb_1_7/io_i_3_in1[7]
+ cb_1_7/io_i_4_ci cb_1_7/io_i_4_in1[0] cb_1_7/io_i_4_in1[1] cb_1_7/io_i_4_in1[2]
+ cb_1_7/io_i_4_in1[3] cb_1_7/io_i_4_in1[4] cb_1_7/io_i_4_in1[5] cb_1_7/io_i_4_in1[6]
+ cb_1_7/io_i_4_in1[7] cb_1_7/io_i_5_ci cb_1_7/io_i_5_in1[0] cb_1_7/io_i_5_in1[1]
+ cb_1_7/io_i_5_in1[2] cb_1_7/io_i_5_in1[3] cb_1_7/io_i_5_in1[4] cb_1_7/io_i_5_in1[5]
+ cb_1_7/io_i_5_in1[6] cb_1_7/io_i_5_in1[7] cb_1_7/io_i_6_ci cb_1_7/io_i_6_in1[0]
+ cb_1_7/io_i_6_in1[1] cb_1_7/io_i_6_in1[2] cb_1_7/io_i_6_in1[3] cb_1_7/io_i_6_in1[4]
+ cb_1_7/io_i_6_in1[5] cb_1_7/io_i_6_in1[6] cb_1_7/io_i_6_in1[7] cb_1_7/io_i_7_ci
+ cb_1_7/io_i_7_in1[0] cb_1_7/io_i_7_in1[1] cb_1_7/io_i_7_in1[2] cb_1_7/io_i_7_in1[3]
+ cb_1_7/io_i_7_in1[4] cb_1_7/io_i_7_in1[5] cb_1_7/io_i_7_in1[6] cb_1_7/io_i_7_in1[7]
+ cb_1_8/io_i_0_ci cb_1_8/io_i_0_in1[0] cb_1_8/io_i_0_in1[1] cb_1_8/io_i_0_in1[2]
+ cb_1_8/io_i_0_in1[3] cb_1_8/io_i_0_in1[4] cb_1_8/io_i_0_in1[5] cb_1_8/io_i_0_in1[6]
+ cb_1_8/io_i_0_in1[7] cb_1_8/io_i_1_ci cb_1_8/io_i_1_in1[0] cb_1_8/io_i_1_in1[1]
+ cb_1_8/io_i_1_in1[2] cb_1_8/io_i_1_in1[3] cb_1_8/io_i_1_in1[4] cb_1_8/io_i_1_in1[5]
+ cb_1_8/io_i_1_in1[6] cb_1_8/io_i_1_in1[7] cb_1_8/io_i_2_ci cb_1_8/io_i_2_in1[0]
+ cb_1_8/io_i_2_in1[1] cb_1_8/io_i_2_in1[2] cb_1_8/io_i_2_in1[3] cb_1_8/io_i_2_in1[4]
+ cb_1_8/io_i_2_in1[5] cb_1_8/io_i_2_in1[6] cb_1_8/io_i_2_in1[7] cb_1_8/io_i_3_ci
+ cb_1_8/io_i_3_in1[0] cb_1_8/io_i_3_in1[1] cb_1_8/io_i_3_in1[2] cb_1_8/io_i_3_in1[3]
+ cb_1_8/io_i_3_in1[4] cb_1_8/io_i_3_in1[5] cb_1_8/io_i_3_in1[6] cb_1_8/io_i_3_in1[7]
+ cb_1_8/io_i_4_ci cb_1_8/io_i_4_in1[0] cb_1_8/io_i_4_in1[1] cb_1_8/io_i_4_in1[2]
+ cb_1_8/io_i_4_in1[3] cb_1_8/io_i_4_in1[4] cb_1_8/io_i_4_in1[5] cb_1_8/io_i_4_in1[6]
+ cb_1_8/io_i_4_in1[7] cb_1_8/io_i_5_ci cb_1_8/io_i_5_in1[0] cb_1_8/io_i_5_in1[1]
+ cb_1_8/io_i_5_in1[2] cb_1_8/io_i_5_in1[3] cb_1_8/io_i_5_in1[4] cb_1_8/io_i_5_in1[5]
+ cb_1_8/io_i_5_in1[6] cb_1_8/io_i_5_in1[7] cb_1_8/io_i_6_ci cb_1_8/io_i_6_in1[0]
+ cb_1_8/io_i_6_in1[1] cb_1_8/io_i_6_in1[2] cb_1_8/io_i_6_in1[3] cb_1_8/io_i_6_in1[4]
+ cb_1_8/io_i_6_in1[5] cb_1_8/io_i_6_in1[6] cb_1_8/io_i_6_in1[7] cb_1_8/io_i_7_ci
+ cb_1_8/io_i_7_in1[0] cb_1_8/io_i_7_in1[1] cb_1_8/io_i_7_in1[2] cb_1_8/io_i_7_in1[3]
+ cb_1_8/io_i_7_in1[4] cb_1_8/io_i_7_in1[5] cb_1_8/io_i_7_in1[6] cb_1_8/io_i_7_in1[7]
+ cb_1_7/io_vci cb_1_8/io_vci cb_1_7/io_vi cb_1_9/io_we_i cb_1_7/io_wo[0] cb_1_7/io_wo[10]
+ cb_1_7/io_wo[11] cb_1_7/io_wo[12] cb_1_7/io_wo[13] cb_1_7/io_wo[14] cb_1_7/io_wo[15]
+ cb_1_7/io_wo[16] cb_1_7/io_wo[17] cb_1_7/io_wo[18] cb_1_7/io_wo[19] cb_1_7/io_wo[1]
+ cb_1_7/io_wo[20] cb_1_7/io_wo[21] cb_1_7/io_wo[22] cb_1_7/io_wo[23] cb_1_7/io_wo[24]
+ cb_1_7/io_wo[25] cb_1_7/io_wo[26] cb_1_7/io_wo[27] cb_1_7/io_wo[28] cb_1_7/io_wo[29]
+ cb_1_7/io_wo[2] cb_1_7/io_wo[30] cb_1_7/io_wo[31] cb_1_7/io_wo[32] cb_1_7/io_wo[33]
+ cb_1_7/io_wo[34] cb_1_7/io_wo[35] cb_1_7/io_wo[36] cb_1_7/io_wo[37] cb_1_7/io_wo[38]
+ cb_1_7/io_wo[39] cb_1_7/io_wo[3] cb_1_7/io_wo[40] cb_1_7/io_wo[41] cb_1_7/io_wo[42]
+ cb_1_7/io_wo[43] cb_1_7/io_wo[44] cb_1_7/io_wo[45] cb_1_7/io_wo[46] cb_1_7/io_wo[47]
+ cb_1_7/io_wo[48] cb_1_7/io_wo[49] cb_1_7/io_wo[4] cb_1_7/io_wo[50] cb_1_7/io_wo[51]
+ cb_1_7/io_wo[52] cb_1_7/io_wo[53] cb_1_7/io_wo[54] cb_1_7/io_wo[55] cb_1_7/io_wo[56]
+ cb_1_7/io_wo[57] cb_1_7/io_wo[58] cb_1_7/io_wo[59] cb_1_7/io_wo[5] cb_1_7/io_wo[60]
+ cb_1_7/io_wo[61] cb_1_7/io_wo[62] cb_1_7/io_wo[63] cb_1_7/io_wo[6] cb_1_7/io_wo[7]
+ cb_1_7/io_wo[8] cb_1_7/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_1_8 cb_1_9/io_adr_i[0] cb_1_9/io_adr_i[1] cb_1_8/io_cs_i cb_1_9/io_dat_i[0] cb_1_9/io_dat_i[10]
+ cb_1_9/io_dat_i[11] cb_1_9/io_dat_i[12] cb_1_9/io_dat_i[13] cb_1_9/io_dat_i[14]
+ cb_1_9/io_dat_i[15] cb_1_9/io_dat_i[1] cb_1_9/io_dat_i[2] cb_1_9/io_dat_i[3] cb_1_9/io_dat_i[4]
+ cb_1_9/io_dat_i[5] cb_1_9/io_dat_i[6] cb_1_9/io_dat_i[7] cb_1_9/io_dat_i[8] cb_1_9/io_dat_i[9]
+ cb_1_8/io_dat_o[0] cb_1_8/io_dat_o[10] cb_1_8/io_dat_o[11] cb_1_8/io_dat_o[12] cb_1_8/io_dat_o[13]
+ cb_1_8/io_dat_o[14] cb_1_8/io_dat_o[15] cb_1_8/io_dat_o[1] cb_1_8/io_dat_o[2] cb_1_8/io_dat_o[3]
+ cb_1_8/io_dat_o[4] cb_1_8/io_dat_o[5] cb_1_8/io_dat_o[6] cb_1_8/io_dat_o[7] cb_1_8/io_dat_o[8]
+ cb_1_8/io_dat_o[9] cb_1_9/io_wo[0] cb_1_9/io_wo[10] cb_1_9/io_wo[11] cb_1_9/io_wo[12]
+ cb_1_9/io_wo[13] cb_1_9/io_wo[14] cb_1_9/io_wo[15] cb_1_9/io_wo[16] cb_1_9/io_wo[17]
+ cb_1_9/io_wo[18] cb_1_9/io_wo[19] cb_1_9/io_wo[1] cb_1_9/io_wo[20] cb_1_9/io_wo[21]
+ cb_1_9/io_wo[22] cb_1_9/io_wo[23] cb_1_9/io_wo[24] cb_1_9/io_wo[25] cb_1_9/io_wo[26]
+ cb_1_9/io_wo[27] cb_1_9/io_wo[28] cb_1_9/io_wo[29] cb_1_9/io_wo[2] cb_1_9/io_wo[30]
+ cb_1_9/io_wo[31] cb_1_9/io_wo[32] cb_1_9/io_wo[33] cb_1_9/io_wo[34] cb_1_9/io_wo[35]
+ cb_1_9/io_wo[36] cb_1_9/io_wo[37] cb_1_9/io_wo[38] cb_1_9/io_wo[39] cb_1_9/io_wo[3]
+ cb_1_9/io_wo[40] cb_1_9/io_wo[41] cb_1_9/io_wo[42] cb_1_9/io_wo[43] cb_1_9/io_wo[44]
+ cb_1_9/io_wo[45] cb_1_9/io_wo[46] cb_1_9/io_wo[47] cb_1_9/io_wo[48] cb_1_9/io_wo[49]
+ cb_1_9/io_wo[4] cb_1_9/io_wo[50] cb_1_9/io_wo[51] cb_1_9/io_wo[52] cb_1_9/io_wo[53]
+ cb_1_9/io_wo[54] cb_1_9/io_wo[55] cb_1_9/io_wo[56] cb_1_9/io_wo[57] cb_1_9/io_wo[58]
+ cb_1_9/io_wo[59] cb_1_9/io_wo[5] cb_1_9/io_wo[60] cb_1_9/io_wo[61] cb_1_9/io_wo[62]
+ cb_1_9/io_wo[63] cb_1_9/io_wo[6] cb_1_9/io_wo[7] cb_1_9/io_wo[8] cb_1_9/io_wo[9]
+ cb_1_8/io_i_0_ci cb_1_8/io_i_0_in1[0] cb_1_8/io_i_0_in1[1] cb_1_8/io_i_0_in1[2]
+ cb_1_8/io_i_0_in1[3] cb_1_8/io_i_0_in1[4] cb_1_8/io_i_0_in1[5] cb_1_8/io_i_0_in1[6]
+ cb_1_8/io_i_0_in1[7] cb_1_8/io_i_1_ci cb_1_8/io_i_1_in1[0] cb_1_8/io_i_1_in1[1]
+ cb_1_8/io_i_1_in1[2] cb_1_8/io_i_1_in1[3] cb_1_8/io_i_1_in1[4] cb_1_8/io_i_1_in1[5]
+ cb_1_8/io_i_1_in1[6] cb_1_8/io_i_1_in1[7] cb_1_8/io_i_2_ci cb_1_8/io_i_2_in1[0]
+ cb_1_8/io_i_2_in1[1] cb_1_8/io_i_2_in1[2] cb_1_8/io_i_2_in1[3] cb_1_8/io_i_2_in1[4]
+ cb_1_8/io_i_2_in1[5] cb_1_8/io_i_2_in1[6] cb_1_8/io_i_2_in1[7] cb_1_8/io_i_3_ci
+ cb_1_8/io_i_3_in1[0] cb_1_8/io_i_3_in1[1] cb_1_8/io_i_3_in1[2] cb_1_8/io_i_3_in1[3]
+ cb_1_8/io_i_3_in1[4] cb_1_8/io_i_3_in1[5] cb_1_8/io_i_3_in1[6] cb_1_8/io_i_3_in1[7]
+ cb_1_8/io_i_4_ci cb_1_8/io_i_4_in1[0] cb_1_8/io_i_4_in1[1] cb_1_8/io_i_4_in1[2]
+ cb_1_8/io_i_4_in1[3] cb_1_8/io_i_4_in1[4] cb_1_8/io_i_4_in1[5] cb_1_8/io_i_4_in1[6]
+ cb_1_8/io_i_4_in1[7] cb_1_8/io_i_5_ci cb_1_8/io_i_5_in1[0] cb_1_8/io_i_5_in1[1]
+ cb_1_8/io_i_5_in1[2] cb_1_8/io_i_5_in1[3] cb_1_8/io_i_5_in1[4] cb_1_8/io_i_5_in1[5]
+ cb_1_8/io_i_5_in1[6] cb_1_8/io_i_5_in1[7] cb_1_8/io_i_6_ci cb_1_8/io_i_6_in1[0]
+ cb_1_8/io_i_6_in1[1] cb_1_8/io_i_6_in1[2] cb_1_8/io_i_6_in1[3] cb_1_8/io_i_6_in1[4]
+ cb_1_8/io_i_6_in1[5] cb_1_8/io_i_6_in1[6] cb_1_8/io_i_6_in1[7] cb_1_8/io_i_7_ci
+ cb_1_8/io_i_7_in1[0] cb_1_8/io_i_7_in1[1] cb_1_8/io_i_7_in1[2] cb_1_8/io_i_7_in1[3]
+ cb_1_8/io_i_7_in1[4] cb_1_8/io_i_7_in1[5] cb_1_8/io_i_7_in1[6] cb_1_8/io_i_7_in1[7]
+ cb_1_9/io_i_0_ci cb_1_9/io_i_0_in1[0] cb_1_9/io_i_0_in1[1] cb_1_9/io_i_0_in1[2]
+ cb_1_9/io_i_0_in1[3] cb_1_9/io_i_0_in1[4] cb_1_9/io_i_0_in1[5] cb_1_9/io_i_0_in1[6]
+ cb_1_9/io_i_0_in1[7] cb_1_9/io_i_1_ci cb_1_9/io_i_1_in1[0] cb_1_9/io_i_1_in1[1]
+ cb_1_9/io_i_1_in1[2] cb_1_9/io_i_1_in1[3] cb_1_9/io_i_1_in1[4] cb_1_9/io_i_1_in1[5]
+ cb_1_9/io_i_1_in1[6] cb_1_9/io_i_1_in1[7] cb_1_9/io_i_2_ci cb_1_9/io_i_2_in1[0]
+ cb_1_9/io_i_2_in1[1] cb_1_9/io_i_2_in1[2] cb_1_9/io_i_2_in1[3] cb_1_9/io_i_2_in1[4]
+ cb_1_9/io_i_2_in1[5] cb_1_9/io_i_2_in1[6] cb_1_9/io_i_2_in1[7] cb_1_9/io_i_3_ci
+ cb_1_9/io_i_3_in1[0] cb_1_9/io_i_3_in1[1] cb_1_9/io_i_3_in1[2] cb_1_9/io_i_3_in1[3]
+ cb_1_9/io_i_3_in1[4] cb_1_9/io_i_3_in1[5] cb_1_9/io_i_3_in1[6] cb_1_9/io_i_3_in1[7]
+ cb_1_9/io_i_4_ci cb_1_9/io_i_4_in1[0] cb_1_9/io_i_4_in1[1] cb_1_9/io_i_4_in1[2]
+ cb_1_9/io_i_4_in1[3] cb_1_9/io_i_4_in1[4] cb_1_9/io_i_4_in1[5] cb_1_9/io_i_4_in1[6]
+ cb_1_9/io_i_4_in1[7] cb_1_9/io_i_5_ci cb_1_9/io_i_5_in1[0] cb_1_9/io_i_5_in1[1]
+ cb_1_9/io_i_5_in1[2] cb_1_9/io_i_5_in1[3] cb_1_9/io_i_5_in1[4] cb_1_9/io_i_5_in1[5]
+ cb_1_9/io_i_5_in1[6] cb_1_9/io_i_5_in1[7] cb_1_9/io_i_6_ci cb_1_9/io_i_6_in1[0]
+ cb_1_9/io_i_6_in1[1] cb_1_9/io_i_6_in1[2] cb_1_9/io_i_6_in1[3] cb_1_9/io_i_6_in1[4]
+ cb_1_9/io_i_6_in1[5] cb_1_9/io_i_6_in1[6] cb_1_9/io_i_6_in1[7] cb_1_9/io_i_7_ci
+ cb_1_9/io_i_7_in1[0] cb_1_9/io_i_7_in1[1] cb_1_9/io_i_7_in1[2] cb_1_9/io_i_7_in1[3]
+ cb_1_9/io_i_7_in1[4] cb_1_9/io_i_7_in1[5] cb_1_9/io_i_7_in1[6] cb_1_9/io_i_7_in1[7]
+ cb_1_8/io_vci cb_1_9/io_vci cb_1_8/io_vi cb_1_9/io_we_i cb_1_8/io_wo[0] cb_1_8/io_wo[10]
+ cb_1_8/io_wo[11] cb_1_8/io_wo[12] cb_1_8/io_wo[13] cb_1_8/io_wo[14] cb_1_8/io_wo[15]
+ cb_1_8/io_wo[16] cb_1_8/io_wo[17] cb_1_8/io_wo[18] cb_1_8/io_wo[19] cb_1_8/io_wo[1]
+ cb_1_8/io_wo[20] cb_1_8/io_wo[21] cb_1_8/io_wo[22] cb_1_8/io_wo[23] cb_1_8/io_wo[24]
+ cb_1_8/io_wo[25] cb_1_8/io_wo[26] cb_1_8/io_wo[27] cb_1_8/io_wo[28] cb_1_8/io_wo[29]
+ cb_1_8/io_wo[2] cb_1_8/io_wo[30] cb_1_8/io_wo[31] cb_1_8/io_wo[32] cb_1_8/io_wo[33]
+ cb_1_8/io_wo[34] cb_1_8/io_wo[35] cb_1_8/io_wo[36] cb_1_8/io_wo[37] cb_1_8/io_wo[38]
+ cb_1_8/io_wo[39] cb_1_8/io_wo[3] cb_1_8/io_wo[40] cb_1_8/io_wo[41] cb_1_8/io_wo[42]
+ cb_1_8/io_wo[43] cb_1_8/io_wo[44] cb_1_8/io_wo[45] cb_1_8/io_wo[46] cb_1_8/io_wo[47]
+ cb_1_8/io_wo[48] cb_1_8/io_wo[49] cb_1_8/io_wo[4] cb_1_8/io_wo[50] cb_1_8/io_wo[51]
+ cb_1_8/io_wo[52] cb_1_8/io_wo[53] cb_1_8/io_wo[54] cb_1_8/io_wo[55] cb_1_8/io_wo[56]
+ cb_1_8/io_wo[57] cb_1_8/io_wo[58] cb_1_8/io_wo[59] cb_1_8/io_wo[5] cb_1_8/io_wo[60]
+ cb_1_8/io_wo[61] cb_1_8/io_wo[62] cb_1_8/io_wo[63] cb_1_8/io_wo[6] cb_1_8/io_wo[7]
+ cb_1_8/io_wo[8] cb_1_8/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_1_9 cb_1_9/io_adr_i[0] cb_1_9/io_adr_i[1] cb_1_9/io_cs_i cb_1_9/io_dat_i[0] cb_1_9/io_dat_i[10]
+ cb_1_9/io_dat_i[11] cb_1_9/io_dat_i[12] cb_1_9/io_dat_i[13] cb_1_9/io_dat_i[14]
+ cb_1_9/io_dat_i[15] cb_1_9/io_dat_i[1] cb_1_9/io_dat_i[2] cb_1_9/io_dat_i[3] cb_1_9/io_dat_i[4]
+ cb_1_9/io_dat_i[5] cb_1_9/io_dat_i[6] cb_1_9/io_dat_i[7] cb_1_9/io_dat_i[8] cb_1_9/io_dat_i[9]
+ cb_1_9/io_dat_o[0] cb_1_9/io_dat_o[10] cb_1_9/io_dat_o[11] cb_1_9/io_dat_o[12] cb_1_9/io_dat_o[13]
+ cb_1_9/io_dat_o[14] cb_1_9/io_dat_o[15] cb_1_9/io_dat_o[1] cb_1_9/io_dat_o[2] cb_1_9/io_dat_o[3]
+ cb_1_9/io_dat_o[4] cb_1_9/io_dat_o[5] cb_1_9/io_dat_o[6] cb_1_9/io_dat_o[7] cb_1_9/io_dat_o[8]
+ cb_1_9/io_dat_o[9] cb_1_9/io_eo[0] cb_1_9/io_eo[10] cb_1_9/io_eo[11] cb_1_9/io_eo[12]
+ cb_1_9/io_eo[13] cb_1_9/io_eo[14] cb_1_9/io_eo[15] cb_1_9/io_eo[16] cb_1_9/io_eo[17]
+ cb_1_9/io_eo[18] cb_1_9/io_eo[19] cb_1_9/io_eo[1] cb_1_9/io_eo[20] cb_1_9/io_eo[21]
+ cb_1_9/io_eo[22] cb_1_9/io_eo[23] cb_1_9/io_eo[24] cb_1_9/io_eo[25] cb_1_9/io_eo[26]
+ cb_1_9/io_eo[27] cb_1_9/io_eo[28] cb_1_9/io_eo[29] cb_1_9/io_eo[2] cb_1_9/io_eo[30]
+ cb_1_9/io_eo[31] cb_1_9/io_eo[32] cb_1_9/io_eo[33] cb_1_9/io_eo[34] cb_1_9/io_eo[35]
+ cb_1_9/io_eo[36] cb_1_9/io_eo[37] cb_1_9/io_eo[38] cb_1_9/io_eo[39] cb_1_9/io_eo[3]
+ cb_1_9/io_eo[40] cb_1_9/io_eo[41] cb_1_9/io_eo[42] cb_1_9/io_eo[43] cb_1_9/io_eo[44]
+ cb_1_9/io_eo[45] cb_1_9/io_eo[46] cb_1_9/io_eo[47] cb_1_9/io_eo[48] cb_1_9/io_eo[49]
+ cb_1_9/io_eo[4] cb_1_9/io_eo[50] cb_1_9/io_eo[51] cb_1_9/io_eo[52] cb_1_9/io_eo[53]
+ cb_1_9/io_eo[54] cb_1_9/io_eo[55] cb_1_9/io_eo[56] cb_1_9/io_eo[57] cb_1_9/io_eo[58]
+ cb_1_9/io_eo[59] cb_1_9/io_eo[5] cb_1_9/io_eo[60] cb_1_9/io_eo[61] cb_1_9/io_eo[62]
+ cb_1_9/io_eo[63] cb_1_9/io_eo[6] cb_1_9/io_eo[7] cb_1_9/io_eo[8] cb_1_9/io_eo[9]
+ cb_1_9/io_i_0_ci cb_1_9/io_i_0_in1[0] cb_1_9/io_i_0_in1[1] cb_1_9/io_i_0_in1[2]
+ cb_1_9/io_i_0_in1[3] cb_1_9/io_i_0_in1[4] cb_1_9/io_i_0_in1[5] cb_1_9/io_i_0_in1[6]
+ cb_1_9/io_i_0_in1[7] cb_1_9/io_i_1_ci cb_1_9/io_i_1_in1[0] cb_1_9/io_i_1_in1[1]
+ cb_1_9/io_i_1_in1[2] cb_1_9/io_i_1_in1[3] cb_1_9/io_i_1_in1[4] cb_1_9/io_i_1_in1[5]
+ cb_1_9/io_i_1_in1[6] cb_1_9/io_i_1_in1[7] cb_1_9/io_i_2_ci cb_1_9/io_i_2_in1[0]
+ cb_1_9/io_i_2_in1[1] cb_1_9/io_i_2_in1[2] cb_1_9/io_i_2_in1[3] cb_1_9/io_i_2_in1[4]
+ cb_1_9/io_i_2_in1[5] cb_1_9/io_i_2_in1[6] cb_1_9/io_i_2_in1[7] cb_1_9/io_i_3_ci
+ cb_1_9/io_i_3_in1[0] cb_1_9/io_i_3_in1[1] cb_1_9/io_i_3_in1[2] cb_1_9/io_i_3_in1[3]
+ cb_1_9/io_i_3_in1[4] cb_1_9/io_i_3_in1[5] cb_1_9/io_i_3_in1[6] cb_1_9/io_i_3_in1[7]
+ cb_1_9/io_i_4_ci cb_1_9/io_i_4_in1[0] cb_1_9/io_i_4_in1[1] cb_1_9/io_i_4_in1[2]
+ cb_1_9/io_i_4_in1[3] cb_1_9/io_i_4_in1[4] cb_1_9/io_i_4_in1[5] cb_1_9/io_i_4_in1[6]
+ cb_1_9/io_i_4_in1[7] cb_1_9/io_i_5_ci cb_1_9/io_i_5_in1[0] cb_1_9/io_i_5_in1[1]
+ cb_1_9/io_i_5_in1[2] cb_1_9/io_i_5_in1[3] cb_1_9/io_i_5_in1[4] cb_1_9/io_i_5_in1[5]
+ cb_1_9/io_i_5_in1[6] cb_1_9/io_i_5_in1[7] cb_1_9/io_i_6_ci cb_1_9/io_i_6_in1[0]
+ cb_1_9/io_i_6_in1[1] cb_1_9/io_i_6_in1[2] cb_1_9/io_i_6_in1[3] cb_1_9/io_i_6_in1[4]
+ cb_1_9/io_i_6_in1[5] cb_1_9/io_i_6_in1[6] cb_1_9/io_i_6_in1[7] cb_1_9/io_i_7_ci
+ cb_1_9/io_i_7_in1[0] cb_1_9/io_i_7_in1[1] cb_1_9/io_i_7_in1[2] cb_1_9/io_i_7_in1[3]
+ cb_1_9/io_i_7_in1[4] cb_1_9/io_i_7_in1[5] cb_1_9/io_i_7_in1[6] cb_1_9/io_i_7_in1[7]
+ cb_1_9/io_o_0_co cb_1_9/io_o_0_out[0] cb_1_9/io_o_0_out[1] cb_1_9/io_o_0_out[2]
+ cb_1_9/io_o_0_out[3] cb_1_9/io_o_0_out[4] cb_1_9/io_o_0_out[5] cb_1_9/io_o_0_out[6]
+ cb_1_9/io_o_0_out[7] cb_1_9/io_o_1_co cb_1_9/io_o_1_out[0] cb_1_9/io_o_1_out[1]
+ cb_1_9/io_o_1_out[2] cb_1_9/io_o_1_out[3] cb_1_9/io_o_1_out[4] cb_1_9/io_o_1_out[5]
+ cb_1_9/io_o_1_out[6] cb_1_9/io_o_1_out[7] cb_1_9/io_o_2_co cb_1_9/io_o_2_out[0]
+ cb_1_9/io_o_2_out[1] cb_1_9/io_o_2_out[2] cb_1_9/io_o_2_out[3] cb_1_9/io_o_2_out[4]
+ cb_1_9/io_o_2_out[5] cb_1_9/io_o_2_out[6] cb_1_9/io_o_2_out[7] cb_1_9/io_o_3_co
+ cb_1_9/io_o_3_out[0] cb_1_9/io_o_3_out[1] cb_1_9/io_o_3_out[2] cb_1_9/io_o_3_out[3]
+ cb_1_9/io_o_3_out[4] cb_1_9/io_o_3_out[5] cb_1_9/io_o_3_out[6] cb_1_9/io_o_3_out[7]
+ cb_1_9/io_o_4_co cb_1_9/io_o_4_out[0] cb_1_9/io_o_4_out[1] cb_1_9/io_o_4_out[2]
+ cb_1_9/io_o_4_out[3] cb_1_9/io_o_4_out[4] cb_1_9/io_o_4_out[5] cb_1_9/io_o_4_out[6]
+ cb_1_9/io_o_4_out[7] cb_1_9/io_o_5_co cb_1_9/io_o_5_out[0] cb_1_9/io_o_5_out[1]
+ cb_1_9/io_o_5_out[2] cb_1_9/io_o_5_out[3] cb_1_9/io_o_5_out[4] cb_1_9/io_o_5_out[5]
+ cb_1_9/io_o_5_out[6] cb_1_9/io_o_5_out[7] cb_1_9/io_o_6_co cb_1_9/io_o_6_out[0]
+ cb_1_9/io_o_6_out[1] cb_1_9/io_o_6_out[2] cb_1_9/io_o_6_out[3] cb_1_9/io_o_6_out[4]
+ cb_1_9/io_o_6_out[5] cb_1_9/io_o_6_out[6] cb_1_9/io_o_6_out[7] cb_1_9/io_o_7_co
+ cb_1_9/io_o_7_out[0] cb_1_9/io_o_7_out[1] cb_1_9/io_o_7_out[2] cb_1_9/io_o_7_out[3]
+ cb_1_9/io_o_7_out[4] cb_1_9/io_o_7_out[5] cb_1_9/io_o_7_out[6] cb_1_9/io_o_7_out[7]
+ cb_1_9/io_vci cb_1_9/io_vco cb_1_9/io_vi cb_1_9/io_we_i cb_1_9/io_wo[0] cb_1_9/io_wo[10]
+ cb_1_9/io_wo[11] cb_1_9/io_wo[12] cb_1_9/io_wo[13] cb_1_9/io_wo[14] cb_1_9/io_wo[15]
+ cb_1_9/io_wo[16] cb_1_9/io_wo[17] cb_1_9/io_wo[18] cb_1_9/io_wo[19] cb_1_9/io_wo[1]
+ cb_1_9/io_wo[20] cb_1_9/io_wo[21] cb_1_9/io_wo[22] cb_1_9/io_wo[23] cb_1_9/io_wo[24]
+ cb_1_9/io_wo[25] cb_1_9/io_wo[26] cb_1_9/io_wo[27] cb_1_9/io_wo[28] cb_1_9/io_wo[29]
+ cb_1_9/io_wo[2] cb_1_9/io_wo[30] cb_1_9/io_wo[31] cb_1_9/io_wo[32] cb_1_9/io_wo[33]
+ cb_1_9/io_wo[34] cb_1_9/io_wo[35] cb_1_9/io_wo[36] cb_1_9/io_wo[37] cb_1_9/io_wo[38]
+ cb_1_9/io_wo[39] cb_1_9/io_wo[3] cb_1_9/io_wo[40] cb_1_9/io_wo[41] cb_1_9/io_wo[42]
+ cb_1_9/io_wo[43] cb_1_9/io_wo[44] cb_1_9/io_wo[45] cb_1_9/io_wo[46] cb_1_9/io_wo[47]
+ cb_1_9/io_wo[48] cb_1_9/io_wo[49] cb_1_9/io_wo[4] cb_1_9/io_wo[50] cb_1_9/io_wo[51]
+ cb_1_9/io_wo[52] cb_1_9/io_wo[53] cb_1_9/io_wo[54] cb_1_9/io_wo[55] cb_1_9/io_wo[56]
+ cb_1_9/io_wo[57] cb_1_9/io_wo[58] cb_1_9/io_wo[59] cb_1_9/io_wo[5] cb_1_9/io_wo[60]
+ cb_1_9/io_wo[61] cb_1_9/io_wo[62] cb_1_9/io_wo[63] cb_1_9/io_wo[6] cb_1_9/io_wo[7]
+ cb_1_9/io_wo[8] cb_1_9/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xcb_6_0 cb_6_9/io_adr_i[0] cb_6_9/io_adr_i[1] cb_6_0/io_cs_i cb_6_9/io_dat_i[0] cb_6_9/io_dat_i[10]
+ cb_6_9/io_dat_i[11] cb_6_9/io_dat_i[12] cb_6_9/io_dat_i[13] cb_6_9/io_dat_i[14]
+ cb_6_9/io_dat_i[15] cb_6_9/io_dat_i[1] cb_6_9/io_dat_i[2] cb_6_9/io_dat_i[3] cb_6_9/io_dat_i[4]
+ cb_6_9/io_dat_i[5] cb_6_9/io_dat_i[6] cb_6_9/io_dat_i[7] cb_6_9/io_dat_i[8] cb_6_9/io_dat_i[9]
+ cb_6_0/io_dat_o[0] cb_6_0/io_dat_o[10] cb_6_0/io_dat_o[11] cb_6_0/io_dat_o[12] cb_6_0/io_dat_o[13]
+ cb_6_0/io_dat_o[14] cb_6_0/io_dat_o[15] cb_6_0/io_dat_o[1] cb_6_0/io_dat_o[2] cb_6_0/io_dat_o[3]
+ cb_6_0/io_dat_o[4] cb_6_0/io_dat_o[5] cb_6_0/io_dat_o[6] cb_6_0/io_dat_o[7] cb_6_0/io_dat_o[8]
+ cb_6_0/io_dat_o[9] cb_6_1/io_wo[0] cb_6_1/io_wo[10] cb_6_1/io_wo[11] cb_6_1/io_wo[12]
+ cb_6_1/io_wo[13] cb_6_1/io_wo[14] cb_6_1/io_wo[15] cb_6_1/io_wo[16] cb_6_1/io_wo[17]
+ cb_6_1/io_wo[18] cb_6_1/io_wo[19] cb_6_1/io_wo[1] cb_6_1/io_wo[20] cb_6_1/io_wo[21]
+ cb_6_1/io_wo[22] cb_6_1/io_wo[23] cb_6_1/io_wo[24] cb_6_1/io_wo[25] cb_6_1/io_wo[26]
+ cb_6_1/io_wo[27] cb_6_1/io_wo[28] cb_6_1/io_wo[29] cb_6_1/io_wo[2] cb_6_1/io_wo[30]
+ cb_6_1/io_wo[31] cb_6_1/io_wo[32] cb_6_1/io_wo[33] cb_6_1/io_wo[34] cb_6_1/io_wo[35]
+ cb_6_1/io_wo[36] cb_6_1/io_wo[37] cb_6_1/io_wo[38] cb_6_1/io_wo[39] cb_6_1/io_wo[3]
+ cb_6_1/io_wo[40] cb_6_1/io_wo[41] cb_6_1/io_wo[42] cb_6_1/io_wo[43] cb_6_1/io_wo[44]
+ cb_6_1/io_wo[45] cb_6_1/io_wo[46] cb_6_1/io_wo[47] cb_6_1/io_wo[48] cb_6_1/io_wo[49]
+ cb_6_1/io_wo[4] cb_6_1/io_wo[50] cb_6_1/io_wo[51] cb_6_1/io_wo[52] cb_6_1/io_wo[53]
+ cb_6_1/io_wo[54] cb_6_1/io_wo[55] cb_6_1/io_wo[56] cb_6_1/io_wo[57] cb_6_1/io_wo[58]
+ cb_6_1/io_wo[59] cb_6_1/io_wo[5] cb_6_1/io_wo[60] cb_6_1/io_wo[61] cb_6_1/io_wo[62]
+ cb_6_1/io_wo[63] cb_6_1/io_wo[6] cb_6_1/io_wo[7] cb_6_1/io_wo[8] cb_6_1/io_wo[9]
+ ccon_6/io_dsi_o cb_6_0/io_i_0_in1[0] cb_6_0/io_i_0_in1[1] cb_6_0/io_i_0_in1[2] cb_6_0/io_i_0_in1[3]
+ cb_6_0/io_i_0_in1[4] cb_6_0/io_i_0_in1[5] cb_6_0/io_i_0_in1[6] cb_6_0/io_i_0_in1[7]
+ cb_6_0/io_i_1_ci cb_6_0/io_i_1_in1[0] cb_6_0/io_i_1_in1[1] cb_6_0/io_i_1_in1[2]
+ cb_6_0/io_i_1_in1[3] cb_6_0/io_i_1_in1[4] cb_6_0/io_i_1_in1[5] cb_6_0/io_i_1_in1[6]
+ cb_6_0/io_i_1_in1[7] cb_6_0/io_i_2_ci cb_6_0/io_i_2_in1[0] cb_6_0/io_i_2_in1[1]
+ cb_6_0/io_i_2_in1[2] cb_6_0/io_i_2_in1[3] cb_6_0/io_i_2_in1[4] cb_6_0/io_i_2_in1[5]
+ cb_6_0/io_i_2_in1[6] cb_6_0/io_i_2_in1[7] cb_6_0/io_i_3_ci cb_6_0/io_i_3_in1[0]
+ cb_6_0/io_i_3_in1[1] cb_6_0/io_i_3_in1[2] cb_6_0/io_i_3_in1[3] cb_6_0/io_i_3_in1[4]
+ cb_6_0/io_i_3_in1[5] cb_6_0/io_i_3_in1[6] cb_6_0/io_i_3_in1[7] cb_6_0/io_i_4_ci
+ cb_6_0/io_i_4_in1[0] cb_6_0/io_i_4_in1[1] cb_6_0/io_i_4_in1[2] cb_6_0/io_i_4_in1[3]
+ cb_6_0/io_i_4_in1[4] cb_6_0/io_i_4_in1[5] cb_6_0/io_i_4_in1[6] cb_6_0/io_i_4_in1[7]
+ cb_6_0/io_i_5_ci cb_6_0/io_i_5_in1[0] cb_6_0/io_i_5_in1[1] cb_6_0/io_i_5_in1[2]
+ cb_6_0/io_i_5_in1[3] cb_6_0/io_i_5_in1[4] cb_6_0/io_i_5_in1[5] cb_6_0/io_i_5_in1[6]
+ cb_6_0/io_i_5_in1[7] cb_6_0/io_i_6_ci cb_6_0/io_i_6_in1[0] cb_6_0/io_i_6_in1[1]
+ cb_6_0/io_i_6_in1[2] cb_6_0/io_i_6_in1[3] cb_6_0/io_i_6_in1[4] cb_6_0/io_i_6_in1[5]
+ cb_6_0/io_i_6_in1[6] cb_6_0/io_i_6_in1[7] cb_6_0/io_i_7_ci cb_6_0/io_i_7_in1[0]
+ cb_6_0/io_i_7_in1[1] cb_6_0/io_i_7_in1[2] cb_6_0/io_i_7_in1[3] cb_6_0/io_i_7_in1[4]
+ cb_6_0/io_i_7_in1[5] cb_6_0/io_i_7_in1[6] cb_6_0/io_i_7_in1[7] cb_6_1/io_i_0_ci
+ cb_6_1/io_i_0_in1[0] cb_6_1/io_i_0_in1[1] cb_6_1/io_i_0_in1[2] cb_6_1/io_i_0_in1[3]
+ cb_6_1/io_i_0_in1[4] cb_6_1/io_i_0_in1[5] cb_6_1/io_i_0_in1[6] cb_6_1/io_i_0_in1[7]
+ cb_6_1/io_i_1_ci cb_6_1/io_i_1_in1[0] cb_6_1/io_i_1_in1[1] cb_6_1/io_i_1_in1[2]
+ cb_6_1/io_i_1_in1[3] cb_6_1/io_i_1_in1[4] cb_6_1/io_i_1_in1[5] cb_6_1/io_i_1_in1[6]
+ cb_6_1/io_i_1_in1[7] cb_6_1/io_i_2_ci cb_6_1/io_i_2_in1[0] cb_6_1/io_i_2_in1[1]
+ cb_6_1/io_i_2_in1[2] cb_6_1/io_i_2_in1[3] cb_6_1/io_i_2_in1[4] cb_6_1/io_i_2_in1[5]
+ cb_6_1/io_i_2_in1[6] cb_6_1/io_i_2_in1[7] cb_6_1/io_i_3_ci cb_6_1/io_i_3_in1[0]
+ cb_6_1/io_i_3_in1[1] cb_6_1/io_i_3_in1[2] cb_6_1/io_i_3_in1[3] cb_6_1/io_i_3_in1[4]
+ cb_6_1/io_i_3_in1[5] cb_6_1/io_i_3_in1[6] cb_6_1/io_i_3_in1[7] cb_6_1/io_i_4_ci
+ cb_6_1/io_i_4_in1[0] cb_6_1/io_i_4_in1[1] cb_6_1/io_i_4_in1[2] cb_6_1/io_i_4_in1[3]
+ cb_6_1/io_i_4_in1[4] cb_6_1/io_i_4_in1[5] cb_6_1/io_i_4_in1[6] cb_6_1/io_i_4_in1[7]
+ cb_6_1/io_i_5_ci cb_6_1/io_i_5_in1[0] cb_6_1/io_i_5_in1[1] cb_6_1/io_i_5_in1[2]
+ cb_6_1/io_i_5_in1[3] cb_6_1/io_i_5_in1[4] cb_6_1/io_i_5_in1[5] cb_6_1/io_i_5_in1[6]
+ cb_6_1/io_i_5_in1[7] cb_6_1/io_i_6_ci cb_6_1/io_i_6_in1[0] cb_6_1/io_i_6_in1[1]
+ cb_6_1/io_i_6_in1[2] cb_6_1/io_i_6_in1[3] cb_6_1/io_i_6_in1[4] cb_6_1/io_i_6_in1[5]
+ cb_6_1/io_i_6_in1[6] cb_6_1/io_i_6_in1[7] cb_6_1/io_i_7_ci cb_6_1/io_i_7_in1[0]
+ cb_6_1/io_i_7_in1[1] cb_6_1/io_i_7_in1[2] cb_6_1/io_i_7_in1[3] cb_6_1/io_i_7_in1[4]
+ cb_6_1/io_i_7_in1[5] cb_6_1/io_i_7_in1[6] cb_6_1/io_i_7_in1[7] cb_6_0/io_vci cb_6_1/io_vci
+ cb_6_0/io_vi cb_6_9/io_we_i cb_6_0/io_wo[0] cb_6_0/io_wo[10] cb_6_0/io_wo[11] cb_6_0/io_wo[12]
+ cb_6_0/io_wo[13] cb_6_0/io_wo[14] cb_6_0/io_wo[15] cb_6_0/io_wo[16] cb_6_0/io_wo[17]
+ cb_6_0/io_wo[18] cb_6_0/io_wo[19] cb_6_0/io_wo[1] cb_6_0/io_wo[20] cb_6_0/io_wo[21]
+ cb_6_0/io_wo[22] cb_6_0/io_wo[23] cb_6_0/io_wo[24] cb_6_0/io_wo[25] cb_6_0/io_wo[26]
+ cb_6_0/io_wo[27] cb_6_0/io_wo[28] cb_6_0/io_wo[29] cb_6_0/io_wo[2] cb_6_0/io_wo[30]
+ cb_6_0/io_wo[31] cb_6_0/io_wo[32] cb_6_0/io_wo[33] cb_6_0/io_wo[34] cb_6_0/io_wo[35]
+ cb_6_0/io_wo[36] cb_6_0/io_wo[37] cb_6_0/io_wo[38] cb_6_0/io_wo[39] cb_6_0/io_wo[3]
+ cb_6_0/io_wo[40] cb_6_0/io_wo[41] cb_6_0/io_wo[42] cb_6_0/io_wo[43] cb_6_0/io_wo[44]
+ cb_6_0/io_wo[45] cb_6_0/io_wo[46] cb_6_0/io_wo[47] cb_6_0/io_wo[48] cb_6_0/io_wo[49]
+ cb_6_0/io_wo[4] cb_6_0/io_wo[50] cb_6_0/io_wo[51] cb_6_0/io_wo[52] cb_6_0/io_wo[53]
+ cb_6_0/io_wo[54] cb_6_0/io_wo[55] cb_6_0/io_wo[56] cb_6_0/io_wo[57] cb_6_0/io_wo[58]
+ cb_6_0/io_wo[59] cb_6_0/io_wo[5] cb_6_0/io_wo[60] cb_6_0/io_wo[61] cb_6_0/io_wo[62]
+ cb_6_0/io_wo[63] cb_6_0/io_wo[6] cb_6_0/io_wo[7] cb_6_0/io_wo[8] cb_6_0/io_wo[9]
+ mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
Xmcons_0 mcons_3/clock icon/mt_QEI_ChA_0 icon/mt_QEI_ChB_0 mcons_0/io_irq icon/mt_pwm_h_0
+ icon/mt_pwm_l_0 mcons_0/io_wb_ack_o ccon_7/io_adr_i[0] ccon_7/io_adr_i[10] ccon_7/io_adr_i[11]
+ ccon_7/io_adr_i[1] ccon_7/io_adr_i[2] ccon_7/io_adr_i[3] ccon_7/io_adr_i[4] ccon_7/io_adr_i[5]
+ ccon_7/io_adr_i[6] ccon_7/io_adr_i[7] ccon_7/io_adr_i[8] ccon_7/io_adr_i[9] mcons_0/io_wb_cs_i
+ ccon_7/io_dat_i[0] ccon_7/io_dat_i[10] ccon_7/io_dat_i[11] ccon_7/io_dat_i[12] ccon_7/io_dat_i[13]
+ ccon_7/io_dat_i[14] ccon_7/io_dat_i[15] ccon_7/io_dat_i[16] ccon_7/io_dat_i[17]
+ ccon_7/io_dat_i[18] ccon_7/io_dat_i[19] ccon_7/io_dat_i[1] ccon_7/io_dat_i[20] ccon_7/io_dat_i[21]
+ ccon_7/io_dat_i[22] ccon_7/io_dat_i[23] ccon_7/io_dat_i[24] ccon_7/io_dat_i[25]
+ ccon_7/io_dat_i[26] ccon_7/io_dat_i[27] ccon_7/io_dat_i[28] ccon_7/io_dat_i[29]
+ ccon_7/io_dat_i[2] ccon_7/io_dat_i[30] ccon_7/io_dat_i[31] ccon_7/io_dat_i[3] ccon_7/io_dat_i[4]
+ ccon_7/io_dat_i[5] ccon_7/io_dat_i[6] ccon_7/io_dat_i[7] ccon_7/io_dat_i[8] ccon_7/io_dat_i[9]
+ icon/m_wbs_dat_o_0[0] icon/m_wbs_dat_o_0[10] icon/m_wbs_dat_o_0[11] icon/m_wbs_dat_o_0[12]
+ icon/m_wbs_dat_o_0[13] icon/m_wbs_dat_o_0[14] icon/m_wbs_dat_o_0[15] icon/m_wbs_dat_o_0[16]
+ icon/m_wbs_dat_o_0[17] icon/m_wbs_dat_o_0[18] icon/m_wbs_dat_o_0[19] icon/m_wbs_dat_o_0[1]
+ icon/m_wbs_dat_o_0[20] icon/m_wbs_dat_o_0[21] icon/m_wbs_dat_o_0[22] icon/m_wbs_dat_o_0[23]
+ icon/m_wbs_dat_o_0[24] icon/m_wbs_dat_o_0[25] icon/m_wbs_dat_o_0[26] icon/m_wbs_dat_o_0[27]
+ icon/m_wbs_dat_o_0[28] icon/m_wbs_dat_o_0[29] icon/m_wbs_dat_o_0[2] icon/m_wbs_dat_o_0[30]
+ icon/m_wbs_dat_o_0[31] icon/m_wbs_dat_o_0[3] icon/m_wbs_dat_o_0[4] icon/m_wbs_dat_o_0[5]
+ icon/m_wbs_dat_o_0[6] icon/m_wbs_dat_o_0[7] icon/m_wbs_dat_o_0[8] icon/m_wbs_dat_o_0[9]
+ ccon_7/io_we_i mcons_3/reset vccd1 vssd1 motor_top
Xcb_6_1 cb_6_9/io_adr_i[0] cb_6_9/io_adr_i[1] cb_6_1/io_cs_i cb_6_9/io_dat_i[0] cb_6_9/io_dat_i[10]
+ cb_6_9/io_dat_i[11] cb_6_9/io_dat_i[12] cb_6_9/io_dat_i[13] cb_6_9/io_dat_i[14]
+ cb_6_9/io_dat_i[15] cb_6_9/io_dat_i[1] cb_6_9/io_dat_i[2] cb_6_9/io_dat_i[3] cb_6_9/io_dat_i[4]
+ cb_6_9/io_dat_i[5] cb_6_9/io_dat_i[6] cb_6_9/io_dat_i[7] cb_6_9/io_dat_i[8] cb_6_9/io_dat_i[9]
+ cb_6_1/io_dat_o[0] cb_6_1/io_dat_o[10] cb_6_1/io_dat_o[11] cb_6_1/io_dat_o[12] cb_6_1/io_dat_o[13]
+ cb_6_1/io_dat_o[14] cb_6_1/io_dat_o[15] cb_6_1/io_dat_o[1] cb_6_1/io_dat_o[2] cb_6_1/io_dat_o[3]
+ cb_6_1/io_dat_o[4] cb_6_1/io_dat_o[5] cb_6_1/io_dat_o[6] cb_6_1/io_dat_o[7] cb_6_1/io_dat_o[8]
+ cb_6_1/io_dat_o[9] cb_6_2/io_wo[0] cb_6_2/io_wo[10] cb_6_2/io_wo[11] cb_6_2/io_wo[12]
+ cb_6_2/io_wo[13] cb_6_2/io_wo[14] cb_6_2/io_wo[15] cb_6_2/io_wo[16] cb_6_2/io_wo[17]
+ cb_6_2/io_wo[18] cb_6_2/io_wo[19] cb_6_2/io_wo[1] cb_6_2/io_wo[20] cb_6_2/io_wo[21]
+ cb_6_2/io_wo[22] cb_6_2/io_wo[23] cb_6_2/io_wo[24] cb_6_2/io_wo[25] cb_6_2/io_wo[26]
+ cb_6_2/io_wo[27] cb_6_2/io_wo[28] cb_6_2/io_wo[29] cb_6_2/io_wo[2] cb_6_2/io_wo[30]
+ cb_6_2/io_wo[31] cb_6_2/io_wo[32] cb_6_2/io_wo[33] cb_6_2/io_wo[34] cb_6_2/io_wo[35]
+ cb_6_2/io_wo[36] cb_6_2/io_wo[37] cb_6_2/io_wo[38] cb_6_2/io_wo[39] cb_6_2/io_wo[3]
+ cb_6_2/io_wo[40] cb_6_2/io_wo[41] cb_6_2/io_wo[42] cb_6_2/io_wo[43] cb_6_2/io_wo[44]
+ cb_6_2/io_wo[45] cb_6_2/io_wo[46] cb_6_2/io_wo[47] cb_6_2/io_wo[48] cb_6_2/io_wo[49]
+ cb_6_2/io_wo[4] cb_6_2/io_wo[50] cb_6_2/io_wo[51] cb_6_2/io_wo[52] cb_6_2/io_wo[53]
+ cb_6_2/io_wo[54] cb_6_2/io_wo[55] cb_6_2/io_wo[56] cb_6_2/io_wo[57] cb_6_2/io_wo[58]
+ cb_6_2/io_wo[59] cb_6_2/io_wo[5] cb_6_2/io_wo[60] cb_6_2/io_wo[61] cb_6_2/io_wo[62]
+ cb_6_2/io_wo[63] cb_6_2/io_wo[6] cb_6_2/io_wo[7] cb_6_2/io_wo[8] cb_6_2/io_wo[9]
+ cb_6_1/io_i_0_ci cb_6_1/io_i_0_in1[0] cb_6_1/io_i_0_in1[1] cb_6_1/io_i_0_in1[2]
+ cb_6_1/io_i_0_in1[3] cb_6_1/io_i_0_in1[4] cb_6_1/io_i_0_in1[5] cb_6_1/io_i_0_in1[6]
+ cb_6_1/io_i_0_in1[7] cb_6_1/io_i_1_ci cb_6_1/io_i_1_in1[0] cb_6_1/io_i_1_in1[1]
+ cb_6_1/io_i_1_in1[2] cb_6_1/io_i_1_in1[3] cb_6_1/io_i_1_in1[4] cb_6_1/io_i_1_in1[5]
+ cb_6_1/io_i_1_in1[6] cb_6_1/io_i_1_in1[7] cb_6_1/io_i_2_ci cb_6_1/io_i_2_in1[0]
+ cb_6_1/io_i_2_in1[1] cb_6_1/io_i_2_in1[2] cb_6_1/io_i_2_in1[3] cb_6_1/io_i_2_in1[4]
+ cb_6_1/io_i_2_in1[5] cb_6_1/io_i_2_in1[6] cb_6_1/io_i_2_in1[7] cb_6_1/io_i_3_ci
+ cb_6_1/io_i_3_in1[0] cb_6_1/io_i_3_in1[1] cb_6_1/io_i_3_in1[2] cb_6_1/io_i_3_in1[3]
+ cb_6_1/io_i_3_in1[4] cb_6_1/io_i_3_in1[5] cb_6_1/io_i_3_in1[6] cb_6_1/io_i_3_in1[7]
+ cb_6_1/io_i_4_ci cb_6_1/io_i_4_in1[0] cb_6_1/io_i_4_in1[1] cb_6_1/io_i_4_in1[2]
+ cb_6_1/io_i_4_in1[3] cb_6_1/io_i_4_in1[4] cb_6_1/io_i_4_in1[5] cb_6_1/io_i_4_in1[6]
+ cb_6_1/io_i_4_in1[7] cb_6_1/io_i_5_ci cb_6_1/io_i_5_in1[0] cb_6_1/io_i_5_in1[1]
+ cb_6_1/io_i_5_in1[2] cb_6_1/io_i_5_in1[3] cb_6_1/io_i_5_in1[4] cb_6_1/io_i_5_in1[5]
+ cb_6_1/io_i_5_in1[6] cb_6_1/io_i_5_in1[7] cb_6_1/io_i_6_ci cb_6_1/io_i_6_in1[0]
+ cb_6_1/io_i_6_in1[1] cb_6_1/io_i_6_in1[2] cb_6_1/io_i_6_in1[3] cb_6_1/io_i_6_in1[4]
+ cb_6_1/io_i_6_in1[5] cb_6_1/io_i_6_in1[6] cb_6_1/io_i_6_in1[7] cb_6_1/io_i_7_ci
+ cb_6_1/io_i_7_in1[0] cb_6_1/io_i_7_in1[1] cb_6_1/io_i_7_in1[2] cb_6_1/io_i_7_in1[3]
+ cb_6_1/io_i_7_in1[4] cb_6_1/io_i_7_in1[5] cb_6_1/io_i_7_in1[6] cb_6_1/io_i_7_in1[7]
+ cb_6_2/io_i_0_ci cb_6_2/io_i_0_in1[0] cb_6_2/io_i_0_in1[1] cb_6_2/io_i_0_in1[2]
+ cb_6_2/io_i_0_in1[3] cb_6_2/io_i_0_in1[4] cb_6_2/io_i_0_in1[5] cb_6_2/io_i_0_in1[6]
+ cb_6_2/io_i_0_in1[7] cb_6_2/io_i_1_ci cb_6_2/io_i_1_in1[0] cb_6_2/io_i_1_in1[1]
+ cb_6_2/io_i_1_in1[2] cb_6_2/io_i_1_in1[3] cb_6_2/io_i_1_in1[4] cb_6_2/io_i_1_in1[5]
+ cb_6_2/io_i_1_in1[6] cb_6_2/io_i_1_in1[7] cb_6_2/io_i_2_ci cb_6_2/io_i_2_in1[0]
+ cb_6_2/io_i_2_in1[1] cb_6_2/io_i_2_in1[2] cb_6_2/io_i_2_in1[3] cb_6_2/io_i_2_in1[4]
+ cb_6_2/io_i_2_in1[5] cb_6_2/io_i_2_in1[6] cb_6_2/io_i_2_in1[7] cb_6_2/io_i_3_ci
+ cb_6_2/io_i_3_in1[0] cb_6_2/io_i_3_in1[1] cb_6_2/io_i_3_in1[2] cb_6_2/io_i_3_in1[3]
+ cb_6_2/io_i_3_in1[4] cb_6_2/io_i_3_in1[5] cb_6_2/io_i_3_in1[6] cb_6_2/io_i_3_in1[7]
+ cb_6_2/io_i_4_ci cb_6_2/io_i_4_in1[0] cb_6_2/io_i_4_in1[1] cb_6_2/io_i_4_in1[2]
+ cb_6_2/io_i_4_in1[3] cb_6_2/io_i_4_in1[4] cb_6_2/io_i_4_in1[5] cb_6_2/io_i_4_in1[6]
+ cb_6_2/io_i_4_in1[7] cb_6_2/io_i_5_ci cb_6_2/io_i_5_in1[0] cb_6_2/io_i_5_in1[1]
+ cb_6_2/io_i_5_in1[2] cb_6_2/io_i_5_in1[3] cb_6_2/io_i_5_in1[4] cb_6_2/io_i_5_in1[5]
+ cb_6_2/io_i_5_in1[6] cb_6_2/io_i_5_in1[7] cb_6_2/io_i_6_ci cb_6_2/io_i_6_in1[0]
+ cb_6_2/io_i_6_in1[1] cb_6_2/io_i_6_in1[2] cb_6_2/io_i_6_in1[3] cb_6_2/io_i_6_in1[4]
+ cb_6_2/io_i_6_in1[5] cb_6_2/io_i_6_in1[6] cb_6_2/io_i_6_in1[7] cb_6_2/io_i_7_ci
+ cb_6_2/io_i_7_in1[0] cb_6_2/io_i_7_in1[1] cb_6_2/io_i_7_in1[2] cb_6_2/io_i_7_in1[3]
+ cb_6_2/io_i_7_in1[4] cb_6_2/io_i_7_in1[5] cb_6_2/io_i_7_in1[6] cb_6_2/io_i_7_in1[7]
+ cb_6_1/io_vci cb_6_2/io_vci cb_6_1/io_vi cb_6_9/io_we_i cb_6_1/io_wo[0] cb_6_1/io_wo[10]
+ cb_6_1/io_wo[11] cb_6_1/io_wo[12] cb_6_1/io_wo[13] cb_6_1/io_wo[14] cb_6_1/io_wo[15]
+ cb_6_1/io_wo[16] cb_6_1/io_wo[17] cb_6_1/io_wo[18] cb_6_1/io_wo[19] cb_6_1/io_wo[1]
+ cb_6_1/io_wo[20] cb_6_1/io_wo[21] cb_6_1/io_wo[22] cb_6_1/io_wo[23] cb_6_1/io_wo[24]
+ cb_6_1/io_wo[25] cb_6_1/io_wo[26] cb_6_1/io_wo[27] cb_6_1/io_wo[28] cb_6_1/io_wo[29]
+ cb_6_1/io_wo[2] cb_6_1/io_wo[30] cb_6_1/io_wo[31] cb_6_1/io_wo[32] cb_6_1/io_wo[33]
+ cb_6_1/io_wo[34] cb_6_1/io_wo[35] cb_6_1/io_wo[36] cb_6_1/io_wo[37] cb_6_1/io_wo[38]
+ cb_6_1/io_wo[39] cb_6_1/io_wo[3] cb_6_1/io_wo[40] cb_6_1/io_wo[41] cb_6_1/io_wo[42]
+ cb_6_1/io_wo[43] cb_6_1/io_wo[44] cb_6_1/io_wo[45] cb_6_1/io_wo[46] cb_6_1/io_wo[47]
+ cb_6_1/io_wo[48] cb_6_1/io_wo[49] cb_6_1/io_wo[4] cb_6_1/io_wo[50] cb_6_1/io_wo[51]
+ cb_6_1/io_wo[52] cb_6_1/io_wo[53] cb_6_1/io_wo[54] cb_6_1/io_wo[55] cb_6_1/io_wo[56]
+ cb_6_1/io_wo[57] cb_6_1/io_wo[58] cb_6_1/io_wo[59] cb_6_1/io_wo[5] cb_6_1/io_wo[60]
+ cb_6_1/io_wo[61] cb_6_1/io_wo[62] cb_6_1/io_wo[63] cb_6_1/io_wo[6] cb_6_1/io_wo[7]
+ cb_6_1/io_wo[8] cb_6_1/io_wo[9] mcons_3/clock mcons_3/reset vccd1 vssd1 cic_block
.ends

