* NGSPICE file created from cic_con.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

.subckt cic_con io_ack_o io_adr_i[0] io_adr_i[10] io_adr_i[11] io_adr_i[1] io_adr_i[2]
+ io_adr_i[3] io_adr_i[4] io_adr_i[5] io_adr_i[6] io_adr_i[7] io_adr_i[8] io_adr_i[9]
+ io_b_adr_i[0] io_b_adr_i[1] io_b_cs_i_0 io_b_cs_i_1 io_b_cs_i_10 io_b_cs_i_2 io_b_cs_i_3
+ io_b_cs_i_4 io_b_cs_i_5 io_b_cs_i_6 io_b_cs_i_7 io_b_cs_i_8 io_b_cs_i_9 io_b_dat_i[0]
+ io_b_dat_i[10] io_b_dat_i[11] io_b_dat_i[12] io_b_dat_i[13] io_b_dat_i[14] io_b_dat_i[15]
+ io_b_dat_i[1] io_b_dat_i[2] io_b_dat_i[3] io_b_dat_i[4] io_b_dat_i[5] io_b_dat_i[6]
+ io_b_dat_i[7] io_b_dat_i[8] io_b_dat_i[9] io_b_dat_o_0[0] io_b_dat_o_0[10] io_b_dat_o_0[11]
+ io_b_dat_o_0[12] io_b_dat_o_0[13] io_b_dat_o_0[14] io_b_dat_o_0[15] io_b_dat_o_0[1]
+ io_b_dat_o_0[2] io_b_dat_o_0[3] io_b_dat_o_0[4] io_b_dat_o_0[5] io_b_dat_o_0[6]
+ io_b_dat_o_0[7] io_b_dat_o_0[8] io_b_dat_o_0[9] io_b_dat_o_10[0] io_b_dat_o_10[10]
+ io_b_dat_o_10[11] io_b_dat_o_10[12] io_b_dat_o_10[13] io_b_dat_o_10[14] io_b_dat_o_10[15]
+ io_b_dat_o_10[1] io_b_dat_o_10[2] io_b_dat_o_10[3] io_b_dat_o_10[4] io_b_dat_o_10[5]
+ io_b_dat_o_10[6] io_b_dat_o_10[7] io_b_dat_o_10[8] io_b_dat_o_10[9] io_b_dat_o_1[0]
+ io_b_dat_o_1[10] io_b_dat_o_1[11] io_b_dat_o_1[12] io_b_dat_o_1[13] io_b_dat_o_1[14]
+ io_b_dat_o_1[15] io_b_dat_o_1[1] io_b_dat_o_1[2] io_b_dat_o_1[3] io_b_dat_o_1[4]
+ io_b_dat_o_1[5] io_b_dat_o_1[6] io_b_dat_o_1[7] io_b_dat_o_1[8] io_b_dat_o_1[9]
+ io_b_dat_o_2[0] io_b_dat_o_2[10] io_b_dat_o_2[11] io_b_dat_o_2[12] io_b_dat_o_2[13]
+ io_b_dat_o_2[14] io_b_dat_o_2[15] io_b_dat_o_2[1] io_b_dat_o_2[2] io_b_dat_o_2[3]
+ io_b_dat_o_2[4] io_b_dat_o_2[5] io_b_dat_o_2[6] io_b_dat_o_2[7] io_b_dat_o_2[8]
+ io_b_dat_o_2[9] io_b_dat_o_3[0] io_b_dat_o_3[10] io_b_dat_o_3[11] io_b_dat_o_3[12]
+ io_b_dat_o_3[13] io_b_dat_o_3[14] io_b_dat_o_3[15] io_b_dat_o_3[1] io_b_dat_o_3[2]
+ io_b_dat_o_3[3] io_b_dat_o_3[4] io_b_dat_o_3[5] io_b_dat_o_3[6] io_b_dat_o_3[7]
+ io_b_dat_o_3[8] io_b_dat_o_3[9] io_b_dat_o_4[0] io_b_dat_o_4[10] io_b_dat_o_4[11]
+ io_b_dat_o_4[12] io_b_dat_o_4[13] io_b_dat_o_4[14] io_b_dat_o_4[15] io_b_dat_o_4[1]
+ io_b_dat_o_4[2] io_b_dat_o_4[3] io_b_dat_o_4[4] io_b_dat_o_4[5] io_b_dat_o_4[6]
+ io_b_dat_o_4[7] io_b_dat_o_4[8] io_b_dat_o_4[9] io_b_dat_o_5[0] io_b_dat_o_5[10]
+ io_b_dat_o_5[11] io_b_dat_o_5[12] io_b_dat_o_5[13] io_b_dat_o_5[14] io_b_dat_o_5[15]
+ io_b_dat_o_5[1] io_b_dat_o_5[2] io_b_dat_o_5[3] io_b_dat_o_5[4] io_b_dat_o_5[5]
+ io_b_dat_o_5[6] io_b_dat_o_5[7] io_b_dat_o_5[8] io_b_dat_o_5[9] io_b_dat_o_6[0]
+ io_b_dat_o_6[10] io_b_dat_o_6[11] io_b_dat_o_6[12] io_b_dat_o_6[13] io_b_dat_o_6[14]
+ io_b_dat_o_6[15] io_b_dat_o_6[1] io_b_dat_o_6[2] io_b_dat_o_6[3] io_b_dat_o_6[4]
+ io_b_dat_o_6[5] io_b_dat_o_6[6] io_b_dat_o_6[7] io_b_dat_o_6[8] io_b_dat_o_6[9]
+ io_b_dat_o_7[0] io_b_dat_o_7[10] io_b_dat_o_7[11] io_b_dat_o_7[12] io_b_dat_o_7[13]
+ io_b_dat_o_7[14] io_b_dat_o_7[15] io_b_dat_o_7[1] io_b_dat_o_7[2] io_b_dat_o_7[3]
+ io_b_dat_o_7[4] io_b_dat_o_7[5] io_b_dat_o_7[6] io_b_dat_o_7[7] io_b_dat_o_7[8]
+ io_b_dat_o_7[9] io_b_dat_o_8[0] io_b_dat_o_8[10] io_b_dat_o_8[11] io_b_dat_o_8[12]
+ io_b_dat_o_8[13] io_b_dat_o_8[14] io_b_dat_o_8[15] io_b_dat_o_8[1] io_b_dat_o_8[2]
+ io_b_dat_o_8[3] io_b_dat_o_8[4] io_b_dat_o_8[5] io_b_dat_o_8[6] io_b_dat_o_8[7]
+ io_b_dat_o_8[8] io_b_dat_o_8[9] io_b_dat_o_9[0] io_b_dat_o_9[10] io_b_dat_o_9[11]
+ io_b_dat_o_9[12] io_b_dat_o_9[13] io_b_dat_o_9[14] io_b_dat_o_9[15] io_b_dat_o_9[1]
+ io_b_dat_o_9[2] io_b_dat_o_9[3] io_b_dat_o_9[4] io_b_dat_o_9[5] io_b_dat_o_9[6]
+ io_b_dat_o_9[7] io_b_dat_o_9[8] io_b_dat_o_9[9] io_b_we_i io_cs_i io_dat_i[0] io_dat_i[10]
+ io_dat_i[11] io_dat_i[12] io_dat_i[13] io_dat_i[14] io_dat_i[15] io_dat_i[16] io_dat_i[17]
+ io_dat_i[18] io_dat_i[19] io_dat_i[1] io_dat_i[20] io_dat_i[21] io_dat_i[22] io_dat_i[23]
+ io_dat_i[24] io_dat_i[25] io_dat_i[26] io_dat_i[27] io_dat_i[28] io_dat_i[29] io_dat_i[2]
+ io_dat_i[30] io_dat_i[31] io_dat_i[3] io_dat_i[4] io_dat_i[5] io_dat_i[6] io_dat_i[7]
+ io_dat_i[8] io_dat_i[9] io_dat_o[0] io_dat_o[10] io_dat_o[11] io_dat_o[12] io_dat_o[13]
+ io_dat_o[14] io_dat_o[15] io_dat_o[16] io_dat_o[17] io_dat_o[18] io_dat_o[19] io_dat_o[1]
+ io_dat_o[20] io_dat_o[21] io_dat_o[22] io_dat_o[23] io_dat_o[24] io_dat_o[25] io_dat_o[26]
+ io_dat_o[27] io_dat_o[28] io_dat_o[29] io_dat_o[2] io_dat_o[30] io_dat_o[31] io_dat_o[3]
+ io_dat_o[4] io_dat_o[5] io_dat_o[6] io_dat_o[7] io_dat_o[8] io_dat_o[9] io_dataLastBlock[0]
+ io_dataLastBlock[10] io_dataLastBlock[11] io_dataLastBlock[12] io_dataLastBlock[13]
+ io_dataLastBlock[14] io_dataLastBlock[15] io_dataLastBlock[16] io_dataLastBlock[17]
+ io_dataLastBlock[18] io_dataLastBlock[19] io_dataLastBlock[1] io_dataLastBlock[20]
+ io_dataLastBlock[21] io_dataLastBlock[22] io_dataLastBlock[23] io_dataLastBlock[24]
+ io_dataLastBlock[25] io_dataLastBlock[26] io_dataLastBlock[27] io_dataLastBlock[28]
+ io_dataLastBlock[29] io_dataLastBlock[2] io_dataLastBlock[30] io_dataLastBlock[31]
+ io_dataLastBlock[32] io_dataLastBlock[33] io_dataLastBlock[34] io_dataLastBlock[35]
+ io_dataLastBlock[36] io_dataLastBlock[37] io_dataLastBlock[38] io_dataLastBlock[39]
+ io_dataLastBlock[3] io_dataLastBlock[40] io_dataLastBlock[41] io_dataLastBlock[42]
+ io_dataLastBlock[43] io_dataLastBlock[44] io_dataLastBlock[45] io_dataLastBlock[46]
+ io_dataLastBlock[47] io_dataLastBlock[48] io_dataLastBlock[49] io_dataLastBlock[4]
+ io_dataLastBlock[50] io_dataLastBlock[51] io_dataLastBlock[52] io_dataLastBlock[53]
+ io_dataLastBlock[54] io_dataLastBlock[55] io_dataLastBlock[56] io_dataLastBlock[57]
+ io_dataLastBlock[58] io_dataLastBlock[59] io_dataLastBlock[5] io_dataLastBlock[60]
+ io_dataLastBlock[61] io_dataLastBlock[62] io_dataLastBlock[63] io_dataLastBlock[6]
+ io_dataLastBlock[7] io_dataLastBlock[8] io_dataLastBlock[9] io_dsi_in[0] io_dsi_in[1]
+ io_dsi_in[2] io_dsi_in[3] io_dsi_in[4] io_dsi_in[5] io_dsi_in[6] io_dsi_in[7] io_dsi_o
+ io_irq io_vout[0] io_vout[10] io_vout[1] io_vout[2] io_vout[3] io_vout[4] io_vout[5]
+ io_vout[6] io_vout[7] io_vout[8] io_vout[9] io_we_i wb_clk_i wb_rst_i vccd1 vssd1
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3155_ _3677_/Q _3661_/Q _3645_/Q _3621_/Q _3370_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3155_/X sky130_fd_sc_hd__mux4_2
X_3086_ _2899_/Y _2900_/Y _2897_/Y _2898_/Y _3102_/S0 _3148_/X vssd1 vssd1 vccd1 vccd1
+ _3086_/X sky130_fd_sc_hd__mux4_2
X_2106_ _3700_/Q _2100_/X _1879_/X _2101_/X vssd1 vssd1 vccd1 vccd1 _3700_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2037_ _3743_/Q _2030_/A _1891_/X _2031_/A vssd1 vssd1 vccd1 vccd1 _3743_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2939_ _3449_/Q vssd1 vssd1 vccd1 vccd1 _2939_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_60_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3859_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_76_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3842_ _3845_/CLK _3842_/D vssd1 vssd1 vccd1 vccd1 _3842_/Q sky130_fd_sc_hd__dfxtp_1
X_3773_ _3773_/CLK _3773_/D vssd1 vssd1 vccd1 vccd1 _3773_/Q sky130_fd_sc_hd__dfxtp_1
X_2724_ _2836_/A _2724_/B vssd1 vssd1 vccd1 vccd1 _2724_/X sky130_fd_sc_hd__and2_1
X_2655_ _2661_/A _2969_/X vssd1 vssd1 vccd1 vccd1 _2655_/X sky130_fd_sc_hd__and2_1
X_2586_ _3403_/Q _2583_/X _2540_/X _2584_/X vssd1 vssd1 vccd1 vccd1 _3403_/D sky130_fd_sc_hd__a22o_1
XFILLER_47_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3207_ _3403_/Q _3395_/Q _3387_/Q _3627_/Q _3860_/Q _3861_/Q vssd1 vssd1 vccd1 vccd1
+ _3207_/X sky130_fd_sc_hd__mux4_2
XFILLER_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3138_ _3134_/X _3135_/X _3136_/X _3137_/X _3862_/Q _3863_/Q vssd1 vssd1 vccd1 vccd1
+ _3138_/X sky130_fd_sc_hd__mux4_2
XFILLER_55_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3069_ _2642_/X _3223_/X _3858_/Q vssd1 vssd1 vccd1 vccd1 _3069_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2440_ _3499_/Q _2435_/X _2328_/X _2437_/X vssd1 vssd1 vccd1 vccd1 _3499_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2371_ _3548_/Q _2367_/X _2326_/X _2369_/X vssd1 vssd1 vccd1 vccd1 _3548_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3825_ _3829_/CLK _3825_/D vssd1 vssd1 vccd1 vccd1 _3825_/Q sky130_fd_sc_hd__dfxtp_1
X_3756_ _3826_/CLK _3756_/D vssd1 vssd1 vccd1 vccd1 _3756_/Q sky130_fd_sc_hd__dfxtp_1
X_2707_ _3800_/Q vssd1 vssd1 vccd1 vccd1 _2707_/Y sky130_fd_sc_hd__inv_2
X_3687_ _3687_/CLK _3687_/D vssd1 vssd1 vccd1 vccd1 _3687_/Q sky130_fd_sc_hd__dfxtp_1
X_2638_ _2638_/A _2975_/X vssd1 vssd1 vccd1 vccd1 _2638_/X sky130_fd_sc_hd__and2_1
X_2569_ _3416_/Q _2563_/X _2546_/X _2564_/X vssd1 vssd1 vccd1 vccd1 _3416_/D sky130_fd_sc_hd__a22o_1
XINSDIODE2_4 _3055_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput297 _2942_/X vssd1 vssd1 vccd1 vccd1 io_b_adr_i[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_67_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1940_ _2583_/A vssd1 vssd1 vccd1 vccd1 _1940_/X sky130_fd_sc_hd__buf_2
XFILLER_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1871_ _3817_/Q _1860_/X _1829_/X _1863_/X vssd1 vssd1 vccd1 vccd1 _3817_/D sky130_fd_sc_hd__a22o_1
X_3610_ _3682_/CLK _3610_/D vssd1 vssd1 vccd1 vccd1 _3610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3541_ _3817_/CLK _3541_/D vssd1 vssd1 vccd1 vccd1 _3541_/Q sky130_fd_sc_hd__dfxtp_1
X_3472_ _3826_/CLK _3472_/D vssd1 vssd1 vccd1 vccd1 _3472_/Q sky130_fd_sc_hd__dfxtp_1
X_2423_ _3510_/Q _2416_/A _2364_/X _2417_/A vssd1 vssd1 vccd1 vccd1 _3510_/D sky130_fd_sc_hd__a22o_1
X_2354_ _2949_/A vssd1 vssd1 vccd1 vccd1 _2354_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2285_ _3597_/Q _2282_/X _2155_/X _2284_/X vssd1 vssd1 vccd1 vccd1 _3597_/D sky130_fd_sc_hd__a22o_1
XFILLER_92_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3808_ _3811_/CLK _3808_/D vssd1 vssd1 vccd1 vccd1 _3808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3739_ _3831_/CLK _3739_/D vssd1 vssd1 vccd1 vccd1 _3739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2070_ _3725_/Q _2067_/X _1861_/X _2069_/X vssd1 vssd1 vccd1 vccd1 _3725_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2972_ _2971_/X _2646_/X _2981_/S vssd1 vssd1 vccd1 vccd1 _2972_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1923_ _1972_/A vssd1 vssd1 vccd1 vccd1 _1923_/X sky130_fd_sc_hd__clkbuf_2
X_1854_ _1905_/B vssd1 vssd1 vccd1 vccd1 _1928_/B sky130_fd_sc_hd__inv_2
X_1785_ _1789_/A _3239_/X vssd1 vssd1 vccd1 vccd1 _3856_/D sky130_fd_sc_hd__and2_1
X_3524_ _3832_/CLK _3524_/D vssd1 vssd1 vccd1 vccd1 _3524_/Q sky130_fd_sc_hd__dfxtp_1
X_3455_ _3726_/CLK _3455_/D vssd1 vssd1 vccd1 vccd1 _3455_/Q sky130_fd_sc_hd__dfxtp_1
X_2406_ _3523_/Q _2401_/X _2328_/X _2403_/X vssd1 vssd1 vccd1 vccd1 _3523_/D sky130_fd_sc_hd__a22o_1
X_3386_ _3746_/CLK _3386_/D vssd1 vssd1 vccd1 vccd1 _3386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2337_ _3566_/Q _2333_/X _2297_/X _2334_/X vssd1 vssd1 vccd1 vccd1 _3566_/D sky130_fd_sc_hd__a22o_1
X_2268_ _3607_/Q _2257_/X _2267_/X _2259_/X vssd1 vssd1 vccd1 vccd1 _3607_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2199_ _3651_/Q _2197_/X _2138_/X _2198_/X vssd1 vssd1 vccd1 vccd1 _3651_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3746_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3240_ input17/X input49/X input65/X input81/X _2971_/S _2981_/S vssd1 vssd1 vccd1
+ vccd1 _3240_/X sky130_fd_sc_hd__mux4_1
X_3171_ _3594_/Q _3818_/Q _3546_/Q _3522_/Q _3292_/S0 _3292_/S1 vssd1 vssd1 vccd1
+ vccd1 _3171_/X sky130_fd_sc_hd__mux4_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2122_ _3690_/Q _2116_/X _1869_/X _2118_/X vssd1 vssd1 vccd1 vccd1 _3690_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2053_ _3735_/Q _2050_/X _2017_/X _2051_/X vssd1 vssd1 vccd1 vccd1 _3735_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2955_ _2955_/A vssd1 vssd1 vccd1 vccd1 _2955_/X sky130_fd_sc_hd__clkbuf_1
X_2886_ _3814_/Q vssd1 vssd1 vccd1 vccd1 _2886_/Y sky130_fd_sc_hd__inv_2
X_1906_ _2476_/A _1977_/B _2065_/A _1915_/D vssd1 vssd1 vccd1 vccd1 _2553_/A sky130_fd_sc_hd__or4_4
X_1837_ _1972_/A vssd1 vssd1 vccd1 vccd1 _1837_/X sky130_fd_sc_hd__clkbuf_2
X_1768_ _1768_/A _3008_/X vssd1 vssd1 vccd1 vccd1 _3870_/D sky130_fd_sc_hd__nor2b_4
X_3507_ _3603_/CLK _3507_/D vssd1 vssd1 vccd1 vccd1 _3507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1699_ _3898_/Q _1680_/B _1681_/A _1707_/B vssd1 vssd1 vccd1 vccd1 _1699_/X sky130_fd_sc_hd__o211a_1
X_3438_ _3812_/CLK _3438_/D vssd1 vssd1 vccd1 vccd1 _3438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3369_ _3558_/Q _3710_/Q _3694_/Q _3678_/Q _3372_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3369_/X sky130_fd_sc_hd__mux4_2
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater372 _3132_/S1 vssd1 vssd1 vccd1 vccd1 _3126_/S1 sky130_fd_sc_hd__buf_8
Xrepeater383 _2613_/A vssd1 vssd1 vccd1 vccd1 _3062_/S sky130_fd_sc_hd__buf_8
XFILLER_72_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater394 _1905_/B vssd1 vssd1 vccd1 vccd1 _3372_/S1 sky130_fd_sc_hd__buf_8
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput120 io_b_dat_o_5[5] vssd1 vssd1 vccd1 vccd1 _3315_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput142 io_b_dat_o_7[10] vssd1 vssd1 vccd1 vccd1 _3260_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput131 io_b_dat_o_6[15] vssd1 vssd1 vccd1 vccd1 _3235_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput153 io_b_dat_o_7[6] vssd1 vssd1 vccd1 vccd1 _3302_/A3 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput175 io_b_dat_o_9[11] vssd1 vssd1 vccd1 vccd1 _2974_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput186 io_b_dat_o_9[7] vssd1 vssd1 vccd1 vccd1 _2982_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput164 io_b_dat_o_8[1] vssd1 vssd1 vccd1 vccd1 _2994_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput197 io_dat_i[16] vssd1 vssd1 vccd1 vccd1 input197/X sky130_fd_sc_hd__buf_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2740_ _3781_/Q vssd1 vssd1 vccd1 vccd1 _2740_/Y sky130_fd_sc_hd__inv_2
XPHY_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2671_ _2671_/A _2682_/B vssd1 vssd1 vccd1 vccd1 _2683_/C sky130_fd_sc_hd__or2_4
X_3223_ _3219_/X _3220_/X _3221_/X _3222_/X _3862_/Q _3863_/Q vssd1 vssd1 vccd1 vccd1
+ _3223_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3154_ _3573_/Q _3725_/Q _3709_/Q _3693_/Q _3372_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3154_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2105_ _3701_/Q _2100_/X _1877_/X _2101_/X vssd1 vssd1 vccd1 vccd1 _3701_/D sky130_fd_sc_hd__a22o_1
X_3085_ _2903_/Y _2904_/Y _2901_/Y _2902_/Y _3102_/S0 _3148_/X vssd1 vssd1 vccd1 vccd1
+ _3085_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2036_ _3744_/Q _2030_/X _1889_/X _2031_/X vssd1 vssd1 vccd1 vccd1 _3744_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2938_ _3473_/Q vssd1 vssd1 vccd1 vccd1 _2938_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2869_ _3718_/Q vssd1 vssd1 vccd1 vccd1 _2869_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3841_ _3841_/CLK _3841_/D vssd1 vssd1 vccd1 vccd1 _3841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3772_ _3799_/CLK _3772_/D vssd1 vssd1 vccd1 vccd1 _3772_/Q sky130_fd_sc_hd__dfxtp_1
X_2723_ _3764_/Q vssd1 vssd1 vccd1 vccd1 _2723_/Y sky130_fd_sc_hd__inv_2
X_2654_ _2654_/A _2654_/B vssd1 vssd1 vccd1 vccd1 _2654_/X sky130_fd_sc_hd__and2_1
X_2585_ _3404_/Q _2583_/X _2537_/X _2584_/X vssd1 vssd1 vccd1 vccd1 _3404_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3206_ _3435_/Q _3747_/Q _3419_/Q _3411_/Q _3860_/Q _3232_/S1 vssd1 vssd1 vccd1 vccd1
+ _3206_/X sky130_fd_sc_hd__mux4_1
X_3137_ _2742_/Y _2743_/Y _2744_/Y _2745_/Y _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3137_/X sky130_fd_sc_hd__mux4_2
XFILLER_82_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3068_ _2633_/X _3218_/X _3858_/Q vssd1 vssd1 vccd1 vccd1 _3068_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2019_ _2952_/A vssd1 vssd1 vccd1 vccd1 _2019_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2370_ _3549_/Q _2367_/X _2322_/X _2369_/X vssd1 vssd1 vccd1 vccd1 _3549_/D sky130_fd_sc_hd__a22o_1
XFILLER_78_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3824_ _3827_/CLK _3824_/D vssd1 vssd1 vccd1 vccd1 _3824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3755_ _3826_/CLK _3755_/D vssd1 vssd1 vccd1 vccd1 _3755_/Q sky130_fd_sc_hd__dfxtp_1
X_3686_ _3687_/CLK _3686_/D vssd1 vssd1 vccd1 vccd1 _3686_/Q sky130_fd_sc_hd__dfxtp_1
X_2706_ _3678_/Q vssd1 vssd1 vccd1 vccd1 _2706_/Y sky130_fd_sc_hd__inv_2
X_2637_ _2637_/A _2637_/B vssd1 vssd1 vccd1 vccd1 _2637_/X sky130_fd_sc_hd__and2_1
X_2568_ _3417_/Q _2563_/X _2544_/X _2564_/X vssd1 vssd1 vccd1 vccd1 _3417_/D sky130_fd_sc_hd__a22o_1
Xoutput298 _2943_/X vssd1 vssd1 vccd1 vccd1 io_b_adr_i[1] sky130_fd_sc_hd__clkbuf_2
X_2499_ _3462_/Q _2492_/A _2464_/X _2493_/A vssd1 vssd1 vccd1 vccd1 _3462_/D sky130_fd_sc_hd__a22o_1
XINSDIODE2_5 _3052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_39_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3700_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1870_ _3818_/Q _1860_/X _1869_/X _1863_/X vssd1 vssd1 vccd1 vccd1 _3818_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3540_ _3812_/CLK _3540_/D vssd1 vssd1 vccd1 vccd1 _3540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3471_ _3816_/CLK _3471_/D vssd1 vssd1 vccd1 vccd1 _3471_/Q sky130_fd_sc_hd__dfxtp_1
X_2422_ _3511_/Q _2416_/X _2362_/X _2417_/X vssd1 vssd1 vccd1 vccd1 _3511_/D sky130_fd_sc_hd__a22o_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2353_ _3556_/Q _2350_/X _2351_/X _2352_/X vssd1 vssd1 vccd1 vccd1 _3556_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2284_ _2302_/A vssd1 vssd1 vccd1 vccd1 _2284_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3807_ _3807_/CLK _3807_/D vssd1 vssd1 vccd1 vccd1 _3807_/Q sky130_fd_sc_hd__dfxtp_1
X_1999_ _3763_/Q _1994_/X _1972_/X _1996_/X vssd1 vssd1 vccd1 vccd1 _3763_/D sky130_fd_sc_hd__a22o_1
X_3738_ _3832_/CLK _3738_/D vssd1 vssd1 vccd1 vccd1 _3738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3669_ _3841_/CLK _3669_/D vssd1 vssd1 vccd1 vccd1 _3669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2971_ _2971_/A0 _2971_/A1 _2971_/S vssd1 vssd1 vccd1 vccd1 _2971_/X sky130_fd_sc_hd__mux2_1
X_1922_ _3796_/Q _1916_/X _1921_/X _1919_/X vssd1 vssd1 vccd1 vccd1 _3796_/D sky130_fd_sc_hd__a22o_1
XFILLER_42_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1853_ _2021_/B vssd1 vssd1 vccd1 vccd1 _2181_/B sky130_fd_sc_hd__buf_1
XFILLER_30_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1784_ _1796_/A vssd1 vssd1 vccd1 vccd1 _1789_/A sky130_fd_sc_hd__buf_1
X_3523_ _3831_/CLK _3523_/D vssd1 vssd1 vccd1 vccd1 _3523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3454_ _3812_/CLK _3454_/D vssd1 vssd1 vccd1 vccd1 _3454_/Q sky130_fd_sc_hd__dfxtp_1
X_2405_ _3524_/Q _2401_/X _2326_/X _2403_/X vssd1 vssd1 vccd1 vccd1 _3524_/D sky130_fd_sc_hd__a22o_1
X_3385_ _3896_/CLK _3385_/D vssd1 vssd1 vccd1 vccd1 _3385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2336_ _3567_/Q _2333_/X _2295_/X _2334_/X vssd1 vssd1 vccd1 vccd1 _3567_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2267_ _2945_/A vssd1 vssd1 vccd1 vccd1 _2267_/X sky130_fd_sc_hd__buf_2
XFILLER_37_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2198_ _2198_/A vssd1 vssd1 vccd1 vccd1 _2198_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_54_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3662_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3170_ _3674_/Q _3658_/Q _3642_/Q _3618_/Q _3370_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3170_/X sky130_fd_sc_hd__mux4_2
XFILLER_66_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2121_ _3691_/Q _2116_/X _1867_/X _2118_/X vssd1 vssd1 vccd1 vccd1 _3691_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2052_ _3736_/Q _2050_/X _2015_/X _2051_/X vssd1 vssd1 vccd1 vccd1 _3736_/D sky130_fd_sc_hd__a22o_1
XFILLER_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2954_ _2954_/A vssd1 vssd1 vccd1 vccd1 _2954_/X sky130_fd_sc_hd__clkbuf_1
X_2885_ _3590_/Q vssd1 vssd1 vccd1 vccd1 _2885_/Y sky130_fd_sc_hd__inv_2
X_1905_ _1905_/A _1905_/B vssd1 vssd1 vccd1 vccd1 _2065_/A sky130_fd_sc_hd__or2_2
XFILLER_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1836_ _2953_/A vssd1 vssd1 vccd1 vccd1 _1972_/A sky130_fd_sc_hd__clkbuf_2
X_1767_ _1768_/A _3007_/X vssd1 vssd1 vccd1 vccd1 _3871_/D sky130_fd_sc_hd__nor2b_4
X_3506_ _3603_/CLK _3506_/D vssd1 vssd1 vccd1 vccd1 _3506_/Q sky130_fd_sc_hd__dfxtp_1
X_1698_ _1700_/A vssd1 vssd1 vccd1 vccd1 _3073_/S sky130_fd_sc_hd__buf_2
XFILLER_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3437_ _3829_/CLK _3437_/D vssd1 vssd1 vccd1 vccd1 _3437_/Q sky130_fd_sc_hd__dfxtp_1
X_3368_ _3055_/X _3057_/X _3058_/X _2843_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3368_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2319_ _2510_/D vssd1 vssd1 vccd1 vccd1 _2476_/D sky130_fd_sc_hd__buf_1
X_3299_ _3404_/Q _3396_/Q _3388_/Q _3628_/Q _3364_/S0 _3338_/S1 vssd1 vssd1 vccd1
+ vccd1 _3299_/X sky130_fd_sc_hd__mux4_2
XFILLER_45_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater384 _3373_/S0 vssd1 vssd1 vccd1 vccd1 _2613_/A sky130_fd_sc_hd__buf_8
Xrepeater373 _3148_/X vssd1 vssd1 vccd1 vccd1 _3132_/S1 sky130_fd_sc_hd__buf_12
Xrepeater395 _3357_/S1 vssd1 vssd1 vccd1 vccd1 _1905_/B sky130_fd_sc_hd__buf_8
XFILLER_82_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput110 io_b_dat_o_5[10] vssd1 vssd1 vccd1 vccd1 _3260_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput121 io_b_dat_o_5[6] vssd1 vssd1 vccd1 vccd1 _3302_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput143 io_b_dat_o_7[11] vssd1 vssd1 vccd1 vccd1 _3252_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput154 io_b_dat_o_7[7] vssd1 vssd1 vccd1 vccd1 _3289_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput132 io_b_dat_o_6[1] vssd1 vssd1 vccd1 vccd1 _3367_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput176 io_b_dat_o_9[12] vssd1 vssd1 vccd1 vccd1 _2971_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput165 io_b_dat_o_8[2] vssd1 vssd1 vccd1 vccd1 _2992_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput187 io_b_dat_o_9[8] vssd1 vssd1 vccd1 vccd1 _2980_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput198 io_dat_i[17] vssd1 vssd1 vccd1 vccd1 input198/X sky130_fd_sc_hd__buf_1
XFILLER_44_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2670_ _2686_/A input3/X input2/X vssd1 vssd1 vccd1 vccd1 _2682_/B sky130_fd_sc_hd__or3b_4
XFILLER_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3222_ _3400_/Q _3392_/Q _3384_/Q _3624_/Q _3860_/Q _3861_/Q vssd1 vssd1 vccd1 vccd1
+ _3222_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3153_ _3149_/X _3150_/X _3151_/X _3152_/X _3862_/Q _3863_/Q vssd1 vssd1 vccd1 vccd1
+ _3153_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2104_ _3702_/Q _2100_/X _2019_/X _2101_/X vssd1 vssd1 vccd1 vccd1 _3702_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3084_ _2907_/Y _2908_/Y _2905_/Y _2906_/Y _3102_/S0 _3148_/X vssd1 vssd1 vccd1 vccd1
+ _3084_/X sky130_fd_sc_hd__mux4_2
X_2035_ _3745_/Q _2030_/X _1887_/X _2031_/X vssd1 vssd1 vccd1 vccd1 _3745_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2937_ _3497_/Q vssd1 vssd1 vccd1 vccd1 _2937_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2868_ _3566_/Q vssd1 vssd1 vccd1 vccd1 _2868_/Y sky130_fd_sc_hd__inv_2
X_2799_ _3465_/Q vssd1 vssd1 vccd1 vccd1 _2799_/Y sky130_fd_sc_hd__inv_2
X_1819_ input1/X vssd1 vssd1 vccd1 vccd1 _2510_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_89_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3840_ _3841_/CLK _3840_/D vssd1 vssd1 vccd1 vccd1 _3840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3771_ _3799_/CLK _3771_/D vssd1 vssd1 vccd1 vccd1 _3771_/Q sky130_fd_sc_hd__dfxtp_1
X_2722_ _3792_/Q vssd1 vssd1 vccd1 vccd1 _2722_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2653_ _2654_/A _2653_/B vssd1 vssd1 vccd1 vccd1 _2653_/X sky130_fd_sc_hd__and2_1
X_2584_ _2584_/A vssd1 vssd1 vccd1 vccd1 _2584_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3205_ _3531_/Q _3507_/Q _3483_/Q _3459_/Q _3860_/Q _3232_/S1 vssd1 vssd1 vccd1 vccd1
+ _3205_/X sky130_fd_sc_hd__mux4_2
X_3136_ _2738_/Y _2739_/Y _2740_/Y _2741_/Y _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3136_/X sky130_fd_sc_hd__mux4_1
X_3067_ _2634_/X _3213_/X _3858_/Q vssd1 vssd1 vccd1 vccd1 _3067_/X sky130_fd_sc_hd__mux2_1
X_2018_ _3755_/Q _2010_/X _2017_/X _2013_/X vssd1 vssd1 vccd1 vccd1 _3755_/D sky130_fd_sc_hd__a22o_1
XFILLER_70_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3823_ _3823_/CLK _3823_/D vssd1 vssd1 vccd1 vccd1 _3823_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_9_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3747_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3754_ _3826_/CLK _3754_/D vssd1 vssd1 vccd1 vccd1 _3754_/Q sky130_fd_sc_hd__dfxtp_1
X_3685_ _3720_/CLK _3685_/D vssd1 vssd1 vccd1 vccd1 _3685_/Q sky130_fd_sc_hd__dfxtp_1
X_2705_ _3694_/Q vssd1 vssd1 vccd1 vccd1 _2705_/Y sky130_fd_sc_hd__inv_2
X_2636_ _2644_/A _3178_/X vssd1 vssd1 vccd1 vccd1 _2636_/X sky130_fd_sc_hd__and2_1
XFILLER_87_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2567_ _3418_/Q _2563_/X _2542_/X _2564_/X vssd1 vssd1 vccd1 vccd1 _3418_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_6 _3866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput299 _2685_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_0 sky130_fd_sc_hd__clkbuf_2
X_2498_ _3463_/Q _2492_/X _2462_/X _2493_/X vssd1 vssd1 vccd1 vccd1 _3463_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3119_ _2784_/Y _2785_/Y _2782_/Y _2783_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3119_/X sky130_fd_sc_hd__mux4_2
XFILLER_82_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3470_ _3816_/CLK _3470_/D vssd1 vssd1 vccd1 vccd1 _3470_/Q sky130_fd_sc_hd__dfxtp_1
X_2421_ _3512_/Q _2416_/X _2360_/X _2417_/X vssd1 vssd1 vccd1 vccd1 _3512_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2352_ _2352_/A vssd1 vssd1 vccd1 vccd1 _2352_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2283_ _2301_/A vssd1 vssd1 vccd1 vccd1 _2302_/A sky130_fd_sc_hd__inv_2
XFILLER_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3806_ _3821_/CLK _3806_/D vssd1 vssd1 vccd1 vccd1 _3806_/Q sky130_fd_sc_hd__dfxtp_1
X_1998_ _3764_/Q _1994_/X _1970_/X _1996_/X vssd1 vssd1 vccd1 vccd1 _3764_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3737_ _3741_/CLK _3737_/D vssd1 vssd1 vccd1 vccd1 _3737_/Q sky130_fd_sc_hd__dfxtp_1
X_3668_ _3672_/CLK _3668_/D vssd1 vssd1 vccd1 vccd1 _3668_/Q sky130_fd_sc_hd__dfxtp_1
X_2619_ _2647_/A vssd1 vssd1 vccd1 vccd1 _2681_/A sky130_fd_sc_hd__buf_4
X_3599_ _3743_/CLK _3599_/D vssd1 vssd1 vccd1 vccd1 _3599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2970_ _2970_/A0 _2970_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _2970_/X sky130_fd_sc_hd__mux2_2
XFILLER_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1921_ _1970_/A vssd1 vssd1 vccd1 vccd1 _1921_/X sky130_fd_sc_hd__clkbuf_2
X_1852_ input4/X vssd1 vssd1 vccd1 vccd1 _2281_/A sky130_fd_sc_hd__buf_1
X_1783_ _1783_/A _3236_/X vssd1 vssd1 vccd1 vccd1 _3857_/D sky130_fd_sc_hd__and2_1
X_3522_ _3832_/CLK _3522_/D vssd1 vssd1 vccd1 vccd1 _3522_/Q sky130_fd_sc_hd__dfxtp_1
X_3453_ _3700_/CLK _3453_/D vssd1 vssd1 vccd1 vccd1 _3453_/Q sky130_fd_sc_hd__dfxtp_1
X_2404_ _3525_/Q _2401_/X _2322_/X _2403_/X vssd1 vssd1 vccd1 vccd1 _3525_/D sky130_fd_sc_hd__a22o_1
X_3384_ _3896_/CLK _3384_/D vssd1 vssd1 vccd1 vccd1 _3384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2335_ _3568_/Q _2333_/X _2292_/X _2334_/X vssd1 vssd1 vccd1 vccd1 _3568_/D sky130_fd_sc_hd__a22o_1
X_2266_ _3608_/Q _2257_/X _2265_/X _2259_/X vssd1 vssd1 vccd1 vccd1 _3608_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2197_ _2197_/A vssd1 vssd1 vccd1 vccd1 _2197_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3748_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2120_ _3692_/Q _2116_/X _1865_/X _2118_/X vssd1 vssd1 vccd1 vccd1 _3692_/D sky130_fd_sc_hd__a22o_1
X_2051_ _2058_/A vssd1 vssd1 vccd1 vccd1 _2051_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2953_ _2953_/A vssd1 vssd1 vccd1 vccd1 _2953_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1904_ input1/X vssd1 vssd1 vccd1 vccd1 _1977_/B sky130_fd_sc_hd__clkbuf_2
X_2884_ _3614_/Q vssd1 vssd1 vccd1 vccd1 _2884_/Y sky130_fd_sc_hd__inv_2
X_1835_ _3828_/Q _1827_/X _1834_/X _1831_/X vssd1 vssd1 vccd1 vccd1 _3828_/D sky130_fd_sc_hd__a22o_1
X_1766_ _1768_/A _3006_/X vssd1 vssd1 vccd1 vccd1 _3872_/D sky130_fd_sc_hd__nor2b_4
X_3505_ _3603_/CLK _3505_/D vssd1 vssd1 vccd1 vccd1 _3505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1697_ _1802_/B _1697_/B vssd1 vssd1 vccd1 vccd1 _1700_/A sky130_fd_sc_hd__or2_2
XFILLER_89_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3436_ _3627_/CLK _3436_/D vssd1 vssd1 vccd1 vccd1 _3436_/Q sky130_fd_sc_hd__dfxtp_1
X_3367_ _3367_/A0 _3367_/A1 _3367_/A2 _3367_/A3 _2996_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3367_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2318_ _3574_/Q _2310_/A _2269_/X _2311_/A vssd1 vssd1 vccd1 vccd1 _3574_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3298_ _3436_/Q _3748_/Q _3420_/Q _3412_/Q _3364_/S0 _3338_/S1 vssd1 vssd1 vccd1
+ vccd1 _3298_/X sky130_fd_sc_hd__mux4_1
XFILLER_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater396 input6/X vssd1 vssd1 vccd1 vccd1 _3357_/S1 sky130_fd_sc_hd__buf_8
X_2249_ _2259_/A vssd1 vssd1 vccd1 vccd1 _2249_/X sky130_fd_sc_hd__clkbuf_2
Xrepeater385 input7/X vssd1 vssd1 vccd1 vccd1 _3373_/S0 sky130_fd_sc_hd__buf_8
Xrepeater374 _3143_/X vssd1 vssd1 vccd1 vccd1 _3133_/S0 sky130_fd_sc_hd__buf_12
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput111 io_b_dat_o_5[11] vssd1 vssd1 vccd1 vccd1 _3252_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput100 io_b_dat_o_4[1] vssd1 vssd1 vccd1 vccd1 _3367_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput122 io_b_dat_o_5[7] vssd1 vssd1 vccd1 vccd1 _3289_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput144 io_b_dat_o_7[12] vssd1 vssd1 vccd1 vccd1 _3244_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput133 io_b_dat_o_6[2] vssd1 vssd1 vccd1 vccd1 _3354_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput155 io_b_dat_o_7[8] vssd1 vssd1 vccd1 vccd1 _3276_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput166 io_b_dat_o_8[3] vssd1 vssd1 vccd1 vccd1 _2990_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput177 io_b_dat_o_9[13] vssd1 vssd1 vccd1 vccd1 _2968_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput188 io_b_dat_o_9[9] vssd1 vssd1 vccd1 vccd1 _2978_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput199 io_dat_i[18] vssd1 vssd1 vccd1 vccd1 input199/X sky130_fd_sc_hd__buf_1
XFILLER_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3221_ _3432_/Q _3744_/Q _3416_/Q _3408_/Q _3860_/Q _3861_/Q vssd1 vssd1 vccd1 vccd1
+ _3221_/X sky130_fd_sc_hd__mux4_1
X_3152_ _3786_/Q _3782_/Q _3790_/Q _3762_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3152_/X sky130_fd_sc_hd__mux4_2
XFILLER_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2103_ _3703_/Q _2100_/X _2017_/X _2101_/X vssd1 vssd1 vccd1 vccd1 _3703_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3083_ _3079_/X _3080_/X _3081_/X _3082_/X _3133_/S0 _3138_/X vssd1 vssd1 vccd1 vccd1
+ _3083_/X sky130_fd_sc_hd__mux4_2
X_2034_ _3746_/Q _2030_/X _1885_/X _2031_/X vssd1 vssd1 vccd1 vccd1 _3746_/D sky130_fd_sc_hd__a22o_1
XFILLER_47_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2936_ _3521_/Q vssd1 vssd1 vccd1 vccd1 _2936_/Y sky130_fd_sc_hd__inv_2
X_2867_ _3733_/Q vssd1 vssd1 vccd1 vccd1 _2867_/Y sky130_fd_sc_hd__inv_2
X_1818_ _2039_/A vssd1 vssd1 vccd1 vccd1 _2510_/A sky130_fd_sc_hd__buf_1
X_2798_ _3489_/Q vssd1 vssd1 vccd1 vccd1 _2798_/Y sky130_fd_sc_hd__inv_2
X_1749_ _3882_/Q _1734_/A _2141_/A _1736_/A _1742_/X vssd1 vssd1 vccd1 vccd1 _3882_/D
+ sky130_fd_sc_hd__o221a_1
X_3419_ _3627_/CLK _3419_/D vssd1 vssd1 vccd1 vccd1 _3419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3770_ _3826_/CLK _3770_/D vssd1 vssd1 vccd1 vccd1 _3770_/Q sky130_fd_sc_hd__dfxtp_1
X_2721_ _2721_/A _3193_/X vssd1 vssd1 vccd1 vccd1 _2721_/X sky130_fd_sc_hd__and2_1
XFILLER_12_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2652_ _2664_/A _2970_/X vssd1 vssd1 vccd1 vccd1 _2652_/X sky130_fd_sc_hd__and2_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2583_ _2583_/A vssd1 vssd1 vccd1 vccd1 _2583_/X sky130_fd_sc_hd__clkbuf_2
X_3204_ _3427_/Q _3603_/Q _3579_/Q _3555_/Q _3860_/Q _3232_/S1 vssd1 vssd1 vccd1 vccd1
+ _3204_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3135_ _2734_/Y _2735_/Y _2736_/Y _2737_/Y _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3135_/X sky130_fd_sc_hd__mux4_2
X_3066_ _2635_/Y _3208_/X _3858_/Q vssd1 vssd1 vccd1 vccd1 _3066_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2017_ _2953_/A vssd1 vssd1 vccd1 vccd1 _2017_/X sky130_fd_sc_hd__clkbuf_2
XPHY_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2919_ _3544_/Q vssd1 vssd1 vccd1 vccd1 _2919_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3899_ _3899_/CLK _3899_/D vssd1 vssd1 vccd1 vccd1 _3899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3822_ _3826_/CLK _3822_/D vssd1 vssd1 vccd1 vccd1 _3822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3753_ _3773_/CLK _3753_/D vssd1 vssd1 vccd1 vccd1 _3753_/Q sky130_fd_sc_hd__dfxtp_1
X_2704_ _3763_/Q vssd1 vssd1 vccd1 vccd1 _2704_/Y sky130_fd_sc_hd__inv_2
X_3684_ _3740_/CLK _3684_/D vssd1 vssd1 vccd1 vccd1 _3684_/Q sky130_fd_sc_hd__dfxtp_1
X_2635_ _1715_/A _1715_/B _1716_/B vssd1 vssd1 vccd1 vccd1 _2635_/Y sky130_fd_sc_hd__o21ai_1
X_2566_ _3419_/Q _2563_/X _2540_/X _2564_/X vssd1 vssd1 vccd1 vccd1 _3419_/D sky130_fd_sc_hd__a22o_1
XINSDIODE2_7 _3872_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2497_ _3464_/Q _2492_/X _2460_/X _2493_/X vssd1 vssd1 vccd1 vccd1 _3464_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3118_ _3114_/X _3115_/X _3116_/X _3117_/X _3133_/S0 _3138_/X vssd1 vssd1 vccd1 vccd1
+ _3118_/X sky130_fd_sc_hd__mux4_2
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3049_ _3339_/X _3048_/X _3053_/S vssd1 vssd1 vccd1 vccd1 _3049_/X sky130_fd_sc_hd__mux2_1
XPHY_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_48_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3831_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2420_ _3513_/Q _2416_/X _2358_/X _2417_/X vssd1 vssd1 vccd1 vccd1 _3513_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2351_ _2950_/A vssd1 vssd1 vccd1 vccd1 _2351_/X sky130_fd_sc_hd__clkbuf_2
X_2282_ _2301_/A vssd1 vssd1 vccd1 vccd1 _2282_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1997_ _3765_/Q _1994_/X _1966_/X _1996_/X vssd1 vssd1 vccd1 vccd1 _3765_/D sky130_fd_sc_hd__a22o_1
X_3805_ _3829_/CLK _3805_/D vssd1 vssd1 vccd1 vccd1 _3805_/Q sky130_fd_sc_hd__dfxtp_1
X_3736_ _3826_/CLK _3736_/D vssd1 vssd1 vccd1 vccd1 _3736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3667_ _3667_/CLK _3667_/D vssd1 vssd1 vccd1 vccd1 _3667_/Q sky130_fd_sc_hd__dfxtp_1
X_2618_ _2637_/A _2618_/B vssd1 vssd1 vccd1 vccd1 _2618_/X sky130_fd_sc_hd__and2_1
X_3598_ _3801_/CLK _3598_/D vssd1 vssd1 vccd1 vccd1 _3598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2549_ _3431_/Q _2536_/A _2548_/X _2538_/A vssd1 vssd1 vccd1 vccd1 _3431_/D sky130_fd_sc_hd__a22o_1
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1920_ _3797_/Q _1916_/X _1917_/X _1919_/X vssd1 vssd1 vccd1 vccd1 _3797_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1851_ _3822_/Q _1845_/X _1840_/X _1847_/X vssd1 vssd1 vccd1 vccd1 _3822_/D sky130_fd_sc_hd__a22o_1
X_1782_ _1802_/A _3073_/S vssd1 vssd1 vccd1 vccd1 _3858_/D sky130_fd_sc_hd__nor2_1
X_3521_ _3832_/CLK _3521_/D vssd1 vssd1 vccd1 vccd1 _3521_/Q sky130_fd_sc_hd__dfxtp_1
X_3452_ _3740_/CLK _3452_/D vssd1 vssd1 vccd1 vccd1 _3452_/Q sky130_fd_sc_hd__dfxtp_1
X_3383_ _3895_/CLK _3383_/D vssd1 vssd1 vccd1 vccd1 _3383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2403_ _2417_/A vssd1 vssd1 vccd1 vccd1 _2403_/X sky130_fd_sc_hd__buf_2
XFILLER_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2334_ _2341_/A vssd1 vssd1 vccd1 vccd1 _2334_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2265_ _2946_/A vssd1 vssd1 vccd1 vccd1 _2265_/X sky130_fd_sc_hd__buf_2
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2196_ _3652_/Q _2190_/X _2135_/X _2191_/X vssd1 vssd1 vccd1 vccd1 _3652_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3719_ _3719_/CLK _3719_/D vssd1 vssd1 vccd1 vccd1 _3719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2050_ _2057_/A vssd1 vssd1 vccd1 vccd1 _2050_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2952_ _2952_/A vssd1 vssd1 vccd1 vccd1 _2952_/X sky130_fd_sc_hd__clkbuf_1
X_1903_ _3802_/Q _1897_/X _1840_/X _1899_/X vssd1 vssd1 vccd1 vccd1 _3802_/D sky130_fd_sc_hd__a22o_1
X_2883_ _3638_/Q vssd1 vssd1 vccd1 vccd1 _2883_/Y sky130_fd_sc_hd__inv_2
X_1834_ _1970_/A vssd1 vssd1 vccd1 vccd1 _1834_/X sky130_fd_sc_hd__clkbuf_2
X_1765_ _1768_/A _3005_/X vssd1 vssd1 vccd1 vccd1 _3873_/D sky130_fd_sc_hd__nor2b_4
XFILLER_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3504_ _3530_/CLK _3504_/D vssd1 vssd1 vccd1 vccd1 _3504_/Q sky130_fd_sc_hd__dfxtp_1
X_1696_ _1691_/X _1692_/X _1693_/X _1695_/X vssd1 vssd1 vccd1 vccd1 _1697_/B sky130_fd_sc_hd__o22a_1
X_3435_ _3747_/CLK _3435_/D vssd1 vssd1 vccd1 vccd1 _3435_/Q sky130_fd_sc_hd__dfxtp_1
X_3366_ input20/X input52/X input68/X input84/X _2996_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3366_/X sky130_fd_sc_hd__mux4_1
X_3297_ _3532_/Q _3508_/Q _3484_/Q _3460_/Q _3364_/S0 _1905_/B vssd1 vssd1 vccd1 vccd1
+ _3297_/X sky130_fd_sc_hd__mux4_2
X_2317_ _3575_/Q _2310_/A _2267_/X _2311_/A vssd1 vssd1 vccd1 vccd1 _3575_/D sky130_fd_sc_hd__a22o_1
X_2248_ _2257_/A vssd1 vssd1 vccd1 vccd1 _2248_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater375 _3132_/S0 vssd1 vssd1 vccd1 vccd1 _3126_/S0 sky130_fd_sc_hd__buf_12
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater386 _3338_/S1 vssd1 vssd1 vccd1 vccd1 _3351_/S1 sky130_fd_sc_hd__buf_4
XFILLER_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2179_ _3663_/Q _2173_/X _2147_/X _2174_/X vssd1 vssd1 vccd1 vccd1 _3663_/D sky130_fd_sc_hd__a22o_1
Xrepeater397 _3372_/S0 vssd1 vssd1 vccd1 vccd1 _3292_/S0 sky130_fd_sc_hd__buf_8
XFILLER_53_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput101 io_b_dat_o_4[2] vssd1 vssd1 vccd1 vccd1 _3354_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput123 io_b_dat_o_5[8] vssd1 vssd1 vccd1 vccd1 _3276_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput134 io_b_dat_o_6[3] vssd1 vssd1 vccd1 vccd1 _3341_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput145 io_b_dat_o_7[13] vssd1 vssd1 vccd1 vccd1 _3241_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput112 io_b_dat_o_5[12] vssd1 vssd1 vccd1 vccd1 _3244_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput156 io_b_dat_o_7[9] vssd1 vssd1 vccd1 vccd1 _3268_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput167 io_b_dat_o_8[4] vssd1 vssd1 vccd1 vccd1 _2988_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput178 io_b_dat_o_9[14] vssd1 vssd1 vccd1 vccd1 _2965_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput189 io_cs_i vssd1 vssd1 vccd1 vccd1 _1729_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3220_ _3528_/Q _3504_/Q _3480_/Q _3456_/Q _3860_/Q _3232_/S1 vssd1 vssd1 vccd1 vccd1
+ _3220_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3151_ _3802_/Q _3750_/Q _3778_/Q _3774_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3151_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2102_ _3704_/Q _2100_/X _2015_/X _2101_/X vssd1 vssd1 vccd1 vccd1 _3704_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3082_ _2911_/Y _2912_/Y _2909_/Y _2910_/Y _3102_/S0 _3148_/X vssd1 vssd1 vccd1 vccd1
+ _3082_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2033_ _3747_/Q _2030_/X _1882_/X _2031_/X vssd1 vssd1 vccd1 vccd1 _3747_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2935_ _3545_/Q vssd1 vssd1 vccd1 vccd1 _2935_/Y sky130_fd_sc_hd__inv_2
X_2866_ _3445_/Q vssd1 vssd1 vccd1 vccd1 _2866_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1817_ input4/X vssd1 vssd1 vccd1 vccd1 _2039_/A sky130_fd_sc_hd__inv_2
XFILLER_7_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2797_ _3513_/Q vssd1 vssd1 vccd1 vccd1 _2797_/Y sky130_fd_sc_hd__inv_2
X_1748_ _2948_/A vssd1 vssd1 vccd1 vccd1 _2141_/A sky130_fd_sc_hd__clkbuf_2
X_1679_ _1679_/A _1707_/A vssd1 vssd1 vccd1 vccd1 _1680_/B sky130_fd_sc_hd__nor2_1
X_3418_ _3867_/CLK _3418_/D vssd1 vssd1 vccd1 vccd1 _3418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3349_ _3528_/Q _3504_/Q _3480_/Q _3456_/Q _3351_/S0 _3351_/S1 vssd1 vssd1 vccd1
+ vccd1 _3349_/X sky130_fd_sc_hd__mux4_2
XFILLER_85_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2720_ _3784_/Q vssd1 vssd1 vccd1 vccd1 _2720_/Y sky130_fd_sc_hd__inv_2
X_2651_ _2664_/A _3168_/X vssd1 vssd1 vccd1 vccd1 _2651_/X sky130_fd_sc_hd__and2_1
X_2582_ _3405_/Q _1940_/X _2534_/X _1942_/X vssd1 vssd1 vccd1 vccd1 _3405_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3203_ _3199_/X _3200_/X _3201_/X _3202_/X _3862_/Q _3863_/Q vssd1 vssd1 vccd1 vccd1
+ _3203_/X sky130_fd_sc_hd__mux4_2
XFILLER_79_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3134_ _2730_/Y _2731_/Y _2732_/Y _2733_/Y _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3134_/X sky130_fd_sc_hd__mux4_1
X_3065_ _2627_/X _3203_/X _3858_/Q vssd1 vssd1 vccd1 vccd1 _3065_/X sky130_fd_sc_hd__mux2_1
X_2016_ _3756_/Q _2010_/X _2015_/X _2013_/X vssd1 vssd1 vccd1 vccd1 _3756_/D sky130_fd_sc_hd__a22o_1
XPHY_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2918_ _3816_/Q vssd1 vssd1 vccd1 vccd1 _2918_/Y sky130_fd_sc_hd__inv_2
X_3898_ _3899_/CLK _3898_/D vssd1 vssd1 vccd1 vccd1 _3898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2849_ _3468_/Q vssd1 vssd1 vccd1 vccd1 _2849_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3821_ _3821_/CLK _3821_/D vssd1 vssd1 vccd1 vccd1 _3821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3752_ _3826_/CLK _3752_/D vssd1 vssd1 vccd1 vccd1 _3752_/Q sky130_fd_sc_hd__dfxtp_1
X_2703_ _3791_/Q vssd1 vssd1 vccd1 vccd1 _2703_/Y sky130_fd_sc_hd__inv_2
X_3683_ _3730_/CLK _3683_/D vssd1 vssd1 vccd1 vccd1 _3683_/Q sky130_fd_sc_hd__dfxtp_1
X_2634_ _3892_/Q _1714_/B _1715_/B vssd1 vssd1 vccd1 vccd1 _2634_/X sky130_fd_sc_hd__a21o_1
X_2565_ _3420_/Q _2563_/X _2537_/X _2564_/X vssd1 vssd1 vccd1 vccd1 _3420_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2496_ _3465_/Q _2492_/X _2458_/X _2493_/X vssd1 vssd1 vccd1 vccd1 _3465_/D sky130_fd_sc_hd__a22o_1
XINSDIODE2_8 _3873_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3117_ _2788_/Y _2789_/Y _2786_/Y _2787_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3117_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3048_ _3048_/A0 _3048_/A1 _3060_/S vssd1 vssd1 vccd1 vccd1 _3048_/X sky130_fd_sc_hd__mux2_2
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_17_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3877_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_69_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2350_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2350_/X sky130_fd_sc_hd__clkbuf_2
X_2281_ _2281_/A _2320_/B _2671_/A _2281_/D vssd1 vssd1 vccd1 vccd1 _2301_/A sky130_fd_sc_hd__or4_4
XFILLER_65_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1996_ _2231_/A vssd1 vssd1 vccd1 vccd1 _1996_/X sky130_fd_sc_hd__clkbuf_2
X_3804_ _3827_/CLK _3804_/D vssd1 vssd1 vccd1 vccd1 _3804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3735_ _3799_/CLK _3735_/D vssd1 vssd1 vccd1 vccd1 _3735_/Q sky130_fd_sc_hd__dfxtp_1
X_3666_ _3859_/CLK _3666_/D vssd1 vssd1 vccd1 vccd1 _3666_/Q sky130_fd_sc_hd__dfxtp_1
X_2617_ _2637_/A _2617_/B vssd1 vssd1 vccd1 vccd1 _2617_/X sky130_fd_sc_hd__and2_1
X_3597_ _3724_/CLK _3597_/D vssd1 vssd1 vccd1 vccd1 _3597_/Q sky130_fd_sc_hd__dfxtp_1
X_2548_ _2945_/A vssd1 vssd1 vccd1 vccd1 _2548_/X sky130_fd_sc_hd__clkbuf_2
X_2479_ _2493_/A vssd1 vssd1 vccd1 vccd1 _2479_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1850_ _3823_/Q _1845_/X _1837_/X _1847_/X vssd1 vssd1 vccd1 vccd1 _3823_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1781_ _1802_/A _2686_/A vssd1 vssd1 vccd1 vccd1 _3859_/D sky130_fd_sc_hd__nor2_1
XFILLER_30_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3520_ _3813_/CLK _3520_/D vssd1 vssd1 vccd1 vccd1 _3520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3451_ _3740_/CLK _3451_/D vssd1 vssd1 vccd1 vccd1 _3451_/Q sky130_fd_sc_hd__dfxtp_1
X_3382_ _3890_/CLK _3382_/D vssd1 vssd1 vccd1 vccd1 _3382_/Q sky130_fd_sc_hd__dfxtp_1
X_2402_ _2416_/A vssd1 vssd1 vccd1 vccd1 _2417_/A sky130_fd_sc_hd__inv_2
X_2333_ _2340_/A vssd1 vssd1 vccd1 vccd1 _2333_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2264_ _3609_/Q _2257_/X _2263_/X _2259_/X vssd1 vssd1 vccd1 vccd1 _3609_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2195_ _3653_/Q _2190_/X _2133_/X _2191_/X vssd1 vssd1 vccd1 vccd1 _3653_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1979_ _2310_/A vssd1 vssd1 vccd1 vccd1 _2311_/A sky130_fd_sc_hd__inv_2
X_3718_ _3719_/CLK _3718_/D vssd1 vssd1 vccd1 vccd1 _3718_/Q sky130_fd_sc_hd__dfxtp_1
X_3649_ _3859_/CLK _3649_/D vssd1 vssd1 vccd1 vccd1 _3649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2951_ _2951_/A vssd1 vssd1 vccd1 vccd1 _2951_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3827_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1902_ _3803_/Q _1897_/X _1837_/X _1899_/X vssd1 vssd1 vccd1 vccd1 _3803_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2882_ _3654_/Q vssd1 vssd1 vccd1 vccd1 _2882_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1833_ _2954_/A vssd1 vssd1 vccd1 vccd1 _1970_/A sky130_fd_sc_hd__clkbuf_2
X_1764_ _1768_/A _3004_/X vssd1 vssd1 vccd1 vccd1 _3874_/D sky130_fd_sc_hd__nor2b_4
X_3503_ _3726_/CLK _3503_/D vssd1 vssd1 vccd1 vccd1 _3503_/Q sky130_fd_sc_hd__dfxtp_1
X_1695_ _3889_/Q _1695_/B _3893_/Q _3892_/Q vssd1 vssd1 vccd1 vccd1 _1695_/X sky130_fd_sc_hd__or4_4
X_3434_ _3851_/CLK _3434_/D vssd1 vssd1 vccd1 vccd1 _3434_/Q sky130_fd_sc_hd__dfxtp_1
X_3365_ _3361_/X _3362_/X _3363_/X _3364_/X _2613_/A _3378_/S1 vssd1 vssd1 vccd1 vccd1
+ _3365_/X sky130_fd_sc_hd__mux4_1
X_2316_ _3576_/Q _2310_/X _2265_/X _2311_/X vssd1 vssd1 vccd1 vccd1 _3576_/D sky130_fd_sc_hd__a22o_1
X_3296_ _3428_/Q _3604_/Q _3580_/Q _3556_/Q _3364_/S0 _3338_/S1 vssd1 vssd1 vccd1
+ vccd1 _3296_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2247_ _3617_/Q _2240_/X _2123_/X _2242_/X vssd1 vssd1 vccd1 vccd1 _3617_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater376 _3102_/S0 vssd1 vssd1 vccd1 vccd1 _3132_/S0 sky130_fd_sc_hd__buf_12
Xrepeater387 _1905_/B vssd1 vssd1 vccd1 vccd1 _3338_/S1 sky130_fd_sc_hd__buf_4
X_2178_ _3664_/Q _2173_/X _2145_/X _2174_/X vssd1 vssd1 vccd1 vccd1 _3664_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater398 _3036_/S vssd1 vssd1 vccd1 vccd1 _3060_/S sky130_fd_sc_hd__buf_8
XFILLER_15_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput102 io_b_dat_o_4[3] vssd1 vssd1 vccd1 vccd1 _3341_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput135 io_b_dat_o_6[4] vssd1 vssd1 vccd1 vccd1 _3328_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput113 io_b_dat_o_5[13] vssd1 vssd1 vccd1 vccd1 _3241_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput124 io_b_dat_o_5[9] vssd1 vssd1 vccd1 vccd1 _3268_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput168 io_b_dat_o_8[5] vssd1 vssd1 vccd1 vccd1 _2986_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput146 io_b_dat_o_7[14] vssd1 vssd1 vccd1 vccd1 _3238_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput157 io_b_dat_o_8[0] vssd1 vssd1 vccd1 vccd1 _2996_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput179 io_b_dat_o_9[15] vssd1 vssd1 vccd1 vccd1 _2962_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3150_ _3758_/Q _3794_/Q _3826_/Q _3822_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3150_/X sky130_fd_sc_hd__mux4_2
X_3081_ _2915_/Y _2916_/Y _2913_/Y _2914_/Y _3102_/S0 _3148_/X vssd1 vssd1 vccd1 vccd1
+ _3081_/X sky130_fd_sc_hd__mux4_1
X_2101_ _2108_/A vssd1 vssd1 vccd1 vccd1 _2101_/X sky130_fd_sc_hd__clkbuf_2
X_2032_ _3748_/Q _2030_/X _1879_/X _2031_/X vssd1 vssd1 vccd1 vccd1 _3748_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2934_ _3817_/Q vssd1 vssd1 vccd1 vccd1 _2934_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2865_ _3469_/Q vssd1 vssd1 vccd1 vccd1 _2865_/Y sky130_fd_sc_hd__inv_2
X_1816_ _3133_/X _1816_/B vssd1 vssd1 vccd1 vccd1 _3830_/D sky130_fd_sc_hd__nor2_2
X_2796_ _3537_/Q vssd1 vssd1 vccd1 vccd1 _2796_/Y sky130_fd_sc_hd__inv_2
X_1747_ _3883_/Q _1734_/X _2138_/A _1736_/X _1742_/X vssd1 vssd1 vccd1 vccd1 _3883_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_89_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1678_ _3896_/Q vssd1 vssd1 vccd1 vccd1 _1707_/A sky130_fd_sc_hd__inv_2
X_3417_ _3746_/CLK _3417_/D vssd1 vssd1 vccd1 vccd1 _3417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3348_ _3424_/Q _3600_/Q _3576_/Q _3552_/Q _3351_/S0 _3351_/S1 vssd1 vssd1 vccd1
+ vccd1 _3348_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3279_ _3669_/Q _3653_/Q _3637_/Q _3613_/Q _3292_/S0 _3292_/S1 vssd1 vssd1 vccd1
+ vccd1 _3279_/X sky130_fd_sc_hd__mux4_2
XFILLER_26_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2650_ _2721_/A vssd1 vssd1 vccd1 vccd1 _2664_/A sky130_fd_sc_hd__buf_1
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2581_ _3406_/Q _2573_/A _2550_/X _2574_/A vssd1 vssd1 vccd1 vccd1 _3406_/D sky130_fd_sc_hd__a22o_1
X_3202_ _3404_/Q _3396_/Q _3388_/Q _3628_/Q _3860_/Q _3232_/S1 vssd1 vssd1 vccd1 vccd1
+ _3202_/X sky130_fd_sc_hd__mux4_1
X_3133_ _3129_/X _3130_/X _3131_/X _3132_/X _3133_/S0 _3138_/X vssd1 vssd1 vccd1 vccd1
+ _3133_/X sky130_fd_sc_hd__mux4_2
XFILLER_82_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3064_ _2628_/X _3198_/X _3858_/Q vssd1 vssd1 vccd1 vccd1 _3064_/X sky130_fd_sc_hd__mux2_1
X_2015_ _2954_/A vssd1 vssd1 vccd1 vccd1 _2015_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2917_ _3592_/Q vssd1 vssd1 vccd1 vccd1 _2917_/Y sky130_fd_sc_hd__inv_2
X_3897_ _3897_/CLK _3897_/D vssd1 vssd1 vccd1 vccd1 _3897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2848_ _3492_/Q vssd1 vssd1 vccd1 vccd1 _2848_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2779_ _3808_/Q vssd1 vssd1 vccd1 vccd1 _2779_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3820_ _3832_/CLK _3820_/D vssd1 vssd1 vccd1 vccd1 _3820_/Q sky130_fd_sc_hd__dfxtp_1
X_3751_ _3826_/CLK _3751_/D vssd1 vssd1 vccd1 vccd1 _3751_/Q sky130_fd_sc_hd__dfxtp_1
X_2702_ _3783_/Q vssd1 vssd1 vccd1 vccd1 _2702_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3682_ _3682_/CLK _3682_/D vssd1 vssd1 vccd1 vccd1 _3682_/Q sky130_fd_sc_hd__dfxtp_1
X_2633_ _3891_/Q _1713_/B _1714_/B vssd1 vssd1 vccd1 vccd1 _2633_/X sky130_fd_sc_hd__a21bo_1
X_2564_ _2564_/A vssd1 vssd1 vccd1 vccd1 _2564_/X sky130_fd_sc_hd__clkbuf_2
X_2495_ _3466_/Q _2492_/X _2456_/X _2493_/X vssd1 vssd1 vccd1 vccd1 _3466_/D sky130_fd_sc_hd__a22o_1
XINSDIODE2_9 _3875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3116_ _2792_/Y _2793_/Y _2790_/Y _2791_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3116_/X sky130_fd_sc_hd__mux4_2
X_3047_ _3881_/Q _3334_/X _3053_/S vssd1 vssd1 vccd1 vccd1 _3047_/X sky130_fd_sc_hd__mux2_1
XPHY_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_57_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3676_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2280_ _3598_/Q _2272_/A _2269_/X _2273_/A vssd1 vssd1 vccd1 vccd1 _3598_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3803_ _3827_/CLK _3803_/D vssd1 vssd1 vccd1 vccd1 _3803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1995_ _2230_/A vssd1 vssd1 vccd1 vccd1 _2231_/A sky130_fd_sc_hd__inv_2
XFILLER_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3734_ _3816_/CLK _3734_/D vssd1 vssd1 vccd1 vccd1 _3734_/Q sky130_fd_sc_hd__dfxtp_1
X_3665_ _3859_/CLK _3665_/D vssd1 vssd1 vccd1 vccd1 _3665_/Q sky130_fd_sc_hd__dfxtp_1
X_2616_ _2659_/A vssd1 vssd1 vccd1 vccd1 _2637_/A sky130_fd_sc_hd__clkbuf_2
X_3596_ _3723_/CLK _3596_/D vssd1 vssd1 vccd1 vccd1 _3596_/Q sky130_fd_sc_hd__dfxtp_1
X_2547_ _3432_/Q _2536_/X _2546_/X _2538_/X vssd1 vssd1 vccd1 vccd1 _3432_/D sky130_fd_sc_hd__a22o_1
X_2478_ _2492_/A vssd1 vssd1 vccd1 vccd1 _2493_/A sky130_fd_sc_hd__inv_2
XFILLER_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1780_ _1783_/A _3073_/X vssd1 vssd1 vccd1 vccd1 _3860_/D sky130_fd_sc_hd__and2_1
XFILLER_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3450_ _3740_/CLK _3450_/D vssd1 vssd1 vccd1 vccd1 _3450_/Q sky130_fd_sc_hd__dfxtp_1
X_3381_ _3059_/X _3061_/X _3062_/X _2725_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3381_/X sky130_fd_sc_hd__mux4_1
X_2401_ _2416_/A vssd1 vssd1 vccd1 vccd1 _2401_/X sky130_fd_sc_hd__buf_2
XFILLER_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2332_ _3569_/Q _2321_/X _2289_/X _2324_/X vssd1 vssd1 vccd1 vccd1 _3569_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2263_ _2947_/A vssd1 vssd1 vccd1 vccd1 _2263_/X sky130_fd_sc_hd__buf_2
X_2194_ _3654_/Q _2190_/X _2131_/X _2191_/X vssd1 vssd1 vccd1 vccd1 _3654_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3717_ _3813_/CLK _3717_/D vssd1 vssd1 vccd1 vccd1 _3717_/Q sky130_fd_sc_hd__dfxtp_1
X_1978_ _2310_/A vssd1 vssd1 vccd1 vccd1 _1978_/X sky130_fd_sc_hd__clkbuf_2
X_3648_ _3682_/CLK _3648_/D vssd1 vssd1 vccd1 vccd1 _3648_/Q sky130_fd_sc_hd__dfxtp_1
X_3579_ _3604_/CLK _3579_/D vssd1 vssd1 vccd1 vccd1 _3579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3714_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2950_ _2950_/A vssd1 vssd1 vccd1 vccd1 _2950_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1901_ _3804_/Q _1897_/X _1834_/X _1899_/X vssd1 vssd1 vccd1 vccd1 _3804_/D sky130_fd_sc_hd__a22o_1
X_2881_ _3670_/Q vssd1 vssd1 vccd1 vccd1 _2881_/Y sky130_fd_sc_hd__inv_2
X_1832_ _3829_/Q _1827_/X _1829_/X _1831_/X vssd1 vssd1 vccd1 vccd1 _3829_/D sky130_fd_sc_hd__a22o_1
XPHY_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1763_ _1775_/A vssd1 vssd1 vccd1 vccd1 _1768_/A sky130_fd_sc_hd__buf_4
X_1694_ _3888_/Q vssd1 vssd1 vccd1 vccd1 _1695_/B sky130_fd_sc_hd__inv_2
X_3502_ _3801_/CLK _3502_/D vssd1 vssd1 vccd1 vccd1 _3502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3433_ _3746_/CLK _3433_/D vssd1 vssd1 vccd1 vccd1 _3433_/Q sky130_fd_sc_hd__dfxtp_1
X_3364_ _3399_/Q _3391_/Q _3383_/Q _3623_/Q _3364_/S0 _1905_/B vssd1 vssd1 vccd1 vccd1
+ _3364_/X sky130_fd_sc_hd__mux4_2
X_3295_ _3291_/X _3292_/X _3293_/X _3294_/X _3295_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3295_/X sky130_fd_sc_hd__mux4_2
X_2315_ _3577_/Q _2310_/X _2263_/X _2311_/X vssd1 vssd1 vccd1 vccd1 _3577_/D sky130_fd_sc_hd__a22o_1
X_2246_ _3618_/Q _2240_/X _2163_/X _2242_/X vssd1 vssd1 vccd1 vccd1 _3618_/D sky130_fd_sc_hd__a22o_1
Xrepeater377 _3153_/X vssd1 vssd1 vccd1 vccd1 _3102_/S0 sky130_fd_sc_hd__buf_12
XFILLER_93_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater399 _3009_/S vssd1 vssd1 vccd1 vccd1 _3036_/S sky130_fd_sc_hd__buf_8
X_2177_ _3665_/Q _2173_/X _2143_/X _2174_/X vssd1 vssd1 vccd1 vccd1 _3665_/D sky130_fd_sc_hd__a22o_1
Xrepeater388 _3292_/S1 vssd1 vssd1 vccd1 vccd1 _3192_/S1 sky130_fd_sc_hd__buf_4
XFILLER_41_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput103 io_b_dat_o_4[4] vssd1 vssd1 vccd1 vccd1 _3328_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput136 io_b_dat_o_6[5] vssd1 vssd1 vccd1 vccd1 _3315_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput114 io_b_dat_o_5[14] vssd1 vssd1 vccd1 vccd1 _3238_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput125 io_b_dat_o_6[0] vssd1 vssd1 vccd1 vccd1 _3380_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput158 io_b_dat_o_8[10] vssd1 vssd1 vccd1 vccd1 _2976_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput169 io_b_dat_o_8[6] vssd1 vssd1 vccd1 vccd1 _2984_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput147 io_b_dat_o_7[15] vssd1 vssd1 vccd1 vccd1 _3235_/A3 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2100_ _2107_/A vssd1 vssd1 vccd1 vccd1 _2100_/X sky130_fd_sc_hd__clkbuf_2
X_3080_ _2919_/Y _2920_/Y _2917_/Y _2918_/Y _3102_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3080_/X sky130_fd_sc_hd__mux4_2
X_2031_ _2031_/A vssd1 vssd1 vccd1 vccd1 _2031_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2933_ _3593_/Q vssd1 vssd1 vccd1 vccd1 _2933_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2864_ _3493_/Q vssd1 vssd1 vccd1 vccd1 _2864_/Y sky130_fd_sc_hd__inv_2
X_1815_ _3128_/X _1816_/B vssd1 vssd1 vccd1 vccd1 _3831_/D sky130_fd_sc_hd__nor2_1
X_2795_ _3809_/Q vssd1 vssd1 vccd1 vccd1 _2795_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1746_ _2949_/A vssd1 vssd1 vccd1 vccd1 _2138_/A sky130_fd_sc_hd__clkbuf_2
X_1677_ _3897_/Q vssd1 vssd1 vccd1 vccd1 _1679_/A sky130_fd_sc_hd__inv_2
X_3416_ _3851_/CLK _3416_/D vssd1 vssd1 vccd1 vccd1 _3416_/Q sky130_fd_sc_hd__dfxtp_1
X_3347_ _3343_/X _3344_/X _3345_/X _3346_/X _3373_/S0 input8/X vssd1 vssd1 vccd1 vccd1
+ _3347_/X sky130_fd_sc_hd__mux4_2
XFILLER_58_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3278_ _3565_/Q _3717_/Q _3701_/Q _3685_/Q _3291_/S0 _3292_/S1 vssd1 vssd1 vccd1
+ vccd1 _3278_/X sky130_fd_sc_hd__mux4_2
XFILLER_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2229_ _3629_/Q _1994_/X _2133_/X _1996_/X vssd1 vssd1 vccd1 vccd1 _3629_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2580_ _3407_/Q _2573_/A _2548_/X _2574_/A vssd1 vssd1 vccd1 vccd1 _3407_/D sky130_fd_sc_hd__a22o_1
X_3201_ _3436_/Q _3748_/Q _3420_/Q _3412_/Q _3860_/Q _3232_/S1 vssd1 vssd1 vccd1 vccd1
+ _3201_/X sky130_fd_sc_hd__mux4_1
X_3132_ _2705_/Y _2706_/Y _2687_/Y _2688_/Y _3132_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3132_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3063_ _1699_/X _3898_/Q _3073_/S vssd1 vssd1 vccd1 vccd1 _3063_/X sky130_fd_sc_hd__mux2_1
X_2014_ _3757_/Q _2010_/X _2011_/X _2013_/X vssd1 vssd1 vccd1 vccd1 _3757_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3896_ _3896_/CLK _3896_/D vssd1 vssd1 vccd1 vccd1 _3896_/Q sky130_fd_sc_hd__dfxtp_1
X_2916_ _3616_/Q vssd1 vssd1 vccd1 vccd1 _2916_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2847_ _3516_/Q vssd1 vssd1 vccd1 vccd1 _2847_/Y sky130_fd_sc_hd__inv_2
X_2778_ _3584_/Q vssd1 vssd1 vccd1 vccd1 _2778_/Y sky130_fd_sc_hd__inv_2
X_1729_ _1729_/A vssd1 vssd1 vccd1 vccd1 _2686_/A sky130_fd_sc_hd__inv_2
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3750_ _3826_/CLK _3750_/D vssd1 vssd1 vccd1 vccd1 _3750_/Q sky130_fd_sc_hd__dfxtp_1
X_2701_ _3787_/Q vssd1 vssd1 vccd1 vccd1 _2701_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3681_ _3730_/CLK _3681_/D vssd1 vssd1 vccd1 vccd1 _3681_/Q sky130_fd_sc_hd__dfxtp_1
X_2632_ _2638_/A _2977_/X vssd1 vssd1 vccd1 vccd1 _2632_/X sky130_fd_sc_hd__and2_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2563_ _2563_/A vssd1 vssd1 vccd1 vccd1 _2563_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2494_ _3467_/Q _2492_/X _2453_/X _2493_/X vssd1 vssd1 vccd1 vccd1 _3467_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3115_ _2796_/Y _2797_/Y _2794_/Y _2795_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3115_/X sky130_fd_sc_hd__mux4_2
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3046_ _3327_/X _3328_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3046_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3879_ _3896_/CLK _3879_/D vssd1 vssd1 vccd1 vccd1 _3879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_26_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3829_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3802_ _3823_/CLK _3802_/D vssd1 vssd1 vccd1 vccd1 _3802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1994_ _2230_/A vssd1 vssd1 vccd1 vccd1 _1994_/X sky130_fd_sc_hd__clkbuf_2
X_3733_ _3773_/CLK _3733_/D vssd1 vssd1 vccd1 vccd1 _3733_/Q sky130_fd_sc_hd__dfxtp_1
X_3664_ _3682_/CLK _3664_/D vssd1 vssd1 vccd1 vccd1 _3664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2615_ _2987_/X _2843_/A vssd1 vssd1 vccd1 vccd1 _2615_/X sky130_fd_sc_hd__and2_1
X_3595_ _3676_/CLK _3595_/D vssd1 vssd1 vccd1 vccd1 _3595_/Q sky130_fd_sc_hd__dfxtp_1
X_2546_ _2946_/A vssd1 vssd1 vccd1 vccd1 _2546_/X sky130_fd_sc_hd__clkbuf_2
X_2477_ _2492_/A vssd1 vssd1 vccd1 vccd1 _2477_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3029_ _3274_/X _3028_/X _3061_/S vssd1 vssd1 vccd1 vccd1 _3029_/X sky130_fd_sc_hd__mux2_2
XFILLER_70_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2400_ _2510_/A _2476_/B _2671_/A _2476_/D vssd1 vssd1 vccd1 vccd1 _2416_/A sky130_fd_sc_hd__or4_4
X_3380_ input93/X _3380_/A1 _3380_/A2 _3380_/A3 _2996_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3380_/X sky130_fd_sc_hd__mux4_1
X_2331_ _3570_/Q _2321_/X _2330_/X _2324_/X vssd1 vssd1 vccd1 vccd1 _3570_/D sky130_fd_sc_hd__a22o_1
X_2262_ _3610_/Q _2257_/X _2261_/X _2259_/X vssd1 vssd1 vccd1 vccd1 _3610_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2193_ _3655_/Q _2190_/X _2129_/X _2191_/X vssd1 vssd1 vccd1 vccd1 _3655_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3716_ _3741_/CLK _3716_/D vssd1 vssd1 vccd1 vccd1 _3716_/Q sky130_fd_sc_hd__dfxtp_1
X_1977_ _1985_/A _1977_/B _2065_/A _2009_/D vssd1 vssd1 vccd1 vccd1 _2310_/A sky130_fd_sc_hd__or4_4
X_3647_ _3667_/CLK _3647_/D vssd1 vssd1 vccd1 vccd1 _3647_/Q sky130_fd_sc_hd__dfxtp_1
X_3578_ _3845_/CLK _3578_/D vssd1 vssd1 vccd1 vccd1 _3578_/Q sky130_fd_sc_hd__dfxtp_1
X_2529_ _3442_/Q _2526_/X _2456_/X _2527_/X vssd1 vssd1 vccd1 vccd1 _3442_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2880_ _2873_/X _2875_/X _2876_/Y _2879_/X vssd1 vssd1 vccd1 vccd1 _2880_/X sky130_fd_sc_hd__a31o_4
XFILLER_70_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1900_ _3805_/Q _1897_/X _1829_/X _1899_/X vssd1 vssd1 vccd1 vccd1 _3805_/D sky130_fd_sc_hd__a22o_1
XPHY_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1831_ _2468_/A vssd1 vssd1 vccd1 vccd1 _1831_/X sky130_fd_sc_hd__buf_2
XPHY_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1762_ _1762_/A _3003_/X vssd1 vssd1 vccd1 vccd1 _3875_/D sky130_fd_sc_hd__nor2b_4
X_1693_ _3895_/Q _3894_/Q _3891_/Q _3890_/Q vssd1 vssd1 vccd1 vccd1 _1693_/X sky130_fd_sc_hd__or4_4
X_3501_ _3741_/CLK _3501_/D vssd1 vssd1 vccd1 vccd1 _3501_/Q sky130_fd_sc_hd__dfxtp_1
X_3432_ _3845_/CLK _3432_/D vssd1 vssd1 vccd1 vccd1 _3432_/Q sky130_fd_sc_hd__dfxtp_1
X_3363_ _3431_/Q _3743_/Q _3415_/Q _3407_/Q _3364_/S0 _1905_/B vssd1 vssd1 vccd1 vccd1
+ _3363_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3816_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3294_ _3492_/Q _3468_/Q _3444_/Q _3732_/Q _3377_/S0 _3294_/S1 vssd1 vssd1 vccd1
+ vccd1 _3294_/X sky130_fd_sc_hd__mux4_1
X_2314_ _3578_/Q _2310_/X _2261_/X _2311_/X vssd1 vssd1 vccd1 vccd1 _3578_/D sky130_fd_sc_hd__a22o_1
X_2245_ _3619_/Q _2240_/X _2161_/X _2242_/X vssd1 vssd1 vccd1 vccd1 _3619_/D sky130_fd_sc_hd__a22o_1
X_2176_ _3666_/Q _2173_/X _2141_/X _2174_/X vssd1 vssd1 vccd1 vccd1 _3666_/D sky130_fd_sc_hd__a22o_1
Xrepeater378 _3861_/Q vssd1 vssd1 vccd1 vccd1 _3232_/S1 sky130_fd_sc_hd__clkbuf_16
Xrepeater389 _2981_/S vssd1 vssd1 vccd1 vccd1 _2997_/S sky130_fd_sc_hd__buf_8
XFILLER_65_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput104 io_b_dat_o_4[5] vssd1 vssd1 vccd1 vccd1 _3315_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput126 io_b_dat_o_6[10] vssd1 vssd1 vccd1 vccd1 _3260_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput115 io_b_dat_o_5[15] vssd1 vssd1 vccd1 vccd1 _3235_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput159 io_b_dat_o_8[11] vssd1 vssd1 vccd1 vccd1 _2974_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput148 io_b_dat_o_7[1] vssd1 vssd1 vccd1 vccd1 _3367_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput137 io_b_dat_o_6[6] vssd1 vssd1 vccd1 vccd1 _3302_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2030_ _2030_/A vssd1 vssd1 vccd1 vccd1 _2030_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2932_ _3617_/Q vssd1 vssd1 vccd1 vccd1 _2932_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2863_ _3517_/Q vssd1 vssd1 vccd1 vccd1 _2863_/Y sky130_fd_sc_hd__inv_2
X_1814_ _3123_/X _1814_/B vssd1 vssd1 vccd1 vccd1 _3832_/D sky130_fd_sc_hd__nor2_1
X_2794_ _3585_/Q vssd1 vssd1 vccd1 vccd1 _2794_/Y sky130_fd_sc_hd__inv_2
X_1745_ _3884_/Q _1734_/X _2135_/A _1736_/X _1742_/X vssd1 vssd1 vccd1 vccd1 _3884_/D
+ sky130_fd_sc_hd__o221a_1
X_3415_ _3743_/CLK _3415_/D vssd1 vssd1 vccd1 vccd1 _3415_/Q sky130_fd_sc_hd__dfxtp_1
X_3346_ _3488_/Q _3464_/Q _3440_/Q _3728_/Q input5/X _3357_/S1 vssd1 vssd1 vccd1 vccd1
+ _3346_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3277_ _2721_/X _3029_/X _3030_/X _2620_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3277_/X sky130_fd_sc_hd__mux4_2
XFILLER_66_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2228_ _3630_/Q _2221_/A _2149_/X _2222_/A vssd1 vssd1 vccd1 vccd1 _3630_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2159_ _2958_/A vssd1 vssd1 vccd1 vccd1 _2159_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3200_ _3532_/Q _3508_/Q _3484_/Q _3460_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3200_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3131_ _2728_/Y _2729_/Y _2726_/Y _2727_/Y _3132_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3131_/X sky130_fd_sc_hd__mux4_2
X_3062_ _3379_/X _3380_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3062_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2013_ _2273_/A vssd1 vssd1 vccd1 vccd1 _2013_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3895_ _3895_/CLK _3895_/D vssd1 vssd1 vccd1 vccd1 _3895_/Q sky130_fd_sc_hd__dfxtp_1
X_2915_ _3640_/Q vssd1 vssd1 vccd1 vccd1 _2915_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2846_ _3540_/Q vssd1 vssd1 vccd1 vccd1 _2846_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2777_ _3608_/Q vssd1 vssd1 vccd1 vccd1 _2777_/Y sky130_fd_sc_hd__inv_2
X_1728_ _3061_/S vssd1 vssd1 vccd1 vccd1 _2721_/A sky130_fd_sc_hd__clkbuf_2
X_3329_ _3043_/X _3045_/X _3046_/X _2656_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3329_/X sky130_fd_sc_hd__mux4_2
XFILLER_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2700_ _3775_/Q vssd1 vssd1 vccd1 vccd1 _2700_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3680_ _3682_/CLK _3680_/D vssd1 vssd1 vccd1 vccd1 _3680_/Q sky130_fd_sc_hd__dfxtp_1
X_2631_ _2637_/A _2631_/B vssd1 vssd1 vccd1 vccd1 _2631_/X sky130_fd_sc_hd__and2_1
X_2562_ _3421_/Q _1957_/X _2534_/X _1959_/X vssd1 vssd1 vccd1 vccd1 _3421_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2493_ _2493_/A vssd1 vssd1 vccd1 vccd1 _2493_/X sky130_fd_sc_hd__buf_2
X_3114_ _2800_/Y _2801_/Y _2798_/Y _2799_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3114_/X sky130_fd_sc_hd__mux4_2
X_3045_ _3326_/X _3044_/X _3053_/S vssd1 vssd1 vccd1 vccd1 _3045_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3878_ _3899_/CLK _3878_/D vssd1 vssd1 vccd1 vccd1 _3878_/Q sky130_fd_sc_hd__dfxtp_1
X_2829_ _3515_/Q vssd1 vssd1 vccd1 vccd1 _2829_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3801_ _3801_/CLK _3801_/D vssd1 vssd1 vccd1 vccd1 _3801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ _2039_/A _2009_/B _2510_/C _2009_/D vssd1 vssd1 vccd1 vccd1 _2230_/A sky130_fd_sc_hd__or4_4
X_3732_ _3773_/CLK _3732_/D vssd1 vssd1 vccd1 vccd1 _3732_/Q sky130_fd_sc_hd__dfxtp_1
X_3663_ _3667_/CLK _3663_/D vssd1 vssd1 vccd1 vccd1 _3663_/Q sky130_fd_sc_hd__dfxtp_1
X_2614_ _2647_/A vssd1 vssd1 vccd1 vccd1 _2843_/A sky130_fd_sc_hd__clkbuf_2
X_3594_ _3723_/CLK _3594_/D vssd1 vssd1 vccd1 vccd1 _3594_/Q sky130_fd_sc_hd__dfxtp_1
X_2545_ _3433_/Q _2536_/X _2544_/X _2538_/X vssd1 vssd1 vccd1 vccd1 _3433_/D sky130_fd_sc_hd__a22o_1
X_2476_ _2476_/A _2476_/B _2682_/A _2476_/D vssd1 vssd1 vccd1 vccd1 _2492_/A sky130_fd_sc_hd__or4_4
XFILLER_18_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3028_ _3028_/A0 _3028_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3028_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2330_ _2956_/A vssd1 vssd1 vccd1 vccd1 _2330_/X sky130_fd_sc_hd__clkbuf_2
X_2261_ _2948_/A vssd1 vssd1 vccd1 vccd1 _2261_/X sky130_fd_sc_hd__buf_2
XFILLER_77_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2192_ _3656_/Q _2190_/X _2126_/X _2191_/X vssd1 vssd1 vccd1 vccd1 _3656_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1976_ _2021_/D vssd1 vssd1 vccd1 vccd1 _2009_/D sky130_fd_sc_hd__buf_1
X_3715_ _3731_/CLK _3715_/D vssd1 vssd1 vccd1 vccd1 _3715_/Q sky130_fd_sc_hd__dfxtp_1
X_3646_ _3662_/CLK _3646_/D vssd1 vssd1 vccd1 vccd1 _3646_/Q sky130_fd_sc_hd__dfxtp_1
X_3577_ _3603_/CLK _3577_/D vssd1 vssd1 vccd1 vccd1 _3577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2528_ _3443_/Q _2526_/X _2453_/X _2527_/X vssd1 vssd1 vccd1 vccd1 _3443_/D sky130_fd_sc_hd__a22o_1
X_2459_ _3489_/Q _2452_/X _2458_/X _2454_/X vssd1 vssd1 vccd1 vccd1 _3489_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ _2467_/A vssd1 vssd1 vccd1 vccd1 _2468_/A sky130_fd_sc_hd__inv_2
XPHY_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1761_ _1762_/A _3002_/X vssd1 vssd1 vccd1 vccd1 _3876_/D sky130_fd_sc_hd__nor2b_4
XFILLER_11_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3500_ _3740_/CLK _3500_/D vssd1 vssd1 vccd1 vccd1 _3500_/Q sky130_fd_sc_hd__dfxtp_1
X_1692_ _3198_/X _3203_/X _3208_/X _3213_/X vssd1 vssd1 vccd1 vccd1 _1692_/X sky130_fd_sc_hd__or4_4
X_3431_ _3748_/CLK _3431_/D vssd1 vssd1 vccd1 vccd1 _3431_/Q sky130_fd_sc_hd__dfxtp_1
X_3362_ _3527_/Q _3503_/Q _3479_/Q _3455_/Q _3364_/S0 _1905_/B vssd1 vssd1 vccd1 vccd1
+ _3362_/X sky130_fd_sc_hd__mux4_2
X_2313_ _3579_/Q _2310_/X _2258_/X _2311_/X vssd1 vssd1 vccd1 vccd1 _3579_/D sky130_fd_sc_hd__a22o_1
X_3293_ _3588_/Q _3812_/Q _3540_/Q _3516_/Q _3377_/S0 _3294_/S1 vssd1 vssd1 vccd1
+ vccd1 _3293_/X sky130_fd_sc_hd__mux4_1
X_2244_ _3620_/Q _2240_/X _2159_/X _2242_/X vssd1 vssd1 vccd1 vccd1 _3620_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2175_ _3667_/Q _2173_/X _2138_/X _2174_/X vssd1 vssd1 vccd1 vccd1 _3667_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_10_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3603_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater379 _3860_/Q vssd1 vssd1 vccd1 vccd1 _3232_/S0 sky130_fd_sc_hd__clkbuf_16
XFILLER_80_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1959_ _2564_/A vssd1 vssd1 vccd1 vccd1 _1959_/X sky130_fd_sc_hd__clkbuf_2
X_3629_ _3796_/CLK _3629_/D vssd1 vssd1 vccd1 vccd1 _3629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput105 io_b_dat_o_4[6] vssd1 vssd1 vccd1 vccd1 _3302_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput127 io_b_dat_o_6[11] vssd1 vssd1 vccd1 vccd1 _3252_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput116 io_b_dat_o_5[1] vssd1 vssd1 vccd1 vccd1 _3367_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput138 io_b_dat_o_6[7] vssd1 vssd1 vccd1 vccd1 _3289_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput149 io_b_dat_o_7[2] vssd1 vssd1 vccd1 vccd1 _3354_/A3 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2931_ _3641_/Q vssd1 vssd1 vccd1 vccd1 _2931_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2862_ _3541_/Q vssd1 vssd1 vccd1 vccd1 _2862_/Y sky130_fd_sc_hd__inv_2
X_2793_ _3609_/Q vssd1 vssd1 vccd1 vccd1 _2793_/Y sky130_fd_sc_hd__inv_2
X_1813_ _3118_/X _1814_/B vssd1 vssd1 vccd1 vccd1 _3833_/D sky130_fd_sc_hd__nor2_1
X_1744_ _2950_/A vssd1 vssd1 vccd1 vccd1 _2135_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3414_ _3829_/CLK _3414_/D vssd1 vssd1 vccd1 vccd1 _3414_/Q sky130_fd_sc_hd__dfxtp_1
X_3345_ _3584_/Q _3808_/Q _3536_/Q _3512_/Q _1905_/A _3357_/S1 vssd1 vssd1 vccd1 vccd1
+ _3345_/X sky130_fd_sc_hd__mux4_2
X_3276_ _3276_/A0 _3276_/A1 _3276_/A2 _3276_/A3 _2984_/S _2981_/S vssd1 vssd1 vccd1
+ vccd1 _3276_/X sky130_fd_sc_hd__mux4_1
X_2227_ _3631_/Q _2221_/X _2147_/X _2222_/X vssd1 vssd1 vccd1 vccd1 _3631_/D sky130_fd_sc_hd__a22o_1
X_2158_ _3677_/Q _2154_/X _2155_/X _2157_/X vssd1 vssd1 vccd1 vccd1 _3677_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2089_ _3710_/Q _2082_/A _1893_/X _2083_/A vssd1 vssd1 vccd1 vccd1 _3710_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3130_ _2748_/Y _2749_/Y _2746_/Y _2747_/Y _3132_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3130_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3061_ _3378_/X _3060_/X _3061_/S vssd1 vssd1 vccd1 vccd1 _3061_/X sky130_fd_sc_hd__mux2_2
XFILLER_82_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2012_ _2272_/A vssd1 vssd1 vccd1 vccd1 _2273_/A sky130_fd_sc_hd__inv_2
XFILLER_90_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3894_ _3895_/CLK _3894_/D vssd1 vssd1 vccd1 vccd1 _3894_/Q sky130_fd_sc_hd__dfxtp_1
X_2914_ _3656_/Q vssd1 vssd1 vccd1 vccd1 _2914_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2845_ _3812_/Q vssd1 vssd1 vccd1 vccd1 _2845_/Y sky130_fd_sc_hd__inv_2
X_2776_ _3632_/Q vssd1 vssd1 vccd1 vccd1 _2776_/Y sky130_fd_sc_hd__inv_2
X_1727_ _1727_/A _3071_/X _1727_/C vssd1 vssd1 vccd1 vccd1 _3888_/D sky130_fd_sc_hd__and3_1
X_3328_ _3328_/A0 _3328_/A1 _3328_/A2 _3328_/A3 _2996_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3328_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3259_ input14/X input46/X input62/X input78/X _2984_/S _2981_/S vssd1 vssd1 vccd1
+ vccd1 _3259_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2630_ _2638_/A _2993_/X vssd1 vssd1 vccd1 vccd1 _2630_/X sky130_fd_sc_hd__and2_1
X_2561_ _3422_/Q _2553_/A _2550_/X _2554_/A vssd1 vssd1 vccd1 vccd1 _3422_/D sky130_fd_sc_hd__a22o_1
X_2492_ _2492_/A vssd1 vssd1 vccd1 vccd1 _2492_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3113_ _3109_/X _3110_/X _3111_/X _3112_/X _3133_/S0 _3138_/X vssd1 vssd1 vccd1 vccd1
+ _3113_/X sky130_fd_sc_hd__mux4_2
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3044_ _3044_/A0 _3044_/A1 _3060_/S vssd1 vssd1 vccd1 vccd1 _3044_/X sky130_fd_sc_hd__mux2_2
XFILLER_82_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3877_ _3877_/CLK _3877_/D vssd1 vssd1 vccd1 vccd1 _3877_/Q sky130_fd_sc_hd__dfxtp_1
X_2828_ _3539_/Q vssd1 vssd1 vccd1 vccd1 _2828_/Y sky130_fd_sc_hd__inv_2
X_2759_ _3647_/Q vssd1 vssd1 vccd1 vccd1 _2759_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3800_ _3827_/CLK _3800_/D vssd1 vssd1 vccd1 vccd1 _3800_/Q sky130_fd_sc_hd__dfxtp_1
X_3731_ _3731_/CLK _3731_/D vssd1 vssd1 vccd1 vccd1 _3731_/Q sky130_fd_sc_hd__dfxtp_1
X_1992_ _3766_/Q _1986_/X _1974_/X _1988_/X vssd1 vssd1 vccd1 vccd1 _3766_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_35_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3823_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3662_ _3662_/CLK _3662_/D vssd1 vssd1 vccd1 vccd1 _3662_/Q sky130_fd_sc_hd__dfxtp_1
X_2613_ _2613_/A vssd1 vssd1 vccd1 vccd1 _2647_/A sky130_fd_sc_hd__inv_2
X_3593_ _3724_/CLK _3593_/D vssd1 vssd1 vccd1 vccd1 _3593_/Q sky130_fd_sc_hd__dfxtp_1
X_2544_ _2947_/A vssd1 vssd1 vccd1 vccd1 _2544_/X sky130_fd_sc_hd__clkbuf_2
X_2475_ _3478_/Q _2467_/A _2464_/X _2468_/A vssd1 vssd1 vccd1 vccd1 _3478_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3027_ _3267_/X _3268_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3027_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2260_ _3611_/Q _2257_/X _2258_/X _2259_/X vssd1 vssd1 vccd1 vccd1 _3611_/D sky130_fd_sc_hd__a22o_1
X_2191_ _2198_/A vssd1 vssd1 vccd1 vccd1 _2191_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1975_ _3774_/Q _1965_/X _1974_/X _1968_/X vssd1 vssd1 vccd1 vccd1 _3774_/D sky130_fd_sc_hd__a22o_1
X_3714_ _3714_/CLK _3714_/D vssd1 vssd1 vccd1 vccd1 _3714_/Q sky130_fd_sc_hd__dfxtp_1
X_3645_ _3677_/CLK _3645_/D vssd1 vssd1 vccd1 vccd1 _3645_/Q sky130_fd_sc_hd__dfxtp_1
X_3576_ _3845_/CLK _3576_/D vssd1 vssd1 vccd1 vccd1 _3576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2527_ _2527_/A vssd1 vssd1 vccd1 vccd1 _2527_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2458_ _2947_/A vssd1 vssd1 vccd1 vccd1 _2458_/X sky130_fd_sc_hd__clkbuf_2
X_2389_ _3534_/Q _2382_/A _2364_/X _2383_/A vssd1 vssd1 vccd1 vccd1 _3534_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1760_ _1762_/A _3001_/X vssd1 vssd1 vccd1 vccd1 _3877_/D sky130_fd_sc_hd__nor2b_4
XPHY_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1691_ _3218_/X _3223_/X _3228_/X _3233_/X vssd1 vssd1 vccd1 vccd1 _1691_/X sky130_fd_sc_hd__or4_4
X_3430_ _3801_/CLK _3430_/D vssd1 vssd1 vccd1 vccd1 _3430_/Q sky130_fd_sc_hd__dfxtp_1
X_3361_ _3423_/Q _3599_/Q _3575_/Q _3551_/Q _3364_/S0 _1905_/B vssd1 vssd1 vccd1 vccd1
+ _3361_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2312_ _3580_/Q _2310_/X _2255_/X _2311_/X vssd1 vssd1 vccd1 vccd1 _3580_/D sky130_fd_sc_hd__a22o_1
X_3292_ _3668_/Q _3652_/Q _3636_/Q _3612_/Q _3292_/S0 _3292_/S1 vssd1 vssd1 vccd1
+ vccd1 _3292_/X sky130_fd_sc_hd__mux4_2
X_2243_ _3621_/Q _2240_/X _2155_/X _2242_/X vssd1 vssd1 vccd1 vccd1 _3621_/D sky130_fd_sc_hd__a22o_1
XFILLER_78_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2174_ _2174_/A vssd1 vssd1 vccd1 vccd1 _2174_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_50_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3740_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1958_ _2563_/A vssd1 vssd1 vccd1 vccd1 _2564_/A sky130_fd_sc_hd__inv_2
X_1889_ _2145_/A vssd1 vssd1 vccd1 vccd1 _1889_/X sky130_fd_sc_hd__clkbuf_2
X_3628_ _3895_/CLK _3628_/D vssd1 vssd1 vccd1 vccd1 _3628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3559_ _3727_/CLK _3559_/D vssd1 vssd1 vccd1 vccd1 _3559_/Q sky130_fd_sc_hd__dfxtp_1
Xinput106 io_b_dat_o_4[7] vssd1 vssd1 vccd1 vccd1 _3289_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput117 io_b_dat_o_5[2] vssd1 vssd1 vccd1 vccd1 _3354_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput128 io_b_dat_o_6[12] vssd1 vssd1 vccd1 vccd1 _3244_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput139 io_b_dat_o_6[8] vssd1 vssd1 vccd1 vccd1 _3276_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2930_ _3657_/Q vssd1 vssd1 vccd1 vccd1 _2930_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2861_ _3813_/Q vssd1 vssd1 vccd1 vccd1 _2861_/Y sky130_fd_sc_hd__inv_2
X_2792_ _3633_/Q vssd1 vssd1 vccd1 vccd1 _2792_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1812_ _3113_/X _1814_/B vssd1 vssd1 vccd1 vccd1 _3834_/D sky130_fd_sc_hd__nor2_1
XPHY_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1743_ _1740_/X _1734_/X _2149_/A _1736_/X _1742_/X vssd1 vssd1 vccd1 vccd1 _3885_/D
+ sky130_fd_sc_hd__o221a_1
X_3413_ _3829_/CLK _3413_/D vssd1 vssd1 vccd1 vccd1 _3413_/Q sky130_fd_sc_hd__dfxtp_1
X_3344_ _3664_/Q _3648_/Q _3632_/Q _3608_/Q input5/X _3357_/S1 vssd1 vssd1 vccd1 vccd1
+ _3344_/X sky130_fd_sc_hd__mux4_2
X_3275_ input27/X input59/X input75/X input91/X _2984_/S _2981_/S vssd1 vssd1 vccd1
+ vccd1 _3275_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2226_ _3632_/Q _2221_/X _2145_/X _2222_/X vssd1 vssd1 vccd1 vccd1 _3632_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2157_ _2174_/A vssd1 vssd1 vccd1 vccd1 _2157_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2088_ _3711_/Q _2082_/X _1891_/X _2083_/X vssd1 vssd1 vccd1 vccd1 _3711_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3060_ _3060_/A0 _3060_/A1 _3060_/S vssd1 vssd1 vccd1 vccd1 _3060_/X sky130_fd_sc_hd__mux2_2
X_2011_ _2955_/A vssd1 vssd1 vccd1 vccd1 _2011_/X sky130_fd_sc_hd__buf_2
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3893_ _3899_/CLK _3893_/D vssd1 vssd1 vccd1 vccd1 _3893_/Q sky130_fd_sc_hd__dfxtp_1
X_2913_ _3672_/Q vssd1 vssd1 vccd1 vccd1 _2913_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2844_ _3588_/Q vssd1 vssd1 vccd1 vccd1 _2844_/Y sky130_fd_sc_hd__inv_2
X_2775_ _3648_/Q vssd1 vssd1 vccd1 vccd1 _2775_/Y sky130_fd_sc_hd__inv_2
X_1726_ _1727_/A _3070_/X _1727_/C vssd1 vssd1 vccd1 vccd1 _3889_/D sky130_fd_sc_hd__and3_1
X_3327_ input23/X input55/X input71/X input87/X _2996_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3327_/X sky130_fd_sc_hd__mux4_1
XFILLER_86_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3258_ _3254_/X _3255_/X _3256_/X _3257_/X _2613_/A _3378_/S1 vssd1 vssd1 vccd1 vccd1
+ _3258_/X sky130_fd_sc_hd__mux4_1
X_2209_ _3645_/Q _2206_/X _2155_/X _2208_/X vssd1 vssd1 vccd1 vccd1 _3645_/D sky130_fd_sc_hd__a22o_1
X_3189_ _3566_/Q _3718_/Q _3702_/Q _3686_/Q _3060_/S _3192_/S1 vssd1 vssd1 vccd1 vccd1
+ _3189_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2560_ _3423_/Q _2553_/A _2548_/X _2554_/A vssd1 vssd1 vccd1 vccd1 _3423_/D sky130_fd_sc_hd__a22o_1
X_2491_ _3468_/Q _2485_/X _2450_/X _2486_/X vssd1 vssd1 vccd1 vccd1 _3468_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3112_ _2804_/Y _2805_/Y _2802_/Y _2803_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3112_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3043_ _3882_/Q _3321_/X _3053_/S vssd1 vssd1 vccd1 vccd1 _3043_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3876_ _3877_/CLK _3876_/D vssd1 vssd1 vccd1 vccd1 _3876_/Q sky130_fd_sc_hd__dfxtp_1
X_2827_ _3811_/Q vssd1 vssd1 vccd1 vccd1 _2827_/Y sky130_fd_sc_hd__inv_2
X_2758_ _3663_/Q vssd1 vssd1 vccd1 vccd1 _2758_/Y sky130_fd_sc_hd__inv_2
X_1709_ _1742_/A vssd1 vssd1 vccd1 vccd1 _1721_/A sky130_fd_sc_hd__buf_1
X_2689_ _3799_/Q vssd1 vssd1 vccd1 vccd1 _2689_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3731_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3730_ _3730_/CLK _3730_/D vssd1 vssd1 vccd1 vccd1 _3730_/Q sky130_fd_sc_hd__dfxtp_1
X_1991_ _3767_/Q _1986_/X _1972_/X _1988_/X vssd1 vssd1 vccd1 vccd1 _3767_/D sky130_fd_sc_hd__a22o_1
X_3661_ _3677_/CLK _3661_/D vssd1 vssd1 vccd1 vccd1 _3661_/Q sky130_fd_sc_hd__dfxtp_1
X_2612_ _2612_/A _2659_/A vssd1 vssd1 vccd1 vccd1 _2612_/X sky130_fd_sc_hd__and2_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3592_ _3813_/CLK _3592_/D vssd1 vssd1 vccd1 vccd1 _3592_/Q sky130_fd_sc_hd__dfxtp_1
X_2543_ _3434_/Q _2536_/X _2542_/X _2538_/X vssd1 vssd1 vccd1 vccd1 _3434_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2474_ _3479_/Q _2467_/A _2462_/X _2468_/A vssd1 vssd1 vccd1 vccd1 _3479_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3026_ _3266_/X _3025_/X _3061_/S vssd1 vssd1 vccd1 vccd1 _3026_/X sky130_fd_sc_hd__mux2_2
XFILLER_36_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3859_ _3859_/CLK _3859_/D vssd1 vssd1 vccd1 vccd1 _3859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2190_ _2197_/A vssd1 vssd1 vccd1 vccd1 _2190_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1974_ _1974_/A vssd1 vssd1 vccd1 vccd1 _1974_/X sky130_fd_sc_hd__clkbuf_2
X_3713_ _3730_/CLK _3713_/D vssd1 vssd1 vccd1 vccd1 _3713_/Q sky130_fd_sc_hd__dfxtp_1
X_3644_ _3676_/CLK _3644_/D vssd1 vssd1 vccd1 vccd1 _3644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3575_ _3743_/CLK _3575_/D vssd1 vssd1 vccd1 vccd1 _3575_/Q sky130_fd_sc_hd__dfxtp_1
X_2526_ _2526_/A vssd1 vssd1 vccd1 vccd1 _2526_/X sky130_fd_sc_hd__clkbuf_2
X_2457_ _3490_/Q _2452_/X _2456_/X _2454_/X vssd1 vssd1 vccd1 vccd1 _3490_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2388_ _3535_/Q _2382_/X _2362_/X _2383_/X vssd1 vssd1 vccd1 vccd1 _3535_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3009_ _3009_/A0 _3009_/A1 _3009_/S vssd1 vssd1 vccd1 vccd1 _3009_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1690_ _3880_/Q vssd1 vssd1 vccd1 vccd1 _1802_/B sky130_fd_sc_hd__inv_2
X_3360_ _3356_/X _3357_/X _3358_/X _3359_/X _3373_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3360_/X sky130_fd_sc_hd__mux4_2
X_2311_ _2311_/A vssd1 vssd1 vccd1 vccd1 _2311_/X sky130_fd_sc_hd__clkbuf_2
X_3291_ _3564_/Q _3716_/Q _3700_/Q _3684_/Q _3291_/S0 _3294_/S1 vssd1 vssd1 vccd1
+ vccd1 _3291_/X sky130_fd_sc_hd__mux4_2
XFILLER_78_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2242_ _2259_/A vssd1 vssd1 vccd1 vccd1 _2242_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2173_ _2173_/A vssd1 vssd1 vccd1 vccd1 _2173_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1957_ _2563_/A vssd1 vssd1 vccd1 vccd1 _1957_/X sky130_fd_sc_hd__clkbuf_2
X_1888_ _3809_/Q _1881_/X _1887_/X _1883_/X vssd1 vssd1 vccd1 vccd1 _3809_/D sky130_fd_sc_hd__a22o_1
X_3627_ _3627_/CLK _3627_/D vssd1 vssd1 vccd1 vccd1 _3627_/Q sky130_fd_sc_hd__dfxtp_1
X_3558_ _3727_/CLK _3558_/D vssd1 vssd1 vccd1 vccd1 _3558_/Q sky130_fd_sc_hd__dfxtp_1
X_2509_ _3454_/Q _2501_/A _2464_/X _2502_/A vssd1 vssd1 vccd1 vccd1 _3454_/D sky130_fd_sc_hd__a22o_1
Xinput107 io_b_dat_o_4[8] vssd1 vssd1 vccd1 vccd1 _3276_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput118 io_b_dat_o_5[3] vssd1 vssd1 vccd1 vccd1 _3341_/A1 sky130_fd_sc_hd__clkbuf_1
X_3489_ _3586_/CLK _3489_/D vssd1 vssd1 vccd1 vccd1 _3489_/Q sky130_fd_sc_hd__dfxtp_1
Xinput129 io_b_dat_o_6[13] vssd1 vssd1 vccd1 vccd1 _3241_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2860_ _3589_/Q vssd1 vssd1 vccd1 vccd1 _2860_/Y sky130_fd_sc_hd__inv_2
X_1811_ _3108_/X _1814_/B vssd1 vssd1 vccd1 vccd1 _3835_/D sky130_fd_sc_hd__nor2_1
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2791_ _3649_/Q vssd1 vssd1 vccd1 vccd1 _2791_/Y sky130_fd_sc_hd__inv_2
XPHY_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1742_ _1742_/A vssd1 vssd1 vccd1 vccd1 _1742_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3412_ _3627_/CLK _3412_/D vssd1 vssd1 vccd1 vccd1 _3412_/Q sky130_fd_sc_hd__dfxtp_1
X_3343_ _3560_/Q _3712_/Q _3696_/Q _3680_/Q input5/X _3357_/S1 vssd1 vssd1 vccd1 vccd1
+ _3343_/X sky130_fd_sc_hd__mux4_2
X_3274_ _3270_/X _3271_/X _3272_/X _3273_/X _2613_/A _3378_/S1 vssd1 vssd1 vccd1 vccd1
+ _3274_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2225_ _3633_/Q _2221_/X _2143_/X _2222_/X vssd1 vssd1 vccd1 vccd1 _3633_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2156_ _2173_/A vssd1 vssd1 vccd1 vccd1 _2174_/A sky130_fd_sc_hd__inv_2
X_2087_ _3712_/Q _2082_/X _1889_/X _2083_/X vssd1 vssd1 vccd1 vccd1 _3712_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2989_ _2988_/X _2653_/X _2997_/S vssd1 vssd1 vccd1 vccd1 _2989_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2010_ _2272_/A vssd1 vssd1 vccd1 vccd1 _2010_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_29_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3796_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2912_ _3688_/Q vssd1 vssd1 vccd1 vccd1 _2912_/Y sky130_fd_sc_hd__inv_2
X_3892_ _3899_/CLK _3892_/D vssd1 vssd1 vccd1 vccd1 _3892_/Q sky130_fd_sc_hd__dfxtp_1
X_2843_ _2843_/A _2995_/X vssd1 vssd1 vccd1 vccd1 _2843_/X sky130_fd_sc_hd__and2_1
X_2774_ _3664_/Q vssd1 vssd1 vccd1 vccd1 _2774_/Y sky130_fd_sc_hd__inv_2
X_1725_ _1727_/A _3069_/X _1727_/C vssd1 vssd1 vccd1 vccd1 _3890_/D sky130_fd_sc_hd__and3_1
XFILLER_86_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3326_ _3322_/X _3323_/X _3324_/X _3325_/X _3373_/S0 _3378_/S1 vssd1 vssd1 vccd1
+ vccd1 _3326_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3257_ _3788_/Q _3784_/Q _3792_/Q _3764_/Q _3009_/S _3286_/S1 vssd1 vssd1 vccd1 vccd1
+ _3257_/X sky130_fd_sc_hd__mux4_1
X_2208_ _2222_/A vssd1 vssd1 vccd1 vccd1 _2208_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3188_ _3184_/X _3185_/X _3186_/X _3187_/X _3295_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3188_/X sky130_fd_sc_hd__mux4_2
X_2139_ _2139_/A vssd1 vssd1 vccd1 vccd1 _2139_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2490_ _3469_/Q _2485_/X _2448_/X _2486_/X vssd1 vssd1 vccd1 vccd1 _3469_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3111_ _2808_/Y _2809_/Y _2806_/Y _2807_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3111_/X sky130_fd_sc_hd__mux4_2
XFILLER_4_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3042_ _3314_/X _3315_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3042_/X sky130_fd_sc_hd__mux2_1
Xinput290 io_dsi_in[4] vssd1 vssd1 vccd1 vccd1 _2877_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_82_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3875_ _3877_/CLK _3875_/D vssd1 vssd1 vccd1 vccd1 _3875_/Q sky130_fd_sc_hd__dfxtp_1
X_2826_ _3587_/Q vssd1 vssd1 vccd1 vccd1 _2826_/Y sky130_fd_sc_hd__inv_2
X_2757_ _3679_/Q vssd1 vssd1 vccd1 vccd1 _2757_/Y sky130_fd_sc_hd__inv_2
X_1708_ _3073_/S _1707_/X _3896_/Q _1700_/Y _1703_/X vssd1 vssd1 vccd1 vccd1 _3896_/D
+ sky130_fd_sc_hd__o221a_1
X_2688_ _3710_/Q vssd1 vssd1 vccd1 vccd1 _2688_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3309_ _3427_/Q _3603_/Q _3579_/Q _3555_/Q _3364_/S0 _3338_/S1 vssd1 vssd1 vccd1
+ vccd1 _3309_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1990_ _3768_/Q _1986_/X _1970_/X _1988_/X vssd1 vssd1 vccd1 vccd1 _3768_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3660_ _3676_/CLK _3660_/D vssd1 vssd1 vccd1 vccd1 _3660_/Q sky130_fd_sc_hd__dfxtp_1
X_2611_ _3382_/Q _2603_/A _2149_/A _2604_/A vssd1 vssd1 vccd1 vccd1 _3382_/D sky130_fd_sc_hd__a22o_1
X_3591_ _3719_/CLK _3591_/D vssd1 vssd1 vccd1 vccd1 _3591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2542_ _2948_/A vssd1 vssd1 vccd1 vccd1 _2542_/X sky130_fd_sc_hd__clkbuf_2
X_2473_ _3480_/Q _2467_/X _2460_/X _2468_/X vssd1 vssd1 vccd1 vccd1 _3480_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_44_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3687_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3025_ _3025_/A0 _3025_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3025_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3858_ _3899_/CLK _3858_/D vssd1 vssd1 vccd1 vccd1 _3858_/Q sky130_fd_sc_hd__dfxtp_2
X_3789_ _3890_/CLK _3789_/D vssd1 vssd1 vccd1 vccd1 _3789_/Q sky130_fd_sc_hd__dfxtp_1
X_2809_ _3610_/Q vssd1 vssd1 vccd1 vccd1 _2809_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1973_ _3775_/Q _1965_/X _1972_/X _1968_/X vssd1 vssd1 vccd1 vccd1 _3775_/D sky130_fd_sc_hd__a22o_1
X_3712_ _3730_/CLK _3712_/D vssd1 vssd1 vccd1 vccd1 _3712_/Q sky130_fd_sc_hd__dfxtp_1
X_3643_ _3676_/CLK _3643_/D vssd1 vssd1 vccd1 vccd1 _3643_/Q sky130_fd_sc_hd__dfxtp_1
X_3574_ _3743_/CLK _3574_/D vssd1 vssd1 vccd1 vccd1 _3574_/Q sky130_fd_sc_hd__dfxtp_1
X_2525_ _3444_/Q _2519_/X _2450_/X _2520_/X vssd1 vssd1 vccd1 vccd1 _3444_/D sky130_fd_sc_hd__a22o_1
X_2456_ _2948_/A vssd1 vssd1 vccd1 vccd1 _2456_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2387_ _3536_/Q _2382_/X _2360_/X _2383_/X vssd1 vssd1 vccd1 vccd1 _3536_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3008_ _3008_/A0 _3008_/A1 _3009_/S vssd1 vssd1 vccd1 vccd1 _3008_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3290_ _3031_/X _3033_/X _3034_/X _2663_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3290_/X sky130_fd_sc_hd__mux4_2
X_2310_ _2310_/A vssd1 vssd1 vccd1 vccd1 _2310_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2241_ _2257_/A vssd1 vssd1 vccd1 vccd1 _2259_/A sky130_fd_sc_hd__inv_2
X_2172_ _3668_/Q _2166_/X _2135_/X _2167_/X vssd1 vssd1 vccd1 vccd1 _3668_/D sky130_fd_sc_hd__a22o_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1956_ _1985_/A _1977_/B _2021_/C _1964_/D vssd1 vssd1 vccd1 vccd1 _2563_/A sky130_fd_sc_hd__or4_4
X_1887_ _2143_/A vssd1 vssd1 vccd1 vccd1 _1887_/X sky130_fd_sc_hd__clkbuf_2
X_3626_ _3746_/CLK _3626_/D vssd1 vssd1 vccd1 vccd1 _3626_/Q sky130_fd_sc_hd__dfxtp_1
X_3557_ _3773_/CLK _3557_/D vssd1 vssd1 vccd1 vccd1 _3557_/Q sky130_fd_sc_hd__dfxtp_1
X_2508_ _3455_/Q _2501_/A _2462_/X _2502_/A vssd1 vssd1 vccd1 vccd1 _3455_/D sky130_fd_sc_hd__a22o_1
Xinput108 io_b_dat_o_4[9] vssd1 vssd1 vccd1 vccd1 _3268_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3488_ _3714_/CLK _3488_/D vssd1 vssd1 vccd1 vccd1 _3488_/Q sky130_fd_sc_hd__dfxtp_1
Xinput119 io_b_dat_o_5[4] vssd1 vssd1 vccd1 vccd1 _3328_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2439_ _3500_/Q _2435_/X _2326_/X _2437_/X vssd1 vssd1 vccd1 vccd1 _3500_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1810_ _3103_/X _1814_/B vssd1 vssd1 vccd1 vccd1 _3836_/D sky130_fd_sc_hd__nor2_1
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2790_ _3665_/Q vssd1 vssd1 vccd1 vccd1 _2790_/Y sky130_fd_sc_hd__inv_2
XPHY_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1741_ _2944_/A vssd1 vssd1 vccd1 vccd1 _2149_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3411_ _3627_/CLK _3411_/D vssd1 vssd1 vccd1 vccd1 _3411_/Q sky130_fd_sc_hd__dfxtp_1
X_3342_ _3047_/X _3049_/X _3050_/X _2622_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3342_/X sky130_fd_sc_hd__mux4_2
XFILLER_3_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3273_ _3786_/Q _3782_/Q _3790_/Q _3762_/Q _2971_/S _3286_/S1 vssd1 vssd1 vccd1 vccd1
+ _3273_/X sky130_fd_sc_hd__mux4_2
X_2224_ _3634_/Q _2221_/X _2141_/X _2222_/X vssd1 vssd1 vccd1 vccd1 _3634_/D sky130_fd_sc_hd__a22o_1
X_2155_ _2959_/A vssd1 vssd1 vccd1 vccd1 _2155_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2086_ _3713_/Q _2082_/X _1887_/X _2083_/X vssd1 vssd1 vccd1 vccd1 _3713_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2988_ _2988_/A0 _2988_/A1 _2996_/S vssd1 vssd1 vccd1 vccd1 _2988_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1939_ _2009_/A _1977_/B _2510_/C _1964_/D vssd1 vssd1 vccd1 vccd1 _2583_/A sky130_fd_sc_hd__or4_4
Xinput90 io_b_dat_o_3[7] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_1
X_3609_ _3682_/CLK _3609_/D vssd1 vssd1 vccd1 vccd1 _3609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2911_ _3704_/Q vssd1 vssd1 vccd1 vccd1 _2911_/Y sky130_fd_sc_hd__inv_2
X_3891_ _3899_/CLK _3891_/D vssd1 vssd1 vccd1 vccd1 _3891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2842_ _3612_/Q vssd1 vssd1 vccd1 vccd1 _2842_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2773_ _3680_/Q vssd1 vssd1 vccd1 vccd1 _2773_/Y sky130_fd_sc_hd__inv_2
X_1724_ _1727_/A _3068_/X _1727_/C vssd1 vssd1 vccd1 vccd1 _3891_/D sky130_fd_sc_hd__and3_1
X_3325_ _3402_/Q _3394_/Q _3386_/Q _3626_/Q _3351_/S0 _3351_/S1 vssd1 vssd1 vccd1
+ vccd1 _3325_/X sky130_fd_sc_hd__mux4_2
X_3256_ _3804_/Q _3752_/Q _3780_/Q _3776_/Q _3036_/S _3294_/S1 vssd1 vssd1 vccd1 vccd1
+ _3256_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2207_ _2221_/A vssd1 vssd1 vccd1 vccd1 _2222_/A sky130_fd_sc_hd__inv_2
XFILLER_37_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3187_ _3495_/Q _3471_/Q _3447_/Q _3735_/Q _3060_/S _3192_/S1 vssd1 vssd1 vccd1 vccd1
+ _3187_/X sky130_fd_sc_hd__mux4_2
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2138_ _2138_/A vssd1 vssd1 vccd1 vccd1 _2138_/X sky130_fd_sc_hd__buf_2
XFILLER_26_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2069_ _2083_/A vssd1 vssd1 vccd1 vccd1 _2069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3110_ _2812_/Y _2813_/Y _2810_/Y _2811_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3110_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput280 io_dataLastBlock[62] vssd1 vssd1 vccd1 vccd1 _3000_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3041_ _3313_/X _3040_/X _3053_/S vssd1 vssd1 vccd1 vccd1 _3041_/X sky130_fd_sc_hd__mux2_1
Xinput291 io_dsi_in[5] vssd1 vssd1 vccd1 vccd1 _2877_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3874_ _3896_/CLK _3874_/D vssd1 vssd1 vccd1 vccd1 _3874_/Q sky130_fd_sc_hd__dfxtp_1
X_2825_ _3611_/Q vssd1 vssd1 vccd1 vccd1 _2825_/Y sky130_fd_sc_hd__inv_2
X_2756_ _3695_/Q vssd1 vssd1 vccd1 vccd1 _2756_/Y sky130_fd_sc_hd__inv_2
X_1707_ _1707_/A _1707_/B vssd1 vssd1 vccd1 vccd1 _1707_/X sky130_fd_sc_hd__and2_1
X_2687_ _3558_/Q vssd1 vssd1 vccd1 vccd1 _2687_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3308_ _3304_/X _3305_/X _3306_/X _3307_/X _3373_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3308_/X sky130_fd_sc_hd__mux4_2
X_3239_ _2657_/X _2658_/X _3016_/X _2661_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3239_/X sky130_fd_sc_hd__mux4_2
XFILLER_73_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2610_ _3383_/Q _2603_/A _2147_/A _2604_/A vssd1 vssd1 vccd1 vccd1 _3383_/D sky130_fd_sc_hd__a22o_1
X_3590_ _3719_/CLK _3590_/D vssd1 vssd1 vccd1 vccd1 _3590_/Q sky130_fd_sc_hd__dfxtp_1
X_2541_ _3435_/Q _2536_/X _2540_/X _2538_/X vssd1 vssd1 vccd1 vccd1 _3435_/D sky130_fd_sc_hd__a22o_1
X_2472_ _3481_/Q _2467_/X _2458_/X _2468_/X vssd1 vssd1 vccd1 vccd1 _3481_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3024_ _3259_/X _3260_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3024_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_13_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3851_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3857_ _3873_/CLK _3857_/D vssd1 vssd1 vccd1 vccd1 _3857_/Q sky130_fd_sc_hd__dfxtp_1
X_3788_ _3828_/CLK _3788_/D vssd1 vssd1 vccd1 vccd1 _3788_/Q sky130_fd_sc_hd__dfxtp_1
X_2808_ _3634_/Q vssd1 vssd1 vccd1 vccd1 _2808_/Y sky130_fd_sc_hd__inv_2
X_2739_ _3753_/Q vssd1 vssd1 vccd1 vccd1 _2739_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1972_ _1972_/A vssd1 vssd1 vccd1 vccd1 _1972_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3711_ _3727_/CLK _3711_/D vssd1 vssd1 vccd1 vccd1 _3711_/Q sky130_fd_sc_hd__dfxtp_1
X_3642_ _3723_/CLK _3642_/D vssd1 vssd1 vccd1 vccd1 _3642_/Q sky130_fd_sc_hd__dfxtp_1
X_3573_ _3741_/CLK _3573_/D vssd1 vssd1 vccd1 vccd1 _3573_/Q sky130_fd_sc_hd__dfxtp_1
X_2524_ _3445_/Q _2519_/X _2448_/X _2520_/X vssd1 vssd1 vccd1 vccd1 _3445_/D sky130_fd_sc_hd__a22o_1
X_2455_ _3491_/Q _2452_/X _2453_/X _2454_/X vssd1 vssd1 vccd1 vccd1 _3491_/D sky130_fd_sc_hd__a22o_1
X_2386_ _3537_/Q _2382_/X _2358_/X _2383_/X vssd1 vssd1 vccd1 vccd1 _3537_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3007_ _3007_/A0 _3007_/A1 _3009_/S vssd1 vssd1 vccd1 vccd1 _3007_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput370 _3838_/Q vssd1 vssd1 vccd1 vccd1 io_vout[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2240_ _2257_/A vssd1 vssd1 vccd1 vccd1 _2240_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2171_ _3669_/Q _2166_/X _2133_/X _2167_/X vssd1 vssd1 vccd1 vccd1 _3669_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1955_ _3782_/Q _1949_/X _1925_/X _1951_/X vssd1 vssd1 vccd1 vccd1 _3782_/D sky130_fd_sc_hd__a22o_1
X_1886_ _3810_/Q _1881_/X _1885_/X _1883_/X vssd1 vssd1 vccd1 vccd1 _3810_/D sky130_fd_sc_hd__a22o_1
X_3625_ _3896_/CLK _3625_/D vssd1 vssd1 vccd1 vccd1 _3625_/Q sky130_fd_sc_hd__dfxtp_1
X_3556_ _3604_/CLK _3556_/D vssd1 vssd1 vccd1 vccd1 _3556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2507_ _3456_/Q _2501_/X _2460_/X _2502_/X vssd1 vssd1 vccd1 vccd1 _3456_/D sky130_fd_sc_hd__a22o_1
Xinput109 io_b_dat_o_5[0] vssd1 vssd1 vccd1 vccd1 _3380_/A1 sky130_fd_sc_hd__clkbuf_1
X_3487_ _3727_/CLK _3487_/D vssd1 vssd1 vccd1 vccd1 _3487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2438_ _3501_/Q _2435_/X _2322_/X _2437_/X vssd1 vssd1 vccd1 vccd1 _3501_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2369_ _2383_/A vssd1 vssd1 vccd1 vccd1 _2369_/X sky130_fd_sc_hd__buf_2
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1740_ _3885_/Q vssd1 vssd1 vccd1 vccd1 _1740_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3410_ _3851_/CLK _3410_/D vssd1 vssd1 vccd1 vccd1 _3410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3341_ _3341_/A0 _3341_/A1 _3341_/A2 _3341_/A3 _2996_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3341_/X sky130_fd_sc_hd__mux4_1
X_3272_ _3802_/Q _3750_/Q _3778_/Q _3774_/Q _3285_/S0 _3294_/S1 vssd1 vssd1 vccd1
+ vccd1 _3272_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2223_ _3635_/Q _2221_/X _2138_/X _2222_/X vssd1 vssd1 vccd1 vccd1 _3635_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2154_ _2173_/A vssd1 vssd1 vccd1 vccd1 _2154_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2085_ _3714_/Q _2082_/X _1885_/X _2083_/X vssd1 vssd1 vccd1 vccd1 _3714_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2987_ _2986_/X _2612_/X _2997_/S vssd1 vssd1 vccd1 vccd1 _2987_/X sky130_fd_sc_hd__mux2_1
X_1938_ _3790_/Q _1932_/X _1925_/X _1934_/X vssd1 vssd1 vccd1 vccd1 _3790_/D sky130_fd_sc_hd__a22o_1
X_1869_ _2956_/A vssd1 vssd1 vccd1 vccd1 _1869_/X sky130_fd_sc_hd__clkbuf_2
Xinput80 io_b_dat_o_3[12] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__clkbuf_1
Xinput91 io_b_dat_o_3[8] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__clkbuf_1
X_3608_ _3682_/CLK _3608_/D vssd1 vssd1 vccd1 vccd1 _3608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3539_ _3731_/CLK _3539_/D vssd1 vssd1 vccd1 vccd1 _3539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2910_ _3720_/Q vssd1 vssd1 vccd1 vccd1 _2910_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3890_ _3890_/CLK _3890_/D vssd1 vssd1 vccd1 vccd1 _3890_/Q sky130_fd_sc_hd__dfxtp_1
X_2841_ _3636_/Q vssd1 vssd1 vccd1 vccd1 _2841_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2772_ _3696_/Q vssd1 vssd1 vccd1 vccd1 _2772_/Y sky130_fd_sc_hd__inv_2
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1723_ _1727_/A _3067_/X _1723_/C vssd1 vssd1 vccd1 vccd1 _3892_/D sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3817_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3324_ _3434_/Q _3746_/Q _3418_/Q _3410_/Q _3351_/S0 _3351_/S1 vssd1 vssd1 vccd1
+ vccd1 _3324_/X sky130_fd_sc_hd__mux4_2
X_3255_ _3760_/Q _3796_/Q _3828_/Q _3824_/Q _2971_/S _3286_/S1 vssd1 vssd1 vccd1 vccd1
+ _3255_/X sky130_fd_sc_hd__mux4_1
X_2206_ _2221_/A vssd1 vssd1 vccd1 vccd1 _2206_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3186_ _3591_/Q _3815_/Q _3543_/Q _3519_/Q _3060_/S _3192_/S1 vssd1 vssd1 vccd1 vccd1
+ _3186_/X sky130_fd_sc_hd__mux4_1
X_2137_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2137_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2068_ _2082_/A vssd1 vssd1 vccd1 vccd1 _2083_/A sky130_fd_sc_hd__inv_2
XFILLER_53_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput281 io_dataLastBlock[63] vssd1 vssd1 vccd1 vccd1 _2999_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput270 io_dataLastBlock[53] vssd1 vssd1 vccd1 vccd1 _3009_/A1 sky130_fd_sc_hd__clkbuf_1
X_3040_ _3040_/A0 _3040_/A1 _3060_/S vssd1 vssd1 vccd1 vccd1 _3040_/X sky130_fd_sc_hd__mux2_2
Xinput292 io_dsi_in[6] vssd1 vssd1 vccd1 vccd1 _2878_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3873_ _3873_/CLK _3873_/D vssd1 vssd1 vccd1 vccd1 _3873_/Q sky130_fd_sc_hd__dfxtp_1
X_2824_ _3635_/Q vssd1 vssd1 vccd1 vccd1 _2824_/Y sky130_fd_sc_hd__inv_2
X_2755_ _3711_/Q vssd1 vssd1 vccd1 vccd1 _2755_/Y sky130_fd_sc_hd__inv_2
X_1706_ _3073_/S _1705_/X _3897_/Q _1700_/Y _1703_/X vssd1 vssd1 vccd1 vccd1 _3897_/D
+ sky130_fd_sc_hd__o221a_1
X_2686_ _2686_/A _3859_/Q vssd1 vssd1 vccd1 vccd1 _2686_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3307_ _3491_/Q _3467_/Q _3443_/Q _3731_/Q _1905_/A _1905_/B vssd1 vssd1 vccd1 vccd1
+ _3307_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3238_ input98/X _3238_/A1 _3238_/A2 _3238_/A3 _3009_/S _3286_/S1 vssd1 vssd1 vccd1
+ vccd1 _3238_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3169_ _3570_/Q _3722_/Q _3706_/Q _3690_/Q _3292_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3169_/X sky130_fd_sc_hd__mux4_2
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2540_ _2949_/A vssd1 vssd1 vccd1 vccd1 _2540_/X sky130_fd_sc_hd__clkbuf_2
X_2471_ _3482_/Q _2467_/X _2456_/X _2468_/X vssd1 vssd1 vccd1 vccd1 _3482_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3023_ _3258_/X _3022_/X _3061_/S vssd1 vssd1 vccd1 vccd1 _3023_/X sky130_fd_sc_hd__mux2_2
XFILLER_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3727_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3856_ _3867_/CLK _3856_/D vssd1 vssd1 vccd1 vccd1 _3856_/Q sky130_fd_sc_hd__dfxtp_1
X_3787_ _3791_/CLK _3787_/D vssd1 vssd1 vccd1 vccd1 _3787_/Q sky130_fd_sc_hd__dfxtp_1
X_2807_ _3650_/Q vssd1 vssd1 vccd1 vccd1 _2807_/Y sky130_fd_sc_hd__inv_2
X_2738_ _3805_/Q vssd1 vssd1 vccd1 vccd1 _2738_/Y sky130_fd_sc_hd__inv_2
X_2669_ input8/X vssd1 vssd1 vccd1 vccd1 _2676_/B sky130_fd_sc_hd__inv_2
XFILLER_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1971_ _3776_/Q _1965_/X _1970_/X _1968_/X vssd1 vssd1 vccd1 vccd1 _3776_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3710_ _3821_/CLK _3710_/D vssd1 vssd1 vccd1 vccd1 _3710_/Q sky130_fd_sc_hd__dfxtp_1
X_3641_ _3723_/CLK _3641_/D vssd1 vssd1 vccd1 vccd1 _3641_/Q sky130_fd_sc_hd__dfxtp_1
X_3572_ _3722_/CLK _3572_/D vssd1 vssd1 vccd1 vccd1 _3572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2523_ _3446_/Q _2519_/X _1974_/A _2520_/X vssd1 vssd1 vccd1 vccd1 _3446_/D sky130_fd_sc_hd__a22o_1
X_2454_ _2454_/A vssd1 vssd1 vccd1 vccd1 _2454_/X sky130_fd_sc_hd__buf_2
XFILLER_68_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2385_ _3538_/Q _2382_/X _2356_/X _2383_/X vssd1 vssd1 vccd1 vccd1 _3538_/D sky130_fd_sc_hd__a22o_1
Xinput1 io_adr_i[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_4
X_3006_ _3006_/A0 _3006_/A1 _3009_/S vssd1 vssd1 vccd1 vccd1 _3006_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3839_ _3841_/CLK _3839_/D vssd1 vssd1 vccd1 vccd1 _3839_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput360 _3841_/Q vssd1 vssd1 vccd1 vccd1 io_irq sky130_fd_sc_hd__clkbuf_2
Xoutput371 _3839_/Q vssd1 vssd1 vccd1 vccd1 io_vout[9] sky130_fd_sc_hd__clkbuf_2
XINSDIODE3_0 _3040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2170_ _3670_/Q _2166_/X _2131_/X _2167_/X vssd1 vssd1 vccd1 vccd1 _3670_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1954_ _3783_/Q _1949_/X _1923_/X _1951_/X vssd1 vssd1 vccd1 vccd1 _3783_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3624_ _3867_/CLK _3624_/D vssd1 vssd1 vccd1 vccd1 _3624_/Q sky130_fd_sc_hd__dfxtp_1
X_1885_ _2141_/A vssd1 vssd1 vccd1 vccd1 _1885_/X sky130_fd_sc_hd__clkbuf_2
X_3555_ _3604_/CLK _3555_/D vssd1 vssd1 vccd1 vccd1 _3555_/Q sky130_fd_sc_hd__dfxtp_1
X_3486_ _3812_/CLK _3486_/D vssd1 vssd1 vccd1 vccd1 _3486_/Q sky130_fd_sc_hd__dfxtp_1
X_2506_ _3457_/Q _2501_/X _2458_/X _2502_/X vssd1 vssd1 vccd1 vccd1 _3457_/D sky130_fd_sc_hd__a22o_1
X_2437_ _2454_/A vssd1 vssd1 vccd1 vccd1 _2437_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2368_ _2382_/A vssd1 vssd1 vccd1 vccd1 _2383_/A sky130_fd_sc_hd__inv_2
X_2299_ _3589_/Q _2291_/X _2253_/X _2293_/X vssd1 vssd1 vccd1 vccd1 _3589_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3340_ input22/X input54/X input70/X input86/X _2996_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3340_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_4_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
X_3271_ _3758_/Q _3794_/Q _3826_/Q _3822_/Q _3285_/S0 _3294_/S1 vssd1 vssd1 vccd1
+ vccd1 _3271_/X sky130_fd_sc_hd__mux4_2
X_2222_ _2222_/A vssd1 vssd1 vccd1 vccd1 _2222_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2153_ _2281_/A _2320_/B _2673_/A _2281_/D vssd1 vssd1 vccd1 vccd1 _2173_/A sky130_fd_sc_hd__or4_4
XFILLER_93_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2084_ _3715_/Q _2082_/X _1882_/X _2083_/X vssd1 vssd1 vccd1 vccd1 _3715_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2986_ _2986_/A0 _2986_/A1 _2996_/S vssd1 vssd1 vccd1 vccd1 _2986_/X sky130_fd_sc_hd__mux2_1
X_1937_ _3791_/Q _1932_/X _1923_/X _1934_/X vssd1 vssd1 vccd1 vccd1 _3791_/D sky130_fd_sc_hd__a22o_1
X_1868_ _3819_/Q _1860_/X _1867_/X _1863_/X vssd1 vssd1 vccd1 vccd1 _3819_/D sky130_fd_sc_hd__a22o_1
Xinput70 io_b_dat_o_2[3] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_1
Xinput81 io_b_dat_o_3[13] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__clkbuf_1
X_3607_ _3662_/CLK _3607_/D vssd1 vssd1 vccd1 vccd1 _3607_/Q sky130_fd_sc_hd__dfxtp_1
Xinput92 io_b_dat_o_3[9] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__clkbuf_1
X_1799_ _1801_/A _3355_/X vssd1 vssd1 vccd1 vccd1 _3844_/D sky130_fd_sc_hd__and2_1
X_3538_ _3586_/CLK _3538_/D vssd1 vssd1 vccd1 vccd1 _3538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3469_ _3812_/CLK _3469_/D vssd1 vssd1 vccd1 vccd1 _3469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3604_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2840_ _3652_/Q vssd1 vssd1 vccd1 vccd1 _2840_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2771_ _3712_/Q vssd1 vssd1 vccd1 vccd1 _2771_/Y sky130_fd_sc_hd__inv_2
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ _1742_/A vssd1 vssd1 vccd1 vccd1 _1727_/A sky130_fd_sc_hd__buf_1
XFILLER_7_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3323_ _3530_/Q _3506_/Q _3482_/Q _3458_/Q _3351_/S0 _3351_/S1 vssd1 vssd1 vccd1
+ vccd1 _3323_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3254_ _3800_/Q _3756_/Q _3772_/Q _3768_/Q _3036_/S _3294_/S1 vssd1 vssd1 vccd1 vccd1
+ _3254_/X sky130_fd_sc_hd__mux4_2
XFILLER_58_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2205_ _2239_/A _2320_/B _2673_/A _2281_/D vssd1 vssd1 vccd1 vccd1 _2221_/A sky130_fd_sc_hd__or4_4
X_3185_ _3671_/Q _3655_/Q _3639_/Q _3615_/Q _3060_/S _3192_/S1 vssd1 vssd1 vccd1 vccd1
+ _3185_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2136_ _3684_/Q _2125_/X _2135_/X _2127_/X vssd1 vssd1 vccd1 vccd1 _3684_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2067_ _2082_/A vssd1 vssd1 vccd1 vccd1 _2067_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2969_ _2968_/X _2654_/X _2981_/S vssd1 vssd1 vccd1 vccd1 _2969_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput271 io_dataLastBlock[54] vssd1 vssd1 vccd1 vccd1 _3008_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput260 io_dataLastBlock[44] vssd1 vssd1 vccd1 vccd1 _2973_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput293 io_dsi_in[7] vssd1 vssd1 vccd1 vccd1 _2878_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput282 io_dataLastBlock[6] vssd1 vssd1 vccd1 vccd1 _3036_/A0 sky130_fd_sc_hd__buf_1
XFILLER_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3872_ _3873_/CLK _3872_/D vssd1 vssd1 vccd1 vccd1 _3872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2823_ _3651_/Q vssd1 vssd1 vccd1 vccd1 _2823_/Y sky130_fd_sc_hd__inv_2
X_2754_ _3559_/Q vssd1 vssd1 vccd1 vccd1 _2754_/Y sky130_fd_sc_hd__inv_2
X_1705_ _1679_/A _1707_/A _3897_/Q _3896_/Q _1707_/B vssd1 vssd1 vccd1 vccd1 _1705_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2685_ input7/X input8/X _2685_/C vssd1 vssd1 vccd1 vccd1 _2685_/Y sky130_fd_sc_hd__nor3_2
X_3306_ _3587_/Q _3811_/Q _3539_/Q _3515_/Q _1905_/A _3357_/S1 vssd1 vssd1 vccd1 vccd1
+ _3306_/X sky130_fd_sc_hd__mux4_2
XFILLER_86_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3237_ input18/X input50/X input66/X input82/X _2971_/S _2981_/S vssd1 vssd1 vccd1
+ vccd1 _3237_/X sky130_fd_sc_hd__mux4_1
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3168_ _3164_/X _3165_/X _3166_/X _3167_/X _3295_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3168_/X sky130_fd_sc_hd__mux4_2
X_2119_ _3693_/Q _2116_/X _1861_/X _2118_/X vssd1 vssd1 vccd1 vccd1 _3693_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3099_ _2850_/Y _2851_/Y _2848_/Y _2849_/Y _3153_/X _3132_/S1 vssd1 vssd1 vccd1 vccd1
+ _3099_/X sky130_fd_sc_hd__mux4_2
XFILLER_50_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2470_ _3483_/Q _2467_/X _2453_/X _2468_/X vssd1 vssd1 vccd1 vccd1 _3483_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3022_ _3022_/A0 _3022_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3022_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3855_ _3873_/CLK _3855_/D vssd1 vssd1 vccd1 vccd1 _3855_/Q sky130_fd_sc_hd__dfxtp_1
X_3786_ _3796_/CLK _3786_/D vssd1 vssd1 vccd1 vccd1 _3786_/Q sky130_fd_sc_hd__dfxtp_1
X_2806_ _3666_/Q vssd1 vssd1 vccd1 vccd1 _2806_/Y sky130_fd_sc_hd__inv_2
X_2737_ _3825_/Q vssd1 vssd1 vccd1 vccd1 _2737_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_22_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3627_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2668_ input7/X vssd1 vssd1 vccd1 vccd1 _2684_/A sky130_fd_sc_hd__clkbuf_4
X_2599_ _3392_/Q _2593_/X _2145_/A _2594_/X vssd1 vssd1 vccd1 vccd1 _3392_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1970_ _1970_/A vssd1 vssd1 vccd1 vccd1 _1970_/X sky130_fd_sc_hd__clkbuf_2
X_3640_ _3672_/CLK _3640_/D vssd1 vssd1 vccd1 vccd1 _3640_/Q sky130_fd_sc_hd__dfxtp_1
X_3571_ _3722_/CLK _3571_/D vssd1 vssd1 vccd1 vccd1 _3571_/Q sky130_fd_sc_hd__dfxtp_1
X_2522_ _3447_/Q _2519_/X _1972_/A _2520_/X vssd1 vssd1 vccd1 vccd1 _3447_/D sky130_fd_sc_hd__a22o_1
X_2453_ _2949_/A vssd1 vssd1 vccd1 vccd1 _2453_/X sky130_fd_sc_hd__clkbuf_2
X_2384_ _3539_/Q _2382_/X _2354_/X _2383_/X vssd1 vssd1 vccd1 vccd1 _3539_/D sky130_fd_sc_hd__a22o_1
Xinput2 io_adr_i[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3005_ _3005_/A0 _3005_/A1 _3009_/S vssd1 vssd1 vccd1 vccd1 _3005_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3838_ _3841_/CLK _3838_/D vssd1 vssd1 vccd1 vccd1 _3838_/Q sky130_fd_sc_hd__dfxtp_1
X_3769_ _3773_/CLK _3769_/D vssd1 vssd1 vccd1 vccd1 _3769_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput350 _3878_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput361 _3830_/Q vssd1 vssd1 vccd1 vccd1 io_vout[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE3_1 _3871_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1953_ _3784_/Q _1949_/X _1921_/X _1951_/X vssd1 vssd1 vccd1 vccd1 _3784_/D sky130_fd_sc_hd__a22o_1
X_1884_ _3811_/Q _1881_/X _1882_/X _1883_/X vssd1 vssd1 vccd1 vccd1 _3811_/D sky130_fd_sc_hd__a22o_1
X_3623_ _3895_/CLK _3623_/D vssd1 vssd1 vccd1 vccd1 _3623_/Q sky130_fd_sc_hd__dfxtp_1
X_3554_ _3845_/CLK _3554_/D vssd1 vssd1 vccd1 vccd1 _3554_/Q sky130_fd_sc_hd__dfxtp_1
X_3485_ _3823_/CLK _3485_/D vssd1 vssd1 vccd1 vccd1 _3485_/Q sky130_fd_sc_hd__dfxtp_1
X_2505_ _3458_/Q _2501_/X _2456_/X _2502_/X vssd1 vssd1 vccd1 vccd1 _3458_/D sky130_fd_sc_hd__a22o_1
X_2436_ _2452_/A vssd1 vssd1 vccd1 vccd1 _2454_/A sky130_fd_sc_hd__inv_2
XFILLER_69_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2367_ _2382_/A vssd1 vssd1 vccd1 vccd1 _2367_/X sky130_fd_sc_hd__buf_2
XFILLER_56_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2298_ _3590_/Q _2291_/X _2297_/X _2293_/X vssd1 vssd1 vccd1 vccd1 _3590_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3270_ _3798_/Q _3754_/Q _3770_/Q _3766_/Q _3285_/S0 _3294_/S1 vssd1 vssd1 vccd1
+ vccd1 _3270_/X sky130_fd_sc_hd__mux4_1
X_2221_ _2221_/A vssd1 vssd1 vccd1 vccd1 _2221_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2152_ _2510_/D vssd1 vssd1 vccd1 vccd1 _2281_/D sky130_fd_sc_hd__buf_1
X_2083_ _2083_/A vssd1 vssd1 vccd1 vccd1 _2083_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2985_ _2984_/X _2645_/X _2997_/S vssd1 vssd1 vccd1 vccd1 _2985_/X sky130_fd_sc_hd__mux2_1
X_1936_ _3792_/Q _1932_/X _1921_/X _1934_/X vssd1 vssd1 vccd1 vccd1 _3792_/D sky130_fd_sc_hd__a22o_1
X_1867_ _2957_/A vssd1 vssd1 vccd1 vccd1 _1867_/X sky130_fd_sc_hd__clkbuf_2
Xinput60 io_b_dat_o_1[9] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_1
Xinput71 io_b_dat_o_2[4] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_1
Xinput82 io_b_dat_o_3[14] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__clkbuf_1
X_1798_ _1801_/A _3342_/X vssd1 vssd1 vccd1 vccd1 _3845_/D sky130_fd_sc_hd__and2_1
X_3606_ _3662_/CLK _3606_/D vssd1 vssd1 vccd1 vccd1 _3606_/Q sky130_fd_sc_hd__dfxtp_1
Xinput93 io_b_dat_o_4[0] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_1
X_3537_ _3811_/CLK _3537_/D vssd1 vssd1 vccd1 vccd1 _3537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3468_ _3812_/CLK _3468_/D vssd1 vssd1 vccd1 vccd1 _3468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3399_ _3895_/CLK _3399_/D vssd1 vssd1 vccd1 vccd1 _3399_/Q sky130_fd_sc_hd__dfxtp_1
X_2419_ _3514_/Q _2416_/X _2356_/X _2417_/X vssd1 vssd1 vccd1 vccd1 _3514_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2770_ _3560_/Q vssd1 vssd1 vccd1 vccd1 _2770_/Y sky130_fd_sc_hd__inv_2
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _1721_/A _3066_/X _1723_/C vssd1 vssd1 vccd1 vccd1 _3893_/D sky130_fd_sc_hd__and3_1
XPHY_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3322_ _3426_/Q _3602_/Q _3578_/Q _3554_/Q _3351_/S0 _3351_/S1 vssd1 vssd1 vccd1
+ vccd1 _3322_/X sky130_fd_sc_hd__mux4_1
XFILLER_86_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3253_ _2636_/X _3020_/X _3021_/X _2638_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3253_/X sky130_fd_sc_hd__mux4_2
XFILLER_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3832_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2204_ _3646_/Q _2197_/A _2149_/X _2198_/A vssd1 vssd1 vccd1 vccd1 _3646_/D sky130_fd_sc_hd__a22o_1
X_3184_ _3567_/Q _3719_/Q _3703_/Q _3687_/Q _3060_/S _3192_/S1 vssd1 vssd1 vccd1 vccd1
+ _3184_/X sky130_fd_sc_hd__mux4_2
X_2135_ _2135_/A vssd1 vssd1 vccd1 vccd1 _2135_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_39_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2066_ _2281_/A _2181_/B _2675_/A _2115_/D vssd1 vssd1 vccd1 vccd1 _2082_/A sky130_fd_sc_hd__or4_4
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2968_ _2968_/A0 _2968_/A1 _2971_/S vssd1 vssd1 vccd1 vccd1 _2968_/X sky130_fd_sc_hd__mux2_1
X_1919_ _2426_/A vssd1 vssd1 vccd1 vccd1 _1919_/X sky130_fd_sc_hd__buf_2
X_2899_ _3639_/Q vssd1 vssd1 vccd1 vccd1 _2899_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput272 io_dataLastBlock[55] vssd1 vssd1 vccd1 vccd1 _3007_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput261 io_dataLastBlock[45] vssd1 vssd1 vccd1 vccd1 _2970_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput250 io_dataLastBlock[35] vssd1 vssd1 vccd1 vccd1 _3048_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput283 io_dataLastBlock[7] vssd1 vssd1 vccd1 vccd1 _3032_/A0 sky130_fd_sc_hd__buf_1
Xinput294 io_we_i vssd1 vssd1 vccd1 vccd1 _2960_/A sky130_fd_sc_hd__buf_1
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3871_ _3873_/CLK _3871_/D vssd1 vssd1 vccd1 vccd1 _3871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2822_ _3667_/Q vssd1 vssd1 vccd1 vccd1 _2822_/Y sky130_fd_sc_hd__inv_2
X_2753_ _3726_/Q vssd1 vssd1 vccd1 vccd1 _2753_/Y sky130_fd_sc_hd__inv_2
X_1704_ _3073_/S _1699_/X _3898_/Q _1700_/Y _1703_/X vssd1 vssd1 vccd1 vccd1 _3898_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2684_ _2684_/A _2684_/B _2684_/C vssd1 vssd1 vccd1 vccd1 _2684_/Y sky130_fd_sc_hd__nor3_4
XFILLER_59_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3305_ _3667_/Q _3651_/Q _3635_/Q _3611_/Q _3370_/S0 _3357_/S1 vssd1 vssd1 vccd1
+ vccd1 _3305_/X sky130_fd_sc_hd__mux4_2
XFILLER_86_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3236_ _2664_/X _2665_/X _3015_/X _2667_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3236_/X sky130_fd_sc_hd__mux4_2
XFILLER_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3167_ _3499_/Q _3475_/Q _3451_/Q _3739_/Q _3292_/S0 _3292_/S1 vssd1 vssd1 vccd1
+ vccd1 _3167_/X sky130_fd_sc_hd__mux4_2
XFILLER_27_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3098_ _3094_/X _3095_/X _3096_/X _3097_/X _3133_/S0 _3138_/X vssd1 vssd1 vccd1 vccd1
+ _3098_/X sky130_fd_sc_hd__mux4_2
X_2118_ _2139_/A vssd1 vssd1 vccd1 vccd1 _2118_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2049_ _3737_/Q _2042_/X _2011_/X _2044_/X vssd1 vssd1 vccd1 vccd1 _3737_/D sky130_fd_sc_hd__a22o_1
XFILLER_42_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3021_ _3251_/X _3252_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3021_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3854_ _3873_/CLK _3854_/D vssd1 vssd1 vccd1 vccd1 _3854_/Q sky130_fd_sc_hd__dfxtp_1
X_2805_ _3682_/Q vssd1 vssd1 vccd1 vccd1 _2805_/Y sky130_fd_sc_hd__inv_2
X_3785_ _3890_/CLK _3785_/D vssd1 vssd1 vccd1 vccd1 _3785_/Q sky130_fd_sc_hd__dfxtp_1
X_2736_ _3829_/Q vssd1 vssd1 vccd1 vccd1 _2736_/Y sky130_fd_sc_hd__inv_2
X_2667_ _2843_/A _2963_/X vssd1 vssd1 vccd1 vccd1 _2667_/X sky130_fd_sc_hd__and2_1
X_2598_ _3393_/Q _2593_/X _2143_/A _2594_/X vssd1 vssd1 vccd1 vccd1 _3393_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3219_ _3424_/Q _3600_/Q _3576_/Q _3552_/Q _3860_/Q _3861_/Q vssd1 vssd1 vccd1 vccd1
+ _3219_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3570_ _3722_/CLK _3570_/D vssd1 vssd1 vccd1 vccd1 _3570_/Q sky130_fd_sc_hd__dfxtp_1
X_2521_ _3448_/Q _2519_/X _1970_/A _2520_/X vssd1 vssd1 vccd1 vccd1 _3448_/D sky130_fd_sc_hd__a22o_1
X_2452_ _2452_/A vssd1 vssd1 vccd1 vccd1 _2452_/X sky130_fd_sc_hd__clkbuf_2
X_2383_ _2383_/A vssd1 vssd1 vccd1 vccd1 _2383_/X sky130_fd_sc_hd__buf_2
X_3004_ _3004_/A0 _3004_/A1 _3009_/S vssd1 vssd1 vccd1 vccd1 _3004_/X sky130_fd_sc_hd__mux2_1
Xinput3 io_adr_i[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3837_ _3841_/CLK _3837_/D vssd1 vssd1 vccd1 vccd1 _3837_/Q sky130_fd_sc_hd__dfxtp_1
X_3768_ _3799_/CLK _3768_/D vssd1 vssd1 vccd1 vccd1 _3768_/Q sky130_fd_sc_hd__dfxtp_1
X_2719_ _3788_/Q vssd1 vssd1 vccd1 vccd1 _2719_/Y sky130_fd_sc_hd__inv_2
X_3699_ _3731_/CLK _3699_/D vssd1 vssd1 vccd1 vccd1 _3699_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput351 _3879_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[31] sky130_fd_sc_hd__clkbuf_2
Xoutput340 _3869_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[21] sky130_fd_sc_hd__clkbuf_2
Xoutput362 _3840_/Q vssd1 vssd1 vccd1 vccd1 io_vout[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE3_2 _3871_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1952_ _3785_/Q _1949_/X _1917_/X _1951_/X vssd1 vssd1 vccd1 vccd1 _3785_/D sky130_fd_sc_hd__a22o_1
X_1883_ _1883_/A vssd1 vssd1 vccd1 vccd1 _1883_/X sky130_fd_sc_hd__clkbuf_2
X_3622_ _3890_/CLK _3622_/D vssd1 vssd1 vccd1 vccd1 _3622_/Q sky130_fd_sc_hd__dfxtp_1
X_3553_ _3603_/CLK _3553_/D vssd1 vssd1 vccd1 vccd1 _3553_/Q sky130_fd_sc_hd__dfxtp_1
X_3484_ _3726_/CLK _3484_/D vssd1 vssd1 vccd1 vccd1 _3484_/Q sky130_fd_sc_hd__dfxtp_1
X_2504_ _3459_/Q _2501_/X _2453_/X _2502_/X vssd1 vssd1 vccd1 vccd1 _3459_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2435_ _2452_/A vssd1 vssd1 vccd1 vccd1 _2435_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2366_ _2510_/A _2510_/B _2671_/A _2476_/D vssd1 vssd1 vccd1 vccd1 _2382_/A sky130_fd_sc_hd__or4_4
XFILLER_84_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2297_ _2952_/A vssd1 vssd1 vccd1 vccd1 _2297_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2220_ _3636_/Q _2214_/X _2135_/X _2215_/X vssd1 vssd1 vccd1 vccd1 _3636_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2151_ _2151_/A vssd1 vssd1 vccd1 vccd1 _2673_/A sky130_fd_sc_hd__buf_2
X_2082_ _2082_/A vssd1 vssd1 vccd1 vccd1 _2082_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2984_ _2984_/A0 _2984_/A1 _2984_/S vssd1 vssd1 vccd1 vccd1 _2984_/X sky130_fd_sc_hd__mux2_1
X_1935_ _3793_/Q _1932_/X _1917_/X _1934_/X vssd1 vssd1 vccd1 vccd1 _3793_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1866_ _3820_/Q _1860_/X _1865_/X _1863_/X vssd1 vssd1 vccd1 vccd1 _3820_/D sky130_fd_sc_hd__a22o_1
Xinput72 io_b_dat_o_2[5] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__clkbuf_1
Xinput50 io_b_dat_o_1[14] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_1
Xinput61 io_b_dat_o_2[0] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_1
X_1797_ _1801_/A _3329_/X vssd1 vssd1 vccd1 vccd1 _3846_/D sky130_fd_sc_hd__and2_1
X_3605_ _3773_/CLK _3605_/D vssd1 vssd1 vccd1 vccd1 _3605_/Q sky130_fd_sc_hd__dfxtp_1
Xinput94 io_b_dat_o_4[10] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__clkbuf_1
Xinput83 io_b_dat_o_3[15] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__clkbuf_1
X_3536_ _3586_/CLK _3536_/D vssd1 vssd1 vccd1 vccd1 _3536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3467_ _3811_/CLK _3467_/D vssd1 vssd1 vccd1 vccd1 _3467_/Q sky130_fd_sc_hd__dfxtp_1
X_3398_ _3890_/CLK _3398_/D vssd1 vssd1 vccd1 vccd1 _3398_/Q sky130_fd_sc_hd__dfxtp_1
X_2418_ _3515_/Q _2416_/X _2354_/X _2417_/X vssd1 vssd1 vccd1 vccd1 _3515_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2349_ _3557_/Q _1986_/X _2348_/X _1988_/X vssd1 vssd1 vccd1 vccd1 _3557_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1720_ _1721_/A _3065_/X _1723_/C vssd1 vssd1 vccd1 vccd1 _3894_/D sky130_fd_sc_hd__and3_1
X_3321_ _3317_/X _3318_/X _3319_/X _3320_/X _3373_/S0 input8/X vssd1 vssd1 vccd1 vccd1
+ _3321_/X sky130_fd_sc_hd__mux4_2
X_3252_ input95/X _3252_/A1 _3252_/A2 _3252_/A3 _2984_/S _2981_/S vssd1 vssd1 vccd1
+ vccd1 _3252_/X sky130_fd_sc_hd__mux4_1
X_2203_ _3647_/Q _2197_/X _2147_/X _2198_/X vssd1 vssd1 vccd1 vccd1 _3647_/D sky130_fd_sc_hd__a22o_1
X_3183_ _3179_/X _3180_/X _3181_/X _3182_/X _3295_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3183_/X sky130_fd_sc_hd__mux4_2
XFILLER_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2134_ _3685_/Q _2125_/X _2133_/X _2127_/X vssd1 vssd1 vccd1 vccd1 _3685_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2065_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2675_/A sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_16_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3873_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2967_ _2967_/A0 _2967_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _2967_/X sky130_fd_sc_hd__mux2_2
X_2898_ _3655_/Q vssd1 vssd1 vccd1 vccd1 _2898_/Y sky130_fd_sc_hd__inv_2
X_1918_ _2425_/A vssd1 vssd1 vccd1 vccd1 _2426_/A sky130_fd_sc_hd__inv_2
X_1849_ _3824_/Q _1845_/X _1834_/X _1847_/X vssd1 vssd1 vccd1 vccd1 _3824_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3519_ _3719_/CLK _3519_/D vssd1 vssd1 vccd1 vccd1 _3519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput262 io_dataLastBlock[46] vssd1 vssd1 vccd1 vccd1 _2967_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput240 io_dataLastBlock[26] vssd1 vssd1 vccd1 vccd1 _3004_/A0 sky130_fd_sc_hd__buf_1
XFILLER_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput251 io_dataLastBlock[36] vssd1 vssd1 vccd1 vccd1 _3044_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput295 wb_rst_i vssd1 vssd1 vccd1 vccd1 _1802_/A sky130_fd_sc_hd__buf_6
XFILLER_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput273 io_dataLastBlock[56] vssd1 vssd1 vccd1 vccd1 _3006_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput284 io_dataLastBlock[8] vssd1 vssd1 vccd1 vccd1 _3028_/A0 sky130_fd_sc_hd__buf_1
XFILLER_84_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3870_ _3896_/CLK _3870_/D vssd1 vssd1 vccd1 vccd1 _3870_/Q sky130_fd_sc_hd__dfxtp_1
X_2821_ _3683_/Q vssd1 vssd1 vccd1 vccd1 _2821_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2752_ _3438_/Q vssd1 vssd1 vccd1 vccd1 _2752_/Y sky130_fd_sc_hd__inv_2
X_1703_ _1796_/A vssd1 vssd1 vccd1 vccd1 _1703_/X sky130_fd_sc_hd__clkbuf_2
X_2683_ _2684_/A _2684_/B _2683_/C vssd1 vssd1 vccd1 vccd1 _2683_/Y sky130_fd_sc_hd__nor3_4
XFILLER_59_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3304_ _3563_/Q _3715_/Q _3699_/Q _3683_/Q _3370_/S0 _3357_/S1 vssd1 vssd1 vccd1
+ vccd1 _3304_/X sky130_fd_sc_hd__mux4_2
X_3235_ input99/X _3235_/A1 _3235_/A2 _3235_/A3 _3009_/S _3286_/S1 vssd1 vssd1 vccd1
+ vccd1 _3235_/X sky130_fd_sc_hd__mux4_1
X_3166_ _3595_/Q _3819_/Q _3547_/Q _3523_/Q _3292_/S0 _3292_/S1 vssd1 vssd1 vccd1
+ vccd1 _3166_/X sky130_fd_sc_hd__mux4_1
X_3097_ _2854_/Y _2855_/Y _2852_/Y _2853_/Y _3102_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3097_/X sky130_fd_sc_hd__mux4_1
X_2117_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2139_/A sky130_fd_sc_hd__inv_2
XFILLER_27_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2048_ _3738_/Q _2042_/X _1869_/X _2044_/X vssd1 vssd1 vccd1 vccd1 _3738_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3020_ _3250_/X _3019_/X _3061_/S vssd1 vssd1 vccd1 vccd1 _3020_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3853_ _3877_/CLK _3853_/D vssd1 vssd1 vccd1 vccd1 _3853_/Q sky130_fd_sc_hd__dfxtp_1
X_2804_ _3698_/Q vssd1 vssd1 vccd1 vccd1 _2804_/Y sky130_fd_sc_hd__inv_2
X_3784_ _3828_/CLK _3784_/D vssd1 vssd1 vccd1 vccd1 _3784_/Q sky130_fd_sc_hd__dfxtp_1
X_2735_ _3797_/Q vssd1 vssd1 vccd1 vccd1 _2735_/Y sky130_fd_sc_hd__inv_2
X_2666_ _2836_/A _2666_/B vssd1 vssd1 vccd1 vccd1 _2666_/X sky130_fd_sc_hd__and2_1
X_2597_ _3394_/Q _2593_/X _2141_/A _2594_/X vssd1 vssd1 vccd1 vccd1 _3394_/D sky130_fd_sc_hd__a22o_1
XFILLER_75_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3828_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3218_ _3214_/X _3215_/X _3216_/X _3217_/X _3862_/Q _3863_/Q vssd1 vssd1 vccd1 vccd1
+ _3218_/X sky130_fd_sc_hd__mux4_2
XFILLER_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3149_ _3798_/Q _3754_/Q _3770_/Q _3766_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3149_/X sky130_fd_sc_hd__mux4_1
XFILLER_42_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2520_ _2527_/A vssd1 vssd1 vccd1 vccd1 _2520_/X sky130_fd_sc_hd__clkbuf_2
X_2451_ _3492_/Q _2443_/X _2450_/X _2444_/X vssd1 vssd1 vccd1 vccd1 _3492_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2382_ _2382_/A vssd1 vssd1 vccd1 vccd1 _2382_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3003_ _3003_/A0 _3003_/A1 _3009_/S vssd1 vssd1 vccd1 vccd1 _3003_/X sky130_fd_sc_hd__mux2_1
Xinput4 io_adr_i[1] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_4
XFILLER_91_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3836_ _3841_/CLK _3836_/D vssd1 vssd1 vccd1 vccd1 _3836_/Q sky130_fd_sc_hd__dfxtp_1
X_3767_ _3799_/CLK _3767_/D vssd1 vssd1 vccd1 vccd1 _3767_/Q sky130_fd_sc_hd__dfxtp_1
X_2718_ _3776_/Q vssd1 vssd1 vccd1 vccd1 _2718_/Y sky130_fd_sc_hd__inv_2
X_3698_ _3714_/CLK _3698_/D vssd1 vssd1 vccd1 vccd1 _3698_/Q sky130_fd_sc_hd__dfxtp_1
X_2649_ _2661_/A _2985_/X vssd1 vssd1 vccd1 vccd1 _2649_/X sky130_fd_sc_hd__and2_1
Xoutput341 _3870_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[22] sky130_fd_sc_hd__clkbuf_2
Xoutput330 _3854_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[12] sky130_fd_sc_hd__clkbuf_2
Xoutput352 _3845_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput363 _3831_/Q vssd1 vssd1 vccd1 vccd1 io_vout[1] sky130_fd_sc_hd__clkbuf_2
XINSDIODE3_3 _3874_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1951_ _2594_/A vssd1 vssd1 vccd1 vccd1 _1951_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1882_ _2138_/A vssd1 vssd1 vccd1 vccd1 _1882_/X sky130_fd_sc_hd__clkbuf_2
X_3621_ _3662_/CLK _3621_/D vssd1 vssd1 vccd1 vccd1 _3621_/Q sky130_fd_sc_hd__dfxtp_1
X_3552_ _3845_/CLK _3552_/D vssd1 vssd1 vccd1 vccd1 _3552_/Q sky130_fd_sc_hd__dfxtp_1
X_2503_ _3460_/Q _2501_/X _2450_/X _2502_/X vssd1 vssd1 vccd1 vccd1 _3460_/D sky130_fd_sc_hd__a22o_1
X_3483_ _3807_/CLK _3483_/D vssd1 vssd1 vccd1 vccd1 _3483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2434_ _2476_/A _2510_/B _2682_/A _2476_/D vssd1 vssd1 vccd1 vccd1 _2452_/A sky130_fd_sc_hd__or4_4
X_2365_ _3550_/Q _2350_/A _2364_/X _2352_/A vssd1 vssd1 vccd1 vccd1 _3550_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2296_ _3591_/Q _2291_/X _2295_/X _2293_/X vssd1 vssd1 vccd1 vccd1 _3591_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3819_ _3831_/CLK _3819_/D vssd1 vssd1 vccd1 vccd1 _3819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2150_ _3678_/Q _2137_/A _2149_/X _2139_/A vssd1 vssd1 vccd1 vccd1 _3678_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2081_ _3716_/Q _2075_/X _1879_/X _2076_/X vssd1 vssd1 vccd1 vccd1 _3716_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2983_ _2982_/X _2662_/X _2997_/S vssd1 vssd1 vccd1 vccd1 _2983_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1934_ _2604_/A vssd1 vssd1 vccd1 vccd1 _1934_/X sky130_fd_sc_hd__clkbuf_2
Xinput40 io_b_dat_o_10[5] vssd1 vssd1 vccd1 vccd1 _2612_/A sky130_fd_sc_hd__clkbuf_1
X_1865_ _2958_/A vssd1 vssd1 vccd1 vccd1 _1865_/X sky130_fd_sc_hd__clkbuf_2
Xinput62 io_b_dat_o_2[10] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_1
Xinput51 io_b_dat_o_1[15] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
Xinput73 io_b_dat_o_2[6] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_1
X_1796_ _1796_/A vssd1 vssd1 vccd1 vccd1 _1801_/A sky130_fd_sc_hd__buf_1
X_3604_ _3604_/CLK _3604_/D vssd1 vssd1 vccd1 vccd1 _3604_/Q sky130_fd_sc_hd__dfxtp_1
Xinput95 io_b_dat_o_4[11] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_1
Xinput84 io_b_dat_o_3[1] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_1
X_3535_ _3726_/CLK _3535_/D vssd1 vssd1 vccd1 vccd1 _3535_/Q sky130_fd_sc_hd__dfxtp_1
X_3466_ _3714_/CLK _3466_/D vssd1 vssd1 vccd1 vccd1 _3466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2417_ _2417_/A vssd1 vssd1 vccd1 vccd1 _2417_/X sky130_fd_sc_hd__clkbuf_2
X_3397_ _3796_/CLK _3397_/D vssd1 vssd1 vccd1 vccd1 _3397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2348_ _2951_/A vssd1 vssd1 vccd1 vccd1 _2348_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2279_ _3599_/Q _2272_/A _2267_/X _2273_/A vssd1 vssd1 vccd1 vccd1 _3599_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3320_ _3490_/Q _3466_/Q _3442_/Q _3730_/Q input5/X _3357_/S1 vssd1 vssd1 vccd1 vccd1
+ _3320_/X sky130_fd_sc_hd__mux4_1
X_3251_ input15/X input47/X input63/X input79/X _2984_/S _2981_/S vssd1 vssd1 vccd1
+ vccd1 _3251_/X sky130_fd_sc_hd__mux4_1
X_2202_ _3648_/Q _2197_/X _2145_/X _2198_/X vssd1 vssd1 vccd1 vccd1 _3648_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3182_ _3496_/Q _3472_/Q _3448_/Q _3736_/Q _3291_/S0 _3294_/S1 vssd1 vssd1 vccd1
+ vccd1 _3182_/X sky130_fd_sc_hd__mux4_2
X_2133_ _2133_/A vssd1 vssd1 vccd1 vccd1 _2133_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_39_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2064_ _3726_/Q _2057_/A _1893_/X _2058_/A vssd1 vssd1 vccd1 vccd1 _3726_/D sky130_fd_sc_hd__a22o_1
XFILLER_62_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2966_ _2965_/X _2660_/X _2981_/S vssd1 vssd1 vccd1 vccd1 _2966_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_56_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3723_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1917_ _1966_/A vssd1 vssd1 vccd1 vccd1 _1917_/X sky130_fd_sc_hd__clkbuf_2
X_2897_ _3671_/Q vssd1 vssd1 vccd1 vccd1 _2897_/Y sky130_fd_sc_hd__inv_2
X_1848_ _3825_/Q _1845_/X _1829_/X _1847_/X vssd1 vssd1 vccd1 vccd1 _3825_/D sky130_fd_sc_hd__a22o_1
X_1779_ _1783_/A _2998_/X vssd1 vssd1 vccd1 vccd1 _3861_/D sky130_fd_sc_hd__and2_1
XFILLER_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3518_ _3719_/CLK _3518_/D vssd1 vssd1 vccd1 vccd1 _3518_/Q sky130_fd_sc_hd__dfxtp_1
X_3449_ _3741_/CLK _3449_/D vssd1 vssd1 vccd1 vccd1 _3449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput263 io_dataLastBlock[47] vssd1 vssd1 vccd1 vccd1 _2964_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput230 io_dataLastBlock[17] vssd1 vssd1 vccd1 vccd1 _3013_/A0 sky130_fd_sc_hd__buf_1
Xinput241 io_dataLastBlock[27] vssd1 vssd1 vccd1 vccd1 _3003_/A0 sky130_fd_sc_hd__buf_1
Xinput252 io_dataLastBlock[37] vssd1 vssd1 vccd1 vccd1 _3040_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput274 io_dataLastBlock[57] vssd1 vssd1 vccd1 vccd1 _3005_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput285 io_dataLastBlock[9] vssd1 vssd1 vccd1 vccd1 _3025_/A0 sky130_fd_sc_hd__buf_1
XFILLER_90_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2820_ _3699_/Q vssd1 vssd1 vccd1 vccd1 _2820_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2751_ _3462_/Q vssd1 vssd1 vccd1 vccd1 _2751_/Y sky130_fd_sc_hd__inv_2
X_1702_ _1742_/A vssd1 vssd1 vccd1 vccd1 _1796_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2682_ _2682_/A _2682_/B input7/X input8/X vssd1 vssd1 vccd1 vccd1 _2682_/Y sky130_fd_sc_hd__nor4_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3303_ _3035_/X _3037_/X _3038_/X _2649_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3303_/X sky130_fd_sc_hd__mux4_2
X_3234_ input19/X input51/X input67/X input83/X _3009_/S _3286_/S1 vssd1 vssd1 vccd1
+ vccd1 _3234_/X sky130_fd_sc_hd__mux4_1
X_3165_ _3675_/Q _3659_/Q _3643_/Q _3619_/Q _3370_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3165_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3096_ _2858_/Y _2859_/Y _2856_/Y _2857_/Y _3102_/S0 _3148_/X vssd1 vssd1 vccd1 vccd1
+ _3096_/X sky130_fd_sc_hd__mux4_2
X_2116_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2116_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2047_ _3739_/Q _2042_/X _1867_/X _2044_/X vssd1 vssd1 vccd1 vccd1 _3739_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2949_ _2949_/A vssd1 vssd1 vccd1 vccd1 _2949_/X sky130_fd_sc_hd__buf_1
XFILLER_1_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_1_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3730_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3852_ _3873_/CLK _3852_/D vssd1 vssd1 vccd1 vccd1 _3852_/Q sky130_fd_sc_hd__dfxtp_1
X_2803_ _3714_/Q vssd1 vssd1 vccd1 vccd1 _2803_/Y sky130_fd_sc_hd__inv_2
X_3783_ _3791_/CLK _3783_/D vssd1 vssd1 vccd1 vccd1 _3783_/Q sky130_fd_sc_hd__dfxtp_1
X_2734_ _3761_/Q vssd1 vssd1 vccd1 vccd1 _2734_/Y sky130_fd_sc_hd__inv_2
X_2665_ _2721_/A _2964_/X vssd1 vssd1 vccd1 vccd1 _2665_/X sky130_fd_sc_hd__and2_1
X_2596_ _3395_/Q _2593_/X _2138_/A _2594_/X vssd1 vssd1 vccd1 vccd1 _3395_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3217_ _3401_/Q _3393_/Q _3385_/Q _3625_/Q _3860_/Q _3861_/Q vssd1 vssd1 vccd1 vccd1
+ _3217_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3148_ _3144_/X _3145_/X _3146_/X _3147_/X _3862_/Q _3863_/Q vssd1 vssd1 vccd1 vccd1
+ _3148_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3079_ _2923_/Y _2924_/Y _2921_/Y _2922_/Y _3153_/X _3132_/S1 vssd1 vssd1 vccd1 vccd1
+ _3079_/X sky130_fd_sc_hd__mux4_2
XFILLER_54_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2450_ _2950_/A vssd1 vssd1 vccd1 vccd1 _2450_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2381_ _3540_/Q _2375_/X _2351_/X _2376_/X vssd1 vssd1 vccd1 vccd1 _3540_/D sky130_fd_sc_hd__a22o_1
X_3002_ _3002_/A0 _3002_/A1 _3009_/S vssd1 vssd1 vccd1 vccd1 _3002_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput5 io_adr_i[2] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_6
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3835_ _3841_/CLK _3835_/D vssd1 vssd1 vccd1 vccd1 _3835_/Q sky130_fd_sc_hd__dfxtp_1
X_3766_ _3823_/CLK _3766_/D vssd1 vssd1 vccd1 vccd1 _3766_/Q sky130_fd_sc_hd__dfxtp_1
X_2717_ _3780_/Q vssd1 vssd1 vccd1 vccd1 _2717_/Y sky130_fd_sc_hd__inv_2
X_3697_ _3730_/CLK _3697_/D vssd1 vssd1 vccd1 vccd1 _3697_/Q sky130_fd_sc_hd__dfxtp_1
X_2648_ _2661_/A _2972_/X vssd1 vssd1 vccd1 vccd1 _2648_/X sky130_fd_sc_hd__and2_1
Xoutput342 _3871_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[23] sky130_fd_sc_hd__clkbuf_2
Xoutput331 _3855_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[13] sky130_fd_sc_hd__clkbuf_2
Xoutput353 _3846_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[4] sky130_fd_sc_hd__clkbuf_2
Xoutput320 _2948_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2579_ _3408_/Q _2573_/X _2546_/X _2574_/X vssd1 vssd1 vccd1 vccd1 _3408_/D sky130_fd_sc_hd__a22o_1
Xoutput364 _3832_/Q vssd1 vssd1 vccd1 vccd1 io_vout[2] sky130_fd_sc_hd__clkbuf_2
XINSDIODE3_4 _3879_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1950_ _2593_/A vssd1 vssd1 vccd1 vccd1 _2594_/A sky130_fd_sc_hd__inv_2
X_1881_ _1881_/A vssd1 vssd1 vccd1 vccd1 _1881_/X sky130_fd_sc_hd__clkbuf_2
X_3620_ _3676_/CLK _3620_/D vssd1 vssd1 vccd1 vccd1 _3620_/Q sky130_fd_sc_hd__dfxtp_1
X_3551_ _3743_/CLK _3551_/D vssd1 vssd1 vccd1 vccd1 _3551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2502_ _2502_/A vssd1 vssd1 vccd1 vccd1 _2502_/X sky130_fd_sc_hd__clkbuf_2
X_3482_ _3603_/CLK _3482_/D vssd1 vssd1 vccd1 vccd1 _3482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2433_ _3502_/Q _2425_/A _2364_/X _2426_/A vssd1 vssd1 vccd1 vccd1 _3502_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2364_ _2944_/A vssd1 vssd1 vccd1 vccd1 _2364_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2295_ _2953_/A vssd1 vssd1 vccd1 vccd1 _2295_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3818_ _3831_/CLK _3818_/D vssd1 vssd1 vccd1 vccd1 _3818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3749_ _3773_/CLK _3749_/D vssd1 vssd1 vccd1 vccd1 _3749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2080_ _3717_/Q _2075_/X _1877_/X _2076_/X vssd1 vssd1 vccd1 vccd1 _3717_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2982_ _2982_/A0 _2982_/A1 _2984_/S vssd1 vssd1 vccd1 vccd1 _2982_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1933_ _2603_/A vssd1 vssd1 vccd1 vccd1 _2604_/A sky130_fd_sc_hd__inv_2
Xinput30 io_b_dat_o_10[10] vssd1 vssd1 vccd1 vccd1 _2631_/B sky130_fd_sc_hd__clkbuf_1
X_1864_ _3821_/Q _1860_/X _1861_/X _1863_/X vssd1 vssd1 vccd1 vccd1 _3821_/D sky130_fd_sc_hd__a22o_1
X_3603_ _3603_/CLK _3603_/D vssd1 vssd1 vccd1 vccd1 _3603_/Q sky130_fd_sc_hd__dfxtp_1
Xinput63 io_b_dat_o_2[11] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
Xinput41 io_b_dat_o_10[6] vssd1 vssd1 vccd1 vccd1 _2645_/B sky130_fd_sc_hd__clkbuf_1
Xinput52 io_b_dat_o_1[1] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
X_1795_ _1795_/A _3316_/X vssd1 vssd1 vccd1 vccd1 _3847_/D sky130_fd_sc_hd__and2_1
Xinput74 io_b_dat_o_2[7] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__clkbuf_1
Xinput96 io_b_dat_o_4[12] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_1
Xinput85 io_b_dat_o_3[2] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__clkbuf_1
X_3534_ _3821_/CLK _3534_/D vssd1 vssd1 vccd1 vccd1 _3534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3465_ _3586_/CLK _3465_/D vssd1 vssd1 vccd1 vccd1 _3465_/Q sky130_fd_sc_hd__dfxtp_1
X_2416_ _2416_/A vssd1 vssd1 vccd1 vccd1 _2416_/X sky130_fd_sc_hd__clkbuf_2
X_3396_ _3895_/CLK _3396_/D vssd1 vssd1 vccd1 vccd1 _3396_/Q sky130_fd_sc_hd__dfxtp_1
X_2347_ _3558_/Q _2340_/A _2269_/X _2341_/A vssd1 vssd1 vccd1 vccd1 _3558_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2278_ _3600_/Q _2272_/X _2265_/X _2273_/X vssd1 vssd1 vccd1 vccd1 _3600_/D sky130_fd_sc_hd__a22o_1
XFILLER_16_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3246_/X _3247_/X _3248_/X _3249_/X _2613_/A _3378_/S1 vssd1 vssd1 vccd1 vccd1
+ _3250_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2201_ _3649_/Q _2197_/X _2143_/X _2198_/X vssd1 vssd1 vccd1 vccd1 _3649_/D sky130_fd_sc_hd__a22o_1
X_3181_ _3592_/Q _3816_/Q _3544_/Q _3520_/Q _3291_/S0 _3292_/S1 vssd1 vssd1 vccd1
+ vccd1 _3181_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2132_ _3686_/Q _2125_/X _2131_/X _2127_/X vssd1 vssd1 vccd1 vccd1 _3686_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2063_ _3727_/Q _2057_/X _1891_/X _2058_/X vssd1 vssd1 vccd1 vccd1 _3727_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2965_ _2965_/A0 _2965_/A1 _3009_/S vssd1 vssd1 vccd1 vccd1 _2965_/X sky130_fd_sc_hd__mux2_1
X_2896_ _3687_/Q vssd1 vssd1 vccd1 vccd1 _2896_/Y sky130_fd_sc_hd__inv_2
X_1916_ _2425_/A vssd1 vssd1 vccd1 vccd1 _1916_/X sky130_fd_sc_hd__buf_2
X_1847_ _2502_/A vssd1 vssd1 vccd1 vccd1 _1847_/X sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_25_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3801_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1778_ _1783_/A _3063_/X vssd1 vssd1 vccd1 vccd1 _3862_/D sky130_fd_sc_hd__and2_1
X_3517_ _3817_/CLK _3517_/D vssd1 vssd1 vccd1 vccd1 _3517_/Q sky130_fd_sc_hd__dfxtp_1
X_3448_ _3816_/CLK _3448_/D vssd1 vssd1 vccd1 vccd1 _3448_/Q sky130_fd_sc_hd__dfxtp_1
X_3379_ input13/X input45/X input61/X input77/X _2996_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3379_/X sky130_fd_sc_hd__mux4_1
XFILLER_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput220 io_dat_i[8] vssd1 vssd1 vccd1 vccd1 _2952_/A sky130_fd_sc_hd__buf_4
Xinput231 io_dataLastBlock[18] vssd1 vssd1 vccd1 vccd1 _3012_/A0 sky130_fd_sc_hd__buf_1
Xinput242 io_dataLastBlock[28] vssd1 vssd1 vccd1 vccd1 _3002_/A0 sky130_fd_sc_hd__buf_1
Xinput253 io_dataLastBlock[38] vssd1 vssd1 vccd1 vccd1 _3036_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput275 io_dataLastBlock[58] vssd1 vssd1 vccd1 vccd1 _3004_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput264 io_dataLastBlock[48] vssd1 vssd1 vccd1 vccd1 _3014_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput286 io_dsi_in[0] vssd1 vssd1 vccd1 vccd1 _2873_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_90_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2750_ _3486_/Q vssd1 vssd1 vccd1 vccd1 _2750_/Y sky130_fd_sc_hd__inv_2
X_1701_ _1802_/A vssd1 vssd1 vccd1 vccd1 _1742_/A sky130_fd_sc_hd__inv_2
X_2681_ _2681_/A _2684_/B _2685_/C vssd1 vssd1 vccd1 vccd1 _2681_/Y sky130_fd_sc_hd__nor3_2
X_3302_ _3302_/A0 _3302_/A1 _3302_/A2 _3302_/A3 _2984_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3302_/X sky130_fd_sc_hd__mux4_1
X_3233_ _3229_/X _3230_/X _3231_/X _3232_/X _3862_/Q _3863_/Q vssd1 vssd1 vccd1 vccd1
+ _3233_/X sky130_fd_sc_hd__mux4_2
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3164_ _3571_/Q _3723_/Q _3707_/Q _3691_/Q _3292_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3164_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2115_ _2239_/A _2181_/B _2675_/A _2115_/D vssd1 vssd1 vccd1 vccd1 _2137_/A sky130_fd_sc_hd__or4_4
X_3095_ _2862_/Y _2863_/Y _2860_/Y _2861_/Y _3153_/X _3132_/S1 vssd1 vssd1 vccd1 vccd1
+ _3095_/X sky130_fd_sc_hd__mux4_2
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2046_ _3740_/Q _2042_/X _1865_/X _2044_/X vssd1 vssd1 vccd1 vccd1 _3740_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2948_ _2948_/A vssd1 vssd1 vccd1 vccd1 _2948_/X sky130_fd_sc_hd__buf_1
X_2879_ _2879_/A _2879_/B _3887_/Q vssd1 vssd1 vccd1 vccd1 _2879_/X sky130_fd_sc_hd__and3_1
XFILLER_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_10 _3876_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3851_ _3851_/CLK _3851_/D vssd1 vssd1 vccd1 vccd1 _3851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3782_ _3791_/CLK _3782_/D vssd1 vssd1 vccd1 vccd1 _3782_/Q sky130_fd_sc_hd__dfxtp_1
X_2802_ _3562_/Q vssd1 vssd1 vccd1 vccd1 _2802_/Y sky130_fd_sc_hd__inv_2
X_2733_ _3769_/Q vssd1 vssd1 vccd1 vccd1 _2733_/Y sky130_fd_sc_hd__inv_2
X_2664_ _2664_/A _3158_/X vssd1 vssd1 vccd1 vccd1 _2664_/X sky130_fd_sc_hd__and2_1
X_2595_ _3396_/Q _2593_/X _2135_/A _2594_/X vssd1 vssd1 vccd1 vccd1 _3396_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3216_ _3433_/Q _3745_/Q _3417_/Q _3409_/Q _3860_/Q _3232_/S1 vssd1 vssd1 vccd1 vccd1
+ _3216_/X sky130_fd_sc_hd__mux4_1
X_3147_ _2701_/Y _2702_/Y _2703_/Y _2704_/Y _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3147_/X sky130_fd_sc_hd__mux4_2
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3078_ _3074_/X _3075_/X _3076_/X _3077_/X _3133_/S0 _3138_/X vssd1 vssd1 vccd1 vccd1
+ _3078_/X sky130_fd_sc_hd__mux4_2
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2029_ _3749_/Q _2022_/X _1877_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _3749_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_40_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3813_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2380_ _3541_/Q _2375_/X _2348_/X _2376_/X vssd1 vssd1 vccd1 vccd1 _3541_/D sky130_fd_sc_hd__a22o_1
X_3001_ _3001_/A0 _3001_/A1 _3009_/S vssd1 vssd1 vccd1 vccd1 _3001_/X sky130_fd_sc_hd__mux2_1
Xinput6 io_adr_i[3] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3834_ _3841_/CLK _3834_/D vssd1 vssd1 vccd1 vccd1 _3834_/Q sky130_fd_sc_hd__dfxtp_1
X_3765_ _3796_/CLK _3765_/D vssd1 vssd1 vccd1 vccd1 _3765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2716_ _3752_/Q vssd1 vssd1 vccd1 vccd1 _2716_/Y sky130_fd_sc_hd__inv_2
X_3696_ _3730_/CLK _3696_/D vssd1 vssd1 vccd1 vccd1 _3696_/Q sky130_fd_sc_hd__dfxtp_1
X_2647_ _2647_/A vssd1 vssd1 vccd1 vccd1 _2661_/A sky130_fd_sc_hd__clkbuf_2
Xoutput310 _2944_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[0] sky130_fd_sc_hd__clkbuf_2
Xoutput343 _3872_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[24] sky130_fd_sc_hd__clkbuf_2
Xoutput332 _3856_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[14] sky130_fd_sc_hd__clkbuf_2
Xoutput321 _2949_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[5] sky130_fd_sc_hd__clkbuf_2
X_2578_ _3409_/Q _2573_/X _2544_/X _2574_/X vssd1 vssd1 vccd1 vccd1 _3409_/D sky130_fd_sc_hd__a22o_1
Xoutput354 _3847_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[5] sky130_fd_sc_hd__clkbuf_2
Xoutput365 _3833_/Q vssd1 vssd1 vccd1 vccd1 io_vout[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_19_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _3812_/Q _1872_/X _1879_/X _1873_/X vssd1 vssd1 vccd1 vccd1 _3812_/D sky130_fd_sc_hd__a22o_1
X_3550_ _3801_/CLK _3550_/D vssd1 vssd1 vccd1 vccd1 _3550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2501_ _2501_/A vssd1 vssd1 vccd1 vccd1 _2501_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3481_ _3603_/CLK _3481_/D vssd1 vssd1 vccd1 vccd1 _3481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2432_ _3503_/Q _2425_/A _2362_/X _2426_/A vssd1 vssd1 vccd1 vccd1 _3503_/D sky130_fd_sc_hd__a22o_1
X_2363_ _3551_/Q _2350_/A _2362_/X _2352_/A vssd1 vssd1 vccd1 vccd1 _3551_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2294_ _3592_/Q _2291_/X _2292_/X _2293_/X vssd1 vssd1 vccd1 vccd1 _3592_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3817_ _3817_/CLK _3817_/D vssd1 vssd1 vccd1 vccd1 _3817_/Q sky130_fd_sc_hd__dfxtp_1
X_3748_ _3748_/CLK _3748_/D vssd1 vssd1 vccd1 vccd1 _3748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3679_ _3727_/CLK _3679_/D vssd1 vssd1 vccd1 vccd1 _3679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2981_ _2980_/X _2618_/X _2981_/S vssd1 vssd1 vccd1 vccd1 _2981_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1932_ _2603_/A vssd1 vssd1 vccd1 vccd1 _1932_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1863_ _1883_/A vssd1 vssd1 vccd1 vccd1 _1863_/X sky130_fd_sc_hd__buf_2
Xinput31 io_b_dat_o_10[11] vssd1 vssd1 vccd1 vccd1 _2637_/B sky130_fd_sc_hd__clkbuf_1
Xinput20 io_b_dat_o_0[1] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_1
X_3602_ _3845_/CLK _3602_/D vssd1 vssd1 vccd1 vccd1 _3602_/Q sky130_fd_sc_hd__dfxtp_1
Xinput64 io_b_dat_o_2[12] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_1
Xinput42 io_b_dat_o_10[7] vssd1 vssd1 vccd1 vccd1 _2662_/B sky130_fd_sc_hd__clkbuf_1
Xinput53 io_b_dat_o_1[2] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_1
X_1794_ _1795_/A _3303_/X vssd1 vssd1 vccd1 vccd1 _3848_/D sky130_fd_sc_hd__and2_1
Xinput86 io_b_dat_o_3[3] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__clkbuf_1
Xinput75 io_b_dat_o_2[8] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__clkbuf_1
Xinput97 io_b_dat_o_4[13] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_1
X_3533_ _3823_/CLK _3533_/D vssd1 vssd1 vccd1 vccd1 _3533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3464_ _3811_/CLK _3464_/D vssd1 vssd1 vccd1 vccd1 _3464_/Q sky130_fd_sc_hd__dfxtp_1
X_2415_ _3516_/Q _2409_/X _2351_/X _2410_/X vssd1 vssd1 vccd1 vccd1 _3516_/D sky130_fd_sc_hd__a22o_1
X_3395_ _3897_/CLK _3395_/D vssd1 vssd1 vccd1 vccd1 _3395_/Q sky130_fd_sc_hd__dfxtp_1
X_2346_ _3559_/Q _2340_/X _2267_/X _2341_/X vssd1 vssd1 vccd1 vccd1 _3559_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2277_ _3601_/Q _2272_/X _2263_/X _2273_/X vssd1 vssd1 vccd1 vccd1 _3601_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2200_ _3650_/Q _2197_/X _2141_/X _2198_/X vssd1 vssd1 vccd1 vccd1 _3650_/D sky130_fd_sc_hd__a22o_1
X_3180_ _3672_/Q _3656_/Q _3640_/Q _3616_/Q _3292_/S0 _3192_/S1 vssd1 vssd1 vccd1
+ vccd1 _3180_/X sky130_fd_sc_hd__mux4_2
X_2131_ _2952_/A vssd1 vssd1 vccd1 vccd1 _2131_/X sky130_fd_sc_hd__clkbuf_2
X_2062_ _3728_/Q _2057_/X _1889_/X _2058_/X vssd1 vssd1 vccd1 vccd1 _3728_/D sky130_fd_sc_hd__a22o_1
X_2964_ _2964_/A0 _2964_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _2964_/X sky130_fd_sc_hd__mux2_2
XFILLER_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1915_ _2009_/A _2476_/B _2151_/A _1915_/D vssd1 vssd1 vccd1 vccd1 _2425_/A sky130_fd_sc_hd__or4_4
X_2895_ _3703_/Q vssd1 vssd1 vccd1 vccd1 _2895_/Y sky130_fd_sc_hd__inv_2
X_1846_ _2501_/A vssd1 vssd1 vccd1 vccd1 _2502_/A sky130_fd_sc_hd__inv_2
X_1777_ _1783_/A _3072_/X vssd1 vssd1 vccd1 vccd1 _3863_/D sky130_fd_sc_hd__and2_1
X_3516_ _3812_/CLK _3516_/D vssd1 vssd1 vccd1 vccd1 _3516_/Q sky130_fd_sc_hd__dfxtp_1
X_3447_ _3826_/CLK _3447_/D vssd1 vssd1 vccd1 vccd1 _3447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3378_ _3374_/X _3375_/X _3376_/X _3377_/X _2613_/A _3378_/S1 vssd1 vssd1 vccd1 vccd1
+ _3378_/X sky130_fd_sc_hd__mux4_1
X_2329_ _3571_/Q _2321_/X _2328_/X _2324_/X vssd1 vssd1 vccd1 vccd1 _3571_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput210 io_dat_i[28] vssd1 vssd1 vccd1 vccd1 input210/X sky130_fd_sc_hd__buf_1
XFILLER_0_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput232 io_dataLastBlock[19] vssd1 vssd1 vccd1 vccd1 _3011_/A0 sky130_fd_sc_hd__buf_1
Xinput221 io_dat_i[9] vssd1 vssd1 vccd1 vccd1 _2953_/A sky130_fd_sc_hd__buf_4
Xinput243 io_dataLastBlock[29] vssd1 vssd1 vccd1 vccd1 _3001_/A0 sky130_fd_sc_hd__buf_1
Xinput254 io_dataLastBlock[39] vssd1 vssd1 vccd1 vccd1 _3032_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput287 io_dsi_in[1] vssd1 vssd1 vccd1 vccd1 _2873_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput276 io_dataLastBlock[59] vssd1 vssd1 vccd1 vccd1 _3003_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput265 io_dataLastBlock[49] vssd1 vssd1 vccd1 vccd1 _3013_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1700_ _1700_/A vssd1 vssd1 vccd1 vccd1 _1700_/Y sky130_fd_sc_hd__inv_2
X_2680_ _2681_/A _2684_/B _2684_/C vssd1 vssd1 vccd1 vccd1 _2680_/Y sky130_fd_sc_hd__nor3_2
XFILLER_8_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3301_ input25/X input57/X input73/X input89/X _2996_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3301_/X sky130_fd_sc_hd__mux4_1
X_3232_ _3398_/Q _3390_/Q _3382_/Q _3622_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3232_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3163_ _3159_/X _3160_/X _3161_/X _3162_/X _3295_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3163_/X sky130_fd_sc_hd__mux4_2
X_2114_ _3694_/Q _2107_/A _1893_/X _2108_/A vssd1 vssd1 vccd1 vccd1 _3694_/D sky130_fd_sc_hd__a22o_1
X_3094_ _2866_/Y _2867_/Y _2864_/Y _2865_/Y _3153_/X _3132_/S1 vssd1 vssd1 vccd1 vccd1
+ _3094_/X sky130_fd_sc_hd__mux4_2
X_2045_ _3741_/Q _2042_/X _1861_/X _2044_/X vssd1 vssd1 vccd1 vccd1 _3741_/D sky130_fd_sc_hd__a22o_1
XFILLER_62_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2947_ _2947_/A vssd1 vssd1 vccd1 vccd1 _2947_/X sky130_fd_sc_hd__buf_1
X_2878_ _2872_/Y _2878_/A2 _1740_/X _2878_/B2 _2874_/Y vssd1 vssd1 vccd1 vccd1 _2879_/B
+ sky130_fd_sc_hd__a221o_1
X_1829_ _1966_/A vssd1 vssd1 vccd1 vccd1 _1829_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_11 _2174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3850_ _3867_/CLK _3850_/D vssd1 vssd1 vccd1 vccd1 _3850_/Q sky130_fd_sc_hd__dfxtp_1
X_3781_ _3829_/CLK _3781_/D vssd1 vssd1 vccd1 vccd1 _3781_/Q sky130_fd_sc_hd__dfxtp_1
X_2801_ _3729_/Q vssd1 vssd1 vccd1 vccd1 _2801_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2732_ _3773_/Q vssd1 vssd1 vccd1 vccd1 _2732_/Y sky130_fd_sc_hd__inv_2
X_2663_ _2843_/A _2983_/X vssd1 vssd1 vccd1 vccd1 _2663_/X sky130_fd_sc_hd__and2_1
X_2594_ _2594_/A vssd1 vssd1 vccd1 vccd1 _2594_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3215_ _3529_/Q _3505_/Q _3481_/Q _3457_/Q _3860_/Q _3232_/S1 vssd1 vssd1 vccd1 vccd1
+ _3215_/X sky130_fd_sc_hd__mux4_2
XFILLER_82_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3146_ _2697_/Y _2698_/Y _2699_/Y _2700_/Y _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3146_/X sky130_fd_sc_hd__mux4_1
X_3077_ _2927_/Y _2928_/Y _2925_/Y _2926_/Y _3132_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3077_/X sky130_fd_sc_hd__mux4_2
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2028_ _3750_/Q _2022_/X _2019_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _3750_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3000_ _3000_/A0 _3000_/A1 _3009_/S vssd1 vssd1 vccd1 vccd1 _3000_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 io_adr_i[4] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_2
XFILLER_36_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3833_ _3841_/CLK _3833_/D vssd1 vssd1 vccd1 vccd1 _3833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3764_ _3828_/CLK _3764_/D vssd1 vssd1 vccd1 vccd1 _3764_/Q sky130_fd_sc_hd__dfxtp_1
X_2715_ _3804_/Q vssd1 vssd1 vccd1 vccd1 _2715_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3695_ _3727_/CLK _3695_/D vssd1 vssd1 vccd1 vccd1 _3695_/Q sky130_fd_sc_hd__dfxtp_1
X_2646_ _2654_/A _2646_/B vssd1 vssd1 vccd1 vccd1 _2646_/X sky130_fd_sc_hd__and2_1
Xoutput300 _2684_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_1 sky130_fd_sc_hd__clkbuf_2
Xoutput344 _3873_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[25] sky130_fd_sc_hd__clkbuf_2
Xoutput333 _3857_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[15] sky130_fd_sc_hd__clkbuf_2
Xoutput322 _2950_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[6] sky130_fd_sc_hd__clkbuf_2
Xoutput311 _2954_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[10] sky130_fd_sc_hd__clkbuf_2
X_2577_ _3410_/Q _2573_/X _2542_/X _2574_/X vssd1 vssd1 vccd1 vccd1 _3410_/D sky130_fd_sc_hd__a22o_1
Xoutput355 _3848_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[6] sky130_fd_sc_hd__clkbuf_2
Xoutput366 _3834_/Q vssd1 vssd1 vccd1 vccd1 io_vout[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3129_ _2752_/Y _2753_/Y _2750_/Y _2751_/Y _3132_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3129_/X sky130_fd_sc_hd__mux4_2
XPHY_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2500_ _3461_/Q _1845_/X _2448_/X _1847_/X vssd1 vssd1 vccd1 vccd1 _3461_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3480_ _3811_/CLK _3480_/D vssd1 vssd1 vccd1 vccd1 _3480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2431_ _3504_/Q _2425_/X _2360_/X _2426_/X vssd1 vssd1 vccd1 vccd1 _3504_/D sky130_fd_sc_hd__a22o_1
X_2362_ _2945_/A vssd1 vssd1 vccd1 vccd1 _2362_/X sky130_fd_sc_hd__clkbuf_2
X_2293_ _2302_/A vssd1 vssd1 vccd1 vccd1 _2293_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3897_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3816_ _3816_/CLK _3816_/D vssd1 vssd1 vccd1 vccd1 _3816_/Q sky130_fd_sc_hd__dfxtp_1
X_3747_ _3747_/CLK _3747_/D vssd1 vssd1 vccd1 vccd1 _3747_/Q sky130_fd_sc_hd__dfxtp_1
X_3678_ _3727_/CLK _3678_/D vssd1 vssd1 vccd1 vccd1 _3678_/Q sky130_fd_sc_hd__dfxtp_1
X_2629_ _2644_/A _3183_/X vssd1 vssd1 vccd1 vccd1 _2629_/X sky130_fd_sc_hd__and2_1
XFILLER_87_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2980_ _2980_/A0 _2980_/A1 _2984_/S vssd1 vssd1 vccd1 vccd1 _2980_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1931_ _1985_/A _1977_/B _2510_/C _1964_/D vssd1 vssd1 vccd1 vccd1 _2603_/A sky130_fd_sc_hd__or4_4
X_1862_ _1881_/A vssd1 vssd1 vccd1 vccd1 _1883_/A sky130_fd_sc_hd__inv_2
Xinput21 io_b_dat_o_0[2] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_1
Xinput10 io_adr_i[7] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
X_3601_ _3747_/CLK _3601_/D vssd1 vssd1 vccd1 vccd1 _3601_/Q sky130_fd_sc_hd__dfxtp_1
Xinput32 io_b_dat_o_10[12] vssd1 vssd1 vccd1 vccd1 _2646_/B sky130_fd_sc_hd__clkbuf_1
Xinput43 io_b_dat_o_10[8] vssd1 vssd1 vccd1 vccd1 _2618_/B sky130_fd_sc_hd__clkbuf_1
Xinput54 io_b_dat_o_1[3] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_1
X_1793_ _1795_/A _3290_/X vssd1 vssd1 vccd1 vccd1 _3849_/D sky130_fd_sc_hd__and2_1
Xinput76 io_b_dat_o_2[9] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_1
Xinput87 io_b_dat_o_3[4] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_1
Xinput65 io_b_dat_o_2[13] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_1
Xinput98 io_b_dat_o_4[14] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_1
X_3532_ _3726_/CLK _3532_/D vssd1 vssd1 vccd1 vccd1 _3532_/Q sky130_fd_sc_hd__dfxtp_1
X_3463_ _3731_/CLK _3463_/D vssd1 vssd1 vccd1 vccd1 _3463_/Q sky130_fd_sc_hd__dfxtp_1
X_2414_ _3517_/Q _2409_/X _2348_/X _2410_/X vssd1 vssd1 vccd1 vccd1 _3517_/D sky130_fd_sc_hd__a22o_1
X_3394_ _3867_/CLK _3394_/D vssd1 vssd1 vccd1 vccd1 _3394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2345_ _3560_/Q _2340_/X _2265_/X _2341_/X vssd1 vssd1 vccd1 vccd1 _3560_/D sky130_fd_sc_hd__a22o_1
X_2276_ _3602_/Q _2272_/X _2261_/X _2273_/X vssd1 vssd1 vccd1 vccd1 _3602_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2130_ _3687_/Q _2125_/X _2129_/X _2127_/X vssd1 vssd1 vccd1 vccd1 _3687_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2061_ _3729_/Q _2057_/X _1887_/X _2058_/X vssd1 vssd1 vccd1 vccd1 _3729_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2963_ _2962_/X _2666_/X _2981_/S vssd1 vssd1 vccd1 vccd1 _2963_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1914_ input4/X vssd1 vssd1 vccd1 vccd1 _2009_/A sky130_fd_sc_hd__buf_1
X_2894_ _3719_/Q vssd1 vssd1 vccd1 vccd1 _2894_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1845_ _2501_/A vssd1 vssd1 vccd1 vccd1 _1845_/X sky130_fd_sc_hd__buf_2
X_1776_ _1796_/A vssd1 vssd1 vccd1 vccd1 _1783_/A sky130_fd_sc_hd__buf_1
X_3515_ _3807_/CLK _3515_/D vssd1 vssd1 vccd1 vccd1 _3515_/Q sky130_fd_sc_hd__dfxtp_1
X_3446_ _3816_/CLK _3446_/D vssd1 vssd1 vccd1 vccd1 _3446_/Q sky130_fd_sc_hd__dfxtp_1
X_3377_ _3398_/Q _3390_/Q _3382_/Q _3622_/Q _3377_/S0 _1905_/B vssd1 vssd1 vccd1 vccd1
+ _3377_/X sky130_fd_sc_hd__mux4_2
X_2328_ _2957_/A vssd1 vssd1 vccd1 vccd1 _2328_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2259_ _2259_/A vssd1 vssd1 vccd1 vccd1 _2259_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_34_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3826_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput200 io_dat_i[19] vssd1 vssd1 vccd1 vccd1 input200/X sky130_fd_sc_hd__buf_1
Xinput211 io_dat_i[29] vssd1 vssd1 vccd1 vccd1 input211/X sky130_fd_sc_hd__buf_1
Xinput233 io_dataLastBlock[1] vssd1 vssd1 vccd1 vccd1 _3056_/A0 sky130_fd_sc_hd__buf_1
Xinput222 io_dataLastBlock[0] vssd1 vssd1 vccd1 vccd1 _3060_/A0 sky130_fd_sc_hd__buf_1
Xinput244 io_dataLastBlock[2] vssd1 vssd1 vccd1 vccd1 _3052_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput277 io_dataLastBlock[5] vssd1 vssd1 vccd1 vccd1 _3040_/A0 sky130_fd_sc_hd__buf_1
Xinput266 io_dataLastBlock[4] vssd1 vssd1 vccd1 vccd1 _3044_/A0 sky130_fd_sc_hd__buf_1
Xinput288 io_dsi_in[2] vssd1 vssd1 vccd1 vccd1 _2875_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput255 io_dataLastBlock[3] vssd1 vssd1 vccd1 vccd1 _3048_/A0 sky130_fd_sc_hd__buf_1
XFILLER_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3300_ _3296_/X _3297_/X _3298_/X _3299_/X _2613_/A _3378_/S1 vssd1 vssd1 vccd1 vccd1
+ _3300_/X sky130_fd_sc_hd__mux4_1
X_3231_ _3430_/Q _3742_/Q _3414_/Q _3406_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3231_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3162_ _3500_/Q _3476_/Q _3452_/Q _3740_/Q _3292_/S0 _3292_/S1 vssd1 vssd1 vccd1
+ vccd1 _3162_/X sky130_fd_sc_hd__mux4_1
X_2113_ _3695_/Q _2107_/X _1891_/X _2108_/X vssd1 vssd1 vccd1 vccd1 _3695_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3093_ _3089_/X _3090_/X _3091_/X _3092_/X _3133_/S0 _3138_/X vssd1 vssd1 vccd1 vccd1
+ _3093_/X sky130_fd_sc_hd__mux4_2
XFILLER_81_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2044_ _2058_/A vssd1 vssd1 vccd1 vccd1 _2044_/X sky130_fd_sc_hd__clkbuf_2
X_2946_ _2946_/A vssd1 vssd1 vccd1 vccd1 _2946_/X sky130_fd_sc_hd__buf_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2877_ _2872_/Y _2877_/A2 _1740_/X _2877_/B2 _3886_/Q vssd1 vssd1 vccd1 vccd1 _2879_/A
+ sky130_fd_sc_hd__a221o_1
X_1828_ _2955_/A vssd1 vssd1 vccd1 vccd1 _1966_/A sky130_fd_sc_hd__clkbuf_2
X_1759_ _1762_/A _3000_/X vssd1 vssd1 vccd1 vccd1 _3878_/D sky130_fd_sc_hd__nor2b_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3429_ _3773_/CLK _3429_/D vssd1 vssd1 vccd1 vccd1 _3429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_12 _2956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3780_ _3828_/CLK _3780_/D vssd1 vssd1 vccd1 vccd1 _3780_/Q sky130_fd_sc_hd__dfxtp_1
X_2800_ _3441_/Q vssd1 vssd1 vccd1 vccd1 _2800_/Y sky130_fd_sc_hd__inv_2
X_2731_ _3757_/Q vssd1 vssd1 vccd1 vccd1 _2731_/Y sky130_fd_sc_hd__inv_2
X_2662_ _2836_/A _2662_/B vssd1 vssd1 vccd1 vccd1 _2662_/X sky130_fd_sc_hd__and2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2593_ _2593_/A vssd1 vssd1 vccd1 vccd1 _2593_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3214_ _3425_/Q _3601_/Q _3577_/Q _3553_/Q _3860_/Q _3232_/S1 vssd1 vssd1 vccd1 vccd1
+ _3214_/X sky130_fd_sc_hd__mux4_2
XFILLER_79_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3145_ _2693_/Y _2694_/Y _2695_/Y _2696_/Y _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3145_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3076_ _2931_/Y _2932_/Y _2929_/Y _2930_/Y _3132_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3076_/X sky130_fd_sc_hd__mux4_2
XFILLER_70_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2027_ _3751_/Q _2022_/X _2017_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _3751_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2929_ _3673_/Q vssd1 vssd1 vccd1 vccd1 _2929_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 io_adr_i[5] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_4
XFILLER_76_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3832_ _3832_/CLK _3832_/D vssd1 vssd1 vccd1 vccd1 _3832_/Q sky130_fd_sc_hd__dfxtp_1
X_3763_ _3791_/CLK _3763_/D vssd1 vssd1 vccd1 vccd1 _3763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2714_ _3824_/Q vssd1 vssd1 vccd1 vccd1 _2714_/Y sky130_fd_sc_hd__inv_2
X_3694_ _3821_/CLK _3694_/D vssd1 vssd1 vccd1 vccd1 _3694_/Q sky130_fd_sc_hd__dfxtp_1
X_2645_ _2654_/A _2645_/B vssd1 vssd1 vccd1 vccd1 _2645_/X sky130_fd_sc_hd__and2_1
XFILLER_10_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput301 _2672_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_10 sky130_fd_sc_hd__clkbuf_2
Xoutput334 _3864_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[16] sky130_fd_sc_hd__clkbuf_2
Xoutput323 _2951_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[7] sky130_fd_sc_hd__clkbuf_2
Xoutput312 _2955_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[11] sky130_fd_sc_hd__clkbuf_2
Xoutput345 _3874_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[26] sky130_fd_sc_hd__clkbuf_2
X_2576_ _3411_/Q _2573_/X _2540_/X _2574_/X vssd1 vssd1 vccd1 vccd1 _3411_/D sky130_fd_sc_hd__a22o_1
Xoutput356 _3849_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[7] sky130_fd_sc_hd__clkbuf_2
Xoutput367 _3835_/Q vssd1 vssd1 vccd1 vccd1 io_vout[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3128_ _3124_/X _3125_/X _3126_/X _3127_/X _3133_/S0 _3138_/X vssd1 vssd1 vccd1 vccd1
+ _3128_/X sky130_fd_sc_hd__mux4_2
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3059_ _3885_/Q _3373_/X _3061_/S vssd1 vssd1 vccd1 vccd1 _3059_/X sky130_fd_sc_hd__mux2_2
XPHY_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2430_ _3505_/Q _2425_/X _2358_/X _2426_/X vssd1 vssd1 vccd1 vccd1 _3505_/D sky130_fd_sc_hd__a22o_1
X_2361_ _3552_/Q _2350_/X _2360_/X _2352_/X vssd1 vssd1 vccd1 vccd1 _3552_/D sky130_fd_sc_hd__a22o_1
X_2292_ _2954_/A vssd1 vssd1 vccd1 vccd1 _2292_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_59_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3667_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3815_ _3816_/CLK _3815_/D vssd1 vssd1 vccd1 vccd1 _3815_/Q sky130_fd_sc_hd__dfxtp_1
X_3746_ _3746_/CLK _3746_/D vssd1 vssd1 vccd1 vccd1 _3746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3677_ _3677_/CLK _3677_/D vssd1 vssd1 vccd1 vccd1 _3677_/Q sky130_fd_sc_hd__dfxtp_1
X_2628_ _3895_/Q _1717_/B _1723_/C vssd1 vssd1 vccd1 vccd1 _2628_/X sky130_fd_sc_hd__a21bo_1
X_2559_ _3424_/Q _2553_/X _2546_/X _2554_/X vssd1 vssd1 vccd1 vccd1 _3424_/D sky130_fd_sc_hd__a22o_1
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1930_ _2021_/D vssd1 vssd1 vccd1 vccd1 _1964_/D sky130_fd_sc_hd__buf_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1861_ _2959_/A vssd1 vssd1 vccd1 vccd1 _1861_/X sky130_fd_sc_hd__clkbuf_2
Xinput22 io_b_dat_o_0[3] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_1
Xinput11 io_adr_i[8] vssd1 vssd1 vccd1 vccd1 _3053_/S sky130_fd_sc_hd__clkbuf_8
X_3600_ _3845_/CLK _3600_/D vssd1 vssd1 vccd1 vccd1 _3600_/Q sky130_fd_sc_hd__dfxtp_1
Xinput44 io_b_dat_o_10[9] vssd1 vssd1 vccd1 vccd1 _2625_/B sky130_fd_sc_hd__clkbuf_1
Xinput55 io_b_dat_o_1[4] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_1
Xinput33 io_b_dat_o_10[13] vssd1 vssd1 vccd1 vccd1 _2654_/B sky130_fd_sc_hd__clkbuf_1
X_1792_ _1795_/A _3277_/X vssd1 vssd1 vccd1 vccd1 _3850_/D sky130_fd_sc_hd__and2_1
X_3531_ _3604_/CLK _3531_/D vssd1 vssd1 vccd1 vccd1 _3531_/Q sky130_fd_sc_hd__dfxtp_1
Xinput88 io_b_dat_o_3[5] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__clkbuf_1
Xinput66 io_b_dat_o_2[14] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_1
Xinput77 io_b_dat_o_3[0] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_1
Xinput99 io_b_dat_o_4[15] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__clkbuf_1
X_3462_ _3812_/CLK _3462_/D vssd1 vssd1 vccd1 vccd1 _3462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3393_ _3896_/CLK _3393_/D vssd1 vssd1 vccd1 vccd1 _3393_/Q sky130_fd_sc_hd__dfxtp_1
X_2413_ _3518_/Q _2409_/X _2297_/X _2410_/X vssd1 vssd1 vccd1 vccd1 _3518_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2344_ _3561_/Q _2340_/X _2263_/X _2341_/X vssd1 vssd1 vccd1 vccd1 _3561_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2275_ _3603_/Q _2272_/X _2258_/X _2273_/X vssd1 vssd1 vccd1 vccd1 _3603_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3729_ _3731_/CLK _3729_/D vssd1 vssd1 vccd1 vccd1 _3729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_4_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3811_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2060_ _3730_/Q _2057_/X _1885_/X _2058_/X vssd1 vssd1 vccd1 vccd1 _3730_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2962_ _2962_/A0 _2962_/A1 _3009_/S vssd1 vssd1 vccd1 vccd1 _2962_/X sky130_fd_sc_hd__mux2_1
X_1913_ _3798_/Q _1907_/X _1840_/X _1909_/X vssd1 vssd1 vccd1 vccd1 _3798_/D sky130_fd_sc_hd__a22o_1
X_2893_ _3567_/Q vssd1 vssd1 vccd1 vccd1 _2893_/Y sky130_fd_sc_hd__inv_2
X_1844_ _2510_/A _2476_/B _2151_/A _1915_/D vssd1 vssd1 vccd1 vccd1 _2501_/A sky130_fd_sc_hd__or4_4
X_1775_ _1775_/A _3014_/X vssd1 vssd1 vccd1 vccd1 _3864_/D sky130_fd_sc_hd__nor2b_4
XFILLER_8_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3514_ _3586_/CLK _3514_/D vssd1 vssd1 vccd1 vccd1 _3514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3445_ _3817_/CLK _3445_/D vssd1 vssd1 vccd1 vccd1 _3445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3376_ _3430_/Q _3742_/Q _3414_/Q _3406_/Q _3377_/S0 _1905_/B vssd1 vssd1 vccd1 vccd1
+ _3376_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2327_ _3572_/Q _2321_/X _2326_/X _2324_/X vssd1 vssd1 vccd1 vccd1 _3572_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2258_ _2949_/A vssd1 vssd1 vccd1 vccd1 _2258_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2189_ _3657_/Q _2182_/X _2123_/X _2184_/X vssd1 vssd1 vccd1 vccd1 _3657_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput201 io_dat_i[1] vssd1 vssd1 vccd1 vccd1 _2945_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput223 io_dataLastBlock[10] vssd1 vssd1 vccd1 vccd1 _3022_/A0 sky130_fd_sc_hd__buf_1
Xinput212 io_dat_i[2] vssd1 vssd1 vccd1 vccd1 _2946_/A sky130_fd_sc_hd__clkbuf_4
Xinput234 io_dataLastBlock[20] vssd1 vssd1 vccd1 vccd1 _3010_/A0 sky130_fd_sc_hd__buf_1
Xinput245 io_dataLastBlock[30] vssd1 vssd1 vccd1 vccd1 _3000_/A0 sky130_fd_sc_hd__buf_1
Xinput278 io_dataLastBlock[60] vssd1 vssd1 vccd1 vccd1 _3002_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput267 io_dataLastBlock[50] vssd1 vssd1 vccd1 vccd1 _3012_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput256 io_dataLastBlock[40] vssd1 vssd1 vccd1 vccd1 _3028_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput289 io_dsi_in[3] vssd1 vssd1 vccd1 vccd1 _2875_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_90_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3230_ _3526_/Q _3502_/Q _3478_/Q _3454_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3230_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3161_ _3596_/Q _3820_/Q _3548_/Q _3524_/Q _3292_/S0 _3292_/S1 vssd1 vssd1 vccd1
+ vccd1 _3161_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2112_ _3696_/Q _2107_/X _1889_/X _2108_/X vssd1 vssd1 vccd1 vccd1 _3696_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3092_ _2870_/Y _2871_/Y _2868_/Y _2869_/Y _3102_/S0 _3148_/X vssd1 vssd1 vccd1 vccd1
+ _3092_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2043_ _2057_/A vssd1 vssd1 vccd1 vccd1 _2058_/A sky130_fd_sc_hd__inv_2
XFILLER_47_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2945_ _2945_/A vssd1 vssd1 vccd1 vccd1 _2945_/X sky130_fd_sc_hd__clkbuf_1
X_2876_ _3887_/Q vssd1 vssd1 vccd1 vccd1 _2876_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1827_ _2467_/A vssd1 vssd1 vccd1 vccd1 _1827_/X sky130_fd_sc_hd__buf_2
X_1758_ _1762_/A _2999_/X vssd1 vssd1 vccd1 vccd1 _3879_/D sky130_fd_sc_hd__nor2b_4
XFILLER_2_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1689_ _3899_/Q _1681_/Y _1682_/Y _1681_/A _1707_/B vssd1 vssd1 vccd1 vccd1 _1689_/X
+ sky130_fd_sc_hd__o221a_1
X_3428_ _3627_/CLK _3428_/D vssd1 vssd1 vccd1 vccd1 _3428_/Q sky130_fd_sc_hd__dfxtp_1
X_3359_ _3487_/Q _3463_/Q _3439_/Q _3727_/Q _3370_/S0 _1905_/B vssd1 vssd1 vccd1 vccd1
+ _3359_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2730_ _3801_/Q vssd1 vssd1 vccd1 vccd1 _2730_/Y sky130_fd_sc_hd__inv_2
X_2661_ _2661_/A _2966_/X vssd1 vssd1 vccd1 vccd1 _2661_/X sky130_fd_sc_hd__and2_1
XFILLER_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2592_ _3397_/Q _1949_/X _2133_/A _1951_/X vssd1 vssd1 vccd1 vccd1 _3397_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3213_ _3209_/X _3210_/X _3211_/X _3212_/X _3862_/Q _3863_/Q vssd1 vssd1 vccd1 vccd1
+ _3213_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3144_ _2689_/Y _2690_/Y _2691_/Y _2692_/Y _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3144_/X sky130_fd_sc_hd__mux4_2
XFILLER_82_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3075_ _2935_/Y _2936_/Y _2933_/Y _2934_/Y _3132_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3075_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2026_ _3752_/Q _2022_/X _2015_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _3752_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2928_ _3689_/Q vssd1 vssd1 vccd1 vccd1 _2928_/Y sky130_fd_sc_hd__inv_2
X_2859_ _3613_/Q vssd1 vssd1 vccd1 vccd1 _2859_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 io_adr_i[6] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_1
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3831_ _3831_/CLK _3831_/D vssd1 vssd1 vccd1 vccd1 _3831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3762_ _3796_/CLK _3762_/D vssd1 vssd1 vccd1 vccd1 _3762_/Q sky130_fd_sc_hd__dfxtp_1
X_2713_ _3828_/Q vssd1 vssd1 vccd1 vccd1 _2713_/Y sky130_fd_sc_hd__inv_2
X_3693_ _3727_/CLK _3693_/D vssd1 vssd1 vccd1 vccd1 _3693_/Q sky130_fd_sc_hd__dfxtp_1
X_2644_ _2644_/A _2973_/X vssd1 vssd1 vccd1 vccd1 _2644_/X sky130_fd_sc_hd__and2_1
Xoutput335 _3865_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[17] sky130_fd_sc_hd__clkbuf_2
X_2575_ _3412_/Q _2573_/X _2537_/X _2574_/X vssd1 vssd1 vccd1 vccd1 _3412_/D sky130_fd_sc_hd__a22o_1
Xoutput302 _2683_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_2 sky130_fd_sc_hd__clkbuf_2
Xoutput324 _2952_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[8] sky130_fd_sc_hd__clkbuf_2
Xoutput313 _2956_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[12] sky130_fd_sc_hd__clkbuf_2
Xoutput346 _3875_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[27] sky130_fd_sc_hd__clkbuf_2
Xoutput357 _3850_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[8] sky130_fd_sc_hd__clkbuf_2
Xoutput368 _3836_/Q vssd1 vssd1 vccd1 vccd1 io_vout[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3127_ _2756_/Y _2757_/Y _2754_/Y _2755_/Y _3132_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3127_/X sky130_fd_sc_hd__mux4_1
X_3058_ _3366_/X _3367_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3058_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2009_ _2009_/A _2009_/B _2065_/A _2009_/D vssd1 vssd1 vccd1 vccd1 _2272_/A sky130_fd_sc_hd__or4_4
XPHY_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2360_ _2946_/A vssd1 vssd1 vccd1 vccd1 _2360_/X sky130_fd_sc_hd__clkbuf_2
X_2291_ _2301_/A vssd1 vssd1 vccd1 vccd1 _2291_/X sky130_fd_sc_hd__buf_2
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3814_ _3816_/CLK _3814_/D vssd1 vssd1 vccd1 vccd1 _3814_/Q sky130_fd_sc_hd__dfxtp_1
X_3745_ _3747_/CLK _3745_/D vssd1 vssd1 vccd1 vccd1 _3745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3676_ _3676_/CLK _3676_/D vssd1 vssd1 vccd1 vccd1 _3676_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_28_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3889_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2627_ _3894_/Q _1716_/B _1717_/B vssd1 vssd1 vccd1 vccd1 _2627_/X sky130_fd_sc_hd__a21bo_1
XFILLER_87_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2558_ _3425_/Q _2553_/X _2544_/X _2554_/X vssd1 vssd1 vccd1 vccd1 _3425_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2489_ _3470_/Q _2485_/X _1974_/A _2486_/X vssd1 vssd1 vccd1 vccd1 _3470_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1860_ _1881_/A vssd1 vssd1 vccd1 vccd1 _1860_/X sky130_fd_sc_hd__buf_2
X_1791_ _1795_/A _3269_/X vssd1 vssd1 vccd1 vccd1 _3851_/D sky130_fd_sc_hd__and2_1
Xinput12 io_adr_i[9] vssd1 vssd1 vccd1 vccd1 _2943_/A sky130_fd_sc_hd__clkbuf_4
Xinput23 io_b_dat_o_0[4] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_1
Xinput34 io_b_dat_o_10[14] vssd1 vssd1 vccd1 vccd1 _2660_/B sky130_fd_sc_hd__clkbuf_1
Xinput45 io_b_dat_o_1[0] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
X_3530_ _3530_/CLK _3530_/D vssd1 vssd1 vccd1 vccd1 _3530_/Q sky130_fd_sc_hd__dfxtp_1
Xinput78 io_b_dat_o_3[10] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__clkbuf_1
Xinput56 io_b_dat_o_1[5] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_1
Xinput89 io_b_dat_o_3[6] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_1
Xinput67 io_b_dat_o_2[15] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_1
X_3461_ _3823_/CLK _3461_/D vssd1 vssd1 vccd1 vccd1 _3461_/Q sky130_fd_sc_hd__dfxtp_1
X_3392_ _3867_/CLK _3392_/D vssd1 vssd1 vccd1 vccd1 _3392_/Q sky130_fd_sc_hd__dfxtp_1
X_2412_ _3519_/Q _2409_/X _2295_/X _2410_/X vssd1 vssd1 vccd1 vccd1 _3519_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2343_ _3562_/Q _2340_/X _2261_/X _2341_/X vssd1 vssd1 vccd1 vccd1 _3562_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2274_ _3604_/Q _2272_/X _2255_/X _2273_/X vssd1 vssd1 vccd1 vccd1 _3604_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1989_ _3769_/Q _1986_/X _1966_/X _1988_/X vssd1 vssd1 vccd1 vccd1 _3769_/D sky130_fd_sc_hd__a22o_1
X_3728_ _3731_/CLK _3728_/D vssd1 vssd1 vccd1 vccd1 _3728_/Q sky130_fd_sc_hd__dfxtp_1
X_3659_ _3677_/CLK _3659_/D vssd1 vssd1 vccd1 vccd1 _3659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2961_ _2943_/A _3378_/S1 _2961_/S vssd1 vssd1 vccd1 vccd1 _2961_/X sky130_fd_sc_hd__mux2_8
XFILLER_15_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1912_ _3799_/Q _1907_/X _1837_/X _1909_/X vssd1 vssd1 vccd1 vccd1 _3799_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2892_ _3734_/Q vssd1 vssd1 vccd1 vccd1 _2892_/Y sky130_fd_sc_hd__inv_2
X_1843_ _2021_/B vssd1 vssd1 vccd1 vccd1 _2476_/B sky130_fd_sc_hd__clkbuf_2
X_1774_ _1774_/A _3013_/X vssd1 vssd1 vccd1 vccd1 _3865_/D sky130_fd_sc_hd__nor2b_4
X_3513_ _3811_/CLK _3513_/D vssd1 vssd1 vccd1 vccd1 _3513_/Q sky130_fd_sc_hd__dfxtp_1
X_3444_ _3812_/CLK _3444_/D vssd1 vssd1 vccd1 vccd1 _3444_/Q sky130_fd_sc_hd__dfxtp_1
X_3375_ _3526_/Q _3502_/Q _3478_/Q _3454_/Q _3377_/S0 _1905_/B vssd1 vssd1 vccd1 vccd1
+ _3375_/X sky130_fd_sc_hd__mux4_2
X_2326_ _2958_/A vssd1 vssd1 vccd1 vccd1 _2326_/X sky130_fd_sc_hd__clkbuf_2
Xrepeater410 _1905_/A vssd1 vssd1 vccd1 vccd1 _3364_/S0 sky130_fd_sc_hd__buf_6
X_2257_ _2257_/A vssd1 vssd1 vccd1 vccd1 _2257_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2188_ _3658_/Q _2182_/X _2163_/X _2184_/X vssd1 vssd1 vccd1 vccd1 _3658_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3720_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput202 io_dat_i[20] vssd1 vssd1 vccd1 vccd1 input202/X sky130_fd_sc_hd__buf_1
XFILLER_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput224 io_dataLastBlock[11] vssd1 vssd1 vccd1 vccd1 _3019_/A0 sky130_fd_sc_hd__buf_1
XFILLER_0_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput235 io_dataLastBlock[21] vssd1 vssd1 vccd1 vccd1 _3009_/A0 sky130_fd_sc_hd__buf_1
Xinput213 io_dat_i[30] vssd1 vssd1 vccd1 vccd1 input213/X sky130_fd_sc_hd__buf_1
XFILLER_88_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput279 io_dataLastBlock[61] vssd1 vssd1 vccd1 vccd1 _3001_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput268 io_dataLastBlock[51] vssd1 vssd1 vccd1 vccd1 _3011_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput257 io_dataLastBlock[41] vssd1 vssd1 vccd1 vccd1 _3025_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput246 io_dataLastBlock[31] vssd1 vssd1 vccd1 vccd1 _2999_/A0 sky130_fd_sc_hd__buf_1
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3160_ _3676_/Q _3660_/Q _3644_/Q _3620_/Q _3370_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3160_/X sky130_fd_sc_hd__mux4_2
X_3091_ _2883_/Y _2884_/Y _2881_/Y _2882_/Y _3102_/S0 _3148_/X vssd1 vssd1 vccd1 vccd1
+ _3091_/X sky130_fd_sc_hd__mux4_2
X_2111_ _3697_/Q _2107_/X _1887_/X _2108_/X vssd1 vssd1 vccd1 vccd1 _3697_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2042_ _2057_/A vssd1 vssd1 vccd1 vccd1 _2042_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2944_ _2944_/A vssd1 vssd1 vccd1 vccd1 _2944_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2875_ _2872_/Y _2875_/A2 _1740_/X _2875_/B2 _2874_/Y vssd1 vssd1 vccd1 vccd1 _2875_/X
+ sky130_fd_sc_hd__a221o_1
X_1826_ _2510_/A _2510_/B _2151_/A _1915_/D vssd1 vssd1 vccd1 vccd1 _2467_/A sky130_fd_sc_hd__or4_4
X_1757_ _1775_/A vssd1 vssd1 vccd1 vccd1 _1762_/A sky130_fd_sc_hd__buf_4
XFILLER_89_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1688_ _1688_/A _1688_/B _1688_/C _1688_/D vssd1 vssd1 vccd1 vccd1 _1707_/B sky130_fd_sc_hd__or4_4
X_3427_ _3747_/CLK _3427_/D vssd1 vssd1 vccd1 vccd1 _3427_/Q sky130_fd_sc_hd__dfxtp_1
X_3358_ _3583_/Q _3807_/Q _3535_/Q _3511_/Q _3372_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3358_/X sky130_fd_sc_hd__mux4_2
X_2309_ _3581_/Q _1978_/X _2253_/X _1980_/X vssd1 vssd1 vccd1 vccd1 _3581_/D sky130_fd_sc_hd__a22o_1
X_3289_ _3289_/A0 _3289_/A1 _3289_/A2 _3289_/A3 _2984_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3289_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2660_ _2836_/A _2660_/B vssd1 vssd1 vccd1 vccd1 _2660_/X sky130_fd_sc_hd__and2_1
XFILLER_12_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2591_ _3398_/Q _2583_/A _2550_/X _2584_/A vssd1 vssd1 vccd1 vccd1 _3398_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3212_ _3402_/Q _3394_/Q _3386_/Q _3626_/Q _3860_/Q _3861_/Q vssd1 vssd1 vccd1 vccd1
+ _3212_/X sky130_fd_sc_hd__mux4_1
X_3143_ _3139_/X _3140_/X _3141_/X _3142_/X _3862_/Q _3863_/Q vssd1 vssd1 vccd1 vccd1
+ _3143_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3074_ _2939_/Y _2940_/Y _2937_/Y _2938_/Y _3132_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3074_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2025_ _3753_/Q _2022_/X _2011_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _3753_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2927_ _3705_/Q vssd1 vssd1 vccd1 vccd1 _2927_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2858_ _3637_/Q vssd1 vssd1 vccd1 vccd1 _2858_/Y sky130_fd_sc_hd__inv_2
X_1809_ _1816_/B vssd1 vssd1 vccd1 vccd1 _1814_/B sky130_fd_sc_hd__buf_1
X_2789_ _3681_/Q vssd1 vssd1 vccd1 vccd1 _2789_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3830_ _3831_/CLK _3830_/D vssd1 vssd1 vccd1 vccd1 _3830_/Q sky130_fd_sc_hd__dfxtp_1
X_3761_ _3890_/CLK _3761_/D vssd1 vssd1 vccd1 vccd1 _3761_/Q sky130_fd_sc_hd__dfxtp_1
X_2712_ _3796_/Q vssd1 vssd1 vccd1 vccd1 _2712_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3692_ _3724_/CLK _3692_/D vssd1 vssd1 vccd1 vccd1 _3692_/Q sky130_fd_sc_hd__dfxtp_1
X_2643_ _2644_/A _3173_/X vssd1 vssd1 vccd1 vccd1 _2643_/X sky130_fd_sc_hd__and2_1
X_2574_ _2574_/A vssd1 vssd1 vccd1 vccd1 _2574_/X sky130_fd_sc_hd__clkbuf_2
Xoutput303 _2682_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_3 sky130_fd_sc_hd__clkbuf_2
Xoutput325 _2953_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[9] sky130_fd_sc_hd__clkbuf_2
Xoutput314 _2957_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[13] sky130_fd_sc_hd__clkbuf_2
Xoutput347 _3876_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[28] sky130_fd_sc_hd__clkbuf_2
Xoutput336 _3866_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[18] sky130_fd_sc_hd__clkbuf_2
Xoutput358 _3851_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[9] sky130_fd_sc_hd__clkbuf_2
Xoutput369 _3837_/Q vssd1 vssd1 vccd1 vccd1 io_vout[7] sky130_fd_sc_hd__clkbuf_2
X_3126_ _2760_/Y _2761_/Y _2758_/Y _2759_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3126_/X sky130_fd_sc_hd__mux4_2
X_3057_ _3365_/X _3056_/X _3061_/S vssd1 vssd1 vccd1 vccd1 _3057_/X sky130_fd_sc_hd__mux2_2
XFILLER_35_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2008_ _3758_/Q _2002_/X _1974_/X _2004_/X vssd1 vssd1 vccd1 vccd1 _3758_/D sky130_fd_sc_hd__a22o_1
XPHY_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2290_ _3593_/Q _2282_/X _2289_/X _2284_/X vssd1 vssd1 vccd1 vccd1 _3593_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3813_ _3813_/CLK _3813_/D vssd1 vssd1 vccd1 vccd1 _3813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3744_ _3746_/CLK _3744_/D vssd1 vssd1 vccd1 vccd1 _3744_/Q sky130_fd_sc_hd__dfxtp_1
X_3675_ _3677_/CLK _3675_/D vssd1 vssd1 vccd1 vccd1 _3675_/Q sky130_fd_sc_hd__dfxtp_1
X_2626_ _2638_/A _2979_/X vssd1 vssd1 vccd1 vccd1 _2626_/X sky130_fd_sc_hd__and2_1
X_2557_ _3426_/Q _2553_/X _2542_/X _2554_/X vssd1 vssd1 vccd1 vccd1 _3426_/D sky130_fd_sc_hd__a22o_1
X_2488_ _3471_/Q _2485_/X _1972_/A _2486_/X vssd1 vssd1 vccd1 vccd1 _3471_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3109_ _2816_/Y _2817_/Y _2814_/Y _2815_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3109_/X sky130_fd_sc_hd__mux4_2
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 io_b_dat_o_0[0] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
X_1790_ _1796_/A vssd1 vssd1 vccd1 vccd1 _1795_/A sky130_fd_sc_hd__buf_1
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput46 io_b_dat_o_1[10] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_1
Xinput24 io_b_dat_o_0[5] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_1
Xinput35 io_b_dat_o_10[15] vssd1 vssd1 vccd1 vccd1 _2666_/B sky130_fd_sc_hd__clkbuf_1
Xinput79 io_b_dat_o_3[11] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_1
Xinput57 io_b_dat_o_1[6] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_1
Xinput68 io_b_dat_o_2[1] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_1
X_3460_ _3726_/CLK _3460_/D vssd1 vssd1 vccd1 vccd1 _3460_/Q sky130_fd_sc_hd__dfxtp_1
X_3391_ _3895_/CLK _3391_/D vssd1 vssd1 vccd1 vccd1 _3391_/Q sky130_fd_sc_hd__dfxtp_1
X_2411_ _3520_/Q _2409_/X _2292_/X _2410_/X vssd1 vssd1 vccd1 vccd1 _3520_/D sky130_fd_sc_hd__a22o_1
X_2342_ _3563_/Q _2340_/X _2258_/X _2341_/X vssd1 vssd1 vccd1 vccd1 _3563_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2273_ _2273_/A vssd1 vssd1 vccd1 vccd1 _2273_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3727_ _3727_/CLK _3727_/D vssd1 vssd1 vccd1 vccd1 _3727_/Q sky130_fd_sc_hd__dfxtp_1
X_1988_ _2352_/A vssd1 vssd1 vccd1 vccd1 _1988_/X sky130_fd_sc_hd__clkbuf_2
X_3658_ _3676_/CLK _3658_/D vssd1 vssd1 vccd1 vccd1 _3658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2609_ _3384_/Q _2603_/X _2145_/A _2604_/X vssd1 vssd1 vccd1 vccd1 _3384_/D sky130_fd_sc_hd__a22o_1
X_3589_ _3813_/CLK _3589_/D vssd1 vssd1 vccd1 vccd1 _3589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2960_ _2960_/A vssd1 vssd1 vccd1 vccd1 _2960_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2891_ _3446_/Q vssd1 vssd1 vccd1 vccd1 _2891_/Y sky130_fd_sc_hd__inv_2
X_1911_ _3800_/Q _1907_/X _1834_/X _1909_/X vssd1 vssd1 vccd1 vccd1 _3800_/D sky130_fd_sc_hd__a22o_1
XPHY_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1842_ input1/X vssd1 vssd1 vccd1 vccd1 _2021_/B sky130_fd_sc_hd__inv_2
X_1773_ _1774_/A _3012_/X vssd1 vssd1 vccd1 vccd1 _3866_/D sky130_fd_sc_hd__nor2b_4
X_3512_ _3586_/CLK _3512_/D vssd1 vssd1 vccd1 vccd1 _3512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3443_ _3731_/CLK _3443_/D vssd1 vssd1 vccd1 vccd1 _3443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3374_ _3422_/Q _3598_/Q _3574_/Q _3550_/Q _3377_/S0 _1905_/B vssd1 vssd1 vccd1 vccd1
+ _3374_/X sky130_fd_sc_hd__mux4_1
Xrepeater400 _2971_/S vssd1 vssd1 vccd1 vccd1 _3009_/S sky130_fd_sc_hd__buf_8
X_2325_ _3573_/Q _2321_/X _2322_/X _2324_/X vssd1 vssd1 vccd1 vccd1 _3573_/D sky130_fd_sc_hd__a22o_1
Xrepeater411 input5/X vssd1 vssd1 vccd1 vccd1 _1905_/A sky130_fd_sc_hd__buf_8
XFILLER_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2256_ _3612_/Q _2248_/X _2255_/X _2249_/X vssd1 vssd1 vccd1 vccd1 _3612_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2187_ _3659_/Q _2182_/X _2161_/X _2184_/X vssd1 vssd1 vccd1 vccd1 _3659_/D sky130_fd_sc_hd__a22o_1
XFILLER_92_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_12_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3845_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput225 io_dataLastBlock[12] vssd1 vssd1 vccd1 vccd1 _2973_/A0 sky130_fd_sc_hd__buf_1
Xinput236 io_dataLastBlock[22] vssd1 vssd1 vccd1 vccd1 _3008_/A0 sky130_fd_sc_hd__buf_1
Xinput203 io_dat_i[21] vssd1 vssd1 vccd1 vccd1 input203/X sky130_fd_sc_hd__buf_1
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput214 io_dat_i[31] vssd1 vssd1 vccd1 vccd1 input214/X sky130_fd_sc_hd__buf_1
Xinput269 io_dataLastBlock[52] vssd1 vssd1 vccd1 vccd1 _3010_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput258 io_dataLastBlock[42] vssd1 vssd1 vccd1 vccd1 _3022_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput247 io_dataLastBlock[32] vssd1 vssd1 vccd1 vccd1 _3060_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2110_ _3698_/Q _2107_/X _1885_/X _2108_/X vssd1 vssd1 vccd1 vccd1 _3698_/D sky130_fd_sc_hd__a22o_1
X_3090_ _2887_/Y _2888_/Y _2885_/Y _2886_/Y _3102_/S0 _3148_/X vssd1 vssd1 vccd1 vccd1
+ _3090_/X sky130_fd_sc_hd__mux4_2
X_2041_ _2239_/A _2181_/B _2682_/A _2115_/D vssd1 vssd1 vccd1 vccd1 _2057_/A sky130_fd_sc_hd__or4_4
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2943_ _2943_/A vssd1 vssd1 vccd1 vccd1 _2943_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2874_ _3886_/Q vssd1 vssd1 vccd1 vccd1 _2874_/Y sky130_fd_sc_hd__inv_2
X_1825_ _2021_/D vssd1 vssd1 vccd1 vccd1 _1915_/D sky130_fd_sc_hd__buf_1
X_1756_ _1857_/A input2/X _1802_/A _1823_/C vssd1 vssd1 vccd1 vccd1 _1775_/A sky130_fd_sc_hd__or4_4
X_1687_ _3898_/Q _3883_/Q _3898_/Q _3883_/Q vssd1 vssd1 vccd1 vccd1 _1688_/D sky130_fd_sc_hd__a2bb2oi_1
X_3426_ _3845_/CLK _3426_/D vssd1 vssd1 vccd1 vccd1 _3426_/Q sky130_fd_sc_hd__dfxtp_1
X_3357_ _3663_/Q _3647_/Q _3631_/Q _3607_/Q _3370_/S0 _3357_/S1 vssd1 vssd1 vccd1
+ vccd1 _3357_/X sky130_fd_sc_hd__mux4_2
X_2308_ _3582_/Q _2301_/A _2269_/X _2302_/A vssd1 vssd1 vccd1 vccd1 _3582_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3288_ input26/X input58/X input74/X input90/X _2984_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3288_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2239_ _2239_/A _2476_/B _2673_/A _2281_/D vssd1 vssd1 vccd1 vccd1 _2257_/A sky130_fd_sc_hd__or4_4
XFILLER_53_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2590_ _3399_/Q _2583_/A _2548_/X _2584_/A vssd1 vssd1 vccd1 vccd1 _3399_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3211_ _3434_/Q _3746_/Q _3418_/Q _3410_/Q _3860_/Q _3861_/Q vssd1 vssd1 vccd1 vccd1
+ _3211_/X sky130_fd_sc_hd__mux4_1
X_3142_ _2719_/Y _2720_/Y _2722_/Y _2723_/Y _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3142_/X sky130_fd_sc_hd__mux4_1
X_3073_ _1707_/X _3896_/Q _3073_/S vssd1 vssd1 vccd1 vccd1 _3073_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2024_ _2031_/A vssd1 vssd1 vccd1 vccd1 _2024_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2926_ _3721_/Q vssd1 vssd1 vccd1 vccd1 _2926_/Y sky130_fd_sc_hd__inv_2
X_2857_ _3653_/Q vssd1 vssd1 vccd1 vccd1 _2857_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1808_ _3098_/X _1808_/B vssd1 vssd1 vccd1 vccd1 _3837_/D sky130_fd_sc_hd__nor2_1
X_2788_ _3697_/Q vssd1 vssd1 vccd1 vccd1 _2788_/Y sky130_fd_sc_hd__inv_2
X_1739_ _3886_/Q _1734_/X _2147_/A _1736_/X _1703_/X vssd1 vssd1 vccd1 vccd1 _3886_/D
+ sky130_fd_sc_hd__o221a_1
X_3409_ _3746_/CLK _3409_/D vssd1 vssd1 vccd1 vccd1 _3409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3760_ _3796_/CLK _3760_/D vssd1 vssd1 vccd1 vccd1 _3760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2711_ _3760_/Q vssd1 vssd1 vccd1 vccd1 _2711_/Y sky130_fd_sc_hd__inv_2
X_3691_ _3723_/CLK _3691_/D vssd1 vssd1 vccd1 vccd1 _3691_/Q sky130_fd_sc_hd__dfxtp_1
X_2642_ _3890_/Q _1712_/B _1713_/B vssd1 vssd1 vccd1 vccd1 _2642_/X sky130_fd_sc_hd__a21bo_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2573_ _2573_/A vssd1 vssd1 vccd1 vccd1 _2573_/X sky130_fd_sc_hd__clkbuf_2
Xoutput326 _2960_/X vssd1 vssd1 vccd1 vccd1 io_b_we_i sky130_fd_sc_hd__clkbuf_2
Xoutput304 _2681_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_4 sky130_fd_sc_hd__clkbuf_2
Xoutput315 _2958_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[14] sky130_fd_sc_hd__clkbuf_2
Xoutput348 _3877_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[29] sky130_fd_sc_hd__clkbuf_2
Xoutput337 _3867_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[19] sky130_fd_sc_hd__clkbuf_2
Xoutput359 _2880_/X vssd1 vssd1 vccd1 vccd1 io_dsi_o sky130_fd_sc_hd__clkbuf_2
XFILLER_67_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3125_ _2764_/Y _2765_/Y _2762_/Y _2763_/Y _3132_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3125_/X sky130_fd_sc_hd__mux4_2
XFILLER_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3056_ _3056_/A0 _3056_/A1 _3060_/S vssd1 vssd1 vccd1 vccd1 _3056_/X sky130_fd_sc_hd__mux2_2
X_2007_ _3759_/Q _2002_/X _1972_/X _2004_/X vssd1 vssd1 vccd1 vccd1 _3759_/D sky130_fd_sc_hd__a22o_1
XFILLER_63_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3889_ _3889_/CLK _3889_/D vssd1 vssd1 vccd1 vccd1 _3889_/Q sky130_fd_sc_hd__dfxtp_1
X_2909_ _3568_/Q vssd1 vssd1 vccd1 vccd1 _2909_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3812_ _3812_/CLK _3812_/D vssd1 vssd1 vccd1 vccd1 _3812_/Q sky130_fd_sc_hd__dfxtp_1
X_3743_ _3743_/CLK _3743_/D vssd1 vssd1 vccd1 vccd1 _3743_/Q sky130_fd_sc_hd__dfxtp_1
X_3674_ _3676_/CLK _3674_/D vssd1 vssd1 vccd1 vccd1 _3674_/Q sky130_fd_sc_hd__dfxtp_1
X_2625_ _2637_/A _2625_/B vssd1 vssd1 vccd1 vccd1 _2625_/X sky130_fd_sc_hd__and2_1
X_2556_ _3427_/Q _2553_/X _2540_/X _2554_/X vssd1 vssd1 vccd1 vccd1 _3427_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2487_ _3472_/Q _2485_/X _1970_/A _2486_/X vssd1 vssd1 vccd1 vccd1 _3472_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3108_ _3104_/X _3105_/X _3106_/X _3107_/X _3133_/S0 _3138_/X vssd1 vssd1 vccd1 vccd1
+ _3108_/X sky130_fd_sc_hd__mux4_2
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3039_ _3883_/Q _3308_/X _3061_/S vssd1 vssd1 vccd1 vccd1 _3039_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_37_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3812_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput14 io_b_dat_o_0[10] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_1
Xinput25 io_b_dat_o_0[6] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_1
Xinput36 io_b_dat_o_10[1] vssd1 vssd1 vccd1 vccd1 _2836_/B sky130_fd_sc_hd__clkbuf_1
Xinput47 io_b_dat_o_1[11] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
Xinput58 io_b_dat_o_1[7] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_1
Xinput69 io_b_dat_o_2[2] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2410_ _2417_/A vssd1 vssd1 vccd1 vccd1 _2410_/X sky130_fd_sc_hd__clkbuf_2
X_3390_ _3890_/CLK _3390_/D vssd1 vssd1 vccd1 vccd1 _3390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2341_ _2341_/A vssd1 vssd1 vccd1 vccd1 _2341_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2272_ _2272_/A vssd1 vssd1 vccd1 vccd1 _2272_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1987_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2352_/A sky130_fd_sc_hd__inv_2
X_3726_ _3726_/CLK _3726_/D vssd1 vssd1 vccd1 vccd1 _3726_/Q sky130_fd_sc_hd__dfxtp_1
X_3657_ _3723_/CLK _3657_/D vssd1 vssd1 vccd1 vccd1 _3657_/Q sky130_fd_sc_hd__dfxtp_1
X_2608_ _3385_/Q _2603_/X _2143_/A _2604_/X vssd1 vssd1 vccd1 vccd1 _3385_/D sky130_fd_sc_hd__a22o_1
X_3588_ _3812_/CLK _3588_/D vssd1 vssd1 vccd1 vccd1 _3588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2539_ _3436_/Q _2536_/X _2537_/X _2538_/X vssd1 vssd1 vccd1 vccd1 _3436_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2890_ _3470_/Q vssd1 vssd1 vccd1 vccd1 _2890_/Y sky130_fd_sc_hd__inv_2
X_1910_ _3801_/Q _1907_/X _1829_/X _1909_/X vssd1 vssd1 vccd1 vccd1 _3801_/D sky130_fd_sc_hd__a22o_1
XPHY_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1841_ _3826_/Q _1827_/X _1840_/X _1831_/X vssd1 vssd1 vccd1 vccd1 _3826_/D sky130_fd_sc_hd__a22o_1
XPHY_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1772_ _1774_/A _3011_/X vssd1 vssd1 vccd1 vccd1 _3867_/D sky130_fd_sc_hd__nor2b_4
X_3511_ _3726_/CLK _3511_/D vssd1 vssd1 vccd1 vccd1 _3511_/Q sky130_fd_sc_hd__dfxtp_1
X_3442_ _3714_/CLK _3442_/D vssd1 vssd1 vccd1 vccd1 _3442_/Q sky130_fd_sc_hd__dfxtp_1
X_3373_ _3369_/X _3370_/X _3371_/X _3372_/X _3373_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3373_/X sky130_fd_sc_hd__mux4_2
XFILLER_69_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2324_ _2341_/A vssd1 vssd1 vccd1 vccd1 _2324_/X sky130_fd_sc_hd__clkbuf_2
Xrepeater401 _2984_/S vssd1 vssd1 vccd1 vccd1 _2996_/S sky130_fd_sc_hd__buf_8
XFILLER_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater412 input2/X vssd1 vssd1 vccd1 vccd1 _2961_/S sky130_fd_sc_hd__buf_8
X_2255_ _2950_/A vssd1 vssd1 vccd1 vccd1 _2255_/X sky130_fd_sc_hd__buf_2
X_2186_ _3660_/Q _2182_/X _2159_/X _2184_/X vssd1 vssd1 vccd1 vccd1 _3660_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3709_ _3741_/CLK _3709_/D vssd1 vssd1 vccd1 vccd1 _3709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput226 io_dataLastBlock[13] vssd1 vssd1 vccd1 vccd1 _2970_/A0 sky130_fd_sc_hd__buf_1
Xinput215 io_dat_i[3] vssd1 vssd1 vccd1 vccd1 _2947_/A sky130_fd_sc_hd__clkbuf_4
Xinput204 io_dat_i[22] vssd1 vssd1 vccd1 vccd1 input204/X sky130_fd_sc_hd__buf_1
Xinput259 io_dataLastBlock[43] vssd1 vssd1 vccd1 vccd1 _3019_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput237 io_dataLastBlock[23] vssd1 vssd1 vccd1 vccd1 _3007_/A0 sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_52_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3821_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput248 io_dataLastBlock[33] vssd1 vssd1 vccd1 vccd1 _3056_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_84_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2040_ _2040_/A vssd1 vssd1 vccd1 vccd1 _2682_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2942_ _3053_/S vssd1 vssd1 vccd1 vccd1 _2942_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2873_ _2872_/Y _2873_/A2 _1740_/X _2873_/B2 _3886_/Q vssd1 vssd1 vccd1 vccd1 _2873_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_30_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1824_ _3053_/S input3/X input2/X _1824_/D vssd1 vssd1 vccd1 vccd1 _2021_/D sky130_fd_sc_hd__or4_4
X_1755_ _2943_/A vssd1 vssd1 vccd1 vccd1 _1823_/C sky130_fd_sc_hd__inv_2
X_1686_ _1682_/Y _3884_/Q _1682_/Y _3884_/Q vssd1 vssd1 vccd1 vccd1 _1688_/C sky130_fd_sc_hd__a2bb2o_1
X_3425_ _3747_/CLK _3425_/D vssd1 vssd1 vccd1 vccd1 _3425_/Q sky130_fd_sc_hd__dfxtp_1
X_3356_ _3559_/Q _3711_/Q _3695_/Q _3679_/Q _3370_/S0 _1905_/B vssd1 vssd1 vccd1 vccd1
+ _3356_/X sky130_fd_sc_hd__mux4_2
X_3287_ _3283_/X _3284_/X _3285_/X _3286_/X _2613_/A _3378_/S1 vssd1 vssd1 vccd1 vccd1
+ _3287_/X sky130_fd_sc_hd__mux4_1
X_2307_ _3583_/Q _2301_/X _2267_/X _2302_/X vssd1 vssd1 vccd1 vccd1 _3583_/D sky130_fd_sc_hd__a22o_1
X_2238_ _3622_/Q _2230_/A _2149_/X _2231_/A vssd1 vssd1 vccd1 vccd1 _3622_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2169_ _3671_/Q _2166_/X _2129_/X _2167_/X vssd1 vssd1 vccd1 vccd1 _3671_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3210_ _3530_/Q _3506_/Q _3482_/Q _3458_/Q _3860_/Q _3232_/S1 vssd1 vssd1 vccd1 vccd1
+ _3210_/X sky130_fd_sc_hd__mux4_2
X_3141_ _2715_/Y _2716_/Y _2717_/Y _2718_/Y _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3141_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3072_ _1689_/X _3899_/Q _3073_/S vssd1 vssd1 vccd1 vccd1 _3072_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2023_ _2030_/A vssd1 vssd1 vccd1 vccd1 _2031_/A sky130_fd_sc_hd__inv_2
XFILLER_47_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2925_ _3569_/Q vssd1 vssd1 vccd1 vccd1 _2925_/Y sky130_fd_sc_hd__inv_2
X_2856_ _3669_/Q vssd1 vssd1 vccd1 vccd1 _2856_/Y sky130_fd_sc_hd__inv_2
X_1807_ _3093_/X _1808_/B vssd1 vssd1 vccd1 vccd1 _3838_/D sky130_fd_sc_hd__nor2_1
X_2787_ _3713_/Q vssd1 vssd1 vccd1 vccd1 _2787_/Y sky130_fd_sc_hd__inv_2
X_1738_ _2945_/A vssd1 vssd1 vccd1 vccd1 _2147_/A sky130_fd_sc_hd__clkbuf_2
X_3408_ _3851_/CLK _3408_/D vssd1 vssd1 vccd1 vccd1 _3408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3339_ _3335_/X _3336_/X _3337_/X _3338_/X _2613_/A _3378_/S1 vssd1 vssd1 vccd1 vccd1
+ _3339_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2710_ _3768_/Q vssd1 vssd1 vccd1 vccd1 _2710_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3690_ _3723_/CLK _3690_/D vssd1 vssd1 vccd1 vccd1 _3690_/Q sky130_fd_sc_hd__dfxtp_1
X_2641_ _3889_/Q _3888_/Q _1712_/B vssd1 vssd1 vccd1 vccd1 _2641_/X sky130_fd_sc_hd__a21bo_1
X_2572_ _3413_/Q _1965_/X _2534_/X _1968_/X vssd1 vssd1 vccd1 vccd1 _3413_/D sky130_fd_sc_hd__a22o_1
Xoutput305 _2680_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_5 sky130_fd_sc_hd__clkbuf_2
Xoutput316 _2959_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput327 _3842_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[0] sky130_fd_sc_hd__clkbuf_2
Xoutput338 _3843_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[1] sky130_fd_sc_hd__clkbuf_2
Xoutput349 _3844_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3124_ _2768_/Y _2769_/Y _2766_/Y _2767_/Y _3132_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3124_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3055_ _3886_/Q _3360_/X _3061_/S vssd1 vssd1 vccd1 vccd1 _3055_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2006_ _3760_/Q _2002_/X _1970_/X _2004_/X vssd1 vssd1 vccd1 vccd1 _3760_/D sky130_fd_sc_hd__a22o_1
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2908_ _3735_/Q vssd1 vssd1 vccd1 vccd1 _2908_/Y sky130_fd_sc_hd__inv_2
X_3888_ _3889_/CLK _3888_/D vssd1 vssd1 vccd1 vccd1 _3888_/Q sky130_fd_sc_hd__dfxtp_1
X_2839_ _3668_/Q vssd1 vssd1 vccd1 vccd1 _2839_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3726_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3811_ _3811_/CLK _3811_/D vssd1 vssd1 vccd1 vccd1 _3811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3742_ _3801_/CLK _3742_/D vssd1 vssd1 vccd1 vccd1 _3742_/Q sky130_fd_sc_hd__dfxtp_1
X_3673_ _3724_/CLK _3673_/D vssd1 vssd1 vccd1 vccd1 _3673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2624_ _2644_/A _3188_/X vssd1 vssd1 vccd1 vccd1 _2624_/X sky130_fd_sc_hd__and2_1
X_2555_ _3428_/Q _2553_/X _2537_/X _2554_/X vssd1 vssd1 vccd1 vccd1 _3428_/D sky130_fd_sc_hd__a22o_1
X_2486_ _2493_/A vssd1 vssd1 vccd1 vccd1 _2486_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3107_ _2820_/Y _2821_/Y _2818_/Y _2819_/Y _3132_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3107_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3038_ _3301_/X _3302_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3038_/X sky130_fd_sc_hd__mux2_1
XPHY_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput15 io_b_dat_o_0[11] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_1
Xinput26 io_b_dat_o_0[7] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_1
Xinput37 io_b_dat_o_10[2] vssd1 vssd1 vccd1 vccd1 _2640_/B sky130_fd_sc_hd__clkbuf_1
Xinput48 io_b_dat_o_1[12] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_1
Xinput59 io_b_dat_o_1[8] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2340_ _2340_/A vssd1 vssd1 vccd1 vccd1 _2340_/X sky130_fd_sc_hd__clkbuf_2
X_2271_ _3605_/Q _2010_/X _2253_/X _2013_/X vssd1 vssd1 vccd1 vccd1 _3605_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1986_ _2350_/A vssd1 vssd1 vccd1 vccd1 _1986_/X sky130_fd_sc_hd__clkbuf_2
X_3725_ _3821_/CLK _3725_/D vssd1 vssd1 vccd1 vccd1 _3725_/Q sky130_fd_sc_hd__dfxtp_1
X_3656_ _3672_/CLK _3656_/D vssd1 vssd1 vccd1 vccd1 _3656_/Q sky130_fd_sc_hd__dfxtp_1
X_2607_ _3386_/Q _2603_/X _2141_/A _2604_/X vssd1 vssd1 vccd1 vccd1 _3386_/D sky130_fd_sc_hd__a22o_1
X_3587_ _3731_/CLK _3587_/D vssd1 vssd1 vccd1 vccd1 _3587_/Q sky130_fd_sc_hd__dfxtp_1
X_2538_ _2538_/A vssd1 vssd1 vccd1 vccd1 _2538_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2469_ _3484_/Q _2467_/X _2450_/X _2468_/X vssd1 vssd1 vccd1 vccd1 _3484_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1840_ _1974_/A vssd1 vssd1 vccd1 vccd1 _1840_/X sky130_fd_sc_hd__clkbuf_2
XPHY_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1771_ _1774_/A _3010_/X vssd1 vssd1 vccd1 vccd1 _3868_/D sky130_fd_sc_hd__nor2b_4
XFILLER_8_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3510_ _3821_/CLK _3510_/D vssd1 vssd1 vccd1 vccd1 _3510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3441_ _3586_/CLK _3441_/D vssd1 vssd1 vccd1 vccd1 _3441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3372_ _3486_/Q _3462_/Q _3438_/Q _3726_/Q _3372_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3372_/X sky130_fd_sc_hd__mux4_2
X_2323_ _2340_/A vssd1 vssd1 vccd1 vccd1 _2341_/A sky130_fd_sc_hd__inv_2
Xrepeater402 _2971_/S vssd1 vssd1 vccd1 vccd1 _2984_/S sky130_fd_sc_hd__buf_8
XFILLER_84_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater413 _3053_/S vssd1 vssd1 vccd1 vccd1 _3061_/S sky130_fd_sc_hd__buf_8
X_2254_ _3613_/Q _2248_/X _2253_/X _2249_/X vssd1 vssd1 vccd1 vccd1 _3613_/D sky130_fd_sc_hd__a22o_1
X_2185_ _3661_/Q _2182_/X _2155_/X _2184_/X vssd1 vssd1 vccd1 vccd1 _3661_/D sky130_fd_sc_hd__a22o_1
XFILLER_92_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1969_ _3777_/Q _1965_/X _1966_/X _1968_/X vssd1 vssd1 vccd1 vccd1 _3777_/D sky130_fd_sc_hd__a22o_1
X_3708_ _3722_/CLK _3708_/D vssd1 vssd1 vccd1 vccd1 _3708_/Q sky130_fd_sc_hd__dfxtp_1
X_3639_ _3687_/CLK _3639_/D vssd1 vssd1 vccd1 vccd1 _3639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput227 io_dataLastBlock[14] vssd1 vssd1 vccd1 vccd1 _2967_/A0 sky130_fd_sc_hd__buf_1
Xinput216 io_dat_i[4] vssd1 vssd1 vccd1 vccd1 _2948_/A sky130_fd_sc_hd__clkbuf_4
Xinput205 io_dat_i[23] vssd1 vssd1 vccd1 vccd1 input205/X sky130_fd_sc_hd__buf_1
Xinput238 io_dataLastBlock[24] vssd1 vssd1 vccd1 vccd1 _3006_/A0 sky130_fd_sc_hd__buf_1
Xinput249 io_dataLastBlock[34] vssd1 vssd1 vccd1 vccd1 _3052_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_84_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3895_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2941_ _1689_/X _1700_/A _3899_/Q _1700_/Y _1721_/A vssd1 vssd1 vccd1 vccd1 _3899_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2872_ _3885_/Q vssd1 vssd1 vccd1 vccd1 _2872_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1823_ _2686_/A _1823_/B _1823_/C vssd1 vssd1 vccd1 vccd1 _1824_/D sky130_fd_sc_hd__or3_1
X_1754_ _3053_/S vssd1 vssd1 vccd1 vccd1 _1857_/A sky130_fd_sc_hd__inv_2
XFILLER_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1685_ _1707_/A _3881_/Q _1707_/A _3881_/Q vssd1 vssd1 vccd1 vccd1 _1688_/B sky130_fd_sc_hd__a2bb2o_1
X_3424_ _3845_/CLK _3424_/D vssd1 vssd1 vccd1 vccd1 _3424_/Q sky130_fd_sc_hd__dfxtp_1
X_3355_ _3051_/X _3053_/X _3054_/X _2630_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3355_/X sky130_fd_sc_hd__mux4_1
X_3286_ _3405_/Q _3397_/Q _3389_/Q _3629_/Q _2971_/S _3286_/S1 vssd1 vssd1 vccd1 vccd1
+ _3286_/X sky130_fd_sc_hd__mux4_2
X_2306_ _3584_/Q _2301_/X _2265_/X _2302_/X vssd1 vssd1 vccd1 vccd1 _3584_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2237_ _3623_/Q _2230_/A _2147_/X _2231_/A vssd1 vssd1 vccd1 vccd1 _3623_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2168_ _3672_/Q _2166_/X _2126_/X _2167_/X vssd1 vssd1 vccd1 vccd1 _3672_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2099_ _3705_/Q _2092_/X _2011_/X _2094_/X vssd1 vssd1 vccd1 vccd1 _3705_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3140_ _2711_/Y _2712_/Y _2713_/Y _2714_/Y _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3140_/X sky130_fd_sc_hd__mux4_2
X_3071_ _1695_/B _3233_/X _3858_/Q vssd1 vssd1 vccd1 vccd1 _3071_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2022_ _2030_/A vssd1 vssd1 vccd1 vccd1 _2022_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2924_ _3736_/Q vssd1 vssd1 vccd1 vccd1 _2924_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2855_ _3685_/Q vssd1 vssd1 vccd1 vccd1 _2855_/Y sky130_fd_sc_hd__inv_2
X_1806_ _3088_/X _1808_/B vssd1 vssd1 vccd1 vccd1 _3839_/D sky130_fd_sc_hd__nor2_1
X_2786_ _3561_/Q vssd1 vssd1 vccd1 vccd1 _2786_/Y sky130_fd_sc_hd__inv_2
X_1737_ _3887_/Q _1734_/X _2145_/A _1736_/X _1703_/X vssd1 vssd1 vccd1 vccd1 _3887_/D
+ sky130_fd_sc_hd__o221a_1
X_3407_ _3743_/CLK _3407_/D vssd1 vssd1 vccd1 vccd1 _3407_/Q sky130_fd_sc_hd__dfxtp_1
X_3338_ _3401_/Q _3393_/Q _3385_/Q _3625_/Q _3351_/S0 _3338_/S1 vssd1 vssd1 vccd1
+ vccd1 _3338_/X sky130_fd_sc_hd__mux4_2
X_3269_ _2624_/X _3026_/X _3027_/X _2626_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3269_/X sky130_fd_sc_hd__mux4_2
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2640_ _2654_/A _2640_/B vssd1 vssd1 vccd1 vccd1 _2640_/X sky130_fd_sc_hd__and2_1
XFILLER_9_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2571_ _3414_/Q _2563_/A _2550_/X _2564_/A vssd1 vssd1 vccd1 vccd1 _3414_/D sky130_fd_sc_hd__a22o_1
Xoutput306 _2679_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_6 sky130_fd_sc_hd__clkbuf_2
Xoutput317 _2945_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[1] sky130_fd_sc_hd__clkbuf_2
Xoutput339 _3868_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[20] sky130_fd_sc_hd__clkbuf_2
Xoutput328 _3852_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3123_ _3119_/X _3120_/X _3121_/X _3122_/X _3133_/S0 _3138_/X vssd1 vssd1 vccd1 vccd1
+ _3123_/X sky130_fd_sc_hd__mux4_2
X_3054_ _3353_/X _3354_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3054_/X sky130_fd_sc_hd__mux2_1
X_2005_ _3761_/Q _2002_/X _1966_/X _2004_/X vssd1 vssd1 vccd1 vccd1 _3761_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2907_ _3447_/Q vssd1 vssd1 vccd1 vccd1 _2907_/Y sky130_fd_sc_hd__inv_2
X_3887_ _3897_/CLK _3887_/D vssd1 vssd1 vccd1 vccd1 _3887_/Q sky130_fd_sc_hd__dfxtp_2
X_2838_ _3684_/Q vssd1 vssd1 vccd1 vccd1 _2838_/Y sky130_fd_sc_hd__inv_2
X_2769_ _3727_/Q vssd1 vssd1 vccd1 vccd1 _2769_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3810_ _3811_/CLK _3810_/D vssd1 vssd1 vccd1 vccd1 _3810_/Q sky130_fd_sc_hd__dfxtp_1
X_3741_ _3741_/CLK _3741_/D vssd1 vssd1 vccd1 vccd1 _3741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3672_ _3672_/CLK _3672_/D vssd1 vssd1 vccd1 vccd1 _3672_/Q sky130_fd_sc_hd__dfxtp_1
X_2623_ _2721_/A vssd1 vssd1 vccd1 vccd1 _2644_/A sky130_fd_sc_hd__buf_1
X_2554_ _2554_/A vssd1 vssd1 vccd1 vccd1 _2554_/X sky130_fd_sc_hd__clkbuf_2
X_2485_ _2492_/A vssd1 vssd1 vccd1 vccd1 _2485_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3106_ _2824_/Y _2825_/Y _2822_/Y _2823_/Y _3132_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3106_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3037_ _3300_/X _3036_/X _3061_/S vssd1 vssd1 vccd1 vccd1 _3037_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3672_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput16 io_b_dat_o_0[12] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
Xinput27 io_b_dat_o_0[8] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
Xinput38 io_b_dat_o_10[3] vssd1 vssd1 vccd1 vccd1 _2617_/B sky130_fd_sc_hd__clkbuf_1
Xinput49 io_b_dat_o_1[13] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2270_ _3606_/Q _2257_/A _2269_/X _2259_/A vssd1 vssd1 vccd1 vccd1 _3606_/D sky130_fd_sc_hd__a22o_1
XFILLER_77_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1985_ _1985_/A _2009_/B _2065_/A _2009_/D vssd1 vssd1 vccd1 vccd1 _2350_/A sky130_fd_sc_hd__or4_4
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3724_ _3724_/CLK _3724_/D vssd1 vssd1 vccd1 vccd1 _3724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3655_ _3687_/CLK _3655_/D vssd1 vssd1 vccd1 vccd1 _3655_/Q sky130_fd_sc_hd__dfxtp_1
X_2606_ _3387_/Q _2603_/X _2138_/A _2604_/X vssd1 vssd1 vccd1 vccd1 _3387_/D sky130_fd_sc_hd__a22o_1
X_3586_ _3586_/CLK _3586_/D vssd1 vssd1 vccd1 vccd1 _3586_/Q sky130_fd_sc_hd__dfxtp_1
X_2537_ _2950_/A vssd1 vssd1 vccd1 vccd1 _2537_/X sky130_fd_sc_hd__clkbuf_2
X_2468_ _2468_/A vssd1 vssd1 vccd1 vccd1 _2468_/X sky130_fd_sc_hd__clkbuf_2
X_2399_ _3526_/Q _2391_/A _2364_/X _2392_/A vssd1 vssd1 vccd1 vccd1 _3526_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1770_ _1774_/A _3009_/X vssd1 vssd1 vccd1 vccd1 _3869_/D sky130_fd_sc_hd__nor2b_4
XPHY_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3440_ _3811_/CLK _3440_/D vssd1 vssd1 vccd1 vccd1 _3440_/Q sky130_fd_sc_hd__dfxtp_1
X_3371_ _3582_/Q _3806_/Q _3534_/Q _3510_/Q _3372_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3371_/X sky130_fd_sc_hd__mux4_1
X_2322_ _2959_/A vssd1 vssd1 vccd1 vccd1 _2322_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater403 _3285_/S0 vssd1 vssd1 vccd1 vccd1 _2971_/S sky130_fd_sc_hd__clkbuf_8
X_2253_ _2951_/A vssd1 vssd1 vccd1 vccd1 _2253_/X sky130_fd_sc_hd__buf_2
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2184_ _2198_/A vssd1 vssd1 vccd1 vccd1 _2184_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1968_ _2574_/A vssd1 vssd1 vccd1 vccd1 _1968_/X sky130_fd_sc_hd__clkbuf_2
X_1899_ _2538_/A vssd1 vssd1 vccd1 vccd1 _1899_/X sky130_fd_sc_hd__clkbuf_2
X_3707_ _3831_/CLK _3707_/D vssd1 vssd1 vccd1 vccd1 _3707_/Q sky130_fd_sc_hd__dfxtp_1
X_3638_ _3687_/CLK _3638_/D vssd1 vssd1 vccd1 vccd1 _3638_/Q sky130_fd_sc_hd__dfxtp_1
X_3569_ _3722_/CLK _3569_/D vssd1 vssd1 vccd1 vccd1 _3569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput217 io_dat_i[5] vssd1 vssd1 vccd1 vccd1 _2949_/A sky130_fd_sc_hd__clkbuf_4
Xinput206 io_dat_i[24] vssd1 vssd1 vccd1 vccd1 input206/X sky130_fd_sc_hd__buf_1
Xinput228 io_dataLastBlock[15] vssd1 vssd1 vccd1 vccd1 _2964_/A0 sky130_fd_sc_hd__buf_1
Xinput239 io_dataLastBlock[25] vssd1 vssd1 vccd1 vccd1 _3005_/A0 sky130_fd_sc_hd__buf_1
XFILLER_84_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2940_ _3737_/Q vssd1 vssd1 vccd1 vccd1 _2940_/Y sky130_fd_sc_hd__inv_2
X_2871_ _3686_/Q vssd1 vssd1 vccd1 vccd1 _2871_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1822_ _2659_/A _1905_/B vssd1 vssd1 vccd1 vccd1 _2151_/A sky130_fd_sc_hd__or2_2
XPHY_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1753_ _3880_/Q _1734_/A _2133_/A _1736_/A _1721_/A vssd1 vssd1 vccd1 vccd1 _3880_/D
+ sky130_fd_sc_hd__o221a_1
X_1684_ _3897_/Q _3882_/Q _1679_/A _1683_/Y vssd1 vssd1 vccd1 vccd1 _1688_/A sky130_fd_sc_hd__o22a_1
XFILLER_89_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3423_ _3743_/CLK _3423_/D vssd1 vssd1 vccd1 vccd1 _3423_/Q sky130_fd_sc_hd__dfxtp_1
X_3354_ _3354_/A0 _3354_/A1 _3354_/A2 _3354_/A3 _2996_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3354_/X sky130_fd_sc_hd__mux4_1
X_3285_ _3437_/Q _3749_/Q _3421_/Q _3413_/Q _3285_/S0 _3286_/S1 vssd1 vssd1 vccd1
+ vccd1 _3285_/X sky130_fd_sc_hd__mux4_1
X_2305_ _3585_/Q _2301_/X _2263_/X _2302_/X vssd1 vssd1 vccd1 vccd1 _3585_/D sky130_fd_sc_hd__a22o_1
X_2236_ _3624_/Q _2230_/X _2145_/X _2231_/X vssd1 vssd1 vccd1 vccd1 _3624_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2167_ _2174_/A vssd1 vssd1 vccd1 vccd1 _2167_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2098_ _3706_/Q _2092_/X _1869_/X _2094_/X vssd1 vssd1 vccd1 vccd1 _3706_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3070_ _2641_/X _3228_/X _3858_/Q vssd1 vssd1 vccd1 vccd1 _3070_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2021_ input4/X _2021_/B _2021_/C _2021_/D vssd1 vssd1 vccd1 vccd1 _2030_/A sky130_fd_sc_hd__or4_4
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2923_ _3448_/Q vssd1 vssd1 vccd1 vccd1 _2923_/Y sky130_fd_sc_hd__inv_2
X_2854_ _3701_/Q vssd1 vssd1 vccd1 vccd1 _2854_/Y sky130_fd_sc_hd__inv_2
X_1805_ _3083_/X _1808_/B vssd1 vssd1 vccd1 vccd1 _3840_/D sky130_fd_sc_hd__nor2_1
X_2785_ _3728_/Q vssd1 vssd1 vccd1 vccd1 _2785_/Y sky130_fd_sc_hd__inv_2
X_1736_ _1736_/A vssd1 vssd1 vccd1 vccd1 _1736_/X sky130_fd_sc_hd__clkbuf_2
X_3406_ _3829_/CLK _3406_/D vssd1 vssd1 vccd1 vccd1 _3406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3337_ _3433_/Q _3745_/Q _3417_/Q _3409_/Q _3351_/S0 _3338_/S1 vssd1 vssd1 vccd1
+ vccd1 _3337_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3268_ _3268_/A0 _3268_/A1 _3268_/A2 _3268_/A3 _2984_/S _2981_/S vssd1 vssd1 vccd1
+ vccd1 _3268_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2219_ _3637_/Q _2214_/X _2133_/X _2215_/X vssd1 vssd1 vccd1 vccd1 _3637_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3199_ _3428_/Q _3604_/Q _3580_/Q _3556_/Q _3860_/Q _3232_/S1 vssd1 vssd1 vccd1 vccd1
+ _3199_/X sky130_fd_sc_hd__mux4_2
XFILLER_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2570_ _3415_/Q _2563_/A _2548_/X _2564_/A vssd1 vssd1 vccd1 vccd1 _3415_/D sky130_fd_sc_hd__a22o_1
Xoutput307 _2677_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_7 sky130_fd_sc_hd__clkbuf_2
Xoutput329 _3853_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[11] sky130_fd_sc_hd__clkbuf_2
Xoutput318 _2946_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3122_ _2772_/Y _2773_/Y _2770_/Y _2771_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3122_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3053_ _3352_/X _3052_/X _3053_/S vssd1 vssd1 vccd1 vccd1 _3053_/X sky130_fd_sc_hd__mux2_1
X_2004_ _2392_/A vssd1 vssd1 vccd1 vccd1 _2004_/X sky130_fd_sc_hd__buf_2
XFILLER_90_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2906_ _3471_/Q vssd1 vssd1 vccd1 vccd1 _2906_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3886_ _3895_/CLK _3886_/D vssd1 vssd1 vccd1 vccd1 _3886_/Q sky130_fd_sc_hd__dfxtp_1
X_2837_ _3700_/Q vssd1 vssd1 vccd1 vccd1 _2837_/Y sky130_fd_sc_hd__inv_2
X_2768_ _3439_/Q vssd1 vssd1 vccd1 vccd1 _2768_/Y sky130_fd_sc_hd__inv_2
X_1719_ _1721_/A _3064_/X _1723_/C vssd1 vssd1 vccd1 vccd1 _3895_/D sky130_fd_sc_hd__and3_1
X_2699_ _3779_/Q vssd1 vssd1 vccd1 vccd1 _2699_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3740_ _3740_/CLK _3740_/D vssd1 vssd1 vccd1 vccd1 _3740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3671_ _3687_/CLK _3671_/D vssd1 vssd1 vccd1 vccd1 _3671_/Q sky130_fd_sc_hd__dfxtp_1
X_2622_ _2638_/A _2991_/X vssd1 vssd1 vccd1 vccd1 _2622_/X sky130_fd_sc_hd__and2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2553_ _2553_/A vssd1 vssd1 vccd1 vccd1 _2553_/X sky130_fd_sc_hd__clkbuf_2
X_2484_ _3473_/Q _2477_/X _1966_/A _2479_/X vssd1 vssd1 vccd1 vccd1 _3473_/D sky130_fd_sc_hd__a22o_1
X_3105_ _2828_/Y _2829_/Y _2826_/Y _2827_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3105_/X sky130_fd_sc_hd__mux4_2
X_3036_ _3036_/A0 _3036_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3036_/X sky130_fd_sc_hd__mux2_2
XFILLER_70_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3869_ _3873_/CLK _3869_/D vssd1 vssd1 vccd1 vccd1 _3869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3867_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 io_b_dat_o_0[13] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_1
Xinput28 io_b_dat_o_0[9] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_1
Xinput39 io_b_dat_o_10[4] vssd1 vssd1 vccd1 vccd1 _2653_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1984_ _3770_/Q _1978_/X _1974_/X _1980_/X vssd1 vssd1 vccd1 vccd1 _3770_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3723_ _3723_/CLK _3723_/D vssd1 vssd1 vccd1 vccd1 _3723_/Q sky130_fd_sc_hd__dfxtp_1
X_3654_ _3687_/CLK _3654_/D vssd1 vssd1 vccd1 vccd1 _3654_/Q sky130_fd_sc_hd__dfxtp_1
X_2605_ _3388_/Q _2603_/X _2135_/A _2604_/X vssd1 vssd1 vccd1 vccd1 _3388_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
X_3585_ _3811_/CLK _3585_/D vssd1 vssd1 vccd1 vccd1 _3585_/Q sky130_fd_sc_hd__dfxtp_1
X_2536_ _2536_/A vssd1 vssd1 vccd1 vccd1 _2536_/X sky130_fd_sc_hd__clkbuf_2
X_2467_ _2467_/A vssd1 vssd1 vccd1 vccd1 _2467_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2398_ _3527_/Q _2391_/A _2362_/X _2392_/A vssd1 vssd1 vccd1 vccd1 _3527_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3019_ _3019_/A0 _3019_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3019_/X sky130_fd_sc_hd__mux2_2
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3370_ _3662_/Q _3646_/Q _3630_/Q _3606_/Q _3370_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3370_/X sky130_fd_sc_hd__mux4_2
X_2321_ _2340_/A vssd1 vssd1 vccd1 vccd1 _2321_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2252_ _3614_/Q _2248_/X _2131_/X _2249_/X vssd1 vssd1 vccd1 vccd1 _3614_/D sky130_fd_sc_hd__a22o_1
Xrepeater404 _3377_/S0 vssd1 vssd1 vccd1 vccd1 _3285_/S0 sky130_fd_sc_hd__buf_6
X_2183_ _2197_/A vssd1 vssd1 vccd1 vccd1 _2198_/A sky130_fd_sc_hd__inv_2
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1967_ _2573_/A vssd1 vssd1 vccd1 vccd1 _2574_/A sky130_fd_sc_hd__inv_2
X_3706_ _3831_/CLK _3706_/D vssd1 vssd1 vccd1 vccd1 _3706_/Q sky130_fd_sc_hd__dfxtp_1
X_1898_ _2536_/A vssd1 vssd1 vccd1 vccd1 _2538_/A sky130_fd_sc_hd__inv_2
X_3637_ _3841_/CLK _3637_/D vssd1 vssd1 vccd1 vccd1 _3637_/Q sky130_fd_sc_hd__dfxtp_1
X_3568_ _3720_/CLK _3568_/D vssd1 vssd1 vccd1 vccd1 _3568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2519_ _2526_/A vssd1 vssd1 vccd1 vccd1 _2519_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3499_ _3722_/CLK _3499_/D vssd1 vssd1 vccd1 vccd1 _3499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput218 io_dat_i[6] vssd1 vssd1 vccd1 vccd1 _2950_/A sky130_fd_sc_hd__clkbuf_4
Xinput207 io_dat_i[25] vssd1 vssd1 vccd1 vccd1 input207/X sky130_fd_sc_hd__buf_1
Xinput229 io_dataLastBlock[16] vssd1 vssd1 vccd1 vccd1 _3014_/A0 sky130_fd_sc_hd__buf_1
XFILLER_29_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3791_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2870_ _3702_/Q vssd1 vssd1 vccd1 vccd1 _2870_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1821_ _1928_/A vssd1 vssd1 vccd1 vccd1 _2659_/A sky130_fd_sc_hd__clkbuf_2
XPHY_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1752_ _2951_/A vssd1 vssd1 vccd1 vccd1 _2133_/A sky130_fd_sc_hd__buf_2
X_1683_ _3882_/Q vssd1 vssd1 vccd1 vccd1 _1683_/Y sky130_fd_sc_hd__inv_2
X_3422_ _3801_/CLK _3422_/D vssd1 vssd1 vccd1 vccd1 _3422_/Q sky130_fd_sc_hd__dfxtp_1
X_3353_ input21/X input53/X input69/X input85/X _2996_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3353_/X sky130_fd_sc_hd__mux4_1
X_3284_ _3533_/Q _3509_/Q _3485_/Q _3461_/Q _3285_/S0 _3286_/S1 vssd1 vssd1 vccd1
+ vccd1 _3284_/X sky130_fd_sc_hd__mux4_1
X_2304_ _3586_/Q _2301_/X _2261_/X _2302_/X vssd1 vssd1 vccd1 vccd1 _3586_/D sky130_fd_sc_hd__a22o_1
X_2235_ _3625_/Q _2230_/X _2143_/X _2231_/X vssd1 vssd1 vccd1 vccd1 _3625_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2166_ _2173_/A vssd1 vssd1 vccd1 vccd1 _2166_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2097_ _3707_/Q _2092_/X _1867_/X _2094_/X vssd1 vssd1 vccd1 vccd1 _3707_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2999_ _2999_/A0 _2999_/A1 _3009_/S vssd1 vssd1 vccd1 vccd1 _2999_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2020_ _3754_/Q _2010_/X _2019_/X _2013_/X vssd1 vssd1 vccd1 vccd1 _3754_/D sky130_fd_sc_hd__a22o_1
XFILLER_63_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2922_ _3472_/Q vssd1 vssd1 vccd1 vccd1 _2922_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2853_ _3717_/Q vssd1 vssd1 vccd1 vccd1 _2853_/Y sky130_fd_sc_hd__inv_2
X_1804_ _3078_/X _1808_/B vssd1 vssd1 vccd1 vccd1 _3841_/D sky130_fd_sc_hd__nor2_1
X_2784_ _3440_/Q vssd1 vssd1 vccd1 vccd1 _2784_/Y sky130_fd_sc_hd__inv_2
X_1735_ _2946_/A vssd1 vssd1 vccd1 vccd1 _2145_/A sky130_fd_sc_hd__clkbuf_2
X_3405_ _3796_/CLK _3405_/D vssd1 vssd1 vccd1 vccd1 _3405_/Q sky130_fd_sc_hd__dfxtp_1
X_3336_ _3529_/Q _3505_/Q _3481_/Q _3457_/Q _3351_/S0 _3351_/S1 vssd1 vssd1 vccd1
+ vccd1 _3336_/X sky130_fd_sc_hd__mux4_2
X_3267_ input28/X input60/X input76/X input92/X _2984_/S _2981_/S vssd1 vssd1 vccd1
+ vccd1 _3267_/X sky130_fd_sc_hd__mux4_1
X_3198_ _3194_/X _3195_/X _3196_/X _3197_/X _3862_/Q _3863_/Q vssd1 vssd1 vccd1 vccd1
+ _3198_/X sky130_fd_sc_hd__mux4_2
X_2218_ _3638_/Q _2214_/X _2131_/X _2215_/X vssd1 vssd1 vccd1 vccd1 _3638_/D sky130_fd_sc_hd__a22o_1
X_2149_ _2149_/A vssd1 vssd1 vccd1 vccd1 _2149_/X sky130_fd_sc_hd__buf_2
XFILLER_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput308 _2676_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_8 sky130_fd_sc_hd__clkbuf_2
Xoutput319 _2947_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[3] sky130_fd_sc_hd__clkbuf_2
X_3121_ _2776_/Y _2777_/Y _2774_/Y _2775_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3121_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3052_ _3052_/A0 _3052_/A1 _3060_/S vssd1 vssd1 vccd1 vccd1 _3052_/X sky130_fd_sc_hd__mux2_4
XFILLER_82_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2003_ _2391_/A vssd1 vssd1 vccd1 vccd1 _2392_/A sky130_fd_sc_hd__inv_2
XFILLER_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3885_ _3895_/CLK _3885_/D vssd1 vssd1 vccd1 vccd1 _3885_/Q sky130_fd_sc_hd__dfxtp_1
X_2905_ _3495_/Q vssd1 vssd1 vccd1 vccd1 _2905_/Y sky130_fd_sc_hd__inv_2
X_2836_ _2836_/A _2836_/B vssd1 vssd1 vccd1 vccd1 _2836_/X sky130_fd_sc_hd__and2_1
X_2767_ _3463_/Q vssd1 vssd1 vccd1 vccd1 _2767_/Y sky130_fd_sc_hd__inv_2
X_1718_ _1727_/C vssd1 vssd1 vccd1 vccd1 _1723_/C sky130_fd_sc_hd__buf_1
X_2698_ _3751_/Q vssd1 vssd1 vccd1 vccd1 _2698_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3319_ _3586_/Q _3810_/Q _3538_/Q _3514_/Q _1905_/A _3357_/S1 vssd1 vssd1 vccd1 vccd1
+ _3319_/X sky130_fd_sc_hd__mux4_2
XFILLER_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3670_ _3687_/CLK _3670_/D vssd1 vssd1 vccd1 vccd1 _3670_/Q sky130_fd_sc_hd__dfxtp_1
X_2621_ _2647_/A vssd1 vssd1 vccd1 vccd1 _2638_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2552_ _3429_/Q _1907_/X _2534_/X _1909_/X vssd1 vssd1 vccd1 vccd1 _3429_/D sky130_fd_sc_hd__a22o_1
X_2483_ _3474_/Q _2477_/X _2330_/X _2479_/X vssd1 vssd1 vccd1 vccd1 _3474_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3104_ _2832_/Y _2833_/Y _2830_/Y _2831_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3104_/X sky130_fd_sc_hd__mux4_2
X_3035_ _3884_/Q _3295_/X _3061_/S vssd1 vssd1 vccd1 vccd1 _3035_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3868_ _3873_/CLK _3868_/D vssd1 vssd1 vccd1 vccd1 _3868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2819_ _3715_/Q vssd1 vssd1 vccd1 vccd1 _2819_/Y sky130_fd_sc_hd__inv_2
X_3799_ _3799_/CLK _3799_/D vssd1 vssd1 vccd1 vccd1 _3799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_55_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3724_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 io_b_dat_o_0[14] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_1
Xinput29 io_b_dat_o_10[0] vssd1 vssd1 vccd1 vccd1 _2724_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1983_ _3771_/Q _1978_/X _1972_/X _1980_/X vssd1 vssd1 vccd1 vccd1 _3771_/D sky130_fd_sc_hd__a22o_1
X_3722_ _3722_/CLK _3722_/D vssd1 vssd1 vccd1 vccd1 _3722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3653_ _3672_/CLK _3653_/D vssd1 vssd1 vccd1 vccd1 _3653_/Q sky130_fd_sc_hd__dfxtp_1
X_2604_ _2604_/A vssd1 vssd1 vccd1 vccd1 _2604_/X sky130_fd_sc_hd__clkbuf_2
X_3584_ _3586_/CLK _3584_/D vssd1 vssd1 vccd1 vccd1 _3584_/Q sky130_fd_sc_hd__dfxtp_1
X_2535_ _3437_/Q _1897_/X _2534_/X _1899_/X vssd1 vssd1 vccd1 vccd1 _3437_/D sky130_fd_sc_hd__a22o_1
X_2466_ _3485_/Q _1827_/X _2448_/X _1831_/X vssd1 vssd1 vccd1 vccd1 _3485_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2397_ _3528_/Q _2391_/X _2360_/X _2392_/X vssd1 vssd1 vccd1 vccd1 _3528_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3018_ _3243_/X _3244_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3018_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2320_ _2476_/A _2320_/B _2675_/A _2476_/D vssd1 vssd1 vccd1 vccd1 _2340_/A sky130_fd_sc_hd__or4_4
X_2251_ _3615_/Q _2248_/X _2129_/X _2249_/X vssd1 vssd1 vccd1 vccd1 _3615_/D sky130_fd_sc_hd__a22o_1
Xrepeater405 _3291_/S0 vssd1 vssd1 vccd1 vccd1 _3377_/S0 sky130_fd_sc_hd__buf_6
X_2182_ _2197_/A vssd1 vssd1 vccd1 vccd1 _2182_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3682_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1966_ _1966_/A vssd1 vssd1 vccd1 vccd1 _1966_/X sky130_fd_sc_hd__clkbuf_2
X_3705_ _3741_/CLK _3705_/D vssd1 vssd1 vccd1 vccd1 _3705_/Q sky130_fd_sc_hd__dfxtp_1
X_1897_ _2536_/A vssd1 vssd1 vccd1 vccd1 _1897_/X sky130_fd_sc_hd__clkbuf_2
X_3636_ _3672_/CLK _3636_/D vssd1 vssd1 vccd1 vccd1 _3636_/Q sky130_fd_sc_hd__dfxtp_1
X_3567_ _3719_/CLK _3567_/D vssd1 vssd1 vccd1 vccd1 _3567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2518_ _3449_/Q _2511_/X _1966_/A _2513_/X vssd1 vssd1 vccd1 vccd1 _3449_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3498_ _3832_/CLK _3498_/D vssd1 vssd1 vccd1 vccd1 _3498_/Q sky130_fd_sc_hd__dfxtp_1
Xinput208 io_dat_i[26] vssd1 vssd1 vccd1 vccd1 input208/X sky130_fd_sc_hd__buf_1
Xinput219 io_dat_i[7] vssd1 vssd1 vccd1 vccd1 _2951_/A sky130_fd_sc_hd__buf_4
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2449_ _3493_/Q _2443_/X _2448_/X _2444_/X vssd1 vssd1 vccd1 vccd1 _3493_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1820_ _1905_/A vssd1 vssd1 vccd1 vccd1 _1928_/A sky130_fd_sc_hd__inv_2
XPHY_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1751_ _3881_/Q _1734_/A _2143_/A _1736_/A _1742_/X vssd1 vssd1 vccd1 vccd1 _3881_/D
+ sky130_fd_sc_hd__o221a_1
X_1682_ _3899_/Q vssd1 vssd1 vccd1 vccd1 _1682_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3421_ _3829_/CLK _3421_/D vssd1 vssd1 vccd1 vccd1 _3421_/Q sky130_fd_sc_hd__dfxtp_1
X_3352_ _3348_/X _3349_/X _3350_/X _3351_/X _3373_/S0 _3378_/S1 vssd1 vssd1 vccd1
+ vccd1 _3352_/X sky130_fd_sc_hd__mux4_1
X_2303_ _3587_/Q _2301_/X _2258_/X _2302_/X vssd1 vssd1 vccd1 vccd1 _3587_/D sky130_fd_sc_hd__a22o_1
X_3283_ _3429_/Q _3605_/Q _3581_/Q _3557_/Q _3285_/S0 _3286_/S1 vssd1 vssd1 vccd1
+ vccd1 _3283_/X sky130_fd_sc_hd__mux4_2
X_2234_ _3626_/Q _2230_/X _2141_/X _2231_/X vssd1 vssd1 vccd1 vccd1 _3626_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2165_ _3673_/Q _2154_/X _2123_/X _2157_/X vssd1 vssd1 vccd1 vccd1 _3673_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2096_ _3708_/Q _2092_/X _1865_/X _2094_/X vssd1 vssd1 vccd1 vccd1 _3708_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2998_ _1705_/X _3897_/Q _3073_/S vssd1 vssd1 vccd1 vccd1 _2998_/X sky130_fd_sc_hd__mux2_1
X_1949_ _2593_/A vssd1 vssd1 vccd1 vccd1 _1949_/X sky130_fd_sc_hd__clkbuf_2
X_3619_ _3676_/CLK _3619_/D vssd1 vssd1 vccd1 vccd1 _3619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2921_ _3496_/Q vssd1 vssd1 vccd1 vccd1 _2921_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2852_ _3565_/Q vssd1 vssd1 vccd1 vccd1 _2852_/Y sky130_fd_sc_hd__inv_2
X_1803_ _1816_/B vssd1 vssd1 vccd1 vccd1 _1808_/B sky130_fd_sc_hd__clkbuf_2
X_2783_ _3464_/Q vssd1 vssd1 vccd1 vccd1 _2783_/Y sky130_fd_sc_hd__inv_2
X_1734_ _1734_/A vssd1 vssd1 vccd1 vccd1 _1734_/X sky130_fd_sc_hd__clkbuf_2
X_3404_ _3627_/CLK _3404_/D vssd1 vssd1 vccd1 vccd1 _3404_/Q sky130_fd_sc_hd__dfxtp_1
X_3335_ _3425_/Q _3601_/Q _3577_/Q _3553_/Q _3351_/S0 _3338_/S1 vssd1 vssd1 vccd1
+ vccd1 _3335_/X sky130_fd_sc_hd__mux4_1
X_3266_ _3262_/X _3263_/X _3264_/X _3265_/X _2613_/A _3378_/S1 vssd1 vssd1 vccd1 vccd1
+ _3266_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2217_ _3639_/Q _2214_/X _2129_/X _2215_/X vssd1 vssd1 vccd1 vccd1 _3639_/D sky130_fd_sc_hd__a22o_1
X_3197_ _3405_/Q _3397_/Q _3389_/Q _3629_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3197_/X sky130_fd_sc_hd__mux4_2
XFILLER_93_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2148_ _3679_/Q _2137_/X _2147_/X _2139_/X vssd1 vssd1 vccd1 vccd1 _3679_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2079_ _3718_/Q _2075_/X _2019_/X _2076_/X vssd1 vssd1 vccd1 vccd1 _3718_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput309 _2674_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_9 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3120_ _2780_/Y _2781_/Y _2778_/Y _2779_/Y _3126_/S0 _3126_/S1 vssd1 vssd1 vccd1
+ vccd1 _3120_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3051_ _3887_/Q _3347_/X _3053_/S vssd1 vssd1 vccd1 vccd1 _3051_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2002_ _2391_/A vssd1 vssd1 vccd1 vccd1 _2002_/X sky130_fd_sc_hd__buf_2
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3884_ _3897_/CLK _3884_/D vssd1 vssd1 vccd1 vccd1 _3884_/Q sky130_fd_sc_hd__dfxtp_1
X_2904_ _3519_/Q vssd1 vssd1 vccd1 vccd1 _2904_/Y sky130_fd_sc_hd__inv_2
X_2835_ _3716_/Q vssd1 vssd1 vccd1 vccd1 _2835_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2766_ _3487_/Q vssd1 vssd1 vccd1 vccd1 _2766_/Y sky130_fd_sc_hd__inv_2
X_1717_ _3895_/Q _1717_/B vssd1 vssd1 vccd1 vccd1 _1727_/C sky130_fd_sc_hd__or2_2
X_2697_ _3803_/Q vssd1 vssd1 vccd1 vccd1 _2697_/Y sky130_fd_sc_hd__inv_2
X_3318_ _3666_/Q _3650_/Q _3634_/Q _3610_/Q input5/X input6/X vssd1 vssd1 vccd1 vccd1
+ _3318_/X sky130_fd_sc_hd__mux4_2
XFILLER_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3249_ _3789_/Q _3785_/Q _3793_/Q _3765_/Q _3285_/S0 _3286_/S1 vssd1 vssd1 vccd1
+ vccd1 _3249_/X sky130_fd_sc_hd__mux4_2
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2620_ _2681_/A _2981_/X vssd1 vssd1 vccd1 vccd1 _2620_/X sky130_fd_sc_hd__and2_1
XFILLER_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2551_ _3430_/Q _2536_/A _2550_/X _2538_/A vssd1 vssd1 vccd1 vccd1 _3430_/D sky130_fd_sc_hd__a22o_1
X_2482_ _3475_/Q _2477_/X _2328_/X _2479_/X vssd1 vssd1 vccd1 vccd1 _3475_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3103_ _3099_/X _3100_/X _3101_/X _3102_/X _3133_/S0 _3138_/X vssd1 vssd1 vccd1 vccd1
+ _3103_/X sky130_fd_sc_hd__mux4_2
X_3034_ _3288_/X _3289_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3034_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3867_ _3867_/CLK _3867_/D vssd1 vssd1 vccd1 vccd1 _3867_/Q sky130_fd_sc_hd__dfxtp_1
X_3798_ _3823_/CLK _3798_/D vssd1 vssd1 vccd1 vccd1 _3798_/Q sky130_fd_sc_hd__dfxtp_1
X_2818_ _3563_/Q vssd1 vssd1 vccd1 vccd1 _2818_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2749_ _3510_/Q vssd1 vssd1 vccd1 vccd1 _2749_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_24_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3743_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput19 io_b_dat_o_0[15] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1982_ _3772_/Q _1978_/X _1970_/X _1980_/X vssd1 vssd1 vccd1 vccd1 _3772_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3721_ _3722_/CLK _3721_/D vssd1 vssd1 vccd1 vccd1 _3721_/Q sky130_fd_sc_hd__dfxtp_1
X_3652_ _3832_/CLK _3652_/D vssd1 vssd1 vccd1 vccd1 _3652_/Q sky130_fd_sc_hd__dfxtp_1
X_2603_ _2603_/A vssd1 vssd1 vccd1 vccd1 _2603_/X sky130_fd_sc_hd__clkbuf_2
X_3583_ _3726_/CLK _3583_/D vssd1 vssd1 vccd1 vccd1 _3583_/Q sky130_fd_sc_hd__dfxtp_1
X_2534_ _2951_/A vssd1 vssd1 vccd1 vccd1 _2534_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2465_ _3486_/Q _2452_/A _2464_/X _2454_/A vssd1 vssd1 vccd1 vccd1 _3486_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2396_ _3529_/Q _2391_/X _2358_/X _2392_/X vssd1 vssd1 vccd1 vccd1 _3529_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3017_ _3240_/X _3241_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3017_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2250_ _3616_/Q _2248_/X _2126_/X _2249_/X vssd1 vssd1 vccd1 vccd1 _3616_/D sky130_fd_sc_hd__a22o_1
Xrepeater406 _3372_/S0 vssd1 vssd1 vccd1 vccd1 _3291_/S0 sky130_fd_sc_hd__buf_4
XFILLER_93_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2181_ _2281_/A _2181_/B _2673_/A _2281_/D vssd1 vssd1 vccd1 vccd1 _2197_/A sky130_fd_sc_hd__or4_4
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1965_ _2573_/A vssd1 vssd1 vccd1 vccd1 _1965_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3704_ _3720_/CLK _3704_/D vssd1 vssd1 vccd1 vccd1 _3704_/Q sky130_fd_sc_hd__dfxtp_1
X_1896_ _2476_/A _2510_/B _2021_/C _1915_/D vssd1 vssd1 vccd1 vccd1 _2536_/A sky130_fd_sc_hd__or4_4
X_3635_ _3667_/CLK _3635_/D vssd1 vssd1 vccd1 vccd1 _3635_/Q sky130_fd_sc_hd__dfxtp_1
X_3566_ _3719_/CLK _3566_/D vssd1 vssd1 vccd1 vccd1 _3566_/Q sky130_fd_sc_hd__dfxtp_1
X_2517_ _3450_/Q _2511_/X _2956_/A _2513_/X vssd1 vssd1 vccd1 vccd1 _3450_/D sky130_fd_sc_hd__a22o_1
X_3497_ _3740_/CLK _3497_/D vssd1 vssd1 vccd1 vccd1 _3497_/Q sky130_fd_sc_hd__dfxtp_1
X_2448_ _2951_/A vssd1 vssd1 vccd1 vccd1 _2448_/X sky130_fd_sc_hd__clkbuf_2
Xinput209 io_dat_i[27] vssd1 vssd1 vccd1 vccd1 input209/X sky130_fd_sc_hd__buf_1
XFILLER_68_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2379_ _3542_/Q _2375_/X _2297_/X _2376_/X vssd1 vssd1 vccd1 vccd1 _3542_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1750_ _2947_/A vssd1 vssd1 vccd1 vccd1 _2143_/A sky130_fd_sc_hd__clkbuf_2
X_1681_ _1681_/A vssd1 vssd1 vccd1 vccd1 _1681_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3420_ _3627_/CLK _3420_/D vssd1 vssd1 vccd1 vccd1 _3420_/Q sky130_fd_sc_hd__dfxtp_1
X_3351_ _3400_/Q _3392_/Q _3384_/Q _3624_/Q _3351_/S0 _3351_/S1 vssd1 vssd1 vccd1
+ vccd1 _3351_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2302_ _2302_/A vssd1 vssd1 vccd1 vccd1 _2302_/X sky130_fd_sc_hd__clkbuf_2
X_3282_ _3278_/X _3279_/X _3280_/X _3281_/X _3295_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3282_/X sky130_fd_sc_hd__mux4_2
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2233_ _3627_/Q _2230_/X _2138_/X _2231_/X vssd1 vssd1 vccd1 vccd1 _3627_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2164_ _3674_/Q _2154_/X _2163_/X _2157_/X vssd1 vssd1 vccd1 vccd1 _3674_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2095_ _3709_/Q _2092_/X _1861_/X _2094_/X vssd1 vssd1 vccd1 vccd1 _3709_/D sky130_fd_sc_hd__a22o_1
XFILLER_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2997_ _2996_/X _2724_/X _2997_/S vssd1 vssd1 vccd1 vccd1 _2997_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1948_ _2009_/A _2009_/B _2510_/C _1964_/D vssd1 vssd1 vccd1 vccd1 _2593_/A sky130_fd_sc_hd__or4_4
X_1879_ _2135_/A vssd1 vssd1 vccd1 vccd1 _1879_/X sky130_fd_sc_hd__buf_2
X_3618_ _3676_/CLK _3618_/D vssd1 vssd1 vccd1 vccd1 _3618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3549_ _3700_/CLK _3549_/D vssd1 vssd1 vccd1 vccd1 _3549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2920_ _3520_/Q vssd1 vssd1 vccd1 vccd1 _2920_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2851_ _3732_/Q vssd1 vssd1 vccd1 vccd1 _2851_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2782_ _3488_/Q vssd1 vssd1 vccd1 vccd1 _2782_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1802_ _1802_/A _1802_/B vssd1 vssd1 vccd1 vccd1 _1816_/B sky130_fd_sc_hd__or2_4
XPHY_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1733_ _1736_/A vssd1 vssd1 vccd1 vccd1 _1734_/A sky130_fd_sc_hd__inv_2
X_3403_ _3897_/CLK _3403_/D vssd1 vssd1 vccd1 vccd1 _3403_/Q sky130_fd_sc_hd__dfxtp_1
X_3334_ _3330_/X _3331_/X _3332_/X _3333_/X _3373_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3334_/X sky130_fd_sc_hd__mux4_2
XFILLER_58_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3265_ _3787_/Q _3783_/Q _3791_/Q _3763_/Q _3009_/S _3286_/S1 vssd1 vssd1 vccd1 vccd1
+ _3265_/X sky130_fd_sc_hd__mux4_2
X_2216_ _3640_/Q _2214_/X _2126_/X _2215_/X vssd1 vssd1 vccd1 vccd1 _3640_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3196_ _3437_/Q _3749_/Q _3421_/Q _3413_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3196_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2147_ _2147_/A vssd1 vssd1 vccd1 vccd1 _2147_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_53_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2078_ _3719_/Q _2075_/X _2017_/X _2076_/X vssd1 vssd1 vccd1 vccd1 _3719_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_49_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3722_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3050_ _3340_/X _3341_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3050_/X sky130_fd_sc_hd__mux2_1
X_2001_ _2009_/A input1/X _2151_/A _2009_/D vssd1 vssd1 vccd1 vccd1 _2391_/A sky130_fd_sc_hd__or4_4
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3883_ _3897_/CLK _3883_/D vssd1 vssd1 vccd1 vccd1 _3883_/Q sky130_fd_sc_hd__dfxtp_1
X_2903_ _3543_/Q vssd1 vssd1 vccd1 vccd1 _2903_/Y sky130_fd_sc_hd__inv_2
X_2834_ _3564_/Q vssd1 vssd1 vccd1 vccd1 _2834_/Y sky130_fd_sc_hd__inv_2
X_2765_ _3511_/Q vssd1 vssd1 vccd1 vccd1 _2765_/Y sky130_fd_sc_hd__inv_2
X_1716_ _3894_/Q _1716_/B vssd1 vssd1 vccd1 vccd1 _1717_/B sky130_fd_sc_hd__or2_1
X_2696_ _3823_/Q vssd1 vssd1 vccd1 vccd1 _2696_/Y sky130_fd_sc_hd__inv_2
X_3317_ _3562_/Q _3714_/Q _3698_/Q _3682_/Q input5/X _3357_/S1 vssd1 vssd1 vccd1 vccd1
+ _3317_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3248_ _3805_/Q _3753_/Q _3781_/Q _3777_/Q _3377_/S0 _3286_/S1 vssd1 vssd1 vccd1
+ vccd1 _3248_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3179_ _3568_/Q _3720_/Q _3704_/Q _3688_/Q _3291_/S0 _3192_/S1 vssd1 vssd1 vccd1
+ vccd1 _3179_/X sky130_fd_sc_hd__mux4_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2550_ _2944_/A vssd1 vssd1 vccd1 vccd1 _2550_/X sky130_fd_sc_hd__clkbuf_2
X_2481_ _3476_/Q _2477_/X _2326_/X _2479_/X vssd1 vssd1 vccd1 vccd1 _3476_/D sky130_fd_sc_hd__a22o_1
X_3102_ _2837_/Y _2838_/Y _2834_/Y _2835_/Y _3102_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3102_/X sky130_fd_sc_hd__mux4_1
X_3033_ _3287_/X _3032_/X _3061_/S vssd1 vssd1 vccd1 vccd1 _3033_/X sky130_fd_sc_hd__mux2_2
XFILLER_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3866_ _3867_/CLK _3866_/D vssd1 vssd1 vccd1 vccd1 _3866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3797_ _3890_/CLK _3797_/D vssd1 vssd1 vccd1 vccd1 _3797_/Q sky130_fd_sc_hd__dfxtp_1
X_2817_ _3730_/Q vssd1 vssd1 vccd1 vccd1 _2817_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2748_ _3534_/Q vssd1 vssd1 vccd1 vccd1 _2748_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2679_ _2681_/A _2684_/B _2683_/C vssd1 vssd1 vccd1 vccd1 _2679_/Y sky130_fd_sc_hd__nor3_2
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3720_ _3720_/CLK _3720_/D vssd1 vssd1 vccd1 vccd1 _3720_/Q sky130_fd_sc_hd__dfxtp_1
X_1981_ _3773_/Q _1978_/X _1966_/X _1980_/X vssd1 vssd1 vccd1 vccd1 _3773_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3651_ _3667_/CLK _3651_/D vssd1 vssd1 vccd1 vccd1 _3651_/Q sky130_fd_sc_hd__dfxtp_1
X_2602_ _3389_/Q _1932_/X _2133_/A _1934_/X vssd1 vssd1 vccd1 vccd1 _3389_/D sky130_fd_sc_hd__a22o_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3582_ _3821_/CLK _3582_/D vssd1 vssd1 vccd1 vccd1 _3582_/Q sky130_fd_sc_hd__dfxtp_1
X_2533_ _3438_/Q _2526_/A _2464_/X _2527_/A vssd1 vssd1 vccd1 vccd1 _3438_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2464_ _2944_/A vssd1 vssd1 vccd1 vccd1 _2464_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2395_ _3530_/Q _2391_/X _2356_/X _2392_/X vssd1 vssd1 vccd1 vccd1 _3530_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3016_ _3237_/X _3238_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3016_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3849_ _3851_/CLK _3849_/D vssd1 vssd1 vccd1 vccd1 _3849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE4_0 _3873_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2180_ _3662_/Q _2173_/A _2149_/X _2174_/A vssd1 vssd1 vccd1 vccd1 _3662_/D sky130_fd_sc_hd__a22o_1
Xrepeater407 _3372_/S0 vssd1 vssd1 vccd1 vccd1 _3370_/S0 sky130_fd_sc_hd__buf_8
XFILLER_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1964_ _1985_/A _2009_/B _2021_/C _1964_/D vssd1 vssd1 vccd1 vccd1 _2573_/A sky130_fd_sc_hd__or4_4
X_3703_ _3719_/CLK _3703_/D vssd1 vssd1 vccd1 vccd1 _3703_/Q sky130_fd_sc_hd__dfxtp_1
X_3634_ _3859_/CLK _3634_/D vssd1 vssd1 vccd1 vccd1 _3634_/Q sky130_fd_sc_hd__dfxtp_1
X_1895_ input4/X vssd1 vssd1 vccd1 vccd1 _2476_/A sky130_fd_sc_hd__clkbuf_2
X_3565_ _3813_/CLK _3565_/D vssd1 vssd1 vccd1 vccd1 _3565_/Q sky130_fd_sc_hd__dfxtp_1
X_2516_ _3451_/Q _2511_/X _2957_/A _2513_/X vssd1 vssd1 vccd1 vccd1 _3451_/D sky130_fd_sc_hd__a22o_1
X_3496_ _3816_/CLK _3496_/D vssd1 vssd1 vccd1 vccd1 _3496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2447_ _3494_/Q _2443_/X _2297_/X _2444_/X vssd1 vssd1 vccd1 vccd1 _3494_/D sky130_fd_sc_hd__a22o_1
X_2378_ _3543_/Q _2375_/X _2295_/X _2376_/X vssd1 vssd1 vccd1 vccd1 _3543_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1680_ _3898_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1681_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3350_ _3432_/Q _3744_/Q _3416_/Q _3408_/Q _3351_/S0 _3351_/S1 vssd1 vssd1 vccd1
+ vccd1 _3350_/X sky130_fd_sc_hd__mux4_1
X_2301_ _2301_/A vssd1 vssd1 vccd1 vccd1 _2301_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3281_ _3493_/Q _3469_/Q _3445_/Q _3733_/Q _3291_/S0 _3294_/S1 vssd1 vssd1 vccd1
+ vccd1 _3281_/X sky130_fd_sc_hd__mux4_1
X_2232_ _3628_/Q _2230_/X _2135_/X _2231_/X vssd1 vssd1 vccd1 vccd1 _3628_/D sky130_fd_sc_hd__a22o_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2163_ _2956_/A vssd1 vssd1 vccd1 vccd1 _2163_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2094_ _2108_/A vssd1 vssd1 vccd1 vccd1 _2094_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2996_ _2996_/A0 _2996_/A1 _2996_/S vssd1 vssd1 vccd1 vccd1 _2996_/X sky130_fd_sc_hd__mux2_1
X_1947_ _2021_/B vssd1 vssd1 vccd1 vccd1 _2009_/B sky130_fd_sc_hd__buf_1
X_1878_ _3813_/Q _1872_/X _1877_/X _1873_/X vssd1 vssd1 vccd1 vccd1 _3813_/D sky130_fd_sc_hd__a22o_1
X_3617_ _3662_/CLK _3617_/D vssd1 vssd1 vccd1 vccd1 _3617_/Q sky130_fd_sc_hd__dfxtp_1
X_3548_ _3832_/CLK _3548_/D vssd1 vssd1 vccd1 vccd1 _3548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3479_ _3801_/CLK _3479_/D vssd1 vssd1 vccd1 vccd1 _3479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2850_ _3444_/Q vssd1 vssd1 vccd1 vccd1 _2850_/Y sky130_fd_sc_hd__inv_2
X_1801_ _1801_/A _3381_/X vssd1 vssd1 vccd1 vccd1 _3842_/D sky130_fd_sc_hd__and2_1
XFILLER_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2781_ _3512_/Q vssd1 vssd1 vccd1 vccd1 _2781_/Y sky130_fd_sc_hd__inv_2
XPHY_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1732_ _2721_/A input3/X _2961_/S _1857_/D vssd1 vssd1 vccd1 vccd1 _1736_/A sky130_fd_sc_hd__or4_4
X_3402_ _3867_/CLK _3402_/D vssd1 vssd1 vccd1 vccd1 _3402_/Q sky130_fd_sc_hd__dfxtp_1
X_3333_ _3489_/Q _3465_/Q _3441_/Q _3729_/Q input5/X _3357_/S1 vssd1 vssd1 vccd1 vccd1
+ _3333_/X sky130_fd_sc_hd__mux4_2
X_3264_ _3803_/Q _3751_/Q _3779_/Q _3775_/Q _3036_/S _3294_/S1 vssd1 vssd1 vccd1 vccd1
+ _3264_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2215_ _2222_/A vssd1 vssd1 vccd1 vccd1 _2215_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3195_ _3533_/Q _3509_/Q _3485_/Q _3461_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3195_/X sky130_fd_sc_hd__mux4_2
XFILLER_38_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2146_ _3680_/Q _2137_/X _2145_/X _2139_/X vssd1 vssd1 vccd1 vccd1 _3680_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2077_ _3720_/Q _2075_/X _2015_/X _2076_/X vssd1 vssd1 vccd1 vccd1 _3720_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2979_ _2978_/X _2625_/X _2981_/S vssd1 vssd1 vccd1 vccd1 _2979_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_18_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3896_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2000_ _3762_/Q _1994_/X _1974_/X _1996_/X vssd1 vssd1 vccd1 vccd1 _3762_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2902_ _3815_/Q vssd1 vssd1 vccd1 vccd1 _2902_/Y sky130_fd_sc_hd__inv_2
X_3882_ _3896_/CLK _3882_/D vssd1 vssd1 vccd1 vccd1 _3882_/Q sky130_fd_sc_hd__dfxtp_1
X_2833_ _3731_/Q vssd1 vssd1 vccd1 vccd1 _2833_/Y sky130_fd_sc_hd__inv_2
X_2764_ _3535_/Q vssd1 vssd1 vccd1 vccd1 _2764_/Y sky130_fd_sc_hd__inv_2
X_1715_ _1715_/A _1715_/B vssd1 vssd1 vccd1 vccd1 _1716_/B sky130_fd_sc_hd__nand2_1
X_2695_ _3827_/Q vssd1 vssd1 vccd1 vccd1 _2695_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3316_ _3039_/X _3041_/X _3042_/X _2615_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3316_/X sky130_fd_sc_hd__mux4_2
X_3247_ _3761_/Q _3797_/Q _3829_/Q _3825_/Q _3285_/S0 _3286_/S1 vssd1 vssd1 vccd1
+ vccd1 _3247_/X sky130_fd_sc_hd__mux4_1
X_3178_ _3174_/X _3175_/X _3176_/X _3177_/X _3295_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3178_/X sky130_fd_sc_hd__mux4_2
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2129_ _2953_/A vssd1 vssd1 vccd1 vccd1 _2129_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2480_ _3477_/Q _2477_/X _2322_/X _2479_/X vssd1 vssd1 vccd1 vccd1 _3477_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3101_ _2841_/Y _2842_/Y _2839_/Y _2840_/Y _3132_/S0 _3132_/S1 vssd1 vssd1 vccd1
+ vccd1 _3101_/X sky130_fd_sc_hd__mux4_2
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput190 io_dat_i[0] vssd1 vssd1 vccd1 vccd1 _2944_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3032_ _3032_/A0 _3032_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3032_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3865_ _3867_/CLK _3865_/D vssd1 vssd1 vccd1 vccd1 _3865_/Q sky130_fd_sc_hd__dfxtp_1
X_2816_ _3442_/Q vssd1 vssd1 vccd1 vccd1 _2816_/Y sky130_fd_sc_hd__inv_2
X_3796_ _3796_/CLK _3796_/D vssd1 vssd1 vccd1 vccd1 _3796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2747_ _3806_/Q vssd1 vssd1 vccd1 vccd1 _2747_/Y sky130_fd_sc_hd__inv_2
X_2678_ input8/X vssd1 vssd1 vccd1 vccd1 _2684_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3799_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1980_ _2311_/A vssd1 vssd1 vccd1 vccd1 _1980_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3650_ _3859_/CLK _3650_/D vssd1 vssd1 vccd1 vccd1 _3650_/Q sky130_fd_sc_hd__dfxtp_1
X_2601_ _3390_/Q _2593_/A _2149_/A _2594_/A vssd1 vssd1 vccd1 vccd1 _3390_/D sky130_fd_sc_hd__a22o_1
X_3581_ _3823_/CLK _3581_/D vssd1 vssd1 vccd1 vccd1 _3581_/Q sky130_fd_sc_hd__dfxtp_1
X_2532_ _3439_/Q _2526_/X _2462_/X _2527_/X vssd1 vssd1 vccd1 vccd1 _3439_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2463_ _3487_/Q _2452_/X _2462_/X _2454_/X vssd1 vssd1 vccd1 vccd1 _3487_/D sky130_fd_sc_hd__a22o_1
X_2394_ _3531_/Q _2391_/X _2354_/X _2392_/X vssd1 vssd1 vccd1 vccd1 _3531_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3015_ _3234_/X _3235_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3015_/X sky130_fd_sc_hd__mux2_2
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3848_ _3867_/CLK _3848_/D vssd1 vssd1 vccd1 vccd1 _3848_/Q sky130_fd_sc_hd__dfxtp_1
X_3779_ _3827_/CLK _3779_/D vssd1 vssd1 vccd1 vccd1 _3779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater408 _1905_/A vssd1 vssd1 vccd1 vccd1 _3372_/S0 sky130_fd_sc_hd__buf_8
XFILLER_92_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1963_ _3778_/Q _1957_/X _1925_/X _1959_/X vssd1 vssd1 vccd1 vccd1 _3778_/D sky130_fd_sc_hd__a22o_1
X_3702_ _3719_/CLK _3702_/D vssd1 vssd1 vccd1 vccd1 _3702_/Q sky130_fd_sc_hd__dfxtp_1
X_1894_ _3806_/Q _1881_/A _1893_/X _1883_/A vssd1 vssd1 vccd1 vccd1 _3806_/D sky130_fd_sc_hd__a22o_1
X_3633_ _3667_/CLK _3633_/D vssd1 vssd1 vccd1 vccd1 _3633_/Q sky130_fd_sc_hd__dfxtp_1
X_3564_ _3741_/CLK _3564_/D vssd1 vssd1 vccd1 vccd1 _3564_/Q sky130_fd_sc_hd__dfxtp_1
X_2515_ _3452_/Q _2511_/X _2958_/A _2513_/X vssd1 vssd1 vccd1 vccd1 _3452_/D sky130_fd_sc_hd__a22o_1
X_3495_ _3816_/CLK _3495_/D vssd1 vssd1 vccd1 vccd1 _3495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2446_ _3495_/Q _2443_/X _2295_/X _2444_/X vssd1 vssd1 vccd1 vccd1 _3495_/D sky130_fd_sc_hd__a22o_1
X_2377_ _3544_/Q _2375_/X _2292_/X _2376_/X vssd1 vssd1 vccd1 vccd1 _3544_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3280_ _3589_/Q _3813_/Q _3541_/Q _3517_/Q _3291_/S0 _3292_/S1 vssd1 vssd1 vccd1
+ vccd1 _3280_/X sky130_fd_sc_hd__mux4_1
X_2300_ _3588_/Q _2291_/X _2255_/X _2293_/X vssd1 vssd1 vccd1 vccd1 _3588_/D sky130_fd_sc_hd__a22o_1
X_2231_ _2231_/A vssd1 vssd1 vccd1 vccd1 _2231_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2162_ _3675_/Q _2154_/X _2161_/X _2157_/X vssd1 vssd1 vccd1 vccd1 _3675_/D sky130_fd_sc_hd__a22o_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2093_ _2107_/A vssd1 vssd1 vccd1 vccd1 _2108_/A sky130_fd_sc_hd__inv_2
XFILLER_93_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2995_ _2994_/X _2836_/X _2997_/S vssd1 vssd1 vccd1 vccd1 _2995_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1946_ _3786_/Q _1940_/X _1925_/X _1942_/X vssd1 vssd1 vccd1 vccd1 _3786_/D sky130_fd_sc_hd__a22o_1
X_1877_ _2133_/A vssd1 vssd1 vccd1 vccd1 _1877_/X sky130_fd_sc_hd__clkbuf_2
X_3616_ _3720_/CLK _3616_/D vssd1 vssd1 vccd1 vccd1 _3616_/Q sky130_fd_sc_hd__dfxtp_1
X_3547_ _3831_/CLK _3547_/D vssd1 vssd1 vccd1 vccd1 _3547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3478_ _3812_/CLK _3478_/D vssd1 vssd1 vccd1 vccd1 _3478_/Q sky130_fd_sc_hd__dfxtp_1
X_2429_ _3506_/Q _2425_/X _2356_/X _2426_/X vssd1 vssd1 vccd1 vccd1 _3506_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1800_ _1801_/A _3368_/X vssd1 vssd1 vccd1 vccd1 _3843_/D sky130_fd_sc_hd__and2_1
XFILLER_34_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2780_ _3536_/Q vssd1 vssd1 vccd1 vccd1 _2780_/Y sky130_fd_sc_hd__inv_2
XPHY_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1731_ _2686_/A _1823_/B _2943_/A vssd1 vssd1 vccd1 vccd1 _1857_/D sky130_fd_sc_hd__or3_4
X_3401_ _3746_/CLK _3401_/D vssd1 vssd1 vccd1 vccd1 _3401_/Q sky130_fd_sc_hd__dfxtp_1
X_3332_ _3585_/Q _3809_/Q _3537_/Q _3513_/Q _1905_/A _3357_/S1 vssd1 vssd1 vccd1 vccd1
+ _3332_/X sky130_fd_sc_hd__mux4_1
X_3263_ _3759_/Q _3795_/Q _3827_/Q _3823_/Q _2971_/S _3286_/S1 vssd1 vssd1 vccd1 vccd1
+ _3263_/X sky130_fd_sc_hd__mux4_2
X_2214_ _2221_/A vssd1 vssd1 vccd1 vccd1 _2214_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3194_ _3429_/Q _3605_/Q _3581_/Q _3557_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3194_/X sky130_fd_sc_hd__mux4_2
X_2145_ _2145_/A vssd1 vssd1 vccd1 vccd1 _2145_/X sky130_fd_sc_hd__buf_2
XFILLER_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2076_ _2083_/A vssd1 vssd1 vccd1 vccd1 _2076_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2978_ _2978_/A0 _2978_/A1 _2984_/S vssd1 vssd1 vccd1 vccd1 _2978_/X sky130_fd_sc_hd__mux2_1
X_1929_ _2040_/A vssd1 vssd1 vccd1 vccd1 _2510_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_30_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_58_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3677_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_17_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2901_ _3591_/Q vssd1 vssd1 vccd1 vccd1 _2901_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3881_ _3896_/CLK _3881_/D vssd1 vssd1 vccd1 vccd1 _3881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2832_ _3443_/Q vssd1 vssd1 vccd1 vccd1 _2832_/Y sky130_fd_sc_hd__inv_2
X_2763_ _3807_/Q vssd1 vssd1 vccd1 vccd1 _2763_/Y sky130_fd_sc_hd__inv_2
X_1714_ _3892_/Q _1714_/B vssd1 vssd1 vccd1 vccd1 _1715_/B sky130_fd_sc_hd__nor2_2
XFILLER_8_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2694_ _3795_/Q vssd1 vssd1 vccd1 vccd1 _2694_/Y sky130_fd_sc_hd__inv_2
X_3315_ _3315_/A0 _3315_/A1 _3315_/A2 _3315_/A3 _2996_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3315_/X sky130_fd_sc_hd__mux4_1
XFILLER_86_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3246_ _3801_/Q _3757_/Q _3773_/Q _3769_/Q _3377_/S0 _3286_/S1 vssd1 vssd1 vccd1
+ vccd1 _3246_/X sky130_fd_sc_hd__mux4_2
XFILLER_86_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3177_ _3497_/Q _3473_/Q _3449_/Q _3737_/Q _3372_/S0 _3292_/S1 vssd1 vssd1 vccd1
+ vccd1 _3177_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2128_ _3688_/Q _2125_/X _2126_/X _2127_/X vssd1 vssd1 vccd1 vccd1 _3688_/D sky130_fd_sc_hd__a22o_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2059_ _3731_/Q _2057_/X _1882_/X _2058_/X vssd1 vssd1 vccd1 vccd1 _3731_/D sky130_fd_sc_hd__a22o_1
XFILLER_42_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3100_ _2846_/Y _2847_/Y _2844_/Y _2845_/Y _3153_/X _3132_/S1 vssd1 vssd1 vccd1 vccd1
+ _3100_/X sky130_fd_sc_hd__mux4_2
Xinput180 io_b_dat_o_9[1] vssd1 vssd1 vccd1 vccd1 _2994_/A1 sky130_fd_sc_hd__clkbuf_1
X_3031_ _3880_/Q _3282_/X _3061_/S vssd1 vssd1 vccd1 vccd1 _3031_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput191 io_dat_i[10] vssd1 vssd1 vccd1 vccd1 _2954_/A sky130_fd_sc_hd__buf_4
XFILLER_36_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3586_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3864_ _3867_/CLK _3864_/D vssd1 vssd1 vccd1 vccd1 _3864_/Q sky130_fd_sc_hd__dfxtp_1
X_2815_ _3466_/Q vssd1 vssd1 vccd1 vccd1 _2815_/Y sky130_fd_sc_hd__inv_2
X_3795_ _3796_/CLK _3795_/D vssd1 vssd1 vccd1 vccd1 _3795_/Q sky130_fd_sc_hd__dfxtp_1
X_2746_ _3582_/Q vssd1 vssd1 vccd1 vccd1 _2746_/Y sky130_fd_sc_hd__inv_2
X_2677_ _2681_/A input8/X _2682_/A _2682_/B vssd1 vssd1 vccd1 vccd1 _2677_/Y sky130_fd_sc_hd__nor4_2
XFILLER_86_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3229_ _3422_/Q _3598_/Q _3574_/Q _3550_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3229_/X sky130_fd_sc_hd__mux4_2
XFILLER_36_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2600_ _3391_/Q _2593_/A _2147_/A _2594_/A vssd1 vssd1 vccd1 vccd1 _3391_/D sky130_fd_sc_hd__a22o_1
X_3580_ _3748_/CLK _3580_/D vssd1 vssd1 vccd1 vccd1 _3580_/Q sky130_fd_sc_hd__dfxtp_1
X_2531_ _3440_/Q _2526_/X _2460_/X _2527_/X vssd1 vssd1 vccd1 vccd1 _3440_/D sky130_fd_sc_hd__a22o_1
X_2462_ _2945_/A vssd1 vssd1 vccd1 vccd1 _2462_/X sky130_fd_sc_hd__clkbuf_2
X_2393_ _3532_/Q _2391_/X _2351_/X _2392_/X vssd1 vssd1 vccd1 vccd1 _3532_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3014_ _3014_/A0 _3014_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3014_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3847_ _3867_/CLK _3847_/D vssd1 vssd1 vccd1 vccd1 _3847_/Q sky130_fd_sc_hd__dfxtp_1
X_3778_ _3827_/CLK _3778_/D vssd1 vssd1 vccd1 vccd1 _3778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2729_ _3606_/Q vssd1 vssd1 vccd1 vccd1 _2729_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater409 _1905_/A vssd1 vssd1 vccd1 vccd1 _3351_/S0 sky130_fd_sc_hd__buf_8
XFILLER_65_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1962_ _3779_/Q _1957_/X _1923_/X _1959_/X vssd1 vssd1 vccd1 vccd1 _3779_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3701_ _3813_/CLK _3701_/D vssd1 vssd1 vccd1 vccd1 _3701_/Q sky130_fd_sc_hd__dfxtp_1
X_1893_ _2149_/A vssd1 vssd1 vccd1 vccd1 _1893_/X sky130_fd_sc_hd__clkbuf_2
X_3632_ _3682_/CLK _3632_/D vssd1 vssd1 vccd1 vccd1 _3632_/Q sky130_fd_sc_hd__dfxtp_1
X_3563_ _3667_/CLK _3563_/D vssd1 vssd1 vccd1 vccd1 _3563_/Q sky130_fd_sc_hd__dfxtp_1
X_2514_ _3453_/Q _2511_/X _2959_/A _2513_/X vssd1 vssd1 vccd1 vccd1 _3453_/D sky130_fd_sc_hd__a22o_1
X_3494_ _3816_/CLK _3494_/D vssd1 vssd1 vccd1 vccd1 _3494_/Q sky130_fd_sc_hd__dfxtp_1
X_2445_ _3496_/Q _2443_/X _2292_/X _2444_/X vssd1 vssd1 vccd1 vccd1 _3496_/D sky130_fd_sc_hd__a22o_1
X_2376_ _2383_/A vssd1 vssd1 vccd1 vccd1 _2376_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _2230_/A vssd1 vssd1 vccd1 vccd1 _2230_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2161_ _2957_/A vssd1 vssd1 vccd1 vccd1 _2161_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2092_ _2107_/A vssd1 vssd1 vccd1 vccd1 _2092_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2994_ _2994_/A0 _2994_/A1 _2996_/S vssd1 vssd1 vccd1 vccd1 _2994_/X sky130_fd_sc_hd__mux2_1
X_1945_ _3787_/Q _1940_/X _1923_/X _1942_/X vssd1 vssd1 vccd1 vccd1 _3787_/D sky130_fd_sc_hd__a22o_1
X_1876_ _3814_/Q _1872_/X _1840_/X _1873_/X vssd1 vssd1 vccd1 vccd1 _3814_/D sky130_fd_sc_hd__a22o_1
X_3615_ _3687_/CLK _3615_/D vssd1 vssd1 vccd1 vccd1 _3615_/Q sky130_fd_sc_hd__dfxtp_1
X_3546_ _3832_/CLK _3546_/D vssd1 vssd1 vccd1 vccd1 _3546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3477_ _3741_/CLK _3477_/D vssd1 vssd1 vccd1 vccd1 _3477_/Q sky130_fd_sc_hd__dfxtp_1
X_2428_ _3507_/Q _2425_/X _2354_/X _2426_/X vssd1 vssd1 vccd1 vccd1 _3507_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2359_ _3553_/Q _2350_/X _2358_/X _2352_/X vssd1 vssd1 vccd1 vccd1 _3553_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1730_ _2960_/A vssd1 vssd1 vccd1 vccd1 _1823_/B sky130_fd_sc_hd__inv_2
X_3400_ _3867_/CLK _3400_/D vssd1 vssd1 vccd1 vccd1 _3400_/Q sky130_fd_sc_hd__dfxtp_1
X_3331_ _3665_/Q _3649_/Q _3633_/Q _3609_/Q input5/X _3357_/S1 vssd1 vssd1 vccd1 vccd1
+ _3331_/X sky130_fd_sc_hd__mux4_2
XFILLER_3_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3262_ _3799_/Q _3755_/Q _3771_/Q _3767_/Q _3060_/S _3294_/S1 vssd1 vssd1 vccd1 vccd1
+ _3262_/X sky130_fd_sc_hd__mux4_2
X_2213_ _3641_/Q _2206_/X _2123_/X _2208_/X vssd1 vssd1 vccd1 vccd1 _3641_/D sky130_fd_sc_hd__a22o_1
X_3193_ _3189_/X _3190_/X _3191_/X _3192_/X _3295_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3193_/X sky130_fd_sc_hd__mux4_2
XFILLER_93_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2144_ _3681_/Q _2137_/X _2143_/X _2139_/X vssd1 vssd1 vccd1 vccd1 _3681_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2075_ _2082_/A vssd1 vssd1 vccd1 vccd1 _2075_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2977_ _2976_/X _2631_/X _2981_/S vssd1 vssd1 vccd1 vccd1 _2977_/X sky130_fd_sc_hd__mux2_1
X_1928_ _1928_/A _1928_/B vssd1 vssd1 vccd1 vccd1 _2040_/A sky130_fd_sc_hd__or2_1
X_1859_ _2281_/A _2181_/B _2671_/A _2115_/D vssd1 vssd1 vccd1 vccd1 _1881_/A sky130_fd_sc_hd__or4_4
X_3529_ _3603_/CLK _3529_/D vssd1 vssd1 vccd1 vccd1 _3529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_27_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3890_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2900_ _3615_/Q vssd1 vssd1 vccd1 vccd1 _2900_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3880_ _3895_/CLK _3880_/D vssd1 vssd1 vccd1 vccd1 _3880_/Q sky130_fd_sc_hd__dfxtp_1
X_2831_ _3467_/Q vssd1 vssd1 vccd1 vccd1 _2831_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2762_ _3583_/Q vssd1 vssd1 vccd1 vccd1 _2762_/Y sky130_fd_sc_hd__inv_2
X_1713_ _3891_/Q _1713_/B vssd1 vssd1 vccd1 vccd1 _1714_/B sky130_fd_sc_hd__or2_2
XFILLER_8_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2693_ _3759_/Q vssd1 vssd1 vccd1 vccd1 _2693_/Y sky130_fd_sc_hd__inv_2
X_3314_ input24/X input56/X input72/X input88/X _2996_/S _2997_/S vssd1 vssd1 vccd1
+ vccd1 _3314_/X sky130_fd_sc_hd__mux4_1
XFILLER_86_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3245_ _2643_/X _2644_/X _3018_/X _2648_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3245_/X sky130_fd_sc_hd__mux4_2
XFILLER_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3176_ _3593_/Q _3817_/Q _3545_/Q _3521_/Q _3372_/S0 _3292_/S1 vssd1 vssd1 vccd1
+ vccd1 _3176_/X sky130_fd_sc_hd__mux4_2
X_2127_ _2139_/A vssd1 vssd1 vccd1 vccd1 _2127_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2058_ _2058_/A vssd1 vssd1 vccd1 vccd1 _2058_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3030_ _3275_/X _3276_/X _3062_/S vssd1 vssd1 vccd1 vccd1 _3030_/X sky130_fd_sc_hd__mux2_1
Xinput181 io_b_dat_o_9[2] vssd1 vssd1 vccd1 vccd1 _2992_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput170 io_b_dat_o_8[7] vssd1 vssd1 vccd1 vccd1 _2982_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput192 io_dat_i[11] vssd1 vssd1 vccd1 vccd1 _2955_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3863_ _3899_/CLK _3863_/D vssd1 vssd1 vccd1 vccd1 _3863_/Q sky130_fd_sc_hd__dfxtp_4
X_2814_ _3490_/Q vssd1 vssd1 vccd1 vccd1 _2814_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3794_ _3826_/CLK _3794_/D vssd1 vssd1 vccd1 vccd1 _3794_/Q sky130_fd_sc_hd__dfxtp_1
X_2745_ _3765_/Q vssd1 vssd1 vccd1 vccd1 _2745_/Y sky130_fd_sc_hd__inv_2
X_2676_ _2684_/A _2676_/B _2685_/C vssd1 vssd1 vccd1 vccd1 _2676_/Y sky130_fd_sc_hd__nor3_2
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3228_ _3224_/X _3225_/X _3226_/X _3227_/X _3862_/Q _3863_/Q vssd1 vssd1 vccd1 vccd1
+ _3228_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3159_ _3572_/Q _3724_/Q _3708_/Q _3692_/Q _3292_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3159_/X sky130_fd_sc_hd__mux4_2
XFILLER_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_42_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3719_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2530_ _3441_/Q _2526_/X _2458_/X _2527_/X vssd1 vssd1 vccd1 vccd1 _3441_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2461_ _3488_/Q _2452_/X _2460_/X _2454_/X vssd1 vssd1 vccd1 vccd1 _3488_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2392_ _2392_/A vssd1 vssd1 vccd1 vccd1 _2392_/X sky130_fd_sc_hd__clkbuf_2
X_3013_ _3013_/A0 _3013_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3013_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3846_ _3867_/CLK _3846_/D vssd1 vssd1 vccd1 vccd1 _3846_/Q sky130_fd_sc_hd__dfxtp_1
X_3777_ _3829_/CLK _3777_/D vssd1 vssd1 vccd1 vccd1 _3777_/Q sky130_fd_sc_hd__dfxtp_1
X_2728_ _3630_/Q vssd1 vssd1 vccd1 vccd1 _2728_/Y sky130_fd_sc_hd__inv_2
X_2659_ _2659_/A vssd1 vssd1 vccd1 vccd1 _2836_/A sky130_fd_sc_hd__buf_2
XFILLER_87_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1961_ _3780_/Q _1957_/X _1921_/X _1959_/X vssd1 vssd1 vccd1 vccd1 _3780_/D sky130_fd_sc_hd__a22o_1
X_3700_ _3700_/CLK _3700_/D vssd1 vssd1 vccd1 vccd1 _3700_/Q sky130_fd_sc_hd__dfxtp_1
X_1892_ _3807_/Q _1881_/X _1891_/X _1883_/X vssd1 vssd1 vccd1 vccd1 _3807_/D sky130_fd_sc_hd__a22o_1
X_3631_ _3667_/CLK _3631_/D vssd1 vssd1 vccd1 vccd1 _3631_/Q sky130_fd_sc_hd__dfxtp_1
X_3562_ _3682_/CLK _3562_/D vssd1 vssd1 vccd1 vccd1 _3562_/Q sky130_fd_sc_hd__dfxtp_1
X_2513_ _2527_/A vssd1 vssd1 vccd1 vccd1 _2513_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3493_ _3812_/CLK _3493_/D vssd1 vssd1 vccd1 vccd1 _3493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2444_ _2454_/A vssd1 vssd1 vccd1 vccd1 _2444_/X sky130_fd_sc_hd__clkbuf_2
X_2375_ _2382_/A vssd1 vssd1 vccd1 vccd1 _2375_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3829_ _3829_/CLK _3829_/D vssd1 vssd1 vccd1 vccd1 _3829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_0 _3261_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2160_ _3676_/Q _2154_/X _2159_/X _2157_/X vssd1 vssd1 vccd1 vccd1 _3676_/D sky130_fd_sc_hd__a22o_1
X_2091_ _2239_/A _2320_/B _2675_/A _2115_/D vssd1 vssd1 vccd1 vccd1 _2107_/A sky130_fd_sc_hd__or4_4
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2993_ _2992_/X _2640_/X _2997_/S vssd1 vssd1 vccd1 vccd1 _2993_/X sky130_fd_sc_hd__mux2_1
X_1944_ _3788_/Q _1940_/X _1921_/X _1942_/X vssd1 vssd1 vccd1 vccd1 _3788_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3614_ _3687_/CLK _3614_/D vssd1 vssd1 vccd1 vccd1 _3614_/Q sky130_fd_sc_hd__dfxtp_1
X_1875_ _3815_/Q _1872_/X _1837_/X _1873_/X vssd1 vssd1 vccd1 vccd1 _3815_/D sky130_fd_sc_hd__a22o_1
X_3545_ _3740_/CLK _3545_/D vssd1 vssd1 vccd1 vccd1 _3545_/Q sky130_fd_sc_hd__dfxtp_1
X_3476_ _3722_/CLK _3476_/D vssd1 vssd1 vccd1 vccd1 _3476_/Q sky130_fd_sc_hd__dfxtp_1
X_2427_ _3508_/Q _2425_/X _2351_/X _2426_/X vssd1 vssd1 vccd1 vccd1 _3508_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2358_ _2947_/A vssd1 vssd1 vccd1 vccd1 _2358_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2289_ _2955_/A vssd1 vssd1 vccd1 vccd1 _2289_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3330_ _3561_/Q _3713_/Q _3697_/Q _3681_/Q input5/X _3357_/S1 vssd1 vssd1 vccd1 vccd1
+ _3330_/X sky130_fd_sc_hd__mux4_2
X_3261_ _2629_/X _3023_/X _3024_/X _2632_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3261_/X sky130_fd_sc_hd__mux4_2
XFILLER_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2212_ _3642_/Q _2206_/X _2163_/X _2208_/X vssd1 vssd1 vccd1 vccd1 _3642_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3192_ _3494_/Q _3470_/Q _3446_/Q _3734_/Q _3060_/S _3192_/S1 vssd1 vssd1 vccd1 vccd1
+ _3192_/X sky130_fd_sc_hd__mux4_1
X_2143_ _2143_/A vssd1 vssd1 vccd1 vccd1 _2143_/X sky130_fd_sc_hd__buf_2
XFILLER_66_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2074_ _3721_/Q _2067_/X _2011_/X _2069_/X vssd1 vssd1 vccd1 vccd1 _3721_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2976_ _2976_/A0 _2976_/A1 _2984_/S vssd1 vssd1 vccd1 vccd1 _2976_/X sky130_fd_sc_hd__mux2_1
X_1927_ _2039_/A vssd1 vssd1 vccd1 vccd1 _1985_/A sky130_fd_sc_hd__buf_1
X_1858_ _2510_/D vssd1 vssd1 vccd1 vccd1 _2115_/D sky130_fd_sc_hd__buf_1
XFILLER_89_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1789_ _1789_/A _3261_/X vssd1 vssd1 vccd1 vccd1 _3852_/D sky130_fd_sc_hd__and2_1
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3528_ _3530_/CLK _3528_/D vssd1 vssd1 vccd1 vccd1 _3528_/Q sky130_fd_sc_hd__dfxtp_1
X_3459_ _3604_/CLK _3459_/D vssd1 vssd1 vccd1 vccd1 _3459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2830_ _3491_/Q vssd1 vssd1 vccd1 vccd1 _2830_/Y sky130_fd_sc_hd__inv_2
XPHY_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2761_ _3607_/Q vssd1 vssd1 vccd1 vccd1 _2761_/Y sky130_fd_sc_hd__inv_2
XPHY_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1712_ _3890_/Q _1712_/B vssd1 vssd1 vccd1 vccd1 _1713_/B sky130_fd_sc_hd__or2_1
XFILLER_8_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2692_ _3767_/Q vssd1 vssd1 vccd1 vccd1 _2692_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3313_ _3309_/X _3310_/X _3311_/X _3312_/X _2613_/A _3378_/S1 vssd1 vssd1 vccd1 vccd1
+ _3313_/X sky130_fd_sc_hd__mux4_1
X_3244_ input96/X _3244_/A1 _3244_/A2 _3244_/A3 _2971_/S _2981_/S vssd1 vssd1 vccd1
+ vccd1 _3244_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3175_ _3673_/Q _3657_/Q _3641_/Q _3617_/Q _3370_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3175_/X sky130_fd_sc_hd__mux4_2
X_2126_ _2954_/A vssd1 vssd1 vccd1 vccd1 _2126_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2057_ _2057_/A vssd1 vssd1 vccd1 vccd1 _2057_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2959_ _2959_/A vssd1 vssd1 vccd1 vccd1 _2959_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater390 _3286_/S1 vssd1 vssd1 vccd1 vccd1 _2981_/S sky130_fd_sc_hd__buf_8
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput171 io_b_dat_o_8[8] vssd1 vssd1 vccd1 vccd1 _2980_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput160 io_b_dat_o_8[12] vssd1 vssd1 vccd1 vccd1 _2971_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput182 io_b_dat_o_9[3] vssd1 vssd1 vccd1 vccd1 _2990_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput193 io_dat_i[12] vssd1 vssd1 vccd1 vccd1 _2956_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3862_ _3897_/CLK _3862_/D vssd1 vssd1 vccd1 vccd1 _3862_/Q sky130_fd_sc_hd__dfxtp_4
X_2813_ _3514_/Q vssd1 vssd1 vccd1 vccd1 _2813_/Y sky130_fd_sc_hd__inv_2
X_3793_ _3890_/CLK _3793_/D vssd1 vssd1 vccd1 vccd1 _3793_/Q sky130_fd_sc_hd__dfxtp_1
X_2744_ _3793_/Q vssd1 vssd1 vccd1 vccd1 _2744_/Y sky130_fd_sc_hd__inv_2
X_2675_ _2675_/A _2682_/B vssd1 vssd1 vccd1 vccd1 _2685_/C sky130_fd_sc_hd__or2_2
XFILLER_86_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3227_ _3399_/Q _3391_/Q _3383_/Q _3623_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3227_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3158_ _3154_/X _3155_/X _3156_/X _3157_/X _3295_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3158_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2109_ _3699_/Q _2107_/X _1882_/X _2108_/X vssd1 vssd1 vccd1 vccd1 _3699_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3089_ _2891_/Y _2892_/Y _2889_/Y _2890_/Y _3102_/S0 _3148_/X vssd1 vssd1 vccd1 vccd1
+ _3089_/X sky130_fd_sc_hd__mux4_2
XFILLER_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_11_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3530_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2460_ _2946_/A vssd1 vssd1 vccd1 vccd1 _2460_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2391_ _2391_/A vssd1 vssd1 vccd1 vccd1 _2391_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3012_ _3012_/A0 _3012_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3012_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3845_ _3845_/CLK _3845_/D vssd1 vssd1 vccd1 vccd1 _3845_/Q sky130_fd_sc_hd__dfxtp_1
X_3776_ _3827_/CLK _3776_/D vssd1 vssd1 vccd1 vccd1 _3776_/Q sky130_fd_sc_hd__dfxtp_1
X_2727_ _3646_/Q vssd1 vssd1 vccd1 vccd1 _2727_/Y sky130_fd_sc_hd__inv_2
X_2658_ _2664_/A _2967_/X vssd1 vssd1 vccd1 vccd1 _2658_/X sky130_fd_sc_hd__and2_1
X_2589_ _3400_/Q _2583_/X _2546_/X _2584_/X vssd1 vssd1 vccd1 vccd1 _3400_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1960_ _3781_/Q _1957_/X _1917_/X _1959_/X vssd1 vssd1 vccd1 vccd1 _3781_/D sky130_fd_sc_hd__a22o_1
XFILLER_61_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1891_ _2147_/A vssd1 vssd1 vccd1 vccd1 _1891_/X sky130_fd_sc_hd__buf_2
X_3630_ _3724_/CLK _3630_/D vssd1 vssd1 vccd1 vccd1 _3630_/Q sky130_fd_sc_hd__dfxtp_1
X_3561_ _3682_/CLK _3561_/D vssd1 vssd1 vccd1 vccd1 _3561_/Q sky130_fd_sc_hd__dfxtp_1
X_2512_ _2526_/A vssd1 vssd1 vccd1 vccd1 _2527_/A sky130_fd_sc_hd__inv_2
X_3492_ _3812_/CLK _3492_/D vssd1 vssd1 vccd1 vccd1 _3492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2443_ _2452_/A vssd1 vssd1 vccd1 vccd1 _2443_/X sky130_fd_sc_hd__clkbuf_2
X_2374_ _3545_/Q _2367_/X _2289_/X _2369_/X vssd1 vssd1 vccd1 vccd1 _3545_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3828_ _3828_/CLK _3828_/D vssd1 vssd1 vccd1 vccd1 _3828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3759_ _3796_/CLK _3759_/D vssd1 vssd1 vccd1 vccd1 _3759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_1 _3316_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2090_ input1/X vssd1 vssd1 vccd1 vccd1 _2320_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_93_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2992_ _2992_/A0 _2992_/A1 _2996_/S vssd1 vssd1 vccd1 vccd1 _2992_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1943_ _3789_/Q _1940_/X _1917_/X _1942_/X vssd1 vssd1 vccd1 vccd1 _3789_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3613_ _3672_/CLK _3613_/D vssd1 vssd1 vccd1 vccd1 _3613_/Q sky130_fd_sc_hd__dfxtp_1
X_1874_ _3816_/Q _1872_/X _1834_/X _1873_/X vssd1 vssd1 vccd1 vccd1 _3816_/D sky130_fd_sc_hd__a22o_1
X_3544_ _3813_/CLK _3544_/D vssd1 vssd1 vccd1 vccd1 _3544_/Q sky130_fd_sc_hd__dfxtp_1
X_3475_ _3722_/CLK _3475_/D vssd1 vssd1 vccd1 vccd1 _3475_/Q sky130_fd_sc_hd__dfxtp_1
X_2426_ _2426_/A vssd1 vssd1 vccd1 vccd1 _2426_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2357_ _3554_/Q _2350_/X _2356_/X _2352_/X vssd1 vssd1 vccd1 vccd1 _3554_/D sky130_fd_sc_hd__a22o_1
X_2288_ _3594_/Q _2282_/X _2163_/X _2284_/X vssd1 vssd1 vccd1 vccd1 _3594_/D sky130_fd_sc_hd__a22o_1
XFILLER_72_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3260_ input94/X _3260_/A1 _3260_/A2 _3260_/A3 _2984_/S _2981_/S vssd1 vssd1 vccd1
+ vccd1 _3260_/X sky130_fd_sc_hd__mux4_1
X_2211_ _3643_/Q _2206_/X _2161_/X _2208_/X vssd1 vssd1 vccd1 vccd1 _3643_/D sky130_fd_sc_hd__a22o_1
X_3191_ _3590_/Q _3814_/Q _3542_/Q _3518_/Q _3060_/S _3192_/S1 vssd1 vssd1 vccd1 vccd1
+ _3191_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2142_ _3682_/Q _2137_/X _2141_/X _2139_/X vssd1 vssd1 vccd1 vccd1 _3682_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2073_ _3722_/Q _2067_/X _1869_/X _2069_/X vssd1 vssd1 vccd1 vccd1 _3722_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2975_ _2974_/X _2637_/X _2981_/S vssd1 vssd1 vccd1 vccd1 _2975_/X sky130_fd_sc_hd__mux2_1
X_1926_ _3794_/Q _1916_/X _1925_/X _1919_/X vssd1 vssd1 vccd1 vccd1 _3794_/D sky130_fd_sc_hd__a22o_1
X_1857_ _1857_/A input2/X input3/X _1857_/D vssd1 vssd1 vccd1 vccd1 _2510_/D sky130_fd_sc_hd__or4_4
X_1788_ _1789_/A _3253_/X vssd1 vssd1 vccd1 vccd1 _3853_/D sky130_fd_sc_hd__and2_1
X_3527_ _3743_/CLK _3527_/D vssd1 vssd1 vccd1 vccd1 _3527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3458_ _3530_/CLK _3458_/D vssd1 vssd1 vccd1 vccd1 _3458_/Q sky130_fd_sc_hd__dfxtp_1
X_3389_ _3796_/CLK _3389_/D vssd1 vssd1 vccd1 vccd1 _3389_/Q sky130_fd_sc_hd__dfxtp_1
X_2409_ _2416_/A vssd1 vssd1 vccd1 vccd1 _2409_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3773_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2760_ _3631_/Q vssd1 vssd1 vccd1 vccd1 _2760_/Y sky130_fd_sc_hd__inv_2
XPHY_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1711_ _3889_/Q _3888_/Q vssd1 vssd1 vccd1 vccd1 _1712_/B sky130_fd_sc_hd__or2_1
X_2691_ _3771_/Q vssd1 vssd1 vccd1 vccd1 _2691_/Y sky130_fd_sc_hd__inv_2
X_3312_ _3403_/Q _3395_/Q _3387_/Q _3627_/Q _3364_/S0 _3338_/S1 vssd1 vssd1 vccd1
+ vccd1 _3312_/X sky130_fd_sc_hd__mux4_2
X_3243_ input16/X input48/X input64/X input80/X _2971_/S _2981_/S vssd1 vssd1 vccd1
+ vccd1 _3243_/X sky130_fd_sc_hd__mux4_1
X_3174_ _3569_/Q _3721_/Q _3705_/Q _3689_/Q _3372_/S0 _3372_/S1 vssd1 vssd1 vccd1
+ vccd1 _3174_/X sky130_fd_sc_hd__mux4_2
XFILLER_27_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2125_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2125_/X sky130_fd_sc_hd__clkbuf_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2056_ _3732_/Q _2050_/X _1879_/X _2051_/X vssd1 vssd1 vccd1 vccd1 _3732_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2958_ _2958_/A vssd1 vssd1 vccd1 vccd1 _2958_/X sky130_fd_sc_hd__clkbuf_1
X_1909_ _2554_/A vssd1 vssd1 vccd1 vccd1 _1909_/X sky130_fd_sc_hd__clkbuf_2
X_2889_ _3494_/Q vssd1 vssd1 vccd1 vccd1 _2889_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater380 _3378_/S1 vssd1 vssd1 vccd1 vccd1 _3373_/S1 sky130_fd_sc_hd__buf_8
XFILLER_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater391 _3294_/S1 vssd1 vssd1 vccd1 vccd1 _3286_/S1 sky130_fd_sc_hd__buf_8
XFILLER_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput150 io_b_dat_o_7[3] vssd1 vssd1 vccd1 vccd1 _3341_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput172 io_b_dat_o_8[9] vssd1 vssd1 vccd1 vccd1 _2978_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput161 io_b_dat_o_8[13] vssd1 vssd1 vccd1 vccd1 _2968_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput183 io_b_dat_o_9[4] vssd1 vssd1 vccd1 vccd1 _2988_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput194 io_dat_i[13] vssd1 vssd1 vccd1 vccd1 _2957_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3861_ _3897_/CLK _3861_/D vssd1 vssd1 vccd1 vccd1 _3861_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3792_ _3828_/CLK _3792_/D vssd1 vssd1 vccd1 vccd1 _3792_/Q sky130_fd_sc_hd__dfxtp_1
X_2812_ _3538_/Q vssd1 vssd1 vccd1 vccd1 _2812_/Y sky130_fd_sc_hd__inv_2
X_2743_ _3785_/Q vssd1 vssd1 vccd1 vccd1 _2743_/Y sky130_fd_sc_hd__inv_2
X_2674_ _2684_/A _2676_/B _2684_/C vssd1 vssd1 vccd1 vccd1 _2674_/Y sky130_fd_sc_hd__nor3_2
X_3226_ _3431_/Q _3743_/Q _3415_/Q _3407_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3226_/X sky130_fd_sc_hd__mux4_1
X_3157_ _3501_/Q _3477_/Q _3453_/Q _3741_/Q _3372_/S0 _3294_/S1 vssd1 vssd1 vccd1
+ vccd1 _3157_/X sky130_fd_sc_hd__mux4_2
XFILLER_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2108_ _2108_/A vssd1 vssd1 vccd1 vccd1 _2108_/X sky130_fd_sc_hd__clkbuf_2
X_3088_ _3084_/X _3085_/X _3086_/X _3087_/X _3133_/S0 _3138_/X vssd1 vssd1 vccd1 vccd1
+ _3088_/X sky130_fd_sc_hd__mux4_2
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2039_ _2039_/A vssd1 vssd1 vccd1 vccd1 _2239_/A sky130_fd_sc_hd__buf_1
XFILLER_50_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_51_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3741_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2390_ _3533_/Q _2002_/X _2348_/X _2004_/X vssd1 vssd1 vccd1 vccd1 _3533_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3011_ _3011_/A0 _3011_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3011_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3844_ _3845_/CLK _3844_/D vssd1 vssd1 vccd1 vccd1 _3844_/Q sky130_fd_sc_hd__dfxtp_1
X_3775_ _3827_/CLK _3775_/D vssd1 vssd1 vccd1 vccd1 _3775_/Q sky130_fd_sc_hd__dfxtp_1
X_2726_ _3662_/Q vssd1 vssd1 vccd1 vccd1 _2726_/Y sky130_fd_sc_hd__inv_2
X_2657_ _2664_/A _3163_/X vssd1 vssd1 vccd1 vccd1 _2657_/X sky130_fd_sc_hd__and2_1
X_2588_ _3401_/Q _2583_/X _2544_/X _2584_/X vssd1 vssd1 vccd1 vccd1 _3401_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3209_ _3426_/Q _3602_/Q _3578_/Q _3554_/Q _3860_/Q _3232_/S1 vssd1 vssd1 vccd1 vccd1
+ _3209_/X sky130_fd_sc_hd__mux4_2
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1890_ _3808_/Q _1881_/X _1889_/X _1883_/X vssd1 vssd1 vccd1 vccd1 _3808_/D sky130_fd_sc_hd__a22o_1
X_3560_ _3682_/CLK _3560_/D vssd1 vssd1 vccd1 vccd1 _3560_/Q sky130_fd_sc_hd__dfxtp_1
X_2511_ _2526_/A vssd1 vssd1 vccd1 vccd1 _2511_/X sky130_fd_sc_hd__clkbuf_2
X_3491_ _3731_/CLK _3491_/D vssd1 vssd1 vccd1 vccd1 _3491_/Q sky130_fd_sc_hd__dfxtp_1
X_2442_ _3497_/Q _2435_/X _2289_/X _2437_/X vssd1 vssd1 vccd1 vccd1 _3497_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2373_ _3546_/Q _2367_/X _2330_/X _2369_/X vssd1 vssd1 vccd1 vccd1 _3546_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3827_ _3827_/CLK _3827_/D vssd1 vssd1 vccd1 vccd1 _3827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3758_ _3823_/CLK _3758_/D vssd1 vssd1 vccd1 vccd1 _3758_/Q sky130_fd_sc_hd__dfxtp_1
X_2709_ _3772_/Q vssd1 vssd1 vccd1 vccd1 _2709_/Y sky130_fd_sc_hd__inv_2
X_3689_ _3724_/CLK _3689_/D vssd1 vssd1 vccd1 vccd1 _3689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_2 _3303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2991_ _2990_/X _2617_/X _2997_/S vssd1 vssd1 vccd1 vccd1 _2991_/X sky130_fd_sc_hd__mux2_1
X_1942_ _2584_/A vssd1 vssd1 vccd1 vccd1 _1942_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1873_ _1883_/A vssd1 vssd1 vccd1 vccd1 _1873_/X sky130_fd_sc_hd__clkbuf_2
X_3612_ _3832_/CLK _3612_/D vssd1 vssd1 vccd1 vccd1 _3612_/Q sky130_fd_sc_hd__dfxtp_1
X_3543_ _3719_/CLK _3543_/D vssd1 vssd1 vccd1 vccd1 _3543_/Q sky130_fd_sc_hd__dfxtp_1
X_3474_ _3722_/CLK _3474_/D vssd1 vssd1 vccd1 vccd1 _3474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2425_ _2425_/A vssd1 vssd1 vccd1 vccd1 _2425_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2356_ _2948_/A vssd1 vssd1 vccd1 vccd1 _2356_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2287_ _3595_/Q _2282_/X _2161_/X _2284_/X vssd1 vssd1 vccd1 vccd1 _3595_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _3644_/Q _2206_/X _2159_/X _2208_/X vssd1 vssd1 vccd1 vccd1 _3644_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3190_ _3670_/Q _3654_/Q _3638_/Q _3614_/Q _3060_/S _3192_/S1 vssd1 vssd1 vccd1 vccd1
+ _3190_/X sky130_fd_sc_hd__mux4_2
X_2141_ _2141_/A vssd1 vssd1 vccd1 vccd1 _2141_/X sky130_fd_sc_hd__buf_2
XFILLER_38_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2072_ _3723_/Q _2067_/X _1867_/X _2069_/X vssd1 vssd1 vccd1 vccd1 _3723_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2974_ _2974_/A0 _2974_/A1 _2984_/S vssd1 vssd1 vccd1 vccd1 _2974_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3807_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1925_ _1974_/A vssd1 vssd1 vccd1 vccd1 _1925_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1856_ _2021_/C vssd1 vssd1 vccd1 vccd1 _2671_/A sky130_fd_sc_hd__buf_2
X_1787_ _1789_/A _3245_/X vssd1 vssd1 vccd1 vccd1 _3854_/D sky130_fd_sc_hd__and2_1
X_3526_ _3801_/CLK _3526_/D vssd1 vssd1 vccd1 vccd1 _3526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3457_ _3603_/CLK _3457_/D vssd1 vssd1 vccd1 vccd1 _3457_/Q sky130_fd_sc_hd__dfxtp_1
X_3388_ _3895_/CLK _3388_/D vssd1 vssd1 vccd1 vccd1 _3388_/Q sky130_fd_sc_hd__dfxtp_1
X_2408_ _3521_/Q _2401_/X _2289_/X _2403_/X vssd1 vssd1 vccd1 vccd1 _3521_/D sky130_fd_sc_hd__a22o_1
X_2339_ _3564_/Q _2333_/X _2255_/X _2334_/X vssd1 vssd1 vccd1 vccd1 _3564_/D sky130_fd_sc_hd__a22o_1
XFILLER_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1710_ _3893_/Q vssd1 vssd1 vccd1 vccd1 _1715_/A sky130_fd_sc_hd__inv_2
X_2690_ _3755_/Q vssd1 vssd1 vccd1 vccd1 _2690_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3311_ _3435_/Q _3747_/Q _3419_/Q _3411_/Q _3364_/S0 _3338_/S1 vssd1 vssd1 vccd1
+ vccd1 _3311_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3242_ _2651_/X _2652_/X _3017_/X _2655_/X _2961_/X _2961_/S vssd1 vssd1 vccd1 vccd1
+ _3242_/X sky130_fd_sc_hd__mux4_2
X_3173_ _3169_/X _3170_/X _3171_/X _3172_/X _3295_/S0 _3373_/S1 vssd1 vssd1 vccd1
+ vccd1 _3173_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2124_ _3689_/Q _2116_/X _2123_/X _2118_/X vssd1 vssd1 vccd1 vccd1 _3689_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2055_ _3733_/Q _2050_/X _1877_/X _2051_/X vssd1 vssd1 vccd1 vccd1 _3733_/D sky130_fd_sc_hd__a22o_1
XFILLER_62_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2957_ _2957_/A vssd1 vssd1 vccd1 vccd1 _2957_/X sky130_fd_sc_hd__clkbuf_1
X_2888_ _3518_/Q vssd1 vssd1 vccd1 vccd1 _2888_/Y sky130_fd_sc_hd__inv_2
X_1908_ _2553_/A vssd1 vssd1 vccd1 vccd1 _2554_/A sky130_fd_sc_hd__inv_2
X_1839_ _2952_/A vssd1 vssd1 vccd1 vccd1 _1974_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3509_ _3773_/CLK _3509_/D vssd1 vssd1 vccd1 vccd1 _3509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater381 input8/X vssd1 vssd1 vccd1 vccd1 _3378_/S1 sky130_fd_sc_hd__buf_8
XFILLER_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater392 _3294_/S1 vssd1 vssd1 vccd1 vccd1 _3292_/S1 sky130_fd_sc_hd__buf_6
XFILLER_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput151 io_b_dat_o_7[4] vssd1 vssd1 vccd1 vccd1 _3328_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput140 io_b_dat_o_6[9] vssd1 vssd1 vccd1 vccd1 _3268_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput162 io_b_dat_o_8[14] vssd1 vssd1 vccd1 vccd1 _2965_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput173 io_b_dat_o_9[0] vssd1 vssd1 vccd1 vccd1 _2996_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput184 io_b_dat_o_9[5] vssd1 vssd1 vccd1 vccd1 _2986_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput195 io_dat_i[14] vssd1 vssd1 vccd1 vccd1 _2958_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3860_ _3896_/CLK _3860_/D vssd1 vssd1 vccd1 vccd1 _3860_/Q sky130_fd_sc_hd__dfxtp_4
X_3791_ _3791_/CLK _3791_/D vssd1 vssd1 vccd1 vccd1 _3791_/Q sky130_fd_sc_hd__dfxtp_1
X_2811_ _3810_/Q vssd1 vssd1 vccd1 vccd1 _2811_/Y sky130_fd_sc_hd__inv_2
X_2742_ _3789_/Q vssd1 vssd1 vccd1 vccd1 _2742_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2673_ _2673_/A _2682_/B vssd1 vssd1 vccd1 vccd1 _2684_/C sky130_fd_sc_hd__or2_4
X_3225_ _3527_/Q _3503_/Q _3479_/Q _3455_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3225_/X sky130_fd_sc_hd__mux4_2
XFILLER_82_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3156_ _3597_/Q _3821_/Q _3549_/Q _3525_/Q _3372_/S0 _3294_/S1 vssd1 vssd1 vccd1
+ vccd1 _3156_/X sky130_fd_sc_hd__mux4_1
X_2107_ _2107_/A vssd1 vssd1 vccd1 vccd1 _2107_/X sky130_fd_sc_hd__clkbuf_2
X_3087_ _2895_/Y _2896_/Y _2893_/Y _2894_/Y _3102_/S0 _3148_/X vssd1 vssd1 vccd1 vccd1
+ _3087_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2038_ _3742_/Q _2030_/A _1893_/X _2031_/A vssd1 vssd1 vccd1 vccd1 _3742_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3899_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3010_ _3010_/A0 _3010_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3010_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3843_ _3845_/CLK _3843_/D vssd1 vssd1 vccd1 vccd1 _3843_/Q sky130_fd_sc_hd__dfxtp_1
X_3774_ _3827_/CLK _3774_/D vssd1 vssd1 vccd1 vccd1 _3774_/Q sky130_fd_sc_hd__dfxtp_1
X_2725_ _2843_/A _2997_/X vssd1 vssd1 vccd1 vccd1 _2725_/X sky130_fd_sc_hd__and2_1
X_2656_ _2661_/A _2989_/X vssd1 vssd1 vccd1 vccd1 _2656_/X sky130_fd_sc_hd__and2_1
XFILLER_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2587_ _3402_/Q _2583_/X _2542_/X _2584_/X vssd1 vssd1 vccd1 vccd1 _3402_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3208_ _3204_/X _3205_/X _3206_/X _3207_/X _3862_/Q _3863_/Q vssd1 vssd1 vccd1 vccd1
+ _3208_/X sky130_fd_sc_hd__mux4_2
X_3139_ _2707_/Y _2708_/Y _2709_/Y _2710_/Y _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3139_/X sky130_fd_sc_hd__mux4_2
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3490_ _3714_/CLK _3490_/D vssd1 vssd1 vccd1 vccd1 _3490_/Q sky130_fd_sc_hd__dfxtp_1
X_2510_ _2510_/A _2510_/B _2510_/C _2510_/D vssd1 vssd1 vccd1 vccd1 _2526_/A sky130_fd_sc_hd__or4_4
X_2441_ _3498_/Q _2435_/X _2330_/X _2437_/X vssd1 vssd1 vccd1 vccd1 _3498_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2372_ _3547_/Q _2367_/X _2328_/X _2369_/X vssd1 vssd1 vccd1 vccd1 _3547_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3826_ _3826_/CLK _3826_/D vssd1 vssd1 vccd1 vccd1 _3826_/Q sky130_fd_sc_hd__dfxtp_1
X_3757_ _3773_/CLK _3757_/D vssd1 vssd1 vccd1 vccd1 _3757_/Q sky130_fd_sc_hd__dfxtp_1
X_2708_ _3756_/Q vssd1 vssd1 vccd1 vccd1 _2708_/Y sky130_fd_sc_hd__inv_2
X_3688_ _3720_/CLK _3688_/D vssd1 vssd1 vccd1 vccd1 _3688_/Q sky130_fd_sc_hd__dfxtp_1
X_2639_ _2659_/A vssd1 vssd1 vccd1 vccd1 _2654_/A sky130_fd_sc_hd__buf_2
XFILLER_87_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_3 _3277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput296 _2686_/Y vssd1 vssd1 vccd1 vccd1 io_ack_o sky130_fd_sc_hd__clkbuf_2
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2990_ _2990_/A0 _2990_/A1 _2996_/S vssd1 vssd1 vccd1 vccd1 _2990_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1941_ _2583_/A vssd1 vssd1 vccd1 vccd1 _2584_/A sky130_fd_sc_hd__inv_2
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1872_ _1881_/A vssd1 vssd1 vccd1 vccd1 _1872_/X sky130_fd_sc_hd__clkbuf_2
X_3611_ _3677_/CLK _3611_/D vssd1 vssd1 vccd1 vccd1 _3611_/Q sky130_fd_sc_hd__dfxtp_1
X_3542_ _3719_/CLK _3542_/D vssd1 vssd1 vccd1 vccd1 _3542_/Q sky130_fd_sc_hd__dfxtp_1
X_3473_ _3741_/CLK _3473_/D vssd1 vssd1 vccd1 vccd1 _3473_/Q sky130_fd_sc_hd__dfxtp_1
X_2424_ _3509_/Q _1916_/X _2348_/X _1919_/X vssd1 vssd1 vccd1 vccd1 _3509_/D sky130_fd_sc_hd__a22o_1
X_2355_ _3555_/Q _2350_/X _2354_/X _2352_/X vssd1 vssd1 vccd1 vccd1 _3555_/D sky130_fd_sc_hd__a22o_1
X_2286_ _3596_/Q _2282_/X _2159_/X _2284_/X vssd1 vssd1 vccd1 vccd1 _3596_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3809_ _3811_/CLK _3809_/D vssd1 vssd1 vccd1 vccd1 _3809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2140_ _3683_/Q _2137_/X _2138_/X _2139_/X vssd1 vssd1 vccd1 vccd1 _3683_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2071_ _3724_/Q _2067_/X _1865_/X _2069_/X vssd1 vssd1 vccd1 vccd1 _3724_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2973_ _2973_/A0 _2973_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _2973_/X sky130_fd_sc_hd__mux2_2
XFILLER_15_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1924_ _3795_/Q _1916_/X _1923_/X _1919_/X vssd1 vssd1 vccd1 vccd1 _3795_/D sky130_fd_sc_hd__a22o_1
XFILLER_15_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1855_ _1905_/A _1928_/B vssd1 vssd1 vccd1 vccd1 _2021_/C sky130_fd_sc_hd__or2_2
X_1786_ _1789_/A _3242_/X vssd1 vssd1 vccd1 vccd1 _3855_/D sky130_fd_sc_hd__and2_1
X_3525_ _3821_/CLK _3525_/D vssd1 vssd1 vccd1 vccd1 _3525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3456_ _3530_/CLK _3456_/D vssd1 vssd1 vccd1 vccd1 _3456_/Q sky130_fd_sc_hd__dfxtp_1
X_3387_ _3897_/CLK _3387_/D vssd1 vssd1 vccd1 vccd1 _3387_/Q sky130_fd_sc_hd__dfxtp_1
X_2407_ _3522_/Q _2401_/X _2330_/X _2403_/X vssd1 vssd1 vccd1 vccd1 _3522_/D sky130_fd_sc_hd__a22o_1
X_2338_ _3565_/Q _2333_/X _2253_/X _2334_/X vssd1 vssd1 vccd1 vccd1 _3565_/D sky130_fd_sc_hd__a22o_1
X_2269_ _2944_/A vssd1 vssd1 vccd1 vccd1 _2269_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_45_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3841_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3310_ _3531_/Q _3507_/Q _3483_/Q _3459_/Q _1905_/A _3351_/S1 vssd1 vssd1 vccd1 vccd1
+ _3310_/X sky130_fd_sc_hd__mux4_2
X_3241_ input97/X _3241_/A1 _3241_/A2 _3241_/A3 _2971_/S _2981_/S vssd1 vssd1 vccd1
+ vccd1 _3241_/X sky130_fd_sc_hd__mux4_1
X_3172_ _3498_/Q _3474_/Q _3450_/Q _3738_/Q _3292_/S0 _3292_/S1 vssd1 vssd1 vccd1
+ vccd1 _3172_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2123_ _2955_/A vssd1 vssd1 vccd1 vccd1 _2123_/X sky130_fd_sc_hd__clkbuf_2
X_2054_ _3734_/Q _2050_/X _2019_/X _2051_/X vssd1 vssd1 vccd1 vccd1 _3734_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2956_ _2956_/A vssd1 vssd1 vccd1 vccd1 _2956_/X sky130_fd_sc_hd__clkbuf_1
X_2887_ _3542_/Q vssd1 vssd1 vccd1 vccd1 _2887_/Y sky130_fd_sc_hd__inv_2
X_1907_ _2553_/A vssd1 vssd1 vccd1 vccd1 _1907_/X sky130_fd_sc_hd__clkbuf_2
X_1838_ _3827_/Q _1827_/X _1837_/X _1831_/X vssd1 vssd1 vccd1 vccd1 _3827_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1769_ _1775_/A vssd1 vssd1 vccd1 vccd1 _1774_/A sky130_fd_sc_hd__buf_4
X_3508_ _3604_/CLK _3508_/D vssd1 vssd1 vccd1 vccd1 _3508_/Q sky130_fd_sc_hd__dfxtp_1
X_3439_ _3727_/CLK _3439_/D vssd1 vssd1 vccd1 vccd1 _3439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater382 _3373_/S0 vssd1 vssd1 vccd1 vccd1 _3295_/S0 sky130_fd_sc_hd__buf_8
Xrepeater393 _3372_/S1 vssd1 vssd1 vccd1 vccd1 _3294_/S1 sky130_fd_sc_hd__buf_8
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput130 io_b_dat_o_6[14] vssd1 vssd1 vccd1 vccd1 _3238_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput141 io_b_dat_o_7[0] vssd1 vssd1 vccd1 vccd1 _3380_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput152 io_b_dat_o_7[5] vssd1 vssd1 vccd1 vccd1 _3315_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput163 io_b_dat_o_8[15] vssd1 vssd1 vccd1 vccd1 _2962_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput174 io_b_dat_o_9[10] vssd1 vssd1 vccd1 vccd1 _2976_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput185 io_b_dat_o_9[6] vssd1 vssd1 vccd1 vccd1 _2984_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput196 io_dat_i[15] vssd1 vssd1 vccd1 vccd1 _2959_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3790_ _3791_/CLK _3790_/D vssd1 vssd1 vccd1 vccd1 _3790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2810_ _3586_/Q vssd1 vssd1 vccd1 vccd1 _2810_/Y sky130_fd_sc_hd__inv_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2741_ _3777_/Q vssd1 vssd1 vccd1 vccd1 _2741_/Y sky130_fd_sc_hd__inv_2
XPHY_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2672_ _2684_/A _2676_/B _2683_/C vssd1 vssd1 vccd1 vccd1 _2672_/Y sky130_fd_sc_hd__nor3_2
X_3224_ _3423_/Q _3599_/Q _3575_/Q _3551_/Q _3232_/S0 _3232_/S1 vssd1 vssd1 vccd1
+ vccd1 _3224_/X sky130_fd_sc_hd__mux4_2
.ends

