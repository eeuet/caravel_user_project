VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sin3
  CLASS BLOCK ;
  FOREIGN sin3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN ao_reg[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 596.000 33.950 604.000 ;
    END
  END ao_reg[0]
  PIN ao_reg[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 596.000 170.110 604.000 ;
    END
  END ao_reg[10]
  PIN ao_reg[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 596.000 183.910 604.000 ;
    END
  END ao_reg[11]
  PIN ao_reg[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 596.000 197.710 604.000 ;
    END
  END ao_reg[12]
  PIN ao_reg[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 596.000 211.050 604.000 ;
    END
  END ao_reg[13]
  PIN ao_reg[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 596.000 224.850 604.000 ;
    END
  END ao_reg[14]
  PIN ao_reg[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 596.000 238.650 604.000 ;
    END
  END ao_reg[15]
  PIN ao_reg[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 596.000 251.990 604.000 ;
    END
  END ao_reg[16]
  PIN ao_reg[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 596.000 265.790 604.000 ;
    END
  END ao_reg[17]
  PIN ao_reg[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 596.000 279.590 604.000 ;
    END
  END ao_reg[18]
  PIN ao_reg[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 596.000 292.930 604.000 ;
    END
  END ao_reg[19]
  PIN ao_reg[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 596.000 47.290 604.000 ;
    END
  END ao_reg[1]
  PIN ao_reg[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 596.000 306.730 604.000 ;
    END
  END ao_reg[20]
  PIN ao_reg[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 596.000 320.070 604.000 ;
    END
  END ao_reg[21]
  PIN ao_reg[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 596.000 333.870 604.000 ;
    END
  END ao_reg[22]
  PIN ao_reg[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 596.000 347.670 604.000 ;
    END
  END ao_reg[23]
  PIN ao_reg[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 596.000 361.010 604.000 ;
    END
  END ao_reg[24]
  PIN ao_reg[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 596.000 374.810 604.000 ;
    END
  END ao_reg[25]
  PIN ao_reg[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 596.000 388.610 604.000 ;
    END
  END ao_reg[26]
  PIN ao_reg[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 596.000 401.950 604.000 ;
    END
  END ao_reg[27]
  PIN ao_reg[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 596.000 415.750 604.000 ;
    END
  END ao_reg[28]
  PIN ao_reg[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 596.000 429.550 604.000 ;
    END
  END ao_reg[29]
  PIN ao_reg[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 596.000 61.090 604.000 ;
    END
  END ao_reg[2]
  PIN ao_reg[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 596.000 442.890 604.000 ;
    END
  END ao_reg[30]
  PIN ao_reg[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 596.000 456.690 604.000 ;
    END
  END ao_reg[31]
  PIN ao_reg[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 596.000 74.890 604.000 ;
    END
  END ao_reg[3]
  PIN ao_reg[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 596.000 88.230 604.000 ;
    END
  END ao_reg[4]
  PIN ao_reg[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 596.000 102.030 604.000 ;
    END
  END ao_reg[5]
  PIN ao_reg[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 596.000 115.830 604.000 ;
    END
  END ao_reg[6]
  PIN ao_reg[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 596.000 129.170 604.000 ;
    END
  END ao_reg[7]
  PIN ao_reg[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 596.000 142.970 604.000 ;
    END
  END ao_reg[8]
  PIN ao_reg[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 596.000 156.770 604.000 ;
    END
  END ao_reg[9]
  PIN asel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 596.000 20.150 604.000 ;
    END
  END asel
  PIN bo_reg[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 596.000 470.490 604.000 ;
    END
  END bo_reg[0]
  PIN bo_reg[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 596.000 606.650 604.000 ;
    END
  END bo_reg[10]
  PIN bo_reg[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 596.000 620.450 604.000 ;
    END
  END bo_reg[11]
  PIN bo_reg[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 596.000 633.790 604.000 ;
    END
  END bo_reg[12]
  PIN bo_reg[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 596.000 647.590 604.000 ;
    END
  END bo_reg[13]
  PIN bo_reg[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 596.000 661.390 604.000 ;
    END
  END bo_reg[14]
  PIN bo_reg[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 596.000 674.730 604.000 ;
    END
  END bo_reg[15]
  PIN bo_reg[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 596.000 688.530 604.000 ;
    END
  END bo_reg[16]
  PIN bo_reg[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 596.000 702.330 604.000 ;
    END
  END bo_reg[17]
  PIN bo_reg[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 596.000 715.670 604.000 ;
    END
  END bo_reg[18]
  PIN bo_reg[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 596.000 729.470 604.000 ;
    END
  END bo_reg[19]
  PIN bo_reg[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 596.000 483.830 604.000 ;
    END
  END bo_reg[1]
  PIN bo_reg[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 596.000 743.270 604.000 ;
    END
  END bo_reg[20]
  PIN bo_reg[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 596.000 756.610 604.000 ;
    END
  END bo_reg[21]
  PIN bo_reg[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 596.000 770.410 604.000 ;
    END
  END bo_reg[22]
  PIN bo_reg[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 596.000 784.210 604.000 ;
    END
  END bo_reg[23]
  PIN bo_reg[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 596.000 797.550 604.000 ;
    END
  END bo_reg[24]
  PIN bo_reg[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 596.000 811.350 604.000 ;
    END
  END bo_reg[25]
  PIN bo_reg[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.870 596.000 825.150 604.000 ;
    END
  END bo_reg[26]
  PIN bo_reg[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 596.000 838.490 604.000 ;
    END
  END bo_reg[27]
  PIN bo_reg[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 596.000 852.290 604.000 ;
    END
  END bo_reg[28]
  PIN bo_reg[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 596.000 866.090 604.000 ;
    END
  END bo_reg[29]
  PIN bo_reg[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 596.000 497.630 604.000 ;
    END
  END bo_reg[2]
  PIN bo_reg[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 596.000 879.430 604.000 ;
    END
  END bo_reg[30]
  PIN bo_reg[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.950 596.000 893.230 604.000 ;
    END
  END bo_reg[31]
  PIN bo_reg[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 596.000 511.430 604.000 ;
    END
  END bo_reg[3]
  PIN bo_reg[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 596.000 524.770 604.000 ;
    END
  END bo_reg[4]
  PIN bo_reg[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 596.000 538.570 604.000 ;
    END
  END bo_reg[5]
  PIN bo_reg[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 596.000 552.370 604.000 ;
    END
  END bo_reg[6]
  PIN bo_reg[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 596.000 565.710 604.000 ;
    END
  END bo_reg[7]
  PIN bo_reg[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 596.000 579.510 604.000 ;
    END
  END bo_reg[8]
  PIN bo_reg[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 596.000 593.310 604.000 ;
    END
  END bo_reg[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 596.000 6.810 604.000 ;
    END
  END clk
  PIN e_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 4.120 904.000 4.720 ;
    END
  END e_i[0]
  PIN e_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 191.120 904.000 191.720 ;
    END
  END e_i[10]
  PIN e_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 210.160 904.000 210.760 ;
    END
  END e_i[11]
  PIN e_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 228.520 904.000 229.120 ;
    END
  END e_i[12]
  PIN e_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 247.560 904.000 248.160 ;
    END
  END e_i[13]
  PIN e_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 265.920 904.000 266.520 ;
    END
  END e_i[14]
  PIN e_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 284.960 904.000 285.560 ;
    END
  END e_i[15]
  PIN e_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 304.000 904.000 304.600 ;
    END
  END e_i[16]
  PIN e_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 322.360 904.000 322.960 ;
    END
  END e_i[17]
  PIN e_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 341.400 904.000 342.000 ;
    END
  END e_i[18]
  PIN e_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 359.760 904.000 360.360 ;
    END
  END e_i[19]
  PIN e_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 22.480 904.000 23.080 ;
    END
  END e_i[1]
  PIN e_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 378.800 904.000 379.400 ;
    END
  END e_i[20]
  PIN e_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 397.160 904.000 397.760 ;
    END
  END e_i[21]
  PIN e_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 416.200 904.000 416.800 ;
    END
  END e_i[22]
  PIN e_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 434.560 904.000 435.160 ;
    END
  END e_i[23]
  PIN e_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 453.600 904.000 454.200 ;
    END
  END e_i[24]
  PIN e_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 472.640 904.000 473.240 ;
    END
  END e_i[25]
  PIN e_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 491.000 904.000 491.600 ;
    END
  END e_i[26]
  PIN e_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 510.040 904.000 510.640 ;
    END
  END e_i[27]
  PIN e_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 528.400 904.000 529.000 ;
    END
  END e_i[28]
  PIN e_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 547.440 904.000 548.040 ;
    END
  END e_i[29]
  PIN e_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 41.520 904.000 42.120 ;
    END
  END e_i[2]
  PIN e_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 565.800 904.000 566.400 ;
    END
  END e_i[30]
  PIN e_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 584.840 904.000 585.440 ;
    END
  END e_i[31]
  PIN e_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 59.880 904.000 60.480 ;
    END
  END e_i[3]
  PIN e_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 78.920 904.000 79.520 ;
    END
  END e_i[4]
  PIN e_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 97.280 904.000 97.880 ;
    END
  END e_i[5]
  PIN e_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 116.320 904.000 116.920 ;
    END
  END e_i[6]
  PIN e_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 134.680 904.000 135.280 ;
    END
  END e_i[7]
  PIN e_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 153.720 904.000 154.320 ;
    END
  END e_i[8]
  PIN e_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 172.760 904.000 173.360 ;
    END
  END e_i[9]
  PIN e_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 12.960 904.000 13.560 ;
    END
  END e_o[0]
  PIN e_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 200.640 904.000 201.240 ;
    END
  END e_o[10]
  PIN e_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 219.000 904.000 219.600 ;
    END
  END e_o[11]
  PIN e_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 238.040 904.000 238.640 ;
    END
  END e_o[12]
  PIN e_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 257.080 904.000 257.680 ;
    END
  END e_o[13]
  PIN e_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 275.440 904.000 276.040 ;
    END
  END e_o[14]
  PIN e_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 294.480 904.000 295.080 ;
    END
  END e_o[15]
  PIN e_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 312.840 904.000 313.440 ;
    END
  END e_o[16]
  PIN e_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 331.880 904.000 332.480 ;
    END
  END e_o[17]
  PIN e_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 350.240 904.000 350.840 ;
    END
  END e_o[18]
  PIN e_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 369.280 904.000 369.880 ;
    END
  END e_o[19]
  PIN e_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 32.000 904.000 32.600 ;
    END
  END e_o[1]
  PIN e_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 388.320 904.000 388.920 ;
    END
  END e_o[20]
  PIN e_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 406.680 904.000 407.280 ;
    END
  END e_o[21]
  PIN e_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 425.720 904.000 426.320 ;
    END
  END e_o[22]
  PIN e_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 444.080 904.000 444.680 ;
    END
  END e_o[23]
  PIN e_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 463.120 904.000 463.720 ;
    END
  END e_o[24]
  PIN e_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 481.480 904.000 482.080 ;
    END
  END e_o[25]
  PIN e_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 500.520 904.000 501.120 ;
    END
  END e_o[26]
  PIN e_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 518.880 904.000 519.480 ;
    END
  END e_o[27]
  PIN e_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 537.920 904.000 538.520 ;
    END
  END e_o[28]
  PIN e_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 556.960 904.000 557.560 ;
    END
  END e_o[29]
  PIN e_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 50.360 904.000 50.960 ;
    END
  END e_o[2]
  PIN e_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 575.320 904.000 575.920 ;
    END
  END e_o[30]
  PIN e_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 594.360 904.000 594.960 ;
    END
  END e_o[31]
  PIN e_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 69.400 904.000 70.000 ;
    END
  END e_o[3]
  PIN e_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 88.440 904.000 89.040 ;
    END
  END e_o[4]
  PIN e_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 106.800 904.000 107.400 ;
    END
  END e_o[5]
  PIN e_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 125.840 904.000 126.440 ;
    END
  END e_o[6]
  PIN e_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 144.200 904.000 144.800 ;
    END
  END e_o[7]
  PIN e_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 163.240 904.000 163.840 ;
    END
  END e_o[8]
  PIN e_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 181.600 904.000 182.200 ;
    END
  END e_o[9]
  PIN se_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 -4.000 453.470 4.000 ;
    END
  END se_i[0]
  PIN se_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 -4.000 594.230 4.000 ;
    END
  END se_i[10]
  PIN se_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.750 -4.000 608.030 4.000 ;
    END
  END se_i[11]
  PIN se_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 -4.000 622.290 4.000 ;
    END
  END se_i[12]
  PIN se_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 -4.000 636.550 4.000 ;
    END
  END se_i[13]
  PIN se_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 -4.000 650.350 4.000 ;
    END
  END se_i[14]
  PIN se_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 -4.000 664.610 4.000 ;
    END
  END se_i[15]
  PIN se_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 -4.000 678.410 4.000 ;
    END
  END se_i[16]
  PIN se_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 -4.000 692.670 4.000 ;
    END
  END se_i[17]
  PIN se_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 -4.000 706.470 4.000 ;
    END
  END se_i[18]
  PIN se_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 -4.000 720.730 4.000 ;
    END
  END se_i[19]
  PIN se_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 -4.000 467.730 4.000 ;
    END
  END se_i[1]
  PIN se_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 -4.000 734.990 4.000 ;
    END
  END se_i[20]
  PIN se_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 -4.000 748.790 4.000 ;
    END
  END se_i[21]
  PIN se_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 -4.000 763.050 4.000 ;
    END
  END se_i[22]
  PIN se_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 -4.000 776.850 4.000 ;
    END
  END se_i[23]
  PIN se_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 -4.000 791.110 4.000 ;
    END
  END se_i[24]
  PIN se_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 -4.000 804.910 4.000 ;
    END
  END se_i[25]
  PIN se_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 -4.000 819.170 4.000 ;
    END
  END se_i[26]
  PIN se_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 -4.000 833.430 4.000 ;
    END
  END se_i[27]
  PIN se_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 -4.000 847.230 4.000 ;
    END
  END se_i[28]
  PIN se_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 -4.000 861.490 4.000 ;
    END
  END se_i[29]
  PIN se_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 -4.000 481.530 4.000 ;
    END
  END se_i[2]
  PIN se_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 -4.000 875.290 4.000 ;
    END
  END se_i[30]
  PIN se_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 -4.000 889.550 4.000 ;
    END
  END se_i[31]
  PIN se_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 -4.000 495.790 4.000 ;
    END
  END se_i[3]
  PIN se_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 -4.000 509.590 4.000 ;
    END
  END se_i[4]
  PIN se_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 -4.000 523.850 4.000 ;
    END
  END se_i[5]
  PIN se_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 -4.000 537.650 4.000 ;
    END
  END se_i[6]
  PIN se_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 -4.000 551.910 4.000 ;
    END
  END se_i[7]
  PIN se_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 -4.000 566.170 4.000 ;
    END
  END se_i[8]
  PIN se_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 -4.000 579.970 4.000 ;
    END
  END se_i[9]
  PIN se_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 -4.000 460.370 4.000 ;
    END
  END se_o[0]
  PIN se_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 -4.000 601.130 4.000 ;
    END
  END se_o[10]
  PIN se_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 -4.000 615.390 4.000 ;
    END
  END se_o[11]
  PIN se_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 -4.000 629.190 4.000 ;
    END
  END se_o[12]
  PIN se_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 -4.000 643.450 4.000 ;
    END
  END se_o[13]
  PIN se_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 -4.000 657.250 4.000 ;
    END
  END se_o[14]
  PIN se_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 -4.000 671.510 4.000 ;
    END
  END se_o[15]
  PIN se_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 -4.000 685.770 4.000 ;
    END
  END se_o[16]
  PIN se_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 -4.000 699.570 4.000 ;
    END
  END se_o[17]
  PIN se_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 -4.000 713.830 4.000 ;
    END
  END se_o[18]
  PIN se_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 -4.000 727.630 4.000 ;
    END
  END se_o[19]
  PIN se_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 -4.000 474.630 4.000 ;
    END
  END se_o[1]
  PIN se_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 -4.000 741.890 4.000 ;
    END
  END se_o[20]
  PIN se_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 -4.000 755.690 4.000 ;
    END
  END se_o[21]
  PIN se_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 -4.000 769.950 4.000 ;
    END
  END se_o[22]
  PIN se_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 -4.000 784.210 4.000 ;
    END
  END se_o[23]
  PIN se_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 -4.000 798.010 4.000 ;
    END
  END se_o[24]
  PIN se_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 -4.000 812.270 4.000 ;
    END
  END se_o[25]
  PIN se_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 -4.000 826.070 4.000 ;
    END
  END se_o[26]
  PIN se_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.050 -4.000 840.330 4.000 ;
    END
  END se_o[27]
  PIN se_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.850 -4.000 854.130 4.000 ;
    END
  END se_o[28]
  PIN se_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 -4.000 868.390 4.000 ;
    END
  END se_o[29]
  PIN se_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 -4.000 488.430 4.000 ;
    END
  END se_o[2]
  PIN se_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 -4.000 882.650 4.000 ;
    END
  END se_o[30]
  PIN se_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.170 -4.000 896.450 4.000 ;
    END
  END se_o[31]
  PIN se_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 -4.000 502.690 4.000 ;
    END
  END se_o[3]
  PIN se_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 -4.000 516.950 4.000 ;
    END
  END se_o[4]
  PIN se_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 -4.000 530.750 4.000 ;
    END
  END se_o[5]
  PIN se_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 -4.000 545.010 4.000 ;
    END
  END se_o[6]
  PIN se_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 -4.000 558.810 4.000 ;
    END
  END se_o[7]
  PIN se_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 -4.000 573.070 4.000 ;
    END
  END se_o[8]
  PIN se_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 -4.000 586.870 4.000 ;
    END
  END se_o[9]
  PIN sw_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 -4.000 3.590 4.000 ;
    END
  END sw_i[0]
  PIN sw_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 -4.000 143.890 4.000 ;
    END
  END sw_i[10]
  PIN sw_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 -4.000 158.150 4.000 ;
    END
  END sw_i[11]
  PIN sw_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 -4.000 171.950 4.000 ;
    END
  END sw_i[12]
  PIN sw_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 -4.000 186.210 4.000 ;
    END
  END sw_i[13]
  PIN sw_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 -4.000 200.470 4.000 ;
    END
  END sw_i[14]
  PIN sw_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 -4.000 214.270 4.000 ;
    END
  END sw_i[15]
  PIN sw_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 -4.000 228.530 4.000 ;
    END
  END sw_i[16]
  PIN sw_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 -4.000 242.330 4.000 ;
    END
  END sw_i[17]
  PIN sw_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 -4.000 256.590 4.000 ;
    END
  END sw_i[18]
  PIN sw_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 -4.000 270.390 4.000 ;
    END
  END sw_i[19]
  PIN sw_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 -4.000 17.390 4.000 ;
    END
  END sw_i[1]
  PIN sw_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 -4.000 284.650 4.000 ;
    END
  END sw_i[20]
  PIN sw_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 -4.000 298.910 4.000 ;
    END
  END sw_i[21]
  PIN sw_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 -4.000 312.710 4.000 ;
    END
  END sw_i[22]
  PIN sw_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 -4.000 326.970 4.000 ;
    END
  END sw_i[23]
  PIN sw_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 -4.000 340.770 4.000 ;
    END
  END sw_i[24]
  PIN sw_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 -4.000 355.030 4.000 ;
    END
  END sw_i[25]
  PIN sw_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 -4.000 369.290 4.000 ;
    END
  END sw_i[26]
  PIN sw_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 -4.000 383.090 4.000 ;
    END
  END sw_i[27]
  PIN sw_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 -4.000 397.350 4.000 ;
    END
  END sw_i[28]
  PIN sw_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 -4.000 411.150 4.000 ;
    END
  END sw_i[29]
  PIN sw_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 -4.000 31.650 4.000 ;
    END
  END sw_i[2]
  PIN sw_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 -4.000 425.410 4.000 ;
    END
  END sw_i[30]
  PIN sw_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 -4.000 439.210 4.000 ;
    END
  END sw_i[31]
  PIN sw_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 -4.000 45.450 4.000 ;
    END
  END sw_i[3]
  PIN sw_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 -4.000 59.710 4.000 ;
    END
  END sw_i[4]
  PIN sw_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 -4.000 73.510 4.000 ;
    END
  END sw_i[5]
  PIN sw_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 -4.000 87.770 4.000 ;
    END
  END sw_i[6]
  PIN sw_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 -4.000 102.030 4.000 ;
    END
  END sw_i[7]
  PIN sw_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 -4.000 115.830 4.000 ;
    END
  END sw_i[8]
  PIN sw_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 -4.000 130.090 4.000 ;
    END
  END sw_i[9]
  PIN sw_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 -4.000 10.490 4.000 ;
    END
  END sw_o[0]
  PIN sw_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 -4.000 151.250 4.000 ;
    END
  END sw_o[10]
  PIN sw_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 -4.000 165.050 4.000 ;
    END
  END sw_o[11]
  PIN sw_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 -4.000 179.310 4.000 ;
    END
  END sw_o[12]
  PIN sw_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 -4.000 193.110 4.000 ;
    END
  END sw_o[13]
  PIN sw_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 -4.000 207.370 4.000 ;
    END
  END sw_o[14]
  PIN sw_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 -4.000 221.170 4.000 ;
    END
  END sw_o[15]
  PIN sw_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 -4.000 235.430 4.000 ;
    END
  END sw_o[16]
  PIN sw_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 -4.000 249.690 4.000 ;
    END
  END sw_o[17]
  PIN sw_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 -4.000 263.490 4.000 ;
    END
  END sw_o[18]
  PIN sw_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 -4.000 277.750 4.000 ;
    END
  END sw_o[19]
  PIN sw_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 -4.000 24.290 4.000 ;
    END
  END sw_o[1]
  PIN sw_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 -4.000 291.550 4.000 ;
    END
  END sw_o[20]
  PIN sw_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 -4.000 305.810 4.000 ;
    END
  END sw_o[21]
  PIN sw_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 -4.000 320.070 4.000 ;
    END
  END sw_o[22]
  PIN sw_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 -4.000 333.870 4.000 ;
    END
  END sw_o[23]
  PIN sw_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 -4.000 348.130 4.000 ;
    END
  END sw_o[24]
  PIN sw_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 -4.000 361.930 4.000 ;
    END
  END sw_o[25]
  PIN sw_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 -4.000 376.190 4.000 ;
    END
  END sw_o[26]
  PIN sw_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 -4.000 389.990 4.000 ;
    END
  END sw_o[27]
  PIN sw_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 -4.000 404.250 4.000 ;
    END
  END sw_o[28]
  PIN sw_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 -4.000 418.510 4.000 ;
    END
  END sw_o[29]
  PIN sw_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 -4.000 38.550 4.000 ;
    END
  END sw_o[2]
  PIN sw_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 -4.000 432.310 4.000 ;
    END
  END sw_o[30]
  PIN sw_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 -4.000 446.570 4.000 ;
    END
  END sw_o[31]
  PIN sw_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 -4.000 52.810 4.000 ;
    END
  END sw_o[3]
  PIN sw_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 -4.000 66.610 4.000 ;
    END
  END sw_o[4]
  PIN sw_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 -4.000 80.870 4.000 ;
    END
  END sw_o[5]
  PIN sw_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 -4.000 94.670 4.000 ;
    END
  END sw_o[6]
  PIN sw_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 -4.000 108.930 4.000 ;
    END
  END sw_o[7]
  PIN sw_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 -4.000 122.730 4.000 ;
    END
  END sw_o[8]
  PIN sw_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 -4.000 136.990 4.000 ;
    END
  END sw_o[9]
  PIN w_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 4.120 4.000 4.720 ;
    END
  END w_i[0]
  PIN w_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 191.120 4.000 191.720 ;
    END
  END w_i[10]
  PIN w_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 210.160 4.000 210.760 ;
    END
  END w_i[11]
  PIN w_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 228.520 4.000 229.120 ;
    END
  END w_i[12]
  PIN w_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 247.560 4.000 248.160 ;
    END
  END w_i[13]
  PIN w_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 265.920 4.000 266.520 ;
    END
  END w_i[14]
  PIN w_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 284.960 4.000 285.560 ;
    END
  END w_i[15]
  PIN w_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 304.000 4.000 304.600 ;
    END
  END w_i[16]
  PIN w_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 322.360 4.000 322.960 ;
    END
  END w_i[17]
  PIN w_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 341.400 4.000 342.000 ;
    END
  END w_i[18]
  PIN w_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 359.760 4.000 360.360 ;
    END
  END w_i[19]
  PIN w_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 22.480 4.000 23.080 ;
    END
  END w_i[1]
  PIN w_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 378.800 4.000 379.400 ;
    END
  END w_i[20]
  PIN w_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 397.160 4.000 397.760 ;
    END
  END w_i[21]
  PIN w_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 416.200 4.000 416.800 ;
    END
  END w_i[22]
  PIN w_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 434.560 4.000 435.160 ;
    END
  END w_i[23]
  PIN w_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 453.600 4.000 454.200 ;
    END
  END w_i[24]
  PIN w_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 472.640 4.000 473.240 ;
    END
  END w_i[25]
  PIN w_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 491.000 4.000 491.600 ;
    END
  END w_i[26]
  PIN w_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 510.040 4.000 510.640 ;
    END
  END w_i[27]
  PIN w_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 528.400 4.000 529.000 ;
    END
  END w_i[28]
  PIN w_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 547.440 4.000 548.040 ;
    END
  END w_i[29]
  PIN w_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 41.520 4.000 42.120 ;
    END
  END w_i[2]
  PIN w_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 565.800 4.000 566.400 ;
    END
  END w_i[30]
  PIN w_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 584.840 4.000 585.440 ;
    END
  END w_i[31]
  PIN w_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 59.880 4.000 60.480 ;
    END
  END w_i[3]
  PIN w_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 78.920 4.000 79.520 ;
    END
  END w_i[4]
  PIN w_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 97.280 4.000 97.880 ;
    END
  END w_i[5]
  PIN w_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 116.320 4.000 116.920 ;
    END
  END w_i[6]
  PIN w_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 134.680 4.000 135.280 ;
    END
  END w_i[7]
  PIN w_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 153.720 4.000 154.320 ;
    END
  END w_i[8]
  PIN w_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 172.760 4.000 173.360 ;
    END
  END w_i[9]
  PIN w_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 12.960 4.000 13.560 ;
    END
  END w_o[0]
  PIN w_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 200.640 4.000 201.240 ;
    END
  END w_o[10]
  PIN w_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 219.000 4.000 219.600 ;
    END
  END w_o[11]
  PIN w_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 238.040 4.000 238.640 ;
    END
  END w_o[12]
  PIN w_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 257.080 4.000 257.680 ;
    END
  END w_o[13]
  PIN w_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 275.440 4.000 276.040 ;
    END
  END w_o[14]
  PIN w_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 294.480 4.000 295.080 ;
    END
  END w_o[15]
  PIN w_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 312.840 4.000 313.440 ;
    END
  END w_o[16]
  PIN w_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 331.880 4.000 332.480 ;
    END
  END w_o[17]
  PIN w_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 350.240 4.000 350.840 ;
    END
  END w_o[18]
  PIN w_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 369.280 4.000 369.880 ;
    END
  END w_o[19]
  PIN w_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 32.000 4.000 32.600 ;
    END
  END w_o[1]
  PIN w_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 388.320 4.000 388.920 ;
    END
  END w_o[20]
  PIN w_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 406.680 4.000 407.280 ;
    END
  END w_o[21]
  PIN w_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 425.720 4.000 426.320 ;
    END
  END w_o[22]
  PIN w_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 444.080 4.000 444.680 ;
    END
  END w_o[23]
  PIN w_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 463.120 4.000 463.720 ;
    END
  END w_o[24]
  PIN w_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 481.480 4.000 482.080 ;
    END
  END w_o[25]
  PIN w_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 500.520 4.000 501.120 ;
    END
  END w_o[26]
  PIN w_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 518.880 4.000 519.480 ;
    END
  END w_o[27]
  PIN w_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 537.920 4.000 538.520 ;
    END
  END w_o[28]
  PIN w_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 556.960 4.000 557.560 ;
    END
  END w_o[29]
  PIN w_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 50.360 4.000 50.960 ;
    END
  END w_o[2]
  PIN w_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 575.320 4.000 575.920 ;
    END
  END w_o[30]
  PIN w_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 594.360 4.000 594.960 ;
    END
  END w_o[31]
  PIN w_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 69.400 4.000 70.000 ;
    END
  END w_o[3]
  PIN w_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 88.440 4.000 89.040 ;
    END
  END w_o[4]
  PIN w_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 106.800 4.000 107.400 ;
    END
  END w_o[5]
  PIN w_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 125.840 4.000 126.440 ;
    END
  END w_o[6]
  PIN w_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 144.200 4.000 144.800 ;
    END
  END w_o[7]
  PIN w_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 163.240 4.000 163.840 ;
    END
  END w_o[8]
  PIN w_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 181.600 4.000 182.200 ;
    END
  END w_o[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 3.290 10.640 896.470 587.760 ;
      LAYER met2 ;
        RECT 3.320 595.720 6.250 596.000 ;
        RECT 7.090 595.720 19.590 596.000 ;
        RECT 20.430 595.720 33.390 596.000 ;
        RECT 34.230 595.720 46.730 596.000 ;
        RECT 47.570 595.720 60.530 596.000 ;
        RECT 61.370 595.720 74.330 596.000 ;
        RECT 75.170 595.720 87.670 596.000 ;
        RECT 88.510 595.720 101.470 596.000 ;
        RECT 102.310 595.720 115.270 596.000 ;
        RECT 116.110 595.720 128.610 596.000 ;
        RECT 129.450 595.720 142.410 596.000 ;
        RECT 143.250 595.720 156.210 596.000 ;
        RECT 157.050 595.720 169.550 596.000 ;
        RECT 170.390 595.720 183.350 596.000 ;
        RECT 184.190 595.720 197.150 596.000 ;
        RECT 197.990 595.720 210.490 596.000 ;
        RECT 211.330 595.720 224.290 596.000 ;
        RECT 225.130 595.720 238.090 596.000 ;
        RECT 238.930 595.720 251.430 596.000 ;
        RECT 252.270 595.720 265.230 596.000 ;
        RECT 266.070 595.720 279.030 596.000 ;
        RECT 279.870 595.720 292.370 596.000 ;
        RECT 293.210 595.720 306.170 596.000 ;
        RECT 307.010 595.720 319.510 596.000 ;
        RECT 320.350 595.720 333.310 596.000 ;
        RECT 334.150 595.720 347.110 596.000 ;
        RECT 347.950 595.720 360.450 596.000 ;
        RECT 361.290 595.720 374.250 596.000 ;
        RECT 375.090 595.720 388.050 596.000 ;
        RECT 388.890 595.720 401.390 596.000 ;
        RECT 402.230 595.720 415.190 596.000 ;
        RECT 416.030 595.720 428.990 596.000 ;
        RECT 429.830 595.720 442.330 596.000 ;
        RECT 443.170 595.720 456.130 596.000 ;
        RECT 456.970 595.720 469.930 596.000 ;
        RECT 470.770 595.720 483.270 596.000 ;
        RECT 484.110 595.720 497.070 596.000 ;
        RECT 497.910 595.720 510.870 596.000 ;
        RECT 511.710 595.720 524.210 596.000 ;
        RECT 525.050 595.720 538.010 596.000 ;
        RECT 538.850 595.720 551.810 596.000 ;
        RECT 552.650 595.720 565.150 596.000 ;
        RECT 565.990 595.720 578.950 596.000 ;
        RECT 579.790 595.720 592.750 596.000 ;
        RECT 593.590 595.720 606.090 596.000 ;
        RECT 606.930 595.720 619.890 596.000 ;
        RECT 620.730 595.720 633.230 596.000 ;
        RECT 634.070 595.720 647.030 596.000 ;
        RECT 647.870 595.720 660.830 596.000 ;
        RECT 661.670 595.720 674.170 596.000 ;
        RECT 675.010 595.720 687.970 596.000 ;
        RECT 688.810 595.720 701.770 596.000 ;
        RECT 702.610 595.720 715.110 596.000 ;
        RECT 715.950 595.720 728.910 596.000 ;
        RECT 729.750 595.720 742.710 596.000 ;
        RECT 743.550 595.720 756.050 596.000 ;
        RECT 756.890 595.720 769.850 596.000 ;
        RECT 770.690 595.720 783.650 596.000 ;
        RECT 784.490 595.720 796.990 596.000 ;
        RECT 797.830 595.720 810.790 596.000 ;
        RECT 811.630 595.720 824.590 596.000 ;
        RECT 825.430 595.720 837.930 596.000 ;
        RECT 838.770 595.720 851.730 596.000 ;
        RECT 852.570 595.720 865.530 596.000 ;
        RECT 866.370 595.720 878.870 596.000 ;
        RECT 879.710 595.720 892.670 596.000 ;
        RECT 893.510 595.720 896.440 596.000 ;
        RECT 3.320 4.280 896.440 595.720 ;
        RECT 3.870 4.000 9.930 4.280 ;
        RECT 10.770 4.000 16.830 4.280 ;
        RECT 17.670 4.000 23.730 4.280 ;
        RECT 24.570 4.000 31.090 4.280 ;
        RECT 31.930 4.000 37.990 4.280 ;
        RECT 38.830 4.000 44.890 4.280 ;
        RECT 45.730 4.000 52.250 4.280 ;
        RECT 53.090 4.000 59.150 4.280 ;
        RECT 59.990 4.000 66.050 4.280 ;
        RECT 66.890 4.000 72.950 4.280 ;
        RECT 73.790 4.000 80.310 4.280 ;
        RECT 81.150 4.000 87.210 4.280 ;
        RECT 88.050 4.000 94.110 4.280 ;
        RECT 94.950 4.000 101.470 4.280 ;
        RECT 102.310 4.000 108.370 4.280 ;
        RECT 109.210 4.000 115.270 4.280 ;
        RECT 116.110 4.000 122.170 4.280 ;
        RECT 123.010 4.000 129.530 4.280 ;
        RECT 130.370 4.000 136.430 4.280 ;
        RECT 137.270 4.000 143.330 4.280 ;
        RECT 144.170 4.000 150.690 4.280 ;
        RECT 151.530 4.000 157.590 4.280 ;
        RECT 158.430 4.000 164.490 4.280 ;
        RECT 165.330 4.000 171.390 4.280 ;
        RECT 172.230 4.000 178.750 4.280 ;
        RECT 179.590 4.000 185.650 4.280 ;
        RECT 186.490 4.000 192.550 4.280 ;
        RECT 193.390 4.000 199.910 4.280 ;
        RECT 200.750 4.000 206.810 4.280 ;
        RECT 207.650 4.000 213.710 4.280 ;
        RECT 214.550 4.000 220.610 4.280 ;
        RECT 221.450 4.000 227.970 4.280 ;
        RECT 228.810 4.000 234.870 4.280 ;
        RECT 235.710 4.000 241.770 4.280 ;
        RECT 242.610 4.000 249.130 4.280 ;
        RECT 249.970 4.000 256.030 4.280 ;
        RECT 256.870 4.000 262.930 4.280 ;
        RECT 263.770 4.000 269.830 4.280 ;
        RECT 270.670 4.000 277.190 4.280 ;
        RECT 278.030 4.000 284.090 4.280 ;
        RECT 284.930 4.000 290.990 4.280 ;
        RECT 291.830 4.000 298.350 4.280 ;
        RECT 299.190 4.000 305.250 4.280 ;
        RECT 306.090 4.000 312.150 4.280 ;
        RECT 312.990 4.000 319.510 4.280 ;
        RECT 320.350 4.000 326.410 4.280 ;
        RECT 327.250 4.000 333.310 4.280 ;
        RECT 334.150 4.000 340.210 4.280 ;
        RECT 341.050 4.000 347.570 4.280 ;
        RECT 348.410 4.000 354.470 4.280 ;
        RECT 355.310 4.000 361.370 4.280 ;
        RECT 362.210 4.000 368.730 4.280 ;
        RECT 369.570 4.000 375.630 4.280 ;
        RECT 376.470 4.000 382.530 4.280 ;
        RECT 383.370 4.000 389.430 4.280 ;
        RECT 390.270 4.000 396.790 4.280 ;
        RECT 397.630 4.000 403.690 4.280 ;
        RECT 404.530 4.000 410.590 4.280 ;
        RECT 411.430 4.000 417.950 4.280 ;
        RECT 418.790 4.000 424.850 4.280 ;
        RECT 425.690 4.000 431.750 4.280 ;
        RECT 432.590 4.000 438.650 4.280 ;
        RECT 439.490 4.000 446.010 4.280 ;
        RECT 446.850 4.000 452.910 4.280 ;
        RECT 453.750 4.000 459.810 4.280 ;
        RECT 460.650 4.000 467.170 4.280 ;
        RECT 468.010 4.000 474.070 4.280 ;
        RECT 474.910 4.000 480.970 4.280 ;
        RECT 481.810 4.000 487.870 4.280 ;
        RECT 488.710 4.000 495.230 4.280 ;
        RECT 496.070 4.000 502.130 4.280 ;
        RECT 502.970 4.000 509.030 4.280 ;
        RECT 509.870 4.000 516.390 4.280 ;
        RECT 517.230 4.000 523.290 4.280 ;
        RECT 524.130 4.000 530.190 4.280 ;
        RECT 531.030 4.000 537.090 4.280 ;
        RECT 537.930 4.000 544.450 4.280 ;
        RECT 545.290 4.000 551.350 4.280 ;
        RECT 552.190 4.000 558.250 4.280 ;
        RECT 559.090 4.000 565.610 4.280 ;
        RECT 566.450 4.000 572.510 4.280 ;
        RECT 573.350 4.000 579.410 4.280 ;
        RECT 580.250 4.000 586.310 4.280 ;
        RECT 587.150 4.000 593.670 4.280 ;
        RECT 594.510 4.000 600.570 4.280 ;
        RECT 601.410 4.000 607.470 4.280 ;
        RECT 608.310 4.000 614.830 4.280 ;
        RECT 615.670 4.000 621.730 4.280 ;
        RECT 622.570 4.000 628.630 4.280 ;
        RECT 629.470 4.000 635.990 4.280 ;
        RECT 636.830 4.000 642.890 4.280 ;
        RECT 643.730 4.000 649.790 4.280 ;
        RECT 650.630 4.000 656.690 4.280 ;
        RECT 657.530 4.000 664.050 4.280 ;
        RECT 664.890 4.000 670.950 4.280 ;
        RECT 671.790 4.000 677.850 4.280 ;
        RECT 678.690 4.000 685.210 4.280 ;
        RECT 686.050 4.000 692.110 4.280 ;
        RECT 692.950 4.000 699.010 4.280 ;
        RECT 699.850 4.000 705.910 4.280 ;
        RECT 706.750 4.000 713.270 4.280 ;
        RECT 714.110 4.000 720.170 4.280 ;
        RECT 721.010 4.000 727.070 4.280 ;
        RECT 727.910 4.000 734.430 4.280 ;
        RECT 735.270 4.000 741.330 4.280 ;
        RECT 742.170 4.000 748.230 4.280 ;
        RECT 749.070 4.000 755.130 4.280 ;
        RECT 755.970 4.000 762.490 4.280 ;
        RECT 763.330 4.000 769.390 4.280 ;
        RECT 770.230 4.000 776.290 4.280 ;
        RECT 777.130 4.000 783.650 4.280 ;
        RECT 784.490 4.000 790.550 4.280 ;
        RECT 791.390 4.000 797.450 4.280 ;
        RECT 798.290 4.000 804.350 4.280 ;
        RECT 805.190 4.000 811.710 4.280 ;
        RECT 812.550 4.000 818.610 4.280 ;
        RECT 819.450 4.000 825.510 4.280 ;
        RECT 826.350 4.000 832.870 4.280 ;
        RECT 833.710 4.000 839.770 4.280 ;
        RECT 840.610 4.000 846.670 4.280 ;
        RECT 847.510 4.000 853.570 4.280 ;
        RECT 854.410 4.000 860.930 4.280 ;
        RECT 861.770 4.000 867.830 4.280 ;
        RECT 868.670 4.000 874.730 4.280 ;
        RECT 875.570 4.000 882.090 4.280 ;
        RECT 882.930 4.000 888.990 4.280 ;
        RECT 889.830 4.000 895.890 4.280 ;
      LAYER met3 ;
        RECT 4.400 593.960 895.600 594.825 ;
        RECT 4.000 585.840 896.000 593.960 ;
        RECT 4.400 584.440 895.600 585.840 ;
        RECT 4.000 576.320 896.000 584.440 ;
        RECT 4.400 574.920 895.600 576.320 ;
        RECT 4.000 566.800 896.000 574.920 ;
        RECT 4.400 565.400 895.600 566.800 ;
        RECT 4.000 557.960 896.000 565.400 ;
        RECT 4.400 556.560 895.600 557.960 ;
        RECT 4.000 548.440 896.000 556.560 ;
        RECT 4.400 547.040 895.600 548.440 ;
        RECT 4.000 538.920 896.000 547.040 ;
        RECT 4.400 537.520 895.600 538.920 ;
        RECT 4.000 529.400 896.000 537.520 ;
        RECT 4.400 528.000 895.600 529.400 ;
        RECT 4.000 519.880 896.000 528.000 ;
        RECT 4.400 518.480 895.600 519.880 ;
        RECT 4.000 511.040 896.000 518.480 ;
        RECT 4.400 509.640 895.600 511.040 ;
        RECT 4.000 501.520 896.000 509.640 ;
        RECT 4.400 500.120 895.600 501.520 ;
        RECT 4.000 492.000 896.000 500.120 ;
        RECT 4.400 490.600 895.600 492.000 ;
        RECT 4.000 482.480 896.000 490.600 ;
        RECT 4.400 481.080 895.600 482.480 ;
        RECT 4.000 473.640 896.000 481.080 ;
        RECT 4.400 472.240 895.600 473.640 ;
        RECT 4.000 464.120 896.000 472.240 ;
        RECT 4.400 462.720 895.600 464.120 ;
        RECT 4.000 454.600 896.000 462.720 ;
        RECT 4.400 453.200 895.600 454.600 ;
        RECT 4.000 445.080 896.000 453.200 ;
        RECT 4.400 443.680 895.600 445.080 ;
        RECT 4.000 435.560 896.000 443.680 ;
        RECT 4.400 434.160 895.600 435.560 ;
        RECT 4.000 426.720 896.000 434.160 ;
        RECT 4.400 425.320 895.600 426.720 ;
        RECT 4.000 417.200 896.000 425.320 ;
        RECT 4.400 415.800 895.600 417.200 ;
        RECT 4.000 407.680 896.000 415.800 ;
        RECT 4.400 406.280 895.600 407.680 ;
        RECT 4.000 398.160 896.000 406.280 ;
        RECT 4.400 396.760 895.600 398.160 ;
        RECT 4.000 389.320 896.000 396.760 ;
        RECT 4.400 387.920 895.600 389.320 ;
        RECT 4.000 379.800 896.000 387.920 ;
        RECT 4.400 378.400 895.600 379.800 ;
        RECT 4.000 370.280 896.000 378.400 ;
        RECT 4.400 368.880 895.600 370.280 ;
        RECT 4.000 360.760 896.000 368.880 ;
        RECT 4.400 359.360 895.600 360.760 ;
        RECT 4.000 351.240 896.000 359.360 ;
        RECT 4.400 349.840 895.600 351.240 ;
        RECT 4.000 342.400 896.000 349.840 ;
        RECT 4.400 341.000 895.600 342.400 ;
        RECT 4.000 332.880 896.000 341.000 ;
        RECT 4.400 331.480 895.600 332.880 ;
        RECT 4.000 323.360 896.000 331.480 ;
        RECT 4.400 321.960 895.600 323.360 ;
        RECT 4.000 313.840 896.000 321.960 ;
        RECT 4.400 312.440 895.600 313.840 ;
        RECT 4.000 305.000 896.000 312.440 ;
        RECT 4.400 303.600 895.600 305.000 ;
        RECT 4.000 295.480 896.000 303.600 ;
        RECT 4.400 294.080 895.600 295.480 ;
        RECT 4.000 285.960 896.000 294.080 ;
        RECT 4.400 284.560 895.600 285.960 ;
        RECT 4.000 276.440 896.000 284.560 ;
        RECT 4.400 275.040 895.600 276.440 ;
        RECT 4.000 266.920 896.000 275.040 ;
        RECT 4.400 265.520 895.600 266.920 ;
        RECT 4.000 258.080 896.000 265.520 ;
        RECT 4.400 256.680 895.600 258.080 ;
        RECT 4.000 248.560 896.000 256.680 ;
        RECT 4.400 247.160 895.600 248.560 ;
        RECT 4.000 239.040 896.000 247.160 ;
        RECT 4.400 237.640 895.600 239.040 ;
        RECT 4.000 229.520 896.000 237.640 ;
        RECT 4.400 228.120 895.600 229.520 ;
        RECT 4.000 220.000 896.000 228.120 ;
        RECT 4.400 218.600 895.600 220.000 ;
        RECT 4.000 211.160 896.000 218.600 ;
        RECT 4.400 209.760 895.600 211.160 ;
        RECT 4.000 201.640 896.000 209.760 ;
        RECT 4.400 200.240 895.600 201.640 ;
        RECT 4.000 192.120 896.000 200.240 ;
        RECT 4.400 190.720 895.600 192.120 ;
        RECT 4.000 182.600 896.000 190.720 ;
        RECT 4.400 181.200 895.600 182.600 ;
        RECT 4.000 173.760 896.000 181.200 ;
        RECT 4.400 172.360 895.600 173.760 ;
        RECT 4.000 164.240 896.000 172.360 ;
        RECT 4.400 162.840 895.600 164.240 ;
        RECT 4.000 154.720 896.000 162.840 ;
        RECT 4.400 153.320 895.600 154.720 ;
        RECT 4.000 145.200 896.000 153.320 ;
        RECT 4.400 143.800 895.600 145.200 ;
        RECT 4.000 135.680 896.000 143.800 ;
        RECT 4.400 134.280 895.600 135.680 ;
        RECT 4.000 126.840 896.000 134.280 ;
        RECT 4.400 125.440 895.600 126.840 ;
        RECT 4.000 117.320 896.000 125.440 ;
        RECT 4.400 115.920 895.600 117.320 ;
        RECT 4.000 107.800 896.000 115.920 ;
        RECT 4.400 106.400 895.600 107.800 ;
        RECT 4.000 98.280 896.000 106.400 ;
        RECT 4.400 96.880 895.600 98.280 ;
        RECT 4.000 89.440 896.000 96.880 ;
        RECT 4.400 88.040 895.600 89.440 ;
        RECT 4.000 79.920 896.000 88.040 ;
        RECT 4.400 78.520 895.600 79.920 ;
        RECT 4.000 70.400 896.000 78.520 ;
        RECT 4.400 69.000 895.600 70.400 ;
        RECT 4.000 60.880 896.000 69.000 ;
        RECT 4.400 59.480 895.600 60.880 ;
        RECT 4.000 51.360 896.000 59.480 ;
        RECT 4.400 49.960 895.600 51.360 ;
        RECT 4.000 42.520 896.000 49.960 ;
        RECT 4.400 41.120 895.600 42.520 ;
        RECT 4.000 33.000 896.000 41.120 ;
        RECT 4.400 31.600 895.600 33.000 ;
        RECT 4.000 23.480 896.000 31.600 ;
        RECT 4.400 22.080 895.600 23.480 ;
        RECT 4.000 13.960 896.000 22.080 ;
        RECT 4.400 12.560 895.600 13.960 ;
        RECT 4.000 5.120 896.000 12.560 ;
        RECT 4.400 4.255 895.600 5.120 ;
  END
END sin3
END LIBRARY

