VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_local
  CLASS BLOCK ;
  FOREIGN wb_local ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 600.000 ;
  PIN dsi[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 596.000 0.830 604.000 ;
    END
  END dsi[0]
  PIN dsi[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 596.000 1.750 604.000 ;
    END
  END dsi[1]
  PIN dsi[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 596.000 3.130 604.000 ;
    END
  END dsi[2]
  PIN dsi[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 596.000 4.050 604.000 ;
    END
  END dsi[3]
  PIN dsi[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 596.000 5.430 604.000 ;
    END
  END dsi[4]
  PIN dsi[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 596.000 6.350 604.000 ;
    END
  END dsi[5]
  PIN dsi[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 596.000 7.730 604.000 ;
    END
  END dsi[6]
  PIN dsi[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 596.000 8.650 604.000 ;
    END
  END dsi[7]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 596.000 10.030 604.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 596.000 44.530 604.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 596.000 48.210 604.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 596.000 51.430 604.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 596.000 55.110 604.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 596.000 58.330 604.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 596.000 62.010 604.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 596.000 65.230 604.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 596.000 68.910 604.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 596.000 72.130 604.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 596.000 75.810 604.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 596.000 13.250 604.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 596.000 79.030 604.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 596.000 82.710 604.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 596.000 86.390 604.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 596.000 89.610 604.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 596.000 93.290 604.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 596.000 96.510 604.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 596.000 100.190 604.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 596.000 103.410 604.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 596.000 107.090 604.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 596.000 110.310 604.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 596.000 16.930 604.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 596.000 113.990 604.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 596.000 117.210 604.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 596.000 120.890 604.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 596.000 124.570 604.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 596.000 127.790 604.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 596.000 131.470 604.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 596.000 134.690 604.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 596.000 138.370 604.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 596.000 20.150 604.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 596.000 23.830 604.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 596.000 27.050 604.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 596.000 30.730 604.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 596.000 33.950 604.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 596.000 37.630 604.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 596.000 41.310 604.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 596.000 10.950 604.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 596.000 45.910 604.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 596.000 49.130 604.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 596.000 52.810 604.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 596.000 56.030 604.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 596.000 59.710 604.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 596.000 62.930 604.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 596.000 66.610 604.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 596.000 69.830 604.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 596.000 73.510 604.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 596.000 76.730 604.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 596.000 14.630 604.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 596.000 80.410 604.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 596.000 84.090 604.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 596.000 87.310 604.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 596.000 90.990 604.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 596.000 94.210 604.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 596.000 97.890 604.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 596.000 101.110 604.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 596.000 104.790 604.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 596.000 108.010 604.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 596.000 111.690 604.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 596.000 17.850 604.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 596.000 114.910 604.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 596.000 118.590 604.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 596.000 122.270 604.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 596.000 125.490 604.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 596.000 129.170 604.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 596.000 132.390 604.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 596.000 136.070 604.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 596.000 139.290 604.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 596.000 21.530 604.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 596.000 24.750 604.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 596.000 28.430 604.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 596.000 31.650 604.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 596.000 35.330 604.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 596.000 38.550 604.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 596.000 42.230 604.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 596.000 12.330 604.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 596.000 46.830 604.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 596.000 50.510 604.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 596.000 53.730 604.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 596.000 57.410 604.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 596.000 60.630 604.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 596.000 64.310 604.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 596.000 67.530 604.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 596.000 71.210 604.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 596.000 74.430 604.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 596.000 78.110 604.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 596.000 15.550 604.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 596.000 81.790 604.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 596.000 85.010 604.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 596.000 88.690 604.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 596.000 91.910 604.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 596.000 95.590 604.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 596.000 98.810 604.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 596.000 102.490 604.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 596.000 105.710 604.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 596.000 109.390 604.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 596.000 112.610 604.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 596.000 19.230 604.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 596.000 116.290 604.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 596.000 119.510 604.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 596.000 123.190 604.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 596.000 126.870 604.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 596.000 130.090 604.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 596.000 133.770 604.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 596.000 136.990 604.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 596.000 140.670 604.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 596.000 22.450 604.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 596.000 26.130 604.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 596.000 29.350 604.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 596.000 33.030 604.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 596.000 36.250 604.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 596.000 39.930 604.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 596.000 43.610 604.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 -4.000 4.050 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 -4.000 5.430 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 -4.000 7.270 4.000 ;
    END
  END irq[2]
  PIN m_irqs[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 596.000 159.990 604.000 ;
    END
  END m_irqs[0]
  PIN m_irqs[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 596.000 171.950 604.000 ;
    END
  END m_irqs[10]
  PIN m_irqs[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 596.000 172.870 604.000 ;
    END
  END m_irqs[11]
  PIN m_irqs[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 596.000 161.370 604.000 ;
    END
  END m_irqs[1]
  PIN m_irqs[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 596.000 162.750 604.000 ;
    END
  END m_irqs[2]
  PIN m_irqs[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 596.000 163.670 604.000 ;
    END
  END m_irqs[3]
  PIN m_irqs[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 596.000 165.050 604.000 ;
    END
  END m_irqs[4]
  PIN m_irqs[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 596.000 165.970 604.000 ;
    END
  END m_irqs[5]
  PIN m_irqs[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 596.000 167.350 604.000 ;
    END
  END m_irqs[6]
  PIN m_irqs[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 596.000 168.270 604.000 ;
    END
  END m_irqs[7]
  PIN m_irqs[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 596.000 169.650 604.000 ;
    END
  END m_irqs[8]
  PIN m_irqs[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 596.000 170.570 604.000 ;
    END
  END m_irqs[9]
  PIN m_wb_clk_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 -4.000 177.930 4.000 ;
    END
  END m_wb_clk_i
  PIN m_wb_rst_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 596.000 174.250 604.000 ;
    END
  END m_wb_rst_i
  PIN m_wbs_ack_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 -4.000 179.770 4.000 ;
    END
  END m_wbs_ack_o[0]
  PIN m_wbs_ack_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 568.520 4.000 569.120 ;
    END
  END m_wbs_ack_o[10]
  PIN m_wbs_ack_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 596.000 192.650 604.000 ;
    END
  END m_wbs_ack_o[11]
  PIN m_wbs_ack_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 520.920 4.000 521.520 ;
    END
  END m_wbs_ack_o[1]
  PIN m_wbs_ack_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 529.080 4.000 529.680 ;
    END
  END m_wbs_ack_o[2]
  PIN m_wbs_ack_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 596.000 177.470 604.000 ;
    END
  END m_wbs_ack_o[3]
  PIN m_wbs_ack_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 544.720 4.000 545.320 ;
    END
  END m_wbs_ack_o[4]
  PIN m_wbs_ack_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 596.000 182.070 604.000 ;
    END
  END m_wbs_ack_o[5]
  PIN m_wbs_ack_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 596.000 185.750 604.000 ;
    END
  END m_wbs_ack_o[6]
  PIN m_wbs_ack_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 596.000 188.050 604.000 ;
    END
  END m_wbs_ack_o[7]
  PIN m_wbs_ack_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 580.080 204.000 580.680 ;
    END
  END m_wbs_ack_o[8]
  PIN m_wbs_ack_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 -4.000 187.590 4.000 ;
    END
  END m_wbs_ack_o[9]
  PIN m_wbs_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 516.840 4.000 517.440 ;
    END
  END m_wbs_adr_i[0]
  PIN m_wbs_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 572.600 4.000 573.200 ;
    END
  END m_wbs_adr_i[10]
  PIN m_wbs_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 -4.000 190.810 4.000 ;
    END
  END m_wbs_adr_i[11]
  PIN m_wbs_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 -4.000 182.990 4.000 ;
    END
  END m_wbs_adr_i[1]
  PIN m_wbs_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 533.160 4.000 533.760 ;
    END
  END m_wbs_adr_i[2]
  PIN m_wbs_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 540.640 4.000 541.240 ;
    END
  END m_wbs_adr_i[3]
  PIN m_wbs_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 548.800 4.000 549.400 ;
    END
  END m_wbs_adr_i[4]
  PIN m_wbs_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 596.000 183.450 604.000 ;
    END
  END m_wbs_adr_i[5]
  PIN m_wbs_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 552.880 4.000 553.480 ;
    END
  END m_wbs_adr_i[6]
  PIN m_wbs_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 575.320 204.000 575.920 ;
    END
  END m_wbs_adr_i[7]
  PIN m_wbs_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 596.000 190.350 604.000 ;
    END
  END m_wbs_adr_i[8]
  PIN m_wbs_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 565.120 4.000 565.720 ;
    END
  END m_wbs_adr_i[9]
  PIN m_wbs_cs_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 -4.000 181.150 4.000 ;
    END
  END m_wbs_cs_i[0]
  PIN m_wbs_cs_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 596.000 191.270 604.000 ;
    END
  END m_wbs_cs_i[10]
  PIN m_wbs_cs_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 -4.000 192.650 4.000 ;
    END
  END m_wbs_cs_i[11]
  PIN m_wbs_cs_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 596.000 176.550 604.000 ;
    END
  END m_wbs_cs_i[1]
  PIN m_wbs_cs_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 573.280 204.000 573.880 ;
    END
  END m_wbs_cs_i[2]
  PIN m_wbs_cs_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 596.000 178.850 604.000 ;
    END
  END m_wbs_cs_i[3]
  PIN m_wbs_cs_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 596.000 181.150 604.000 ;
    END
  END m_wbs_cs_i[4]
  PIN m_wbs_cs_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 596.000 184.370 604.000 ;
    END
  END m_wbs_cs_i[5]
  PIN m_wbs_cs_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 596.000 186.670 604.000 ;
    END
  END m_wbs_cs_i[6]
  PIN m_wbs_cs_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 596.000 188.970 604.000 ;
    END
  END m_wbs_cs_i[7]
  PIN m_wbs_cs_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 582.120 204.000 582.720 ;
    END
  END m_wbs_cs_i[8]
  PIN m_wbs_cs_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 584.160 204.000 584.760 ;
    END
  END m_wbs_cs_i[9]
  PIN m_wbs_dat_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 596.000 175.170 604.000 ;
    END
  END m_wbs_dat_i[0]
  PIN m_wbs_dat_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 -4.000 189.430 4.000 ;
    END
  END m_wbs_dat_i[10]
  PIN m_wbs_dat_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 576.680 4.000 577.280 ;
    END
  END m_wbs_dat_i[11]
  PIN m_wbs_dat_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 596.000 193.570 604.000 ;
    END
  END m_wbs_dat_i[12]
  PIN m_wbs_dat_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 588.920 204.000 589.520 ;
    END
  END m_wbs_dat_i[13]
  PIN m_wbs_dat_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 580.760 4.000 581.360 ;
    END
  END m_wbs_dat_i[14]
  PIN m_wbs_dat_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 596.000 194.950 604.000 ;
    END
  END m_wbs_dat_i[15]
  PIN m_wbs_dat_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 584.840 4.000 585.440 ;
    END
  END m_wbs_dat_i[16]
  PIN m_wbs_dat_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 590.960 204.000 591.560 ;
    END
  END m_wbs_dat_i[17]
  PIN m_wbs_dat_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 593.680 204.000 594.280 ;
    END
  END m_wbs_dat_i[18]
  PIN m_wbs_dat_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 -4.000 194.030 4.000 ;
    END
  END m_wbs_dat_i[19]
  PIN m_wbs_dat_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 525.000 4.000 525.600 ;
    END
  END m_wbs_dat_i[1]
  PIN m_wbs_dat_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 -4.000 195.870 4.000 ;
    END
  END m_wbs_dat_i[20]
  PIN m_wbs_dat_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 596.000 195.870 604.000 ;
    END
  END m_wbs_dat_i[21]
  PIN m_wbs_dat_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 588.920 4.000 589.520 ;
    END
  END m_wbs_dat_i[22]
  PIN m_wbs_dat_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 596.000 197.250 604.000 ;
    END
  END m_wbs_dat_i[23]
  PIN m_wbs_dat_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 596.000 198.170 604.000 ;
    END
  END m_wbs_dat_i[24]
  PIN m_wbs_dat_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 -4.000 197.250 4.000 ;
    END
  END m_wbs_dat_i[25]
  PIN m_wbs_dat_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 593.000 4.000 593.600 ;
    END
  END m_wbs_dat_i[26]
  PIN m_wbs_dat_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 597.080 4.000 597.680 ;
    END
  END m_wbs_dat_i[27]
  PIN m_wbs_dat_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 -4.000 199.090 4.000 ;
    END
  END m_wbs_dat_i[28]
  PIN m_wbs_dat_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 595.720 204.000 596.320 ;
    END
  END m_wbs_dat_i[29]
  PIN m_wbs_dat_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 536.560 4.000 537.160 ;
    END
  END m_wbs_dat_i[2]
  PIN m_wbs_dat_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 597.760 204.000 598.360 ;
    END
  END m_wbs_dat_i[30]
  PIN m_wbs_dat_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 596.000 199.550 604.000 ;
    END
  END m_wbs_dat_i[31]
  PIN m_wbs_dat_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 596.000 179.770 604.000 ;
    END
  END m_wbs_dat_i[3]
  PIN m_wbs_dat_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 -4.000 184.370 4.000 ;
    END
  END m_wbs_dat_i[4]
  PIN m_wbs_dat_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 -4.000 186.210 4.000 ;
    END
  END m_wbs_dat_i[5]
  PIN m_wbs_dat_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 556.960 4.000 557.560 ;
    END
  END m_wbs_dat_i[6]
  PIN m_wbs_dat_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 578.040 204.000 578.640 ;
    END
  END m_wbs_dat_i[7]
  PIN m_wbs_dat_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 561.040 4.000 561.640 ;
    END
  END m_wbs_dat_i[8]
  PIN m_wbs_dat_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 586.880 204.000 587.480 ;
    END
  END m_wbs_dat_i[9]
  PIN m_wbs_dat_o_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 0.720 204.000 1.320 ;
    END
  END m_wbs_dat_o_0[0]
  PIN m_wbs_dat_o_0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 22.480 204.000 23.080 ;
    END
  END m_wbs_dat_o_0[10]
  PIN m_wbs_dat_o_0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 25.200 204.000 25.800 ;
    END
  END m_wbs_dat_o_0[11]
  PIN m_wbs_dat_o_0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 27.240 204.000 27.840 ;
    END
  END m_wbs_dat_o_0[12]
  PIN m_wbs_dat_o_0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 29.280 204.000 29.880 ;
    END
  END m_wbs_dat_o_0[13]
  PIN m_wbs_dat_o_0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 32.000 204.000 32.600 ;
    END
  END m_wbs_dat_o_0[14]
  PIN m_wbs_dat_o_0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 34.040 204.000 34.640 ;
    END
  END m_wbs_dat_o_0[15]
  PIN m_wbs_dat_o_0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 36.080 204.000 36.680 ;
    END
  END m_wbs_dat_o_0[16]
  PIN m_wbs_dat_o_0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 38.120 204.000 38.720 ;
    END
  END m_wbs_dat_o_0[17]
  PIN m_wbs_dat_o_0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 40.840 204.000 41.440 ;
    END
  END m_wbs_dat_o_0[18]
  PIN m_wbs_dat_o_0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 42.880 204.000 43.480 ;
    END
  END m_wbs_dat_o_0[19]
  PIN m_wbs_dat_o_0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2.760 204.000 3.360 ;
    END
  END m_wbs_dat_o_0[1]
  PIN m_wbs_dat_o_0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 44.920 204.000 45.520 ;
    END
  END m_wbs_dat_o_0[20]
  PIN m_wbs_dat_o_0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 47.640 204.000 48.240 ;
    END
  END m_wbs_dat_o_0[21]
  PIN m_wbs_dat_o_0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 49.680 204.000 50.280 ;
    END
  END m_wbs_dat_o_0[22]
  PIN m_wbs_dat_o_0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 51.720 204.000 52.320 ;
    END
  END m_wbs_dat_o_0[23]
  PIN m_wbs_dat_o_0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 53.760 204.000 54.360 ;
    END
  END m_wbs_dat_o_0[24]
  PIN m_wbs_dat_o_0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 56.480 204.000 57.080 ;
    END
  END m_wbs_dat_o_0[25]
  PIN m_wbs_dat_o_0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 58.520 204.000 59.120 ;
    END
  END m_wbs_dat_o_0[26]
  PIN m_wbs_dat_o_0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 60.560 204.000 61.160 ;
    END
  END m_wbs_dat_o_0[27]
  PIN m_wbs_dat_o_0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 63.280 204.000 63.880 ;
    END
  END m_wbs_dat_o_0[28]
  PIN m_wbs_dat_o_0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 65.320 204.000 65.920 ;
    END
  END m_wbs_dat_o_0[29]
  PIN m_wbs_dat_o_0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 4.800 204.000 5.400 ;
    END
  END m_wbs_dat_o_0[2]
  PIN m_wbs_dat_o_0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 67.360 204.000 67.960 ;
    END
  END m_wbs_dat_o_0[30]
  PIN m_wbs_dat_o_0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 70.080 204.000 70.680 ;
    END
  END m_wbs_dat_o_0[31]
  PIN m_wbs_dat_o_0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 6.840 204.000 7.440 ;
    END
  END m_wbs_dat_o_0[3]
  PIN m_wbs_dat_o_0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 9.560 204.000 10.160 ;
    END
  END m_wbs_dat_o_0[4]
  PIN m_wbs_dat_o_0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 11.600 204.000 12.200 ;
    END
  END m_wbs_dat_o_0[5]
  PIN m_wbs_dat_o_0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 13.640 204.000 14.240 ;
    END
  END m_wbs_dat_o_0[6]
  PIN m_wbs_dat_o_0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 16.360 204.000 16.960 ;
    END
  END m_wbs_dat_o_0[7]
  PIN m_wbs_dat_o_0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 18.400 204.000 19.000 ;
    END
  END m_wbs_dat_o_0[8]
  PIN m_wbs_dat_o_0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 20.440 204.000 21.040 ;
    END
  END m_wbs_dat_o_0[9]
  PIN m_wbs_dat_o_10[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 74.160 204.000 74.760 ;
    END
  END m_wbs_dat_o_10[0]
  PIN m_wbs_dat_o_10[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 141.480 204.000 142.080 ;
    END
  END m_wbs_dat_o_10[10]
  PIN m_wbs_dat_o_10[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 148.280 204.000 148.880 ;
    END
  END m_wbs_dat_o_10[11]
  PIN m_wbs_dat_o_10[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 155.080 204.000 155.680 ;
    END
  END m_wbs_dat_o_10[12]
  PIN m_wbs_dat_o_10[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 161.200 204.000 161.800 ;
    END
  END m_wbs_dat_o_10[13]
  PIN m_wbs_dat_o_10[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 168.000 204.000 168.600 ;
    END
  END m_wbs_dat_o_10[14]
  PIN m_wbs_dat_o_10[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 174.800 204.000 175.400 ;
    END
  END m_wbs_dat_o_10[15]
  PIN m_wbs_dat_o_10[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 181.600 204.000 182.200 ;
    END
  END m_wbs_dat_o_10[16]
  PIN m_wbs_dat_o_10[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 188.400 204.000 189.000 ;
    END
  END m_wbs_dat_o_10[17]
  PIN m_wbs_dat_o_10[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 195.200 204.000 195.800 ;
    END
  END m_wbs_dat_o_10[18]
  PIN m_wbs_dat_o_10[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 202.000 204.000 202.600 ;
    END
  END m_wbs_dat_o_10[19]
  PIN m_wbs_dat_o_10[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 80.960 204.000 81.560 ;
    END
  END m_wbs_dat_o_10[1]
  PIN m_wbs_dat_o_10[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 208.800 204.000 209.400 ;
    END
  END m_wbs_dat_o_10[20]
  PIN m_wbs_dat_o_10[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 214.920 204.000 215.520 ;
    END
  END m_wbs_dat_o_10[21]
  PIN m_wbs_dat_o_10[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 221.720 204.000 222.320 ;
    END
  END m_wbs_dat_o_10[22]
  PIN m_wbs_dat_o_10[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 228.520 204.000 229.120 ;
    END
  END m_wbs_dat_o_10[23]
  PIN m_wbs_dat_o_10[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 235.320 204.000 235.920 ;
    END
  END m_wbs_dat_o_10[24]
  PIN m_wbs_dat_o_10[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 242.120 204.000 242.720 ;
    END
  END m_wbs_dat_o_10[25]
  PIN m_wbs_dat_o_10[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 248.920 204.000 249.520 ;
    END
  END m_wbs_dat_o_10[26]
  PIN m_wbs_dat_o_10[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 255.720 204.000 256.320 ;
    END
  END m_wbs_dat_o_10[27]
  PIN m_wbs_dat_o_10[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 262.520 204.000 263.120 ;
    END
  END m_wbs_dat_o_10[28]
  PIN m_wbs_dat_o_10[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 268.640 204.000 269.240 ;
    END
  END m_wbs_dat_o_10[29]
  PIN m_wbs_dat_o_10[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 87.760 204.000 88.360 ;
    END
  END m_wbs_dat_o_10[2]
  PIN m_wbs_dat_o_10[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 275.440 204.000 276.040 ;
    END
  END m_wbs_dat_o_10[30]
  PIN m_wbs_dat_o_10[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 282.240 204.000 282.840 ;
    END
  END m_wbs_dat_o_10[31]
  PIN m_wbs_dat_o_10[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 94.560 204.000 95.160 ;
    END
  END m_wbs_dat_o_10[3]
  PIN m_wbs_dat_o_10[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 101.360 204.000 101.960 ;
    END
  END m_wbs_dat_o_10[4]
  PIN m_wbs_dat_o_10[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 107.480 204.000 108.080 ;
    END
  END m_wbs_dat_o_10[5]
  PIN m_wbs_dat_o_10[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 114.280 204.000 114.880 ;
    END
  END m_wbs_dat_o_10[6]
  PIN m_wbs_dat_o_10[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 121.080 204.000 121.680 ;
    END
  END m_wbs_dat_o_10[7]
  PIN m_wbs_dat_o_10[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 127.880 204.000 128.480 ;
    END
  END m_wbs_dat_o_10[8]
  PIN m_wbs_dat_o_10[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 134.680 204.000 135.280 ;
    END
  END m_wbs_dat_o_10[9]
  PIN m_wbs_dat_o_11[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 76.200 204.000 76.800 ;
    END
  END m_wbs_dat_o_11[0]
  PIN m_wbs_dat_o_11[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 143.520 204.000 144.120 ;
    END
  END m_wbs_dat_o_11[10]
  PIN m_wbs_dat_o_11[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 150.320 204.000 150.920 ;
    END
  END m_wbs_dat_o_11[11]
  PIN m_wbs_dat_o_11[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 157.120 204.000 157.720 ;
    END
  END m_wbs_dat_o_11[12]
  PIN m_wbs_dat_o_11[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 163.920 204.000 164.520 ;
    END
  END m_wbs_dat_o_11[13]
  PIN m_wbs_dat_o_11[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 170.720 204.000 171.320 ;
    END
  END m_wbs_dat_o_11[14]
  PIN m_wbs_dat_o_11[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 176.840 204.000 177.440 ;
    END
  END m_wbs_dat_o_11[15]
  PIN m_wbs_dat_o_11[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 183.640 204.000 184.240 ;
    END
  END m_wbs_dat_o_11[16]
  PIN m_wbs_dat_o_11[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 190.440 204.000 191.040 ;
    END
  END m_wbs_dat_o_11[17]
  PIN m_wbs_dat_o_11[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 197.240 204.000 197.840 ;
    END
  END m_wbs_dat_o_11[18]
  PIN m_wbs_dat_o_11[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 204.040 204.000 204.640 ;
    END
  END m_wbs_dat_o_11[19]
  PIN m_wbs_dat_o_11[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 83.000 204.000 83.600 ;
    END
  END m_wbs_dat_o_11[1]
  PIN m_wbs_dat_o_11[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 210.840 204.000 211.440 ;
    END
  END m_wbs_dat_o_11[20]
  PIN m_wbs_dat_o_11[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 217.640 204.000 218.240 ;
    END
  END m_wbs_dat_o_11[21]
  PIN m_wbs_dat_o_11[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 224.440 204.000 225.040 ;
    END
  END m_wbs_dat_o_11[22]
  PIN m_wbs_dat_o_11[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 230.560 204.000 231.160 ;
    END
  END m_wbs_dat_o_11[23]
  PIN m_wbs_dat_o_11[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 237.360 204.000 237.960 ;
    END
  END m_wbs_dat_o_11[24]
  PIN m_wbs_dat_o_11[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 244.160 204.000 244.760 ;
    END
  END m_wbs_dat_o_11[25]
  PIN m_wbs_dat_o_11[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 250.960 204.000 251.560 ;
    END
  END m_wbs_dat_o_11[26]
  PIN m_wbs_dat_o_11[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 257.760 204.000 258.360 ;
    END
  END m_wbs_dat_o_11[27]
  PIN m_wbs_dat_o_11[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 264.560 204.000 265.160 ;
    END
  END m_wbs_dat_o_11[28]
  PIN m_wbs_dat_o_11[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 271.360 204.000 271.960 ;
    END
  END m_wbs_dat_o_11[29]
  PIN m_wbs_dat_o_11[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 89.800 204.000 90.400 ;
    END
  END m_wbs_dat_o_11[2]
  PIN m_wbs_dat_o_11[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 278.160 204.000 278.760 ;
    END
  END m_wbs_dat_o_11[30]
  PIN m_wbs_dat_o_11[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 284.280 204.000 284.880 ;
    END
  END m_wbs_dat_o_11[31]
  PIN m_wbs_dat_o_11[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 96.600 204.000 97.200 ;
    END
  END m_wbs_dat_o_11[3]
  PIN m_wbs_dat_o_11[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 103.400 204.000 104.000 ;
    END
  END m_wbs_dat_o_11[4]
  PIN m_wbs_dat_o_11[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 110.200 204.000 110.800 ;
    END
  END m_wbs_dat_o_11[5]
  PIN m_wbs_dat_o_11[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 117.000 204.000 117.600 ;
    END
  END m_wbs_dat_o_11[6]
  PIN m_wbs_dat_o_11[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 123.800 204.000 124.400 ;
    END
  END m_wbs_dat_o_11[7]
  PIN m_wbs_dat_o_11[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 129.920 204.000 130.520 ;
    END
  END m_wbs_dat_o_11[8]
  PIN m_wbs_dat_o_11[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 136.720 204.000 137.320 ;
    END
  END m_wbs_dat_o_11[9]
  PIN m_wbs_dat_o_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 72.120 204.000 72.720 ;
    END
  END m_wbs_dat_o_1[0]
  PIN m_wbs_dat_o_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 139.440 204.000 140.040 ;
    END
  END m_wbs_dat_o_1[10]
  PIN m_wbs_dat_o_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 145.560 204.000 146.160 ;
    END
  END m_wbs_dat_o_1[11]
  PIN m_wbs_dat_o_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 152.360 204.000 152.960 ;
    END
  END m_wbs_dat_o_1[12]
  PIN m_wbs_dat_o_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 159.160 204.000 159.760 ;
    END
  END m_wbs_dat_o_1[13]
  PIN m_wbs_dat_o_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 165.960 204.000 166.560 ;
    END
  END m_wbs_dat_o_1[14]
  PIN m_wbs_dat_o_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 172.760 204.000 173.360 ;
    END
  END m_wbs_dat_o_1[15]
  PIN m_wbs_dat_o_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 179.560 204.000 180.160 ;
    END
  END m_wbs_dat_o_1[16]
  PIN m_wbs_dat_o_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 186.360 204.000 186.960 ;
    END
  END m_wbs_dat_o_1[17]
  PIN m_wbs_dat_o_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 193.160 204.000 193.760 ;
    END
  END m_wbs_dat_o_1[18]
  PIN m_wbs_dat_o_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 199.280 204.000 199.880 ;
    END
  END m_wbs_dat_o_1[19]
  PIN m_wbs_dat_o_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 78.920 204.000 79.520 ;
    END
  END m_wbs_dat_o_1[1]
  PIN m_wbs_dat_o_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 206.080 204.000 206.680 ;
    END
  END m_wbs_dat_o_1[20]
  PIN m_wbs_dat_o_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 212.880 204.000 213.480 ;
    END
  END m_wbs_dat_o_1[21]
  PIN m_wbs_dat_o_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 219.680 204.000 220.280 ;
    END
  END m_wbs_dat_o_1[22]
  PIN m_wbs_dat_o_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 226.480 204.000 227.080 ;
    END
  END m_wbs_dat_o_1[23]
  PIN m_wbs_dat_o_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 233.280 204.000 233.880 ;
    END
  END m_wbs_dat_o_1[24]
  PIN m_wbs_dat_o_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 240.080 204.000 240.680 ;
    END
  END m_wbs_dat_o_1[25]
  PIN m_wbs_dat_o_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 246.880 204.000 247.480 ;
    END
  END m_wbs_dat_o_1[26]
  PIN m_wbs_dat_o_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 253.000 204.000 253.600 ;
    END
  END m_wbs_dat_o_1[27]
  PIN m_wbs_dat_o_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 259.800 204.000 260.400 ;
    END
  END m_wbs_dat_o_1[28]
  PIN m_wbs_dat_o_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 266.600 204.000 267.200 ;
    END
  END m_wbs_dat_o_1[29]
  PIN m_wbs_dat_o_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 85.720 204.000 86.320 ;
    END
  END m_wbs_dat_o_1[2]
  PIN m_wbs_dat_o_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 273.400 204.000 274.000 ;
    END
  END m_wbs_dat_o_1[30]
  PIN m_wbs_dat_o_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 280.200 204.000 280.800 ;
    END
  END m_wbs_dat_o_1[31]
  PIN m_wbs_dat_o_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 91.840 204.000 92.440 ;
    END
  END m_wbs_dat_o_1[3]
  PIN m_wbs_dat_o_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 98.640 204.000 99.240 ;
    END
  END m_wbs_dat_o_1[4]
  PIN m_wbs_dat_o_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 105.440 204.000 106.040 ;
    END
  END m_wbs_dat_o_1[5]
  PIN m_wbs_dat_o_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 112.240 204.000 112.840 ;
    END
  END m_wbs_dat_o_1[6]
  PIN m_wbs_dat_o_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 119.040 204.000 119.640 ;
    END
  END m_wbs_dat_o_1[7]
  PIN m_wbs_dat_o_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 125.840 204.000 126.440 ;
    END
  END m_wbs_dat_o_1[8]
  PIN m_wbs_dat_o_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 132.640 204.000 133.240 ;
    END
  END m_wbs_dat_o_1[9]
  PIN m_wbs_dat_o_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 287.000 204.000 287.600 ;
    END
  END m_wbs_dat_o_2[0]
  PIN m_wbs_dat_o_2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 309.440 204.000 310.040 ;
    END
  END m_wbs_dat_o_2[10]
  PIN m_wbs_dat_o_2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 311.480 204.000 312.080 ;
    END
  END m_wbs_dat_o_2[11]
  PIN m_wbs_dat_o_2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 313.520 204.000 314.120 ;
    END
  END m_wbs_dat_o_2[12]
  PIN m_wbs_dat_o_2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 316.240 204.000 316.840 ;
    END
  END m_wbs_dat_o_2[13]
  PIN m_wbs_dat_o_2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 318.280 204.000 318.880 ;
    END
  END m_wbs_dat_o_2[14]
  PIN m_wbs_dat_o_2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 320.320 204.000 320.920 ;
    END
  END m_wbs_dat_o_2[15]
  PIN m_wbs_dat_o_2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 322.360 204.000 322.960 ;
    END
  END m_wbs_dat_o_2[16]
  PIN m_wbs_dat_o_2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 325.080 204.000 325.680 ;
    END
  END m_wbs_dat_o_2[17]
  PIN m_wbs_dat_o_2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 327.120 204.000 327.720 ;
    END
  END m_wbs_dat_o_2[18]
  PIN m_wbs_dat_o_2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 329.160 204.000 329.760 ;
    END
  END m_wbs_dat_o_2[19]
  PIN m_wbs_dat_o_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 289.040 204.000 289.640 ;
    END
  END m_wbs_dat_o_2[1]
  PIN m_wbs_dat_o_2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 331.880 204.000 332.480 ;
    END
  END m_wbs_dat_o_2[20]
  PIN m_wbs_dat_o_2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 333.920 204.000 334.520 ;
    END
  END m_wbs_dat_o_2[21]
  PIN m_wbs_dat_o_2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 335.960 204.000 336.560 ;
    END
  END m_wbs_dat_o_2[22]
  PIN m_wbs_dat_o_2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 338.000 204.000 338.600 ;
    END
  END m_wbs_dat_o_2[23]
  PIN m_wbs_dat_o_2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 340.720 204.000 341.320 ;
    END
  END m_wbs_dat_o_2[24]
  PIN m_wbs_dat_o_2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 342.760 204.000 343.360 ;
    END
  END m_wbs_dat_o_2[25]
  PIN m_wbs_dat_o_2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 344.800 204.000 345.400 ;
    END
  END m_wbs_dat_o_2[26]
  PIN m_wbs_dat_o_2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 347.520 204.000 348.120 ;
    END
  END m_wbs_dat_o_2[27]
  PIN m_wbs_dat_o_2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 349.560 204.000 350.160 ;
    END
  END m_wbs_dat_o_2[28]
  PIN m_wbs_dat_o_2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 351.600 204.000 352.200 ;
    END
  END m_wbs_dat_o_2[29]
  PIN m_wbs_dat_o_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 291.080 204.000 291.680 ;
    END
  END m_wbs_dat_o_2[2]
  PIN m_wbs_dat_o_2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 353.640 204.000 354.240 ;
    END
  END m_wbs_dat_o_2[30]
  PIN m_wbs_dat_o_2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 356.360 204.000 356.960 ;
    END
  END m_wbs_dat_o_2[31]
  PIN m_wbs_dat_o_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 293.800 204.000 294.400 ;
    END
  END m_wbs_dat_o_2[3]
  PIN m_wbs_dat_o_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 295.840 204.000 296.440 ;
    END
  END m_wbs_dat_o_2[4]
  PIN m_wbs_dat_o_2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 297.880 204.000 298.480 ;
    END
  END m_wbs_dat_o_2[5]
  PIN m_wbs_dat_o_2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 300.600 204.000 301.200 ;
    END
  END m_wbs_dat_o_2[6]
  PIN m_wbs_dat_o_2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 302.640 204.000 303.240 ;
    END
  END m_wbs_dat_o_2[7]
  PIN m_wbs_dat_o_2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 304.680 204.000 305.280 ;
    END
  END m_wbs_dat_o_2[8]
  PIN m_wbs_dat_o_2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 306.720 204.000 307.320 ;
    END
  END m_wbs_dat_o_2[9]
  PIN m_wbs_dat_o_3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 358.400 204.000 359.000 ;
    END
  END m_wbs_dat_o_3[0]
  PIN m_wbs_dat_o_3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 380.840 204.000 381.440 ;
    END
  END m_wbs_dat_o_3[10]
  PIN m_wbs_dat_o_3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 382.880 204.000 383.480 ;
    END
  END m_wbs_dat_o_3[11]
  PIN m_wbs_dat_o_3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 385.600 204.000 386.200 ;
    END
  END m_wbs_dat_o_3[12]
  PIN m_wbs_dat_o_3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 387.640 204.000 388.240 ;
    END
  END m_wbs_dat_o_3[13]
  PIN m_wbs_dat_o_3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 389.680 204.000 390.280 ;
    END
  END m_wbs_dat_o_3[14]
  PIN m_wbs_dat_o_3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 391.720 204.000 392.320 ;
    END
  END m_wbs_dat_o_3[15]
  PIN m_wbs_dat_o_3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 394.440 204.000 395.040 ;
    END
  END m_wbs_dat_o_3[16]
  PIN m_wbs_dat_o_3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 396.480 204.000 397.080 ;
    END
  END m_wbs_dat_o_3[17]
  PIN m_wbs_dat_o_3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 398.520 204.000 399.120 ;
    END
  END m_wbs_dat_o_3[18]
  PIN m_wbs_dat_o_3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 401.240 204.000 401.840 ;
    END
  END m_wbs_dat_o_3[19]
  PIN m_wbs_dat_o_3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 360.440 204.000 361.040 ;
    END
  END m_wbs_dat_o_3[1]
  PIN m_wbs_dat_o_3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 403.280 204.000 403.880 ;
    END
  END m_wbs_dat_o_3[20]
  PIN m_wbs_dat_o_3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 405.320 204.000 405.920 ;
    END
  END m_wbs_dat_o_3[21]
  PIN m_wbs_dat_o_3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 407.360 204.000 407.960 ;
    END
  END m_wbs_dat_o_3[22]
  PIN m_wbs_dat_o_3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 410.080 204.000 410.680 ;
    END
  END m_wbs_dat_o_3[23]
  PIN m_wbs_dat_o_3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 412.120 204.000 412.720 ;
    END
  END m_wbs_dat_o_3[24]
  PIN m_wbs_dat_o_3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 414.160 204.000 414.760 ;
    END
  END m_wbs_dat_o_3[25]
  PIN m_wbs_dat_o_3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 416.880 204.000 417.480 ;
    END
  END m_wbs_dat_o_3[26]
  PIN m_wbs_dat_o_3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 418.920 204.000 419.520 ;
    END
  END m_wbs_dat_o_3[27]
  PIN m_wbs_dat_o_3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 420.960 204.000 421.560 ;
    END
  END m_wbs_dat_o_3[28]
  PIN m_wbs_dat_o_3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 423.680 204.000 424.280 ;
    END
  END m_wbs_dat_o_3[29]
  PIN m_wbs_dat_o_3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 363.160 204.000 363.760 ;
    END
  END m_wbs_dat_o_3[2]
  PIN m_wbs_dat_o_3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 425.720 204.000 426.320 ;
    END
  END m_wbs_dat_o_3[30]
  PIN m_wbs_dat_o_3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 427.760 204.000 428.360 ;
    END
  END m_wbs_dat_o_3[31]
  PIN m_wbs_dat_o_3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 365.200 204.000 365.800 ;
    END
  END m_wbs_dat_o_3[3]
  PIN m_wbs_dat_o_3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 367.240 204.000 367.840 ;
    END
  END m_wbs_dat_o_3[4]
  PIN m_wbs_dat_o_3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 369.960 204.000 370.560 ;
    END
  END m_wbs_dat_o_3[5]
  PIN m_wbs_dat_o_3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 372.000 204.000 372.600 ;
    END
  END m_wbs_dat_o_3[6]
  PIN m_wbs_dat_o_3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 374.040 204.000 374.640 ;
    END
  END m_wbs_dat_o_3[7]
  PIN m_wbs_dat_o_3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 376.080 204.000 376.680 ;
    END
  END m_wbs_dat_o_3[8]
  PIN m_wbs_dat_o_3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 378.800 204.000 379.400 ;
    END
  END m_wbs_dat_o_3[9]
  PIN m_wbs_dat_o_4[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 429.800 204.000 430.400 ;
    END
  END m_wbs_dat_o_4[0]
  PIN m_wbs_dat_o_4[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 452.240 204.000 452.840 ;
    END
  END m_wbs_dat_o_4[10]
  PIN m_wbs_dat_o_4[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 454.960 204.000 455.560 ;
    END
  END m_wbs_dat_o_4[11]
  PIN m_wbs_dat_o_4[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 457.000 204.000 457.600 ;
    END
  END m_wbs_dat_o_4[12]
  PIN m_wbs_dat_o_4[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 459.040 204.000 459.640 ;
    END
  END m_wbs_dat_o_4[13]
  PIN m_wbs_dat_o_4[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 461.080 204.000 461.680 ;
    END
  END m_wbs_dat_o_4[14]
  PIN m_wbs_dat_o_4[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 463.800 204.000 464.400 ;
    END
  END m_wbs_dat_o_4[15]
  PIN m_wbs_dat_o_4[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 465.840 204.000 466.440 ;
    END
  END m_wbs_dat_o_4[16]
  PIN m_wbs_dat_o_4[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 467.880 204.000 468.480 ;
    END
  END m_wbs_dat_o_4[17]
  PIN m_wbs_dat_o_4[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 470.600 204.000 471.200 ;
    END
  END m_wbs_dat_o_4[18]
  PIN m_wbs_dat_o_4[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 472.640 204.000 473.240 ;
    END
  END m_wbs_dat_o_4[19]
  PIN m_wbs_dat_o_4[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 432.520 204.000 433.120 ;
    END
  END m_wbs_dat_o_4[1]
  PIN m_wbs_dat_o_4[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 474.680 204.000 475.280 ;
    END
  END m_wbs_dat_o_4[20]
  PIN m_wbs_dat_o_4[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 476.720 204.000 477.320 ;
    END
  END m_wbs_dat_o_4[21]
  PIN m_wbs_dat_o_4[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 479.440 204.000 480.040 ;
    END
  END m_wbs_dat_o_4[22]
  PIN m_wbs_dat_o_4[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 481.480 204.000 482.080 ;
    END
  END m_wbs_dat_o_4[23]
  PIN m_wbs_dat_o_4[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 483.520 204.000 484.120 ;
    END
  END m_wbs_dat_o_4[24]
  PIN m_wbs_dat_o_4[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 486.240 204.000 486.840 ;
    END
  END m_wbs_dat_o_4[25]
  PIN m_wbs_dat_o_4[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 488.280 204.000 488.880 ;
    END
  END m_wbs_dat_o_4[26]
  PIN m_wbs_dat_o_4[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 490.320 204.000 490.920 ;
    END
  END m_wbs_dat_o_4[27]
  PIN m_wbs_dat_o_4[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 493.040 204.000 493.640 ;
    END
  END m_wbs_dat_o_4[28]
  PIN m_wbs_dat_o_4[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 495.080 204.000 495.680 ;
    END
  END m_wbs_dat_o_4[29]
  PIN m_wbs_dat_o_4[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 434.560 204.000 435.160 ;
    END
  END m_wbs_dat_o_4[2]
  PIN m_wbs_dat_o_4[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 497.120 204.000 497.720 ;
    END
  END m_wbs_dat_o_4[30]
  PIN m_wbs_dat_o_4[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 499.160 204.000 499.760 ;
    END
  END m_wbs_dat_o_4[31]
  PIN m_wbs_dat_o_4[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 436.600 204.000 437.200 ;
    END
  END m_wbs_dat_o_4[3]
  PIN m_wbs_dat_o_4[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 439.320 204.000 439.920 ;
    END
  END m_wbs_dat_o_4[4]
  PIN m_wbs_dat_o_4[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 441.360 204.000 441.960 ;
    END
  END m_wbs_dat_o_4[5]
  PIN m_wbs_dat_o_4[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 443.400 204.000 444.000 ;
    END
  END m_wbs_dat_o_4[6]
  PIN m_wbs_dat_o_4[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 445.440 204.000 446.040 ;
    END
  END m_wbs_dat_o_4[7]
  PIN m_wbs_dat_o_4[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 448.160 204.000 448.760 ;
    END
  END m_wbs_dat_o_4[8]
  PIN m_wbs_dat_o_4[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 450.200 204.000 450.800 ;
    END
  END m_wbs_dat_o_4[9]
  PIN m_wbs_dat_o_5[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 501.880 204.000 502.480 ;
    END
  END m_wbs_dat_o_5[0]
  PIN m_wbs_dat_o_5[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 524.320 204.000 524.920 ;
    END
  END m_wbs_dat_o_5[10]
  PIN m_wbs_dat_o_5[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 526.360 204.000 526.960 ;
    END
  END m_wbs_dat_o_5[11]
  PIN m_wbs_dat_o_5[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 528.400 204.000 529.000 ;
    END
  END m_wbs_dat_o_5[12]
  PIN m_wbs_dat_o_5[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 530.440 204.000 531.040 ;
    END
  END m_wbs_dat_o_5[13]
  PIN m_wbs_dat_o_5[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 533.160 204.000 533.760 ;
    END
  END m_wbs_dat_o_5[14]
  PIN m_wbs_dat_o_5[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 535.200 204.000 535.800 ;
    END
  END m_wbs_dat_o_5[15]
  PIN m_wbs_dat_o_5[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 537.240 204.000 537.840 ;
    END
  END m_wbs_dat_o_5[16]
  PIN m_wbs_dat_o_5[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 539.960 204.000 540.560 ;
    END
  END m_wbs_dat_o_5[17]
  PIN m_wbs_dat_o_5[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 542.000 204.000 542.600 ;
    END
  END m_wbs_dat_o_5[18]
  PIN m_wbs_dat_o_5[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 544.040 204.000 544.640 ;
    END
  END m_wbs_dat_o_5[19]
  PIN m_wbs_dat_o_5[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 503.920 204.000 504.520 ;
    END
  END m_wbs_dat_o_5[1]
  PIN m_wbs_dat_o_5[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 546.760 204.000 547.360 ;
    END
  END m_wbs_dat_o_5[20]
  PIN m_wbs_dat_o_5[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 548.800 204.000 549.400 ;
    END
  END m_wbs_dat_o_5[21]
  PIN m_wbs_dat_o_5[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 550.840 204.000 551.440 ;
    END
  END m_wbs_dat_o_5[22]
  PIN m_wbs_dat_o_5[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 552.880 204.000 553.480 ;
    END
  END m_wbs_dat_o_5[23]
  PIN m_wbs_dat_o_5[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 555.600 204.000 556.200 ;
    END
  END m_wbs_dat_o_5[24]
  PIN m_wbs_dat_o_5[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 557.640 204.000 558.240 ;
    END
  END m_wbs_dat_o_5[25]
  PIN m_wbs_dat_o_5[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 559.680 204.000 560.280 ;
    END
  END m_wbs_dat_o_5[26]
  PIN m_wbs_dat_o_5[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 562.400 204.000 563.000 ;
    END
  END m_wbs_dat_o_5[27]
  PIN m_wbs_dat_o_5[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 564.440 204.000 565.040 ;
    END
  END m_wbs_dat_o_5[28]
  PIN m_wbs_dat_o_5[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 566.480 204.000 567.080 ;
    END
  END m_wbs_dat_o_5[29]
  PIN m_wbs_dat_o_5[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 505.960 204.000 506.560 ;
    END
  END m_wbs_dat_o_5[2]
  PIN m_wbs_dat_o_5[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 568.520 204.000 569.120 ;
    END
  END m_wbs_dat_o_5[30]
  PIN m_wbs_dat_o_5[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 571.240 204.000 571.840 ;
    END
  END m_wbs_dat_o_5[31]
  PIN m_wbs_dat_o_5[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 508.680 204.000 509.280 ;
    END
  END m_wbs_dat_o_5[3]
  PIN m_wbs_dat_o_5[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 510.720 204.000 511.320 ;
    END
  END m_wbs_dat_o_5[4]
  PIN m_wbs_dat_o_5[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 512.760 204.000 513.360 ;
    END
  END m_wbs_dat_o_5[5]
  PIN m_wbs_dat_o_5[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 514.800 204.000 515.400 ;
    END
  END m_wbs_dat_o_5[6]
  PIN m_wbs_dat_o_5[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 517.520 204.000 518.120 ;
    END
  END m_wbs_dat_o_5[7]
  PIN m_wbs_dat_o_5[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 519.560 204.000 520.160 ;
    END
  END m_wbs_dat_o_5[8]
  PIN m_wbs_dat_o_5[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 521.600 204.000 522.200 ;
    END
  END m_wbs_dat_o_5[9]
  PIN m_wbs_dat_o_6[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1.400 4.000 2.000 ;
    END
  END m_wbs_dat_o_6[0]
  PIN m_wbs_dat_o_6[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 40.840 4.000 41.440 ;
    END
  END m_wbs_dat_o_6[10]
  PIN m_wbs_dat_o_6[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 44.920 4.000 45.520 ;
    END
  END m_wbs_dat_o_6[11]
  PIN m_wbs_dat_o_6[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 49.000 4.000 49.600 ;
    END
  END m_wbs_dat_o_6[12]
  PIN m_wbs_dat_o_6[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 53.080 4.000 53.680 ;
    END
  END m_wbs_dat_o_6[13]
  PIN m_wbs_dat_o_6[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 57.160 4.000 57.760 ;
    END
  END m_wbs_dat_o_6[14]
  PIN m_wbs_dat_o_6[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 61.240 4.000 61.840 ;
    END
  END m_wbs_dat_o_6[15]
  PIN m_wbs_dat_o_6[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 65.320 4.000 65.920 ;
    END
  END m_wbs_dat_o_6[16]
  PIN m_wbs_dat_o_6[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 68.720 4.000 69.320 ;
    END
  END m_wbs_dat_o_6[17]
  PIN m_wbs_dat_o_6[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 72.800 4.000 73.400 ;
    END
  END m_wbs_dat_o_6[18]
  PIN m_wbs_dat_o_6[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 76.880 4.000 77.480 ;
    END
  END m_wbs_dat_o_6[19]
  PIN m_wbs_dat_o_6[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 4.800 4.000 5.400 ;
    END
  END m_wbs_dat_o_6[1]
  PIN m_wbs_dat_o_6[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 80.960 4.000 81.560 ;
    END
  END m_wbs_dat_o_6[20]
  PIN m_wbs_dat_o_6[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 85.040 4.000 85.640 ;
    END
  END m_wbs_dat_o_6[21]
  PIN m_wbs_dat_o_6[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 89.120 4.000 89.720 ;
    END
  END m_wbs_dat_o_6[22]
  PIN m_wbs_dat_o_6[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 93.200 4.000 93.800 ;
    END
  END m_wbs_dat_o_6[23]
  PIN m_wbs_dat_o_6[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 97.280 4.000 97.880 ;
    END
  END m_wbs_dat_o_6[24]
  PIN m_wbs_dat_o_6[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 101.360 4.000 101.960 ;
    END
  END m_wbs_dat_o_6[25]
  PIN m_wbs_dat_o_6[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 104.760 4.000 105.360 ;
    END
  END m_wbs_dat_o_6[26]
  PIN m_wbs_dat_o_6[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 108.840 4.000 109.440 ;
    END
  END m_wbs_dat_o_6[27]
  PIN m_wbs_dat_o_6[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 112.920 4.000 113.520 ;
    END
  END m_wbs_dat_o_6[28]
  PIN m_wbs_dat_o_6[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 117.000 4.000 117.600 ;
    END
  END m_wbs_dat_o_6[29]
  PIN m_wbs_dat_o_6[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 8.880 4.000 9.480 ;
    END
  END m_wbs_dat_o_6[2]
  PIN m_wbs_dat_o_6[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 121.080 4.000 121.680 ;
    END
  END m_wbs_dat_o_6[30]
  PIN m_wbs_dat_o_6[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 125.160 4.000 125.760 ;
    END
  END m_wbs_dat_o_6[31]
  PIN m_wbs_dat_o_6[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 12.960 4.000 13.560 ;
    END
  END m_wbs_dat_o_6[3]
  PIN m_wbs_dat_o_6[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 17.040 4.000 17.640 ;
    END
  END m_wbs_dat_o_6[4]
  PIN m_wbs_dat_o_6[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 21.120 4.000 21.720 ;
    END
  END m_wbs_dat_o_6[5]
  PIN m_wbs_dat_o_6[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 25.200 4.000 25.800 ;
    END
  END m_wbs_dat_o_6[6]
  PIN m_wbs_dat_o_6[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 29.280 4.000 29.880 ;
    END
  END m_wbs_dat_o_6[7]
  PIN m_wbs_dat_o_6[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 33.360 4.000 33.960 ;
    END
  END m_wbs_dat_o_6[8]
  PIN m_wbs_dat_o_6[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 36.760 4.000 37.360 ;
    END
  END m_wbs_dat_o_6[9]
  PIN m_wbs_dat_o_7[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 129.240 4.000 129.840 ;
    END
  END m_wbs_dat_o_7[0]
  PIN m_wbs_dat_o_7[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 168.680 4.000 169.280 ;
    END
  END m_wbs_dat_o_7[10]
  PIN m_wbs_dat_o_7[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 172.760 4.000 173.360 ;
    END
  END m_wbs_dat_o_7[11]
  PIN m_wbs_dat_o_7[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 176.840 4.000 177.440 ;
    END
  END m_wbs_dat_o_7[12]
  PIN m_wbs_dat_o_7[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 180.920 4.000 181.520 ;
    END
  END m_wbs_dat_o_7[13]
  PIN m_wbs_dat_o_7[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 185.000 4.000 185.600 ;
    END
  END m_wbs_dat_o_7[14]
  PIN m_wbs_dat_o_7[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 189.080 4.000 189.680 ;
    END
  END m_wbs_dat_o_7[15]
  PIN m_wbs_dat_o_7[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 193.160 4.000 193.760 ;
    END
  END m_wbs_dat_o_7[16]
  PIN m_wbs_dat_o_7[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 197.240 4.000 197.840 ;
    END
  END m_wbs_dat_o_7[17]
  PIN m_wbs_dat_o_7[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 201.320 4.000 201.920 ;
    END
  END m_wbs_dat_o_7[18]
  PIN m_wbs_dat_o_7[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 204.720 4.000 205.320 ;
    END
  END m_wbs_dat_o_7[19]
  PIN m_wbs_dat_o_7[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 133.320 4.000 133.920 ;
    END
  END m_wbs_dat_o_7[1]
  PIN m_wbs_dat_o_7[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 208.800 4.000 209.400 ;
    END
  END m_wbs_dat_o_7[20]
  PIN m_wbs_dat_o_7[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 212.880 4.000 213.480 ;
    END
  END m_wbs_dat_o_7[21]
  PIN m_wbs_dat_o_7[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 216.960 4.000 217.560 ;
    END
  END m_wbs_dat_o_7[22]
  PIN m_wbs_dat_o_7[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 221.040 4.000 221.640 ;
    END
  END m_wbs_dat_o_7[23]
  PIN m_wbs_dat_o_7[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 225.120 4.000 225.720 ;
    END
  END m_wbs_dat_o_7[24]
  PIN m_wbs_dat_o_7[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 229.200 4.000 229.800 ;
    END
  END m_wbs_dat_o_7[25]
  PIN m_wbs_dat_o_7[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 233.280 4.000 233.880 ;
    END
  END m_wbs_dat_o_7[26]
  PIN m_wbs_dat_o_7[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 236.680 4.000 237.280 ;
    END
  END m_wbs_dat_o_7[27]
  PIN m_wbs_dat_o_7[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 240.760 4.000 241.360 ;
    END
  END m_wbs_dat_o_7[28]
  PIN m_wbs_dat_o_7[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 244.840 4.000 245.440 ;
    END
  END m_wbs_dat_o_7[29]
  PIN m_wbs_dat_o_7[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 136.720 4.000 137.320 ;
    END
  END m_wbs_dat_o_7[2]
  PIN m_wbs_dat_o_7[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 248.920 4.000 249.520 ;
    END
  END m_wbs_dat_o_7[30]
  PIN m_wbs_dat_o_7[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 253.000 4.000 253.600 ;
    END
  END m_wbs_dat_o_7[31]
  PIN m_wbs_dat_o_7[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 140.800 4.000 141.400 ;
    END
  END m_wbs_dat_o_7[3]
  PIN m_wbs_dat_o_7[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 144.880 4.000 145.480 ;
    END
  END m_wbs_dat_o_7[4]
  PIN m_wbs_dat_o_7[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 148.960 4.000 149.560 ;
    END
  END m_wbs_dat_o_7[5]
  PIN m_wbs_dat_o_7[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 153.040 4.000 153.640 ;
    END
  END m_wbs_dat_o_7[6]
  PIN m_wbs_dat_o_7[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 157.120 4.000 157.720 ;
    END
  END m_wbs_dat_o_7[7]
  PIN m_wbs_dat_o_7[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 161.200 4.000 161.800 ;
    END
  END m_wbs_dat_o_7[8]
  PIN m_wbs_dat_o_7[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 165.280 4.000 165.880 ;
    END
  END m_wbs_dat_o_7[9]
  PIN m_wbs_dat_o_8[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 257.080 4.000 257.680 ;
    END
  END m_wbs_dat_o_8[0]
  PIN m_wbs_dat_o_8[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 297.200 4.000 297.800 ;
    END
  END m_wbs_dat_o_8[10]
  PIN m_wbs_dat_o_8[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 301.280 4.000 301.880 ;
    END
  END m_wbs_dat_o_8[11]
  PIN m_wbs_dat_o_8[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 304.680 4.000 305.280 ;
    END
  END m_wbs_dat_o_8[12]
  PIN m_wbs_dat_o_8[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 308.760 4.000 309.360 ;
    END
  END m_wbs_dat_o_8[13]
  PIN m_wbs_dat_o_8[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 312.840 4.000 313.440 ;
    END
  END m_wbs_dat_o_8[14]
  PIN m_wbs_dat_o_8[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 316.920 4.000 317.520 ;
    END
  END m_wbs_dat_o_8[15]
  PIN m_wbs_dat_o_8[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 321.000 4.000 321.600 ;
    END
  END m_wbs_dat_o_8[16]
  PIN m_wbs_dat_o_8[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 325.080 4.000 325.680 ;
    END
  END m_wbs_dat_o_8[17]
  PIN m_wbs_dat_o_8[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 329.160 4.000 329.760 ;
    END
  END m_wbs_dat_o_8[18]
  PIN m_wbs_dat_o_8[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 333.240 4.000 333.840 ;
    END
  END m_wbs_dat_o_8[19]
  PIN m_wbs_dat_o_8[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 261.160 4.000 261.760 ;
    END
  END m_wbs_dat_o_8[1]
  PIN m_wbs_dat_o_8[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 336.640 4.000 337.240 ;
    END
  END m_wbs_dat_o_8[20]
  PIN m_wbs_dat_o_8[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 340.720 4.000 341.320 ;
    END
  END m_wbs_dat_o_8[21]
  PIN m_wbs_dat_o_8[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 344.800 4.000 345.400 ;
    END
  END m_wbs_dat_o_8[22]
  PIN m_wbs_dat_o_8[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 348.880 4.000 349.480 ;
    END
  END m_wbs_dat_o_8[23]
  PIN m_wbs_dat_o_8[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 352.960 4.000 353.560 ;
    END
  END m_wbs_dat_o_8[24]
  PIN m_wbs_dat_o_8[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 357.040 4.000 357.640 ;
    END
  END m_wbs_dat_o_8[25]
  PIN m_wbs_dat_o_8[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 361.120 4.000 361.720 ;
    END
  END m_wbs_dat_o_8[26]
  PIN m_wbs_dat_o_8[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 365.200 4.000 365.800 ;
    END
  END m_wbs_dat_o_8[27]
  PIN m_wbs_dat_o_8[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 368.600 4.000 369.200 ;
    END
  END m_wbs_dat_o_8[28]
  PIN m_wbs_dat_o_8[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 372.680 4.000 373.280 ;
    END
  END m_wbs_dat_o_8[29]
  PIN m_wbs_dat_o_8[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 265.240 4.000 265.840 ;
    END
  END m_wbs_dat_o_8[2]
  PIN m_wbs_dat_o_8[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 376.760 4.000 377.360 ;
    END
  END m_wbs_dat_o_8[30]
  PIN m_wbs_dat_o_8[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 380.840 4.000 381.440 ;
    END
  END m_wbs_dat_o_8[31]
  PIN m_wbs_dat_o_8[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 268.640 4.000 269.240 ;
    END
  END m_wbs_dat_o_8[3]
  PIN m_wbs_dat_o_8[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 272.720 4.000 273.320 ;
    END
  END m_wbs_dat_o_8[4]
  PIN m_wbs_dat_o_8[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 276.800 4.000 277.400 ;
    END
  END m_wbs_dat_o_8[5]
  PIN m_wbs_dat_o_8[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 280.880 4.000 281.480 ;
    END
  END m_wbs_dat_o_8[6]
  PIN m_wbs_dat_o_8[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 284.960 4.000 285.560 ;
    END
  END m_wbs_dat_o_8[7]
  PIN m_wbs_dat_o_8[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 289.040 4.000 289.640 ;
    END
  END m_wbs_dat_o_8[8]
  PIN m_wbs_dat_o_8[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 293.120 4.000 293.720 ;
    END
  END m_wbs_dat_o_8[9]
  PIN m_wbs_dat_o_9[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 384.920 4.000 385.520 ;
    END
  END m_wbs_dat_o_9[0]
  PIN m_wbs_dat_o_9[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 425.040 4.000 425.640 ;
    END
  END m_wbs_dat_o_9[10]
  PIN m_wbs_dat_o_9[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 429.120 4.000 429.720 ;
    END
  END m_wbs_dat_o_9[11]
  PIN m_wbs_dat_o_9[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 433.200 4.000 433.800 ;
    END
  END m_wbs_dat_o_9[12]
  PIN m_wbs_dat_o_9[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 436.600 4.000 437.200 ;
    END
  END m_wbs_dat_o_9[13]
  PIN m_wbs_dat_o_9[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 440.680 4.000 441.280 ;
    END
  END m_wbs_dat_o_9[14]
  PIN m_wbs_dat_o_9[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 444.760 4.000 445.360 ;
    END
  END m_wbs_dat_o_9[15]
  PIN m_wbs_dat_o_9[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 448.840 4.000 449.440 ;
    END
  END m_wbs_dat_o_9[16]
  PIN m_wbs_dat_o_9[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 452.920 4.000 453.520 ;
    END
  END m_wbs_dat_o_9[17]
  PIN m_wbs_dat_o_9[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 457.000 4.000 457.600 ;
    END
  END m_wbs_dat_o_9[18]
  PIN m_wbs_dat_o_9[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 461.080 4.000 461.680 ;
    END
  END m_wbs_dat_o_9[19]
  PIN m_wbs_dat_o_9[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 389.000 4.000 389.600 ;
    END
  END m_wbs_dat_o_9[1]
  PIN m_wbs_dat_o_9[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 465.160 4.000 465.760 ;
    END
  END m_wbs_dat_o_9[20]
  PIN m_wbs_dat_o_9[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 468.560 4.000 469.160 ;
    END
  END m_wbs_dat_o_9[21]
  PIN m_wbs_dat_o_9[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 472.640 4.000 473.240 ;
    END
  END m_wbs_dat_o_9[22]
  PIN m_wbs_dat_o_9[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 476.720 4.000 477.320 ;
    END
  END m_wbs_dat_o_9[23]
  PIN m_wbs_dat_o_9[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 480.800 4.000 481.400 ;
    END
  END m_wbs_dat_o_9[24]
  PIN m_wbs_dat_o_9[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 484.880 4.000 485.480 ;
    END
  END m_wbs_dat_o_9[25]
  PIN m_wbs_dat_o_9[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 488.960 4.000 489.560 ;
    END
  END m_wbs_dat_o_9[26]
  PIN m_wbs_dat_o_9[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 493.040 4.000 493.640 ;
    END
  END m_wbs_dat_o_9[27]
  PIN m_wbs_dat_o_9[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 497.120 4.000 497.720 ;
    END
  END m_wbs_dat_o_9[28]
  PIN m_wbs_dat_o_9[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 501.200 4.000 501.800 ;
    END
  END m_wbs_dat_o_9[29]
  PIN m_wbs_dat_o_9[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 393.080 4.000 393.680 ;
    END
  END m_wbs_dat_o_9[2]
  PIN m_wbs_dat_o_9[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 504.600 4.000 505.200 ;
    END
  END m_wbs_dat_o_9[30]
  PIN m_wbs_dat_o_9[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 508.680 4.000 509.280 ;
    END
  END m_wbs_dat_o_9[31]
  PIN m_wbs_dat_o_9[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 397.160 4.000 397.760 ;
    END
  END m_wbs_dat_o_9[3]
  PIN m_wbs_dat_o_9[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 401.240 4.000 401.840 ;
    END
  END m_wbs_dat_o_9[4]
  PIN m_wbs_dat_o_9[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 404.640 4.000 405.240 ;
    END
  END m_wbs_dat_o_9[5]
  PIN m_wbs_dat_o_9[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 408.720 4.000 409.320 ;
    END
  END m_wbs_dat_o_9[6]
  PIN m_wbs_dat_o_9[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 412.800 4.000 413.400 ;
    END
  END m_wbs_dat_o_9[7]
  PIN m_wbs_dat_o_9[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 416.880 4.000 417.480 ;
    END
  END m_wbs_dat_o_9[8]
  PIN m_wbs_dat_o_9[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 420.960 4.000 421.560 ;
    END
  END m_wbs_dat_o_9[9]
  PIN m_wbs_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 512.760 4.000 513.360 ;
    END
  END m_wbs_we_i
  PIN mt_QEI_ChA_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 596.000 141.590 604.000 ;
    END
  END mt_QEI_ChA_0
  PIN mt_QEI_ChA_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 596.000 142.970 604.000 ;
    END
  END mt_QEI_ChA_1
  PIN mt_QEI_ChA_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 596.000 143.890 604.000 ;
    END
  END mt_QEI_ChA_2
  PIN mt_QEI_ChA_3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 596.000 145.270 604.000 ;
    END
  END mt_QEI_ChA_3
  PIN mt_QEI_ChB_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 596.000 146.190 604.000 ;
    END
  END mt_QEI_ChB_0
  PIN mt_QEI_ChB_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 596.000 147.570 604.000 ;
    END
  END mt_QEI_ChB_1
  PIN mt_QEI_ChB_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 596.000 148.490 604.000 ;
    END
  END mt_QEI_ChB_2
  PIN mt_QEI_ChB_3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 596.000 149.870 604.000 ;
    END
  END mt_QEI_ChB_3
  PIN mt_pwm_h_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 596.000 150.790 604.000 ;
    END
  END mt_pwm_h_0
  PIN mt_pwm_h_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 596.000 152.170 604.000 ;
    END
  END mt_pwm_h_1
  PIN mt_pwm_h_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 596.000 153.090 604.000 ;
    END
  END mt_pwm_h_2
  PIN mt_pwm_h_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 596.000 154.470 604.000 ;
    END
  END mt_pwm_h_3
  PIN mt_pwm_l_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 596.000 155.390 604.000 ;
    END
  END mt_pwm_l_0
  PIN mt_pwm_l_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 596.000 156.770 604.000 ;
    END
  END mt_pwm_l_1
  PIN mt_pwm_l_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 596.000 157.690 604.000 ;
    END
  END mt_pwm_l_2
  PIN mt_pwm_l_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 596.000 159.070 604.000 ;
    END
  END mt_pwm_l_3
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 -4.000 0.830 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 -4.000 2.210 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 -4.000 8.650 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 -4.000 15.090 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 -4.000 70.750 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 -4.000 75.350 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 -4.000 80.410 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 -4.000 85.010 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 -4.000 90.070 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 -4.000 95.130 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 -4.000 99.730 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 -4.000 104.790 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 -4.000 109.390 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 -4.000 114.450 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 -4.000 21.530 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 -4.000 119.510 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 -4.000 124.110 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 -4.000 129.170 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 -4.000 134.230 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 -4.000 138.830 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 -4.000 143.890 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 -4.000 148.490 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 -4.000 153.550 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 -4.000 158.610 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 -4.000 163.210 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 -4.000 28.430 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 -4.000 168.270 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 -4.000 172.870 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 -4.000 34.870 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 -4.000 41.310 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 -4.000 46.370 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 -4.000 50.970 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 -4.000 56.030 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 -4.000 60.630 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 -4.000 65.690 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 -4.000 10.490 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 -4.000 16.930 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 -4.000 72.130 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 -4.000 77.190 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 -4.000 81.790 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 -4.000 86.850 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 -4.000 91.910 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 -4.000 96.510 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 -4.000 101.570 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 -4.000 106.170 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 -4.000 111.230 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 -4.000 116.290 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 -4.000 23.370 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 -4.000 120.890 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 -4.000 125.950 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 -4.000 130.550 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 -4.000 135.610 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 -4.000 140.670 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 -4.000 145.270 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 -4.000 150.330 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 -4.000 154.930 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 -4.000 159.990 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 -4.000 165.050 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 -4.000 29.810 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 -4.000 169.650 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 -4.000 174.710 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 -4.000 36.250 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 -4.000 42.690 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 -4.000 47.750 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 -4.000 52.810 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 -4.000 57.410 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 -4.000 62.470 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 -4.000 67.530 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 -4.000 18.310 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 -4.000 73.970 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 -4.000 78.570 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 -4.000 83.630 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 -4.000 88.230 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 -4.000 93.290 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 -4.000 98.350 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 -4.000 102.950 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 -4.000 108.010 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 -4.000 113.070 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 -4.000 117.670 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 -4.000 25.210 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 -4.000 122.730 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 -4.000 127.330 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 -4.000 132.390 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 -4.000 137.450 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 -4.000 142.050 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 -4.000 147.110 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 -4.000 151.710 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 -4.000 156.770 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 -4.000 161.830 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 -4.000 166.430 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 -4.000 31.650 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 -4.000 171.490 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 -4.000 176.090 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 -4.000 38.090 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 -4.000 44.530 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 -4.000 49.590 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 -4.000 54.190 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 -4.000 59.250 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 -4.000 63.850 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 -4.000 68.910 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 -4.000 20.150 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 -4.000 26.590 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 -4.000 33.030 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 -4.000 39.470 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 -4.000 11.870 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 -4.000 13.710 4.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 199.035 587.605 ;
      LAYER met1 ;
        RECT 0.530 411.360 200.000 591.220 ;
        RECT 0.530 411.100 200.030 411.360 ;
        RECT 0.530 325.340 200.000 411.100 ;
        RECT 0.530 325.080 200.030 325.340 ;
        RECT 0.530 7.520 200.000 325.080 ;
      LAYER met2 ;
        RECT 1.110 595.720 1.190 598.245 ;
        RECT 2.030 595.720 2.570 598.245 ;
        RECT 3.410 595.720 3.490 598.245 ;
        RECT 4.330 595.720 4.870 598.245 ;
        RECT 5.710 595.720 5.790 598.245 ;
        RECT 6.630 595.720 7.170 598.245 ;
        RECT 8.010 595.720 8.090 598.245 ;
        RECT 8.930 595.720 9.470 598.245 ;
        RECT 10.310 595.720 10.390 598.245 ;
        RECT 11.230 595.720 11.770 598.245 ;
        RECT 12.610 595.720 12.690 598.245 ;
        RECT 13.530 595.720 14.070 598.245 ;
        RECT 14.910 595.720 14.990 598.245 ;
        RECT 15.830 595.720 16.370 598.245 ;
        RECT 17.210 595.720 17.290 598.245 ;
        RECT 18.130 595.720 18.670 598.245 ;
        RECT 19.510 595.720 19.590 598.245 ;
        RECT 20.430 595.720 20.970 598.245 ;
        RECT 21.810 595.720 21.890 598.245 ;
        RECT 22.730 595.720 23.270 598.245 ;
        RECT 24.110 595.720 24.190 598.245 ;
        RECT 25.030 595.720 25.570 598.245 ;
        RECT 26.410 595.720 26.490 598.245 ;
        RECT 27.330 595.720 27.870 598.245 ;
        RECT 28.710 595.720 28.790 598.245 ;
        RECT 29.630 595.720 30.170 598.245 ;
        RECT 31.010 595.720 31.090 598.245 ;
        RECT 31.930 595.720 32.470 598.245 ;
        RECT 33.310 595.720 33.390 598.245 ;
        RECT 34.230 595.720 34.770 598.245 ;
        RECT 35.610 595.720 35.690 598.245 ;
        RECT 36.530 595.720 37.070 598.245 ;
        RECT 37.910 595.720 37.990 598.245 ;
        RECT 38.830 595.720 39.370 598.245 ;
        RECT 40.210 595.720 40.750 598.245 ;
        RECT 41.590 595.720 41.670 598.245 ;
        RECT 42.510 595.720 43.050 598.245 ;
        RECT 43.890 595.720 43.970 598.245 ;
        RECT 44.810 595.720 45.350 598.245 ;
        RECT 46.190 595.720 46.270 598.245 ;
        RECT 47.110 595.720 47.650 598.245 ;
        RECT 48.490 595.720 48.570 598.245 ;
        RECT 49.410 595.720 49.950 598.245 ;
        RECT 50.790 595.720 50.870 598.245 ;
        RECT 51.710 595.720 52.250 598.245 ;
        RECT 53.090 595.720 53.170 598.245 ;
        RECT 54.010 595.720 54.550 598.245 ;
        RECT 55.390 595.720 55.470 598.245 ;
        RECT 56.310 595.720 56.850 598.245 ;
        RECT 57.690 595.720 57.770 598.245 ;
        RECT 58.610 595.720 59.150 598.245 ;
        RECT 59.990 595.720 60.070 598.245 ;
        RECT 60.910 595.720 61.450 598.245 ;
        RECT 62.290 595.720 62.370 598.245 ;
        RECT 63.210 595.720 63.750 598.245 ;
        RECT 64.590 595.720 64.670 598.245 ;
        RECT 65.510 595.720 66.050 598.245 ;
        RECT 66.890 595.720 66.970 598.245 ;
        RECT 67.810 595.720 68.350 598.245 ;
        RECT 69.190 595.720 69.270 598.245 ;
        RECT 70.110 595.720 70.650 598.245 ;
        RECT 71.490 595.720 71.570 598.245 ;
        RECT 72.410 595.720 72.950 598.245 ;
        RECT 73.790 595.720 73.870 598.245 ;
        RECT 74.710 595.720 75.250 598.245 ;
        RECT 76.090 595.720 76.170 598.245 ;
        RECT 77.010 595.720 77.550 598.245 ;
        RECT 78.390 595.720 78.470 598.245 ;
        RECT 79.310 595.720 79.850 598.245 ;
        RECT 80.690 595.720 81.230 598.245 ;
        RECT 82.070 595.720 82.150 598.245 ;
        RECT 82.990 595.720 83.530 598.245 ;
        RECT 84.370 595.720 84.450 598.245 ;
        RECT 85.290 595.720 85.830 598.245 ;
        RECT 86.670 595.720 86.750 598.245 ;
        RECT 87.590 595.720 88.130 598.245 ;
        RECT 88.970 595.720 89.050 598.245 ;
        RECT 89.890 595.720 90.430 598.245 ;
        RECT 91.270 595.720 91.350 598.245 ;
        RECT 92.190 595.720 92.730 598.245 ;
        RECT 93.570 595.720 93.650 598.245 ;
        RECT 94.490 595.720 95.030 598.245 ;
        RECT 95.870 595.720 95.950 598.245 ;
        RECT 96.790 595.720 97.330 598.245 ;
        RECT 98.170 595.720 98.250 598.245 ;
        RECT 99.090 595.720 99.630 598.245 ;
        RECT 100.470 595.720 100.550 598.245 ;
        RECT 101.390 595.720 101.930 598.245 ;
        RECT 102.770 595.720 102.850 598.245 ;
        RECT 103.690 595.720 104.230 598.245 ;
        RECT 105.070 595.720 105.150 598.245 ;
        RECT 105.990 595.720 106.530 598.245 ;
        RECT 107.370 595.720 107.450 598.245 ;
        RECT 108.290 595.720 108.830 598.245 ;
        RECT 109.670 595.720 109.750 598.245 ;
        RECT 110.590 595.720 111.130 598.245 ;
        RECT 111.970 595.720 112.050 598.245 ;
        RECT 112.890 595.720 113.430 598.245 ;
        RECT 114.270 595.720 114.350 598.245 ;
        RECT 115.190 595.720 115.730 598.245 ;
        RECT 116.570 595.720 116.650 598.245 ;
        RECT 117.490 595.720 118.030 598.245 ;
        RECT 118.870 595.720 118.950 598.245 ;
        RECT 119.790 595.720 120.330 598.245 ;
        RECT 121.170 595.720 121.710 598.245 ;
        RECT 122.550 595.720 122.630 598.245 ;
        RECT 123.470 595.720 124.010 598.245 ;
        RECT 124.850 595.720 124.930 598.245 ;
        RECT 125.770 595.720 126.310 598.245 ;
        RECT 127.150 595.720 127.230 598.245 ;
        RECT 128.070 595.720 128.610 598.245 ;
        RECT 129.450 595.720 129.530 598.245 ;
        RECT 130.370 595.720 130.910 598.245 ;
        RECT 131.750 595.720 131.830 598.245 ;
        RECT 132.670 595.720 133.210 598.245 ;
        RECT 134.050 595.720 134.130 598.245 ;
        RECT 134.970 595.720 135.510 598.245 ;
        RECT 136.350 595.720 136.430 598.245 ;
        RECT 137.270 595.720 137.810 598.245 ;
        RECT 138.650 595.720 138.730 598.245 ;
        RECT 139.570 595.720 140.110 598.245 ;
        RECT 140.950 595.720 141.030 598.245 ;
        RECT 141.870 595.720 142.410 598.245 ;
        RECT 143.250 595.720 143.330 598.245 ;
        RECT 144.170 595.720 144.710 598.245 ;
        RECT 145.550 595.720 145.630 598.245 ;
        RECT 146.470 595.720 147.010 598.245 ;
        RECT 147.850 595.720 147.930 598.245 ;
        RECT 148.770 595.720 149.310 598.245 ;
        RECT 150.150 595.720 150.230 598.245 ;
        RECT 151.070 595.720 151.610 598.245 ;
        RECT 152.450 595.720 152.530 598.245 ;
        RECT 153.370 595.720 153.910 598.245 ;
        RECT 154.750 595.720 154.830 598.245 ;
        RECT 155.670 595.720 156.210 598.245 ;
        RECT 157.050 595.720 157.130 598.245 ;
        RECT 157.970 595.720 158.510 598.245 ;
        RECT 159.350 595.720 159.430 598.245 ;
        RECT 160.270 595.720 160.810 598.245 ;
        RECT 161.650 595.720 162.190 598.245 ;
        RECT 163.030 595.720 163.110 598.245 ;
        RECT 163.950 595.720 164.490 598.245 ;
        RECT 165.330 595.720 165.410 598.245 ;
        RECT 166.250 595.720 166.790 598.245 ;
        RECT 167.630 595.720 167.710 598.245 ;
        RECT 168.550 595.720 169.090 598.245 ;
        RECT 169.930 595.720 170.010 598.245 ;
        RECT 170.850 595.720 171.390 598.245 ;
        RECT 172.230 595.720 172.310 598.245 ;
        RECT 173.150 595.720 173.690 598.245 ;
        RECT 174.530 595.720 174.610 598.245 ;
        RECT 175.450 595.720 175.990 598.245 ;
        RECT 176.830 595.720 176.910 598.245 ;
        RECT 177.750 595.720 178.290 598.245 ;
        RECT 179.130 595.720 179.210 598.245 ;
        RECT 180.050 595.720 180.590 598.245 ;
        RECT 181.430 595.720 181.510 598.245 ;
        RECT 182.350 595.720 182.890 598.245 ;
        RECT 183.730 595.720 183.810 598.245 ;
        RECT 184.650 595.720 185.190 598.245 ;
        RECT 186.030 595.720 186.110 598.245 ;
        RECT 186.950 595.720 187.490 598.245 ;
        RECT 188.330 595.720 188.410 598.245 ;
        RECT 189.250 595.720 189.790 598.245 ;
        RECT 190.630 595.720 190.710 598.245 ;
        RECT 191.550 595.720 192.090 598.245 ;
        RECT 192.930 595.720 193.010 598.245 ;
        RECT 193.850 595.720 194.390 598.245 ;
        RECT 195.230 595.720 195.310 598.245 ;
        RECT 196.150 595.720 196.690 598.245 ;
        RECT 197.530 595.720 197.610 598.245 ;
        RECT 198.450 595.720 198.990 598.245 ;
        RECT 199.830 595.720 200.000 598.245 ;
        RECT 0.560 4.280 200.000 595.720 ;
        RECT 1.110 0.835 1.650 4.280 ;
        RECT 2.490 0.835 3.490 4.280 ;
        RECT 4.330 0.835 4.870 4.280 ;
        RECT 5.710 0.835 6.710 4.280 ;
        RECT 7.550 0.835 8.090 4.280 ;
        RECT 8.930 0.835 9.930 4.280 ;
        RECT 10.770 0.835 11.310 4.280 ;
        RECT 12.150 0.835 13.150 4.280 ;
        RECT 13.990 0.835 14.530 4.280 ;
        RECT 15.370 0.835 16.370 4.280 ;
        RECT 17.210 0.835 17.750 4.280 ;
        RECT 18.590 0.835 19.590 4.280 ;
        RECT 20.430 0.835 20.970 4.280 ;
        RECT 21.810 0.835 22.810 4.280 ;
        RECT 23.650 0.835 24.650 4.280 ;
        RECT 25.490 0.835 26.030 4.280 ;
        RECT 26.870 0.835 27.870 4.280 ;
        RECT 28.710 0.835 29.250 4.280 ;
        RECT 30.090 0.835 31.090 4.280 ;
        RECT 31.930 0.835 32.470 4.280 ;
        RECT 33.310 0.835 34.310 4.280 ;
        RECT 35.150 0.835 35.690 4.280 ;
        RECT 36.530 0.835 37.530 4.280 ;
        RECT 38.370 0.835 38.910 4.280 ;
        RECT 39.750 0.835 40.750 4.280 ;
        RECT 41.590 0.835 42.130 4.280 ;
        RECT 42.970 0.835 43.970 4.280 ;
        RECT 44.810 0.835 45.810 4.280 ;
        RECT 46.650 0.835 47.190 4.280 ;
        RECT 48.030 0.835 49.030 4.280 ;
        RECT 49.870 0.835 50.410 4.280 ;
        RECT 51.250 0.835 52.250 4.280 ;
        RECT 53.090 0.835 53.630 4.280 ;
        RECT 54.470 0.835 55.470 4.280 ;
        RECT 56.310 0.835 56.850 4.280 ;
        RECT 57.690 0.835 58.690 4.280 ;
        RECT 59.530 0.835 60.070 4.280 ;
        RECT 60.910 0.835 61.910 4.280 ;
        RECT 62.750 0.835 63.290 4.280 ;
        RECT 64.130 0.835 65.130 4.280 ;
        RECT 65.970 0.835 66.970 4.280 ;
        RECT 67.810 0.835 68.350 4.280 ;
        RECT 69.190 0.835 70.190 4.280 ;
        RECT 71.030 0.835 71.570 4.280 ;
        RECT 72.410 0.835 73.410 4.280 ;
        RECT 74.250 0.835 74.790 4.280 ;
        RECT 75.630 0.835 76.630 4.280 ;
        RECT 77.470 0.835 78.010 4.280 ;
        RECT 78.850 0.835 79.850 4.280 ;
        RECT 80.690 0.835 81.230 4.280 ;
        RECT 82.070 0.835 83.070 4.280 ;
        RECT 83.910 0.835 84.450 4.280 ;
        RECT 85.290 0.835 86.290 4.280 ;
        RECT 87.130 0.835 87.670 4.280 ;
        RECT 88.510 0.835 89.510 4.280 ;
        RECT 90.350 0.835 91.350 4.280 ;
        RECT 92.190 0.835 92.730 4.280 ;
        RECT 93.570 0.835 94.570 4.280 ;
        RECT 95.410 0.835 95.950 4.280 ;
        RECT 96.790 0.835 97.790 4.280 ;
        RECT 98.630 0.835 99.170 4.280 ;
        RECT 100.010 0.835 101.010 4.280 ;
        RECT 101.850 0.835 102.390 4.280 ;
        RECT 103.230 0.835 104.230 4.280 ;
        RECT 105.070 0.835 105.610 4.280 ;
        RECT 106.450 0.835 107.450 4.280 ;
        RECT 108.290 0.835 108.830 4.280 ;
        RECT 109.670 0.835 110.670 4.280 ;
        RECT 111.510 0.835 112.510 4.280 ;
        RECT 113.350 0.835 113.890 4.280 ;
        RECT 114.730 0.835 115.730 4.280 ;
        RECT 116.570 0.835 117.110 4.280 ;
        RECT 117.950 0.835 118.950 4.280 ;
        RECT 119.790 0.835 120.330 4.280 ;
        RECT 121.170 0.835 122.170 4.280 ;
        RECT 123.010 0.835 123.550 4.280 ;
        RECT 124.390 0.835 125.390 4.280 ;
        RECT 126.230 0.835 126.770 4.280 ;
        RECT 127.610 0.835 128.610 4.280 ;
        RECT 129.450 0.835 129.990 4.280 ;
        RECT 130.830 0.835 131.830 4.280 ;
        RECT 132.670 0.835 133.670 4.280 ;
        RECT 134.510 0.835 135.050 4.280 ;
        RECT 135.890 0.835 136.890 4.280 ;
        RECT 137.730 0.835 138.270 4.280 ;
        RECT 139.110 0.835 140.110 4.280 ;
        RECT 140.950 0.835 141.490 4.280 ;
        RECT 142.330 0.835 143.330 4.280 ;
        RECT 144.170 0.835 144.710 4.280 ;
        RECT 145.550 0.835 146.550 4.280 ;
        RECT 147.390 0.835 147.930 4.280 ;
        RECT 148.770 0.835 149.770 4.280 ;
        RECT 150.610 0.835 151.150 4.280 ;
        RECT 151.990 0.835 152.990 4.280 ;
        RECT 153.830 0.835 154.370 4.280 ;
        RECT 155.210 0.835 156.210 4.280 ;
        RECT 157.050 0.835 158.050 4.280 ;
        RECT 158.890 0.835 159.430 4.280 ;
        RECT 160.270 0.835 161.270 4.280 ;
        RECT 162.110 0.835 162.650 4.280 ;
        RECT 163.490 0.835 164.490 4.280 ;
        RECT 165.330 0.835 165.870 4.280 ;
        RECT 166.710 0.835 167.710 4.280 ;
        RECT 168.550 0.835 169.090 4.280 ;
        RECT 169.930 0.835 170.930 4.280 ;
        RECT 171.770 0.835 172.310 4.280 ;
        RECT 173.150 0.835 174.150 4.280 ;
        RECT 174.990 0.835 175.530 4.280 ;
        RECT 176.370 0.835 177.370 4.280 ;
        RECT 178.210 0.835 179.210 4.280 ;
        RECT 180.050 0.835 180.590 4.280 ;
        RECT 181.430 0.835 182.430 4.280 ;
        RECT 183.270 0.835 183.810 4.280 ;
        RECT 184.650 0.835 185.650 4.280 ;
        RECT 186.490 0.835 187.030 4.280 ;
        RECT 187.870 0.835 188.870 4.280 ;
        RECT 189.710 0.835 190.250 4.280 ;
        RECT 191.090 0.835 192.090 4.280 ;
        RECT 192.930 0.835 193.470 4.280 ;
        RECT 194.310 0.835 195.310 4.280 ;
        RECT 196.150 0.835 196.690 4.280 ;
        RECT 197.530 0.835 198.530 4.280 ;
        RECT 199.370 0.835 200.000 4.280 ;
      LAYER met3 ;
        RECT 4.000 598.080 195.600 598.225 ;
        RECT 4.400 597.360 195.600 598.080 ;
        RECT 4.400 596.720 199.115 597.360 ;
        RECT 4.400 596.680 195.600 596.720 ;
        RECT 4.000 595.320 195.600 596.680 ;
        RECT 4.000 594.680 199.115 595.320 ;
        RECT 4.000 594.000 195.600 594.680 ;
        RECT 4.400 593.280 195.600 594.000 ;
        RECT 4.400 592.600 199.115 593.280 ;
        RECT 4.000 591.960 199.115 592.600 ;
        RECT 4.000 590.560 195.600 591.960 ;
        RECT 4.000 589.920 199.115 590.560 ;
        RECT 4.400 588.520 195.600 589.920 ;
        RECT 4.000 587.880 199.115 588.520 ;
        RECT 4.000 586.480 195.600 587.880 ;
        RECT 4.000 585.840 199.115 586.480 ;
        RECT 4.400 585.160 199.115 585.840 ;
        RECT 4.400 584.440 195.600 585.160 ;
        RECT 4.000 583.760 195.600 584.440 ;
        RECT 4.000 583.120 199.115 583.760 ;
        RECT 4.000 581.760 195.600 583.120 ;
        RECT 4.400 581.720 195.600 581.760 ;
        RECT 4.400 581.080 199.115 581.720 ;
        RECT 4.400 580.360 195.600 581.080 ;
        RECT 4.000 579.680 195.600 580.360 ;
        RECT 4.000 579.040 199.115 579.680 ;
        RECT 4.000 577.680 195.600 579.040 ;
        RECT 4.400 577.640 195.600 577.680 ;
        RECT 4.400 576.320 199.115 577.640 ;
        RECT 4.400 576.280 195.600 576.320 ;
        RECT 4.000 574.920 195.600 576.280 ;
        RECT 4.000 574.280 199.115 574.920 ;
        RECT 4.000 573.600 195.600 574.280 ;
        RECT 4.400 572.880 195.600 573.600 ;
        RECT 4.400 572.240 199.115 572.880 ;
        RECT 4.400 572.200 195.600 572.240 ;
        RECT 4.000 570.840 195.600 572.200 ;
        RECT 4.000 569.520 199.115 570.840 ;
        RECT 4.400 568.120 195.600 569.520 ;
        RECT 4.000 567.480 199.115 568.120 ;
        RECT 4.000 566.120 195.600 567.480 ;
        RECT 4.400 566.080 195.600 566.120 ;
        RECT 4.400 565.440 199.115 566.080 ;
        RECT 4.400 564.720 195.600 565.440 ;
        RECT 4.000 564.040 195.600 564.720 ;
        RECT 4.000 563.400 199.115 564.040 ;
        RECT 4.000 562.040 195.600 563.400 ;
        RECT 4.400 562.000 195.600 562.040 ;
        RECT 4.400 560.680 199.115 562.000 ;
        RECT 4.400 560.640 195.600 560.680 ;
        RECT 4.000 559.280 195.600 560.640 ;
        RECT 4.000 558.640 199.115 559.280 ;
        RECT 4.000 557.960 195.600 558.640 ;
        RECT 4.400 557.240 195.600 557.960 ;
        RECT 4.400 556.600 199.115 557.240 ;
        RECT 4.400 556.560 195.600 556.600 ;
        RECT 4.000 555.200 195.600 556.560 ;
        RECT 4.000 553.880 199.115 555.200 ;
        RECT 4.400 552.480 195.600 553.880 ;
        RECT 4.000 551.840 199.115 552.480 ;
        RECT 4.000 550.440 195.600 551.840 ;
        RECT 4.000 549.800 199.115 550.440 ;
        RECT 4.400 548.400 195.600 549.800 ;
        RECT 4.000 547.760 199.115 548.400 ;
        RECT 4.000 546.360 195.600 547.760 ;
        RECT 4.000 545.720 199.115 546.360 ;
        RECT 4.400 545.040 199.115 545.720 ;
        RECT 4.400 544.320 195.600 545.040 ;
        RECT 4.000 543.640 195.600 544.320 ;
        RECT 4.000 543.000 199.115 543.640 ;
        RECT 4.000 541.640 195.600 543.000 ;
        RECT 4.400 541.600 195.600 541.640 ;
        RECT 4.400 540.960 199.115 541.600 ;
        RECT 4.400 540.240 195.600 540.960 ;
        RECT 4.000 539.560 195.600 540.240 ;
        RECT 4.000 538.240 199.115 539.560 ;
        RECT 4.000 537.560 195.600 538.240 ;
        RECT 4.400 536.840 195.600 537.560 ;
        RECT 4.400 536.200 199.115 536.840 ;
        RECT 4.400 536.160 195.600 536.200 ;
        RECT 4.000 534.800 195.600 536.160 ;
        RECT 4.000 534.160 199.115 534.800 ;
        RECT 4.400 532.760 195.600 534.160 ;
        RECT 4.000 531.440 199.115 532.760 ;
        RECT 4.000 530.080 195.600 531.440 ;
        RECT 4.400 530.040 195.600 530.080 ;
        RECT 4.400 529.400 199.115 530.040 ;
        RECT 4.400 528.680 195.600 529.400 ;
        RECT 4.000 528.000 195.600 528.680 ;
        RECT 4.000 527.360 199.115 528.000 ;
        RECT 4.000 526.000 195.600 527.360 ;
        RECT 4.400 525.960 195.600 526.000 ;
        RECT 4.400 525.320 199.115 525.960 ;
        RECT 4.400 524.600 195.600 525.320 ;
        RECT 4.000 523.920 195.600 524.600 ;
        RECT 4.000 522.600 199.115 523.920 ;
        RECT 4.000 521.920 195.600 522.600 ;
        RECT 4.400 521.200 195.600 521.920 ;
        RECT 4.400 520.560 199.115 521.200 ;
        RECT 4.400 520.520 195.600 520.560 ;
        RECT 4.000 519.160 195.600 520.520 ;
        RECT 4.000 518.520 199.115 519.160 ;
        RECT 4.000 517.840 195.600 518.520 ;
        RECT 4.400 517.120 195.600 517.840 ;
        RECT 4.400 516.440 199.115 517.120 ;
        RECT 4.000 515.800 199.115 516.440 ;
        RECT 4.000 514.400 195.600 515.800 ;
        RECT 4.000 513.760 199.115 514.400 ;
        RECT 4.400 512.360 195.600 513.760 ;
        RECT 4.000 511.720 199.115 512.360 ;
        RECT 4.000 510.320 195.600 511.720 ;
        RECT 4.000 509.680 199.115 510.320 ;
        RECT 4.400 508.280 195.600 509.680 ;
        RECT 4.000 506.960 199.115 508.280 ;
        RECT 4.000 505.600 195.600 506.960 ;
        RECT 4.400 505.560 195.600 505.600 ;
        RECT 4.400 504.920 199.115 505.560 ;
        RECT 4.400 504.200 195.600 504.920 ;
        RECT 4.000 503.520 195.600 504.200 ;
        RECT 4.000 502.880 199.115 503.520 ;
        RECT 4.000 502.200 195.600 502.880 ;
        RECT 4.400 501.480 195.600 502.200 ;
        RECT 4.400 500.800 199.115 501.480 ;
        RECT 4.000 500.160 199.115 500.800 ;
        RECT 4.000 498.760 195.600 500.160 ;
        RECT 4.000 498.120 199.115 498.760 ;
        RECT 4.400 496.720 195.600 498.120 ;
        RECT 4.000 496.080 199.115 496.720 ;
        RECT 4.000 494.680 195.600 496.080 ;
        RECT 4.000 494.040 199.115 494.680 ;
        RECT 4.400 492.640 195.600 494.040 ;
        RECT 4.000 491.320 199.115 492.640 ;
        RECT 4.000 489.960 195.600 491.320 ;
        RECT 4.400 489.920 195.600 489.960 ;
        RECT 4.400 489.280 199.115 489.920 ;
        RECT 4.400 488.560 195.600 489.280 ;
        RECT 4.000 487.880 195.600 488.560 ;
        RECT 4.000 487.240 199.115 487.880 ;
        RECT 4.000 485.880 195.600 487.240 ;
        RECT 4.400 485.840 195.600 485.880 ;
        RECT 4.400 484.520 199.115 485.840 ;
        RECT 4.400 484.480 195.600 484.520 ;
        RECT 4.000 483.120 195.600 484.480 ;
        RECT 4.000 482.480 199.115 483.120 ;
        RECT 4.000 481.800 195.600 482.480 ;
        RECT 4.400 481.080 195.600 481.800 ;
        RECT 4.400 480.440 199.115 481.080 ;
        RECT 4.400 480.400 195.600 480.440 ;
        RECT 4.000 479.040 195.600 480.400 ;
        RECT 4.000 477.720 199.115 479.040 ;
        RECT 4.400 476.320 195.600 477.720 ;
        RECT 4.000 475.680 199.115 476.320 ;
        RECT 4.000 474.280 195.600 475.680 ;
        RECT 4.000 473.640 199.115 474.280 ;
        RECT 4.400 472.240 195.600 473.640 ;
        RECT 4.000 471.600 199.115 472.240 ;
        RECT 4.000 470.200 195.600 471.600 ;
        RECT 4.000 469.560 199.115 470.200 ;
        RECT 4.400 468.880 199.115 469.560 ;
        RECT 4.400 468.160 195.600 468.880 ;
        RECT 4.000 467.480 195.600 468.160 ;
        RECT 4.000 466.840 199.115 467.480 ;
        RECT 4.000 466.160 195.600 466.840 ;
        RECT 4.400 465.440 195.600 466.160 ;
        RECT 4.400 464.800 199.115 465.440 ;
        RECT 4.400 464.760 195.600 464.800 ;
        RECT 4.000 463.400 195.600 464.760 ;
        RECT 4.000 462.080 199.115 463.400 ;
        RECT 4.400 460.680 195.600 462.080 ;
        RECT 4.000 460.040 199.115 460.680 ;
        RECT 4.000 458.640 195.600 460.040 ;
        RECT 4.000 458.000 199.115 458.640 ;
        RECT 4.400 456.600 195.600 458.000 ;
        RECT 4.000 455.960 199.115 456.600 ;
        RECT 4.000 454.560 195.600 455.960 ;
        RECT 4.000 453.920 199.115 454.560 ;
        RECT 4.400 453.240 199.115 453.920 ;
        RECT 4.400 452.520 195.600 453.240 ;
        RECT 4.000 451.840 195.600 452.520 ;
        RECT 4.000 451.200 199.115 451.840 ;
        RECT 4.000 449.840 195.600 451.200 ;
        RECT 4.400 449.800 195.600 449.840 ;
        RECT 4.400 449.160 199.115 449.800 ;
        RECT 4.400 448.440 195.600 449.160 ;
        RECT 4.000 447.760 195.600 448.440 ;
        RECT 4.000 446.440 199.115 447.760 ;
        RECT 4.000 445.760 195.600 446.440 ;
        RECT 4.400 445.040 195.600 445.760 ;
        RECT 4.400 444.400 199.115 445.040 ;
        RECT 4.400 444.360 195.600 444.400 ;
        RECT 4.000 443.000 195.600 444.360 ;
        RECT 4.000 442.360 199.115 443.000 ;
        RECT 4.000 441.680 195.600 442.360 ;
        RECT 4.400 440.960 195.600 441.680 ;
        RECT 4.400 440.320 199.115 440.960 ;
        RECT 4.400 440.280 195.600 440.320 ;
        RECT 4.000 438.920 195.600 440.280 ;
        RECT 4.000 437.600 199.115 438.920 ;
        RECT 4.400 436.200 195.600 437.600 ;
        RECT 4.000 435.560 199.115 436.200 ;
        RECT 4.000 434.200 195.600 435.560 ;
        RECT 4.400 434.160 195.600 434.200 ;
        RECT 4.400 433.520 199.115 434.160 ;
        RECT 4.400 432.800 195.600 433.520 ;
        RECT 4.000 432.120 195.600 432.800 ;
        RECT 4.000 430.800 199.115 432.120 ;
        RECT 4.000 430.120 195.600 430.800 ;
        RECT 4.400 429.400 195.600 430.120 ;
        RECT 4.400 428.760 199.115 429.400 ;
        RECT 4.400 428.720 195.600 428.760 ;
        RECT 4.000 427.360 195.600 428.720 ;
        RECT 4.000 426.720 199.115 427.360 ;
        RECT 4.000 426.040 195.600 426.720 ;
        RECT 4.400 425.320 195.600 426.040 ;
        RECT 4.400 424.680 199.115 425.320 ;
        RECT 4.400 424.640 195.600 424.680 ;
        RECT 4.000 423.280 195.600 424.640 ;
        RECT 4.000 421.960 199.115 423.280 ;
        RECT 4.400 420.560 195.600 421.960 ;
        RECT 4.000 419.920 199.115 420.560 ;
        RECT 4.000 418.520 195.600 419.920 ;
        RECT 4.000 417.880 199.115 418.520 ;
        RECT 4.400 416.480 195.600 417.880 ;
        RECT 4.000 415.160 199.115 416.480 ;
        RECT 4.000 413.800 195.600 415.160 ;
        RECT 4.400 413.760 195.600 413.800 ;
        RECT 4.400 413.120 199.115 413.760 ;
        RECT 4.400 412.400 195.600 413.120 ;
        RECT 4.000 411.720 195.600 412.400 ;
        RECT 4.000 411.080 199.115 411.720 ;
        RECT 4.000 409.720 195.600 411.080 ;
        RECT 4.400 409.680 195.600 409.720 ;
        RECT 4.400 408.360 199.115 409.680 ;
        RECT 4.400 408.320 195.600 408.360 ;
        RECT 4.000 406.960 195.600 408.320 ;
        RECT 4.000 406.320 199.115 406.960 ;
        RECT 4.000 405.640 195.600 406.320 ;
        RECT 4.400 404.920 195.600 405.640 ;
        RECT 4.400 404.280 199.115 404.920 ;
        RECT 4.400 404.240 195.600 404.280 ;
        RECT 4.000 402.880 195.600 404.240 ;
        RECT 4.000 402.240 199.115 402.880 ;
        RECT 4.400 400.840 195.600 402.240 ;
        RECT 4.000 399.520 199.115 400.840 ;
        RECT 4.000 398.160 195.600 399.520 ;
        RECT 4.400 398.120 195.600 398.160 ;
        RECT 4.400 397.480 199.115 398.120 ;
        RECT 4.400 396.760 195.600 397.480 ;
        RECT 4.000 396.080 195.600 396.760 ;
        RECT 4.000 395.440 199.115 396.080 ;
        RECT 4.000 394.080 195.600 395.440 ;
        RECT 4.400 394.040 195.600 394.080 ;
        RECT 4.400 392.720 199.115 394.040 ;
        RECT 4.400 392.680 195.600 392.720 ;
        RECT 4.000 391.320 195.600 392.680 ;
        RECT 4.000 390.680 199.115 391.320 ;
        RECT 4.000 390.000 195.600 390.680 ;
        RECT 4.400 389.280 195.600 390.000 ;
        RECT 4.400 388.640 199.115 389.280 ;
        RECT 4.400 388.600 195.600 388.640 ;
        RECT 4.000 387.240 195.600 388.600 ;
        RECT 4.000 386.600 199.115 387.240 ;
        RECT 4.000 385.920 195.600 386.600 ;
        RECT 4.400 385.200 195.600 385.920 ;
        RECT 4.400 384.520 199.115 385.200 ;
        RECT 4.000 383.880 199.115 384.520 ;
        RECT 4.000 382.480 195.600 383.880 ;
        RECT 4.000 381.840 199.115 382.480 ;
        RECT 4.400 380.440 195.600 381.840 ;
        RECT 4.000 379.800 199.115 380.440 ;
        RECT 4.000 378.400 195.600 379.800 ;
        RECT 4.000 377.760 199.115 378.400 ;
        RECT 4.400 377.080 199.115 377.760 ;
        RECT 4.400 376.360 195.600 377.080 ;
        RECT 4.000 375.680 195.600 376.360 ;
        RECT 4.000 375.040 199.115 375.680 ;
        RECT 4.000 373.680 195.600 375.040 ;
        RECT 4.400 373.640 195.600 373.680 ;
        RECT 4.400 373.000 199.115 373.640 ;
        RECT 4.400 372.280 195.600 373.000 ;
        RECT 4.000 371.600 195.600 372.280 ;
        RECT 4.000 370.960 199.115 371.600 ;
        RECT 4.000 369.600 195.600 370.960 ;
        RECT 4.400 369.560 195.600 369.600 ;
        RECT 4.400 368.240 199.115 369.560 ;
        RECT 4.400 368.200 195.600 368.240 ;
        RECT 4.000 366.840 195.600 368.200 ;
        RECT 4.000 366.200 199.115 366.840 ;
        RECT 4.400 364.800 195.600 366.200 ;
        RECT 4.000 364.160 199.115 364.800 ;
        RECT 4.000 362.760 195.600 364.160 ;
        RECT 4.000 362.120 199.115 362.760 ;
        RECT 4.400 361.440 199.115 362.120 ;
        RECT 4.400 360.720 195.600 361.440 ;
        RECT 4.000 360.040 195.600 360.720 ;
        RECT 4.000 359.400 199.115 360.040 ;
        RECT 4.000 358.040 195.600 359.400 ;
        RECT 4.400 358.000 195.600 358.040 ;
        RECT 4.400 357.360 199.115 358.000 ;
        RECT 4.400 356.640 195.600 357.360 ;
        RECT 4.000 355.960 195.600 356.640 ;
        RECT 4.000 354.640 199.115 355.960 ;
        RECT 4.000 353.960 195.600 354.640 ;
        RECT 4.400 353.240 195.600 353.960 ;
        RECT 4.400 352.600 199.115 353.240 ;
        RECT 4.400 352.560 195.600 352.600 ;
        RECT 4.000 351.200 195.600 352.560 ;
        RECT 4.000 350.560 199.115 351.200 ;
        RECT 4.000 349.880 195.600 350.560 ;
        RECT 4.400 349.160 195.600 349.880 ;
        RECT 4.400 348.520 199.115 349.160 ;
        RECT 4.400 348.480 195.600 348.520 ;
        RECT 4.000 347.120 195.600 348.480 ;
        RECT 4.000 345.800 199.115 347.120 ;
        RECT 4.400 344.400 195.600 345.800 ;
        RECT 4.000 343.760 199.115 344.400 ;
        RECT 4.000 342.360 195.600 343.760 ;
        RECT 4.000 341.720 199.115 342.360 ;
        RECT 4.400 340.320 195.600 341.720 ;
        RECT 4.000 339.000 199.115 340.320 ;
        RECT 4.000 337.640 195.600 339.000 ;
        RECT 4.400 337.600 195.600 337.640 ;
        RECT 4.400 336.960 199.115 337.600 ;
        RECT 4.400 336.240 195.600 336.960 ;
        RECT 4.000 335.560 195.600 336.240 ;
        RECT 4.000 334.920 199.115 335.560 ;
        RECT 4.000 334.240 195.600 334.920 ;
        RECT 4.400 333.520 195.600 334.240 ;
        RECT 4.400 332.880 199.115 333.520 ;
        RECT 4.400 332.840 195.600 332.880 ;
        RECT 4.000 331.480 195.600 332.840 ;
        RECT 4.000 330.160 199.115 331.480 ;
        RECT 4.400 328.760 195.600 330.160 ;
        RECT 4.000 328.120 199.115 328.760 ;
        RECT 4.000 326.720 195.600 328.120 ;
        RECT 4.000 326.080 199.115 326.720 ;
        RECT 4.400 324.680 195.600 326.080 ;
        RECT 4.000 323.360 199.115 324.680 ;
        RECT 4.000 322.000 195.600 323.360 ;
        RECT 4.400 321.960 195.600 322.000 ;
        RECT 4.400 321.320 199.115 321.960 ;
        RECT 4.400 320.600 195.600 321.320 ;
        RECT 4.000 319.920 195.600 320.600 ;
        RECT 4.000 319.280 199.115 319.920 ;
        RECT 4.000 317.920 195.600 319.280 ;
        RECT 4.400 317.880 195.600 317.920 ;
        RECT 4.400 317.240 199.115 317.880 ;
        RECT 4.400 316.520 195.600 317.240 ;
        RECT 4.000 315.840 195.600 316.520 ;
        RECT 4.000 314.520 199.115 315.840 ;
        RECT 4.000 313.840 195.600 314.520 ;
        RECT 4.400 313.120 195.600 313.840 ;
        RECT 4.400 312.480 199.115 313.120 ;
        RECT 4.400 312.440 195.600 312.480 ;
        RECT 4.000 311.080 195.600 312.440 ;
        RECT 4.000 310.440 199.115 311.080 ;
        RECT 4.000 309.760 195.600 310.440 ;
        RECT 4.400 309.040 195.600 309.760 ;
        RECT 4.400 308.360 199.115 309.040 ;
        RECT 4.000 307.720 199.115 308.360 ;
        RECT 4.000 306.320 195.600 307.720 ;
        RECT 4.000 305.680 199.115 306.320 ;
        RECT 4.400 304.280 195.600 305.680 ;
        RECT 4.000 303.640 199.115 304.280 ;
        RECT 4.000 302.280 195.600 303.640 ;
        RECT 4.400 302.240 195.600 302.280 ;
        RECT 4.400 301.600 199.115 302.240 ;
        RECT 4.400 300.880 195.600 301.600 ;
        RECT 4.000 300.200 195.600 300.880 ;
        RECT 4.000 298.880 199.115 300.200 ;
        RECT 4.000 298.200 195.600 298.880 ;
        RECT 4.400 297.480 195.600 298.200 ;
        RECT 4.400 296.840 199.115 297.480 ;
        RECT 4.400 296.800 195.600 296.840 ;
        RECT 4.000 295.440 195.600 296.800 ;
        RECT 4.000 294.800 199.115 295.440 ;
        RECT 4.000 294.120 195.600 294.800 ;
        RECT 4.400 293.400 195.600 294.120 ;
        RECT 4.400 292.720 199.115 293.400 ;
        RECT 4.000 292.080 199.115 292.720 ;
        RECT 4.000 290.680 195.600 292.080 ;
        RECT 4.000 290.040 199.115 290.680 ;
        RECT 4.400 288.640 195.600 290.040 ;
        RECT 4.000 288.000 199.115 288.640 ;
        RECT 4.000 286.600 195.600 288.000 ;
        RECT 4.000 285.960 199.115 286.600 ;
        RECT 4.400 285.280 199.115 285.960 ;
        RECT 4.400 284.560 195.600 285.280 ;
        RECT 4.000 283.880 195.600 284.560 ;
        RECT 4.000 283.240 199.115 283.880 ;
        RECT 4.000 281.880 195.600 283.240 ;
        RECT 4.400 281.840 195.600 281.880 ;
        RECT 4.400 281.200 199.115 281.840 ;
        RECT 4.400 280.480 195.600 281.200 ;
        RECT 4.000 279.800 195.600 280.480 ;
        RECT 4.000 279.160 199.115 279.800 ;
        RECT 4.000 277.800 195.600 279.160 ;
        RECT 4.400 277.760 195.600 277.800 ;
        RECT 4.400 276.440 199.115 277.760 ;
        RECT 4.400 276.400 195.600 276.440 ;
        RECT 4.000 275.040 195.600 276.400 ;
        RECT 4.000 274.400 199.115 275.040 ;
        RECT 4.000 273.720 195.600 274.400 ;
        RECT 4.400 273.000 195.600 273.720 ;
        RECT 4.400 272.360 199.115 273.000 ;
        RECT 4.400 272.320 195.600 272.360 ;
        RECT 4.000 270.960 195.600 272.320 ;
        RECT 4.000 269.640 199.115 270.960 ;
        RECT 4.400 268.240 195.600 269.640 ;
        RECT 4.000 267.600 199.115 268.240 ;
        RECT 4.000 266.240 195.600 267.600 ;
        RECT 4.400 266.200 195.600 266.240 ;
        RECT 4.400 265.560 199.115 266.200 ;
        RECT 4.400 264.840 195.600 265.560 ;
        RECT 4.000 264.160 195.600 264.840 ;
        RECT 4.000 263.520 199.115 264.160 ;
        RECT 4.000 262.160 195.600 263.520 ;
        RECT 4.400 262.120 195.600 262.160 ;
        RECT 4.400 260.800 199.115 262.120 ;
        RECT 4.400 260.760 195.600 260.800 ;
        RECT 4.000 259.400 195.600 260.760 ;
        RECT 4.000 258.760 199.115 259.400 ;
        RECT 4.000 258.080 195.600 258.760 ;
        RECT 4.400 257.360 195.600 258.080 ;
        RECT 4.400 256.720 199.115 257.360 ;
        RECT 4.400 256.680 195.600 256.720 ;
        RECT 4.000 255.320 195.600 256.680 ;
        RECT 4.000 254.000 199.115 255.320 ;
        RECT 4.400 252.600 195.600 254.000 ;
        RECT 4.000 251.960 199.115 252.600 ;
        RECT 4.000 250.560 195.600 251.960 ;
        RECT 4.000 249.920 199.115 250.560 ;
        RECT 4.400 248.520 195.600 249.920 ;
        RECT 4.000 247.880 199.115 248.520 ;
        RECT 4.000 246.480 195.600 247.880 ;
        RECT 4.000 245.840 199.115 246.480 ;
        RECT 4.400 245.160 199.115 245.840 ;
        RECT 4.400 244.440 195.600 245.160 ;
        RECT 4.000 243.760 195.600 244.440 ;
        RECT 4.000 243.120 199.115 243.760 ;
        RECT 4.000 241.760 195.600 243.120 ;
        RECT 4.400 241.720 195.600 241.760 ;
        RECT 4.400 241.080 199.115 241.720 ;
        RECT 4.400 240.360 195.600 241.080 ;
        RECT 4.000 239.680 195.600 240.360 ;
        RECT 4.000 238.360 199.115 239.680 ;
        RECT 4.000 237.680 195.600 238.360 ;
        RECT 4.400 236.960 195.600 237.680 ;
        RECT 4.400 236.320 199.115 236.960 ;
        RECT 4.400 236.280 195.600 236.320 ;
        RECT 4.000 234.920 195.600 236.280 ;
        RECT 4.000 234.280 199.115 234.920 ;
        RECT 4.400 232.880 195.600 234.280 ;
        RECT 4.000 231.560 199.115 232.880 ;
        RECT 4.000 230.200 195.600 231.560 ;
        RECT 4.400 230.160 195.600 230.200 ;
        RECT 4.400 229.520 199.115 230.160 ;
        RECT 4.400 228.800 195.600 229.520 ;
        RECT 4.000 228.120 195.600 228.800 ;
        RECT 4.000 227.480 199.115 228.120 ;
        RECT 4.000 226.120 195.600 227.480 ;
        RECT 4.400 226.080 195.600 226.120 ;
        RECT 4.400 225.440 199.115 226.080 ;
        RECT 4.400 224.720 195.600 225.440 ;
        RECT 4.000 224.040 195.600 224.720 ;
        RECT 4.000 222.720 199.115 224.040 ;
        RECT 4.000 222.040 195.600 222.720 ;
        RECT 4.400 221.320 195.600 222.040 ;
        RECT 4.400 220.680 199.115 221.320 ;
        RECT 4.400 220.640 195.600 220.680 ;
        RECT 4.000 219.280 195.600 220.640 ;
        RECT 4.000 218.640 199.115 219.280 ;
        RECT 4.000 217.960 195.600 218.640 ;
        RECT 4.400 217.240 195.600 217.960 ;
        RECT 4.400 216.560 199.115 217.240 ;
        RECT 4.000 215.920 199.115 216.560 ;
        RECT 4.000 214.520 195.600 215.920 ;
        RECT 4.000 213.880 199.115 214.520 ;
        RECT 4.400 212.480 195.600 213.880 ;
        RECT 4.000 211.840 199.115 212.480 ;
        RECT 4.000 210.440 195.600 211.840 ;
        RECT 4.000 209.800 199.115 210.440 ;
        RECT 4.400 208.400 195.600 209.800 ;
        RECT 4.000 207.080 199.115 208.400 ;
        RECT 4.000 205.720 195.600 207.080 ;
        RECT 4.400 205.680 195.600 205.720 ;
        RECT 4.400 205.040 199.115 205.680 ;
        RECT 4.400 204.320 195.600 205.040 ;
        RECT 4.000 203.640 195.600 204.320 ;
        RECT 4.000 203.000 199.115 203.640 ;
        RECT 4.000 202.320 195.600 203.000 ;
        RECT 4.400 201.600 195.600 202.320 ;
        RECT 4.400 200.920 199.115 201.600 ;
        RECT 4.000 200.280 199.115 200.920 ;
        RECT 4.000 198.880 195.600 200.280 ;
        RECT 4.000 198.240 199.115 198.880 ;
        RECT 4.400 196.840 195.600 198.240 ;
        RECT 4.000 196.200 199.115 196.840 ;
        RECT 4.000 194.800 195.600 196.200 ;
        RECT 4.000 194.160 199.115 194.800 ;
        RECT 4.400 192.760 195.600 194.160 ;
        RECT 4.000 191.440 199.115 192.760 ;
        RECT 4.000 190.080 195.600 191.440 ;
        RECT 4.400 190.040 195.600 190.080 ;
        RECT 4.400 189.400 199.115 190.040 ;
        RECT 4.400 188.680 195.600 189.400 ;
        RECT 4.000 188.000 195.600 188.680 ;
        RECT 4.000 187.360 199.115 188.000 ;
        RECT 4.000 186.000 195.600 187.360 ;
        RECT 4.400 185.960 195.600 186.000 ;
        RECT 4.400 184.640 199.115 185.960 ;
        RECT 4.400 184.600 195.600 184.640 ;
        RECT 4.000 183.240 195.600 184.600 ;
        RECT 4.000 182.600 199.115 183.240 ;
        RECT 4.000 181.920 195.600 182.600 ;
        RECT 4.400 181.200 195.600 181.920 ;
        RECT 4.400 180.560 199.115 181.200 ;
        RECT 4.400 180.520 195.600 180.560 ;
        RECT 4.000 179.160 195.600 180.520 ;
        RECT 4.000 177.840 199.115 179.160 ;
        RECT 4.400 176.440 195.600 177.840 ;
        RECT 4.000 175.800 199.115 176.440 ;
        RECT 4.000 174.400 195.600 175.800 ;
        RECT 4.000 173.760 199.115 174.400 ;
        RECT 4.400 172.360 195.600 173.760 ;
        RECT 4.000 171.720 199.115 172.360 ;
        RECT 4.000 170.320 195.600 171.720 ;
        RECT 4.000 169.680 199.115 170.320 ;
        RECT 4.400 169.000 199.115 169.680 ;
        RECT 4.400 168.280 195.600 169.000 ;
        RECT 4.000 167.600 195.600 168.280 ;
        RECT 4.000 166.960 199.115 167.600 ;
        RECT 4.000 166.280 195.600 166.960 ;
        RECT 4.400 165.560 195.600 166.280 ;
        RECT 4.400 164.920 199.115 165.560 ;
        RECT 4.400 164.880 195.600 164.920 ;
        RECT 4.000 163.520 195.600 164.880 ;
        RECT 4.000 162.200 199.115 163.520 ;
        RECT 4.400 160.800 195.600 162.200 ;
        RECT 4.000 160.160 199.115 160.800 ;
        RECT 4.000 158.760 195.600 160.160 ;
        RECT 4.000 158.120 199.115 158.760 ;
        RECT 4.400 156.720 195.600 158.120 ;
        RECT 4.000 156.080 199.115 156.720 ;
        RECT 4.000 154.680 195.600 156.080 ;
        RECT 4.000 154.040 199.115 154.680 ;
        RECT 4.400 153.360 199.115 154.040 ;
        RECT 4.400 152.640 195.600 153.360 ;
        RECT 4.000 151.960 195.600 152.640 ;
        RECT 4.000 151.320 199.115 151.960 ;
        RECT 4.000 149.960 195.600 151.320 ;
        RECT 4.400 149.920 195.600 149.960 ;
        RECT 4.400 149.280 199.115 149.920 ;
        RECT 4.400 148.560 195.600 149.280 ;
        RECT 4.000 147.880 195.600 148.560 ;
        RECT 4.000 146.560 199.115 147.880 ;
        RECT 4.000 145.880 195.600 146.560 ;
        RECT 4.400 145.160 195.600 145.880 ;
        RECT 4.400 144.520 199.115 145.160 ;
        RECT 4.400 144.480 195.600 144.520 ;
        RECT 4.000 143.120 195.600 144.480 ;
        RECT 4.000 142.480 199.115 143.120 ;
        RECT 4.000 141.800 195.600 142.480 ;
        RECT 4.400 141.080 195.600 141.800 ;
        RECT 4.400 140.440 199.115 141.080 ;
        RECT 4.400 140.400 195.600 140.440 ;
        RECT 4.000 139.040 195.600 140.400 ;
        RECT 4.000 137.720 199.115 139.040 ;
        RECT 4.400 136.320 195.600 137.720 ;
        RECT 4.000 135.680 199.115 136.320 ;
        RECT 4.000 134.320 195.600 135.680 ;
        RECT 4.400 134.280 195.600 134.320 ;
        RECT 4.400 133.640 199.115 134.280 ;
        RECT 4.400 132.920 195.600 133.640 ;
        RECT 4.000 132.240 195.600 132.920 ;
        RECT 4.000 130.920 199.115 132.240 ;
        RECT 4.000 130.240 195.600 130.920 ;
        RECT 4.400 129.520 195.600 130.240 ;
        RECT 4.400 128.880 199.115 129.520 ;
        RECT 4.400 128.840 195.600 128.880 ;
        RECT 4.000 127.480 195.600 128.840 ;
        RECT 4.000 126.840 199.115 127.480 ;
        RECT 4.000 126.160 195.600 126.840 ;
        RECT 4.400 125.440 195.600 126.160 ;
        RECT 4.400 124.800 199.115 125.440 ;
        RECT 4.400 124.760 195.600 124.800 ;
        RECT 4.000 123.400 195.600 124.760 ;
        RECT 4.000 122.080 199.115 123.400 ;
        RECT 4.400 120.680 195.600 122.080 ;
        RECT 4.000 120.040 199.115 120.680 ;
        RECT 4.000 118.640 195.600 120.040 ;
        RECT 4.000 118.000 199.115 118.640 ;
        RECT 4.400 116.600 195.600 118.000 ;
        RECT 4.000 115.280 199.115 116.600 ;
        RECT 4.000 113.920 195.600 115.280 ;
        RECT 4.400 113.880 195.600 113.920 ;
        RECT 4.400 113.240 199.115 113.880 ;
        RECT 4.400 112.520 195.600 113.240 ;
        RECT 4.000 111.840 195.600 112.520 ;
        RECT 4.000 111.200 199.115 111.840 ;
        RECT 4.000 109.840 195.600 111.200 ;
        RECT 4.400 109.800 195.600 109.840 ;
        RECT 4.400 108.480 199.115 109.800 ;
        RECT 4.400 108.440 195.600 108.480 ;
        RECT 4.000 107.080 195.600 108.440 ;
        RECT 4.000 106.440 199.115 107.080 ;
        RECT 4.000 105.760 195.600 106.440 ;
        RECT 4.400 105.040 195.600 105.760 ;
        RECT 4.400 104.400 199.115 105.040 ;
        RECT 4.400 104.360 195.600 104.400 ;
        RECT 4.000 103.000 195.600 104.360 ;
        RECT 4.000 102.360 199.115 103.000 ;
        RECT 4.400 100.960 195.600 102.360 ;
        RECT 4.000 99.640 199.115 100.960 ;
        RECT 4.000 98.280 195.600 99.640 ;
        RECT 4.400 98.240 195.600 98.280 ;
        RECT 4.400 97.600 199.115 98.240 ;
        RECT 4.400 96.880 195.600 97.600 ;
        RECT 4.000 96.200 195.600 96.880 ;
        RECT 4.000 95.560 199.115 96.200 ;
        RECT 4.000 94.200 195.600 95.560 ;
        RECT 4.400 94.160 195.600 94.200 ;
        RECT 4.400 92.840 199.115 94.160 ;
        RECT 4.400 92.800 195.600 92.840 ;
        RECT 4.000 91.440 195.600 92.800 ;
        RECT 4.000 90.800 199.115 91.440 ;
        RECT 4.000 90.120 195.600 90.800 ;
        RECT 4.400 89.400 195.600 90.120 ;
        RECT 4.400 88.760 199.115 89.400 ;
        RECT 4.400 88.720 195.600 88.760 ;
        RECT 4.000 87.360 195.600 88.720 ;
        RECT 4.000 86.720 199.115 87.360 ;
        RECT 4.000 86.040 195.600 86.720 ;
        RECT 4.400 85.320 195.600 86.040 ;
        RECT 4.400 84.640 199.115 85.320 ;
        RECT 4.000 84.000 199.115 84.640 ;
        RECT 4.000 82.600 195.600 84.000 ;
        RECT 4.000 81.960 199.115 82.600 ;
        RECT 4.400 80.560 195.600 81.960 ;
        RECT 4.000 79.920 199.115 80.560 ;
        RECT 4.000 78.520 195.600 79.920 ;
        RECT 4.000 77.880 199.115 78.520 ;
        RECT 4.400 77.200 199.115 77.880 ;
        RECT 4.400 76.480 195.600 77.200 ;
        RECT 4.000 75.800 195.600 76.480 ;
        RECT 4.000 75.160 199.115 75.800 ;
        RECT 4.000 73.800 195.600 75.160 ;
        RECT 4.400 73.760 195.600 73.800 ;
        RECT 4.400 73.120 199.115 73.760 ;
        RECT 4.400 72.400 195.600 73.120 ;
        RECT 4.000 71.720 195.600 72.400 ;
        RECT 4.000 71.080 199.115 71.720 ;
        RECT 4.000 69.720 195.600 71.080 ;
        RECT 4.400 69.680 195.600 69.720 ;
        RECT 4.400 68.360 199.115 69.680 ;
        RECT 4.400 68.320 195.600 68.360 ;
        RECT 4.000 66.960 195.600 68.320 ;
        RECT 4.000 66.320 199.115 66.960 ;
        RECT 4.400 64.920 195.600 66.320 ;
        RECT 4.000 64.280 199.115 64.920 ;
        RECT 4.000 62.880 195.600 64.280 ;
        RECT 4.000 62.240 199.115 62.880 ;
        RECT 4.400 61.560 199.115 62.240 ;
        RECT 4.400 60.840 195.600 61.560 ;
        RECT 4.000 60.160 195.600 60.840 ;
        RECT 4.000 59.520 199.115 60.160 ;
        RECT 4.000 58.160 195.600 59.520 ;
        RECT 4.400 58.120 195.600 58.160 ;
        RECT 4.400 57.480 199.115 58.120 ;
        RECT 4.400 56.760 195.600 57.480 ;
        RECT 4.000 56.080 195.600 56.760 ;
        RECT 4.000 54.760 199.115 56.080 ;
        RECT 4.000 54.080 195.600 54.760 ;
        RECT 4.400 53.360 195.600 54.080 ;
        RECT 4.400 52.720 199.115 53.360 ;
        RECT 4.400 52.680 195.600 52.720 ;
        RECT 4.000 51.320 195.600 52.680 ;
        RECT 4.000 50.680 199.115 51.320 ;
        RECT 4.000 50.000 195.600 50.680 ;
        RECT 4.400 49.280 195.600 50.000 ;
        RECT 4.400 48.640 199.115 49.280 ;
        RECT 4.400 48.600 195.600 48.640 ;
        RECT 4.000 47.240 195.600 48.600 ;
        RECT 4.000 45.920 199.115 47.240 ;
        RECT 4.400 44.520 195.600 45.920 ;
        RECT 4.000 43.880 199.115 44.520 ;
        RECT 4.000 42.480 195.600 43.880 ;
        RECT 4.000 41.840 199.115 42.480 ;
        RECT 4.400 40.440 195.600 41.840 ;
        RECT 4.000 39.120 199.115 40.440 ;
        RECT 4.000 37.760 195.600 39.120 ;
        RECT 4.400 37.720 195.600 37.760 ;
        RECT 4.400 37.080 199.115 37.720 ;
        RECT 4.400 36.360 195.600 37.080 ;
        RECT 4.000 35.680 195.600 36.360 ;
        RECT 4.000 35.040 199.115 35.680 ;
        RECT 4.000 34.360 195.600 35.040 ;
        RECT 4.400 33.640 195.600 34.360 ;
        RECT 4.400 33.000 199.115 33.640 ;
        RECT 4.400 32.960 195.600 33.000 ;
        RECT 4.000 31.600 195.600 32.960 ;
        RECT 4.000 30.280 199.115 31.600 ;
        RECT 4.400 28.880 195.600 30.280 ;
        RECT 4.000 28.240 199.115 28.880 ;
        RECT 4.000 26.840 195.600 28.240 ;
        RECT 4.000 26.200 199.115 26.840 ;
        RECT 4.400 24.800 195.600 26.200 ;
        RECT 4.000 23.480 199.115 24.800 ;
        RECT 4.000 22.120 195.600 23.480 ;
        RECT 4.400 22.080 195.600 22.120 ;
        RECT 4.400 21.440 199.115 22.080 ;
        RECT 4.400 20.720 195.600 21.440 ;
        RECT 4.000 20.040 195.600 20.720 ;
        RECT 4.000 19.400 199.115 20.040 ;
        RECT 4.000 18.040 195.600 19.400 ;
        RECT 4.400 18.000 195.600 18.040 ;
        RECT 4.400 17.360 199.115 18.000 ;
        RECT 4.400 16.640 195.600 17.360 ;
        RECT 4.000 15.960 195.600 16.640 ;
        RECT 4.000 14.640 199.115 15.960 ;
        RECT 4.000 13.960 195.600 14.640 ;
        RECT 4.400 13.240 195.600 13.960 ;
        RECT 4.400 12.600 199.115 13.240 ;
        RECT 4.400 12.560 195.600 12.600 ;
        RECT 4.000 11.200 195.600 12.560 ;
        RECT 4.000 10.560 199.115 11.200 ;
        RECT 4.000 9.880 195.600 10.560 ;
        RECT 4.400 9.160 195.600 9.880 ;
        RECT 4.400 8.480 199.115 9.160 ;
        RECT 4.000 7.840 199.115 8.480 ;
        RECT 4.000 6.440 195.600 7.840 ;
        RECT 4.000 5.800 199.115 6.440 ;
        RECT 4.400 4.400 195.600 5.800 ;
        RECT 4.000 3.760 199.115 4.400 ;
        RECT 4.000 2.400 195.600 3.760 ;
        RECT 4.400 2.360 195.600 2.400 ;
        RECT 4.400 1.720 199.115 2.360 ;
        RECT 4.400 1.000 195.600 1.720 ;
        RECT 4.000 0.855 195.600 1.000 ;
  END
END wb_local
END LIBRARY

