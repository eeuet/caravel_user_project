magic
tech sky130A
magscale 1 2
timestamp 1623880163
<< obsli1 >>
rect 1104 2159 29043 53329
<< obsm1 >>
rect 658 1028 29334 54052
<< metal2 >>
rect 846 55200 902 56800
rect 2594 55200 2650 56800
rect 4342 55200 4398 56800
rect 6090 55200 6146 56800
rect 7838 55200 7894 56800
rect 9586 55200 9642 56800
rect 11426 55200 11482 56800
rect 13174 55200 13230 56800
rect 14922 55200 14978 56800
rect 16670 55200 16726 56800
rect 18418 55200 18474 56800
rect 20166 55200 20222 56800
rect 22006 55200 22062 56800
rect 23754 55200 23810 56800
rect 25502 55200 25558 56800
rect 27250 55200 27306 56800
rect 28998 55200 29054 56800
rect 662 -800 718 800
rect 1950 -800 2006 800
rect 3330 -800 3386 800
rect 4710 -800 4766 800
rect 6090 -800 6146 800
rect 7470 -800 7526 800
rect 8758 -800 8814 800
rect 10138 -800 10194 800
rect 11518 -800 11574 800
rect 12898 -800 12954 800
rect 14278 -800 14334 800
rect 15658 -800 15714 800
rect 16946 -800 17002 800
rect 18326 -800 18382 800
rect 19706 -800 19762 800
rect 21086 -800 21142 800
rect 22466 -800 22522 800
rect 23754 -800 23810 800
rect 25134 -800 25190 800
rect 26514 -800 26570 800
rect 27894 -800 27950 800
rect 29274 -800 29330 800
<< obsm2 >>
rect 664 55144 790 55729
rect 958 55144 2538 55729
rect 2706 55144 4286 55729
rect 4454 55144 6034 55729
rect 6202 55144 7782 55729
rect 7950 55144 9530 55729
rect 9698 55144 11370 55729
rect 11538 55144 13118 55729
rect 13286 55144 14866 55729
rect 15034 55144 16614 55729
rect 16782 55144 18362 55729
rect 18530 55144 20110 55729
rect 20278 55144 21950 55729
rect 22118 55144 23698 55729
rect 23866 55144 25446 55729
rect 25614 55144 27194 55729
rect 27362 55144 28942 55729
rect 29110 55144 29328 55729
rect 664 856 29328 55144
rect 774 167 1894 856
rect 2062 167 3274 856
rect 3442 167 4654 856
rect 4822 167 6034 856
rect 6202 167 7414 856
rect 7582 167 8702 856
rect 8870 167 10082 856
rect 10250 167 11462 856
rect 11630 167 12842 856
rect 13010 167 14222 856
rect 14390 167 15602 856
rect 15770 167 16890 856
rect 17058 167 18270 856
rect 18438 167 19650 856
rect 19818 167 21030 856
rect 21198 167 22410 856
rect 22578 167 23698 856
rect 23866 167 25078 856
rect 25246 167 26458 856
rect 26626 167 27838 856
rect 28006 167 29218 856
<< metal3 >>
rect -800 55632 800 55752
rect 29200 55632 30800 55752
rect -800 55224 800 55344
rect 29200 55224 30800 55344
rect -800 54816 800 54936
rect 29200 54816 30800 54936
rect -800 54408 800 54528
rect 29200 54408 30800 54528
rect -800 54000 800 54120
rect 29200 54000 30800 54120
rect -800 53592 800 53712
rect 29200 53592 30800 53712
rect -800 53184 800 53304
rect 29200 53184 30800 53304
rect -800 52776 800 52896
rect 29200 52776 30800 52896
rect -800 52368 800 52488
rect 29200 52368 30800 52488
rect -800 51960 800 52080
rect 29200 51960 30800 52080
rect -800 51552 800 51672
rect 29200 51552 30800 51672
rect -800 51144 800 51264
rect 29200 51144 30800 51264
rect -800 50736 800 50856
rect 29200 50736 30800 50856
rect -800 50328 800 50448
rect 29200 50328 30800 50448
rect -800 49920 800 50040
rect 29200 49920 30800 50040
rect -800 49512 800 49632
rect 29200 49512 30800 49632
rect -800 49104 800 49224
rect 29200 49104 30800 49224
rect -800 48696 800 48816
rect 29200 48696 30800 48816
rect -800 48288 800 48408
rect 29200 48288 30800 48408
rect -800 47880 800 48000
rect 29200 47880 30800 48000
rect -800 47472 800 47592
rect 29200 47472 30800 47592
rect -800 47064 800 47184
rect 29200 47064 30800 47184
rect -800 46656 800 46776
rect 29200 46656 30800 46776
rect -800 46248 800 46368
rect 29200 46248 30800 46368
rect -800 45840 800 45960
rect 29200 45840 30800 45960
rect -800 45432 800 45552
rect 29200 45432 30800 45552
rect -800 45024 800 45144
rect 29200 45024 30800 45144
rect -800 44616 800 44736
rect 29200 44616 30800 44736
rect -800 44208 800 44328
rect 29200 44208 30800 44328
rect -800 43800 800 43920
rect 29200 43800 30800 43920
rect -800 43392 800 43512
rect 29200 43392 30800 43512
rect -800 42984 800 43104
rect 29200 42984 30800 43104
rect -800 42576 800 42696
rect 29200 42576 30800 42696
rect -800 42168 800 42288
rect 29200 42168 30800 42288
rect -800 41760 800 41880
rect 29200 41760 30800 41880
rect -800 41352 800 41472
rect 29200 41352 30800 41472
rect -800 40944 800 41064
rect 29200 40944 30800 41064
rect -800 40536 800 40656
rect 29200 40536 30800 40656
rect -800 40128 800 40248
rect 29200 40128 30800 40248
rect -800 39720 800 39840
rect 29200 39720 30800 39840
rect -800 39312 800 39432
rect 29200 39312 30800 39432
rect -800 38904 800 39024
rect 29200 38904 30800 39024
rect -800 38496 800 38616
rect 29200 38496 30800 38616
rect -800 38088 800 38208
rect 29200 38088 30800 38208
rect -800 37680 800 37800
rect 29200 37680 30800 37800
rect -800 37272 800 37392
rect 29200 37272 30800 37392
rect -800 36864 800 36984
rect 29200 36864 30800 36984
rect -800 36456 800 36576
rect 29200 36456 30800 36576
rect -800 36048 800 36168
rect 29200 36048 30800 36168
rect -800 35640 800 35760
rect 29200 35640 30800 35760
rect -800 35232 800 35352
rect 29200 35232 30800 35352
rect -800 34824 800 34944
rect 29200 34824 30800 34944
rect -800 34416 800 34536
rect 29200 34416 30800 34536
rect -800 34008 800 34128
rect 29200 34008 30800 34128
rect -800 33600 800 33720
rect 29200 33600 30800 33720
rect -800 33192 800 33312
rect 29200 33192 30800 33312
rect -800 32784 800 32904
rect 29200 32784 30800 32904
rect -800 32376 800 32496
rect 29200 32376 30800 32496
rect -800 31968 800 32088
rect 29200 31968 30800 32088
rect -800 31560 800 31680
rect 29200 31560 30800 31680
rect -800 31152 800 31272
rect 29200 31152 30800 31272
rect -800 30744 800 30864
rect 29200 30744 30800 30864
rect -800 30336 800 30456
rect 29200 30336 30800 30456
rect -800 29928 800 30048
rect 29200 29928 30800 30048
rect -800 29520 800 29640
rect 29200 29520 30800 29640
rect -800 29112 800 29232
rect 29200 29112 30800 29232
rect -800 28704 800 28824
rect 29200 28704 30800 28824
rect -800 28296 800 28416
rect 29200 28296 30800 28416
rect -800 27888 800 28008
rect 29200 27888 30800 28008
rect -800 27480 800 27600
rect 29200 27480 30800 27600
rect -800 27072 800 27192
rect 29200 27072 30800 27192
rect -800 26664 800 26784
rect 29200 26664 30800 26784
rect -800 26256 800 26376
rect 29200 26256 30800 26376
rect -800 25848 800 25968
rect 29200 25848 30800 25968
rect -800 25440 800 25560
rect 29200 25440 30800 25560
rect -800 25032 800 25152
rect 29200 25032 30800 25152
rect -800 24624 800 24744
rect 29200 24624 30800 24744
rect -800 24216 800 24336
rect 29200 24216 30800 24336
rect -800 23808 800 23928
rect 29200 23808 30800 23928
rect -800 23400 800 23520
rect 29200 23400 30800 23520
rect -800 22992 800 23112
rect 29200 22992 30800 23112
rect -800 22584 800 22704
rect 29200 22584 30800 22704
rect -800 22176 800 22296
rect 29200 22176 30800 22296
rect -800 21768 800 21888
rect 29200 21768 30800 21888
rect -800 21360 800 21480
rect 29200 21360 30800 21480
rect -800 20952 800 21072
rect 29200 20952 30800 21072
rect -800 20544 800 20664
rect 29200 20544 30800 20664
rect -800 20136 800 20256
rect 29200 20136 30800 20256
rect -800 19728 800 19848
rect 29200 19728 30800 19848
rect -800 19320 800 19440
rect 29200 19320 30800 19440
rect -800 18912 800 19032
rect 29200 18912 30800 19032
rect -800 18504 800 18624
rect 29200 18504 30800 18624
rect -800 18096 800 18216
rect 29200 18096 30800 18216
rect -800 17688 800 17808
rect 29200 17688 30800 17808
rect -800 17280 800 17400
rect 29200 17280 30800 17400
rect -800 16872 800 16992
rect 29200 16872 30800 16992
rect -800 16464 800 16584
rect 29200 16464 30800 16584
rect -800 16056 800 16176
rect 29200 16056 30800 16176
rect -800 15648 800 15768
rect 29200 15648 30800 15768
rect -800 15240 800 15360
rect 29200 15240 30800 15360
rect -800 14832 800 14952
rect 29200 14832 30800 14952
rect -800 14424 800 14544
rect 29200 14424 30800 14544
rect -800 14016 800 14136
rect 29200 14016 30800 14136
rect -800 13608 800 13728
rect 29200 13608 30800 13728
rect -800 13200 800 13320
rect 29200 13200 30800 13320
rect -800 12792 800 12912
rect 29200 12792 30800 12912
rect -800 12384 800 12504
rect 29200 12384 30800 12504
rect -800 11976 800 12096
rect 29200 11976 30800 12096
rect -800 11568 800 11688
rect 29200 11568 30800 11688
rect -800 11160 800 11280
rect 29200 11160 30800 11280
rect -800 10752 800 10872
rect 29200 10752 30800 10872
rect -800 10344 800 10464
rect 29200 10344 30800 10464
rect -800 9936 800 10056
rect 29200 9936 30800 10056
rect -800 9528 800 9648
rect 29200 9528 30800 9648
rect -800 9120 800 9240
rect 29200 9120 30800 9240
rect -800 8712 800 8832
rect 29200 8712 30800 8832
rect -800 8304 800 8424
rect 29200 8304 30800 8424
rect -800 7896 800 8016
rect 29200 7896 30800 8016
rect -800 7488 800 7608
rect 29200 7488 30800 7608
rect -800 7080 800 7200
rect 29200 7080 30800 7200
rect -800 6672 800 6792
rect 29200 6672 30800 6792
rect -800 6264 800 6384
rect 29200 6264 30800 6384
rect -800 5856 800 5976
rect 29200 5856 30800 5976
rect -800 5448 800 5568
rect 29200 5448 30800 5568
rect -800 5040 800 5160
rect 29200 5040 30800 5160
rect -800 4632 800 4752
rect 29200 4632 30800 4752
rect -800 4224 800 4344
rect 29200 4224 30800 4344
rect -800 3816 800 3936
rect 29200 3816 30800 3936
rect -800 3408 800 3528
rect 29200 3408 30800 3528
rect -800 3000 800 3120
rect 29200 3000 30800 3120
rect -800 2592 800 2712
rect 29200 2592 30800 2712
rect -800 2184 800 2304
rect 29200 2184 30800 2304
rect -800 1776 800 1896
rect 29200 1776 30800 1896
rect -800 1368 800 1488
rect 29200 1368 30800 1488
rect -800 960 800 1080
rect 29200 960 30800 1080
rect -800 552 800 672
rect 29200 552 30800 672
rect -800 144 800 264
rect 29200 144 30800 264
<< obsm3 >>
rect 880 55552 29120 55725
rect 800 55424 29200 55552
rect 880 55144 29120 55424
rect 800 55016 29200 55144
rect 880 54736 29120 55016
rect 800 54608 29200 54736
rect 880 54328 29120 54608
rect 800 54200 29200 54328
rect 880 53920 29120 54200
rect 800 53792 29200 53920
rect 880 53512 29120 53792
rect 800 53384 29200 53512
rect 880 53104 29120 53384
rect 800 52976 29200 53104
rect 880 52696 29120 52976
rect 800 52568 29200 52696
rect 880 52288 29120 52568
rect 800 52160 29200 52288
rect 880 51880 29120 52160
rect 800 51752 29200 51880
rect 880 51472 29120 51752
rect 800 51344 29200 51472
rect 880 51064 29120 51344
rect 800 50936 29200 51064
rect 880 50656 29120 50936
rect 800 50528 29200 50656
rect 880 50248 29120 50528
rect 800 50120 29200 50248
rect 880 49840 29120 50120
rect 800 49712 29200 49840
rect 880 49432 29120 49712
rect 800 49304 29200 49432
rect 880 49024 29120 49304
rect 800 48896 29200 49024
rect 880 48616 29120 48896
rect 800 48488 29200 48616
rect 880 48208 29120 48488
rect 800 48080 29200 48208
rect 880 47800 29120 48080
rect 800 47672 29200 47800
rect 880 47392 29120 47672
rect 800 47264 29200 47392
rect 880 46984 29120 47264
rect 800 46856 29200 46984
rect 880 46576 29120 46856
rect 800 46448 29200 46576
rect 880 46168 29120 46448
rect 800 46040 29200 46168
rect 880 45760 29120 46040
rect 800 45632 29200 45760
rect 880 45352 29120 45632
rect 800 45224 29200 45352
rect 880 44944 29120 45224
rect 800 44816 29200 44944
rect 880 44536 29120 44816
rect 800 44408 29200 44536
rect 880 44128 29120 44408
rect 800 44000 29200 44128
rect 880 43720 29120 44000
rect 800 43592 29200 43720
rect 880 43312 29120 43592
rect 800 43184 29200 43312
rect 880 42904 29120 43184
rect 800 42776 29200 42904
rect 880 42496 29120 42776
rect 800 42368 29200 42496
rect 880 42088 29120 42368
rect 800 41960 29200 42088
rect 880 41680 29120 41960
rect 800 41552 29200 41680
rect 880 41272 29120 41552
rect 800 41144 29200 41272
rect 880 40864 29120 41144
rect 800 40736 29200 40864
rect 880 40456 29120 40736
rect 800 40328 29200 40456
rect 880 40048 29120 40328
rect 800 39920 29200 40048
rect 880 39640 29120 39920
rect 800 39512 29200 39640
rect 880 39232 29120 39512
rect 800 39104 29200 39232
rect 880 38824 29120 39104
rect 800 38696 29200 38824
rect 880 38416 29120 38696
rect 800 38288 29200 38416
rect 880 38008 29120 38288
rect 800 37880 29200 38008
rect 880 37600 29120 37880
rect 800 37472 29200 37600
rect 880 37192 29120 37472
rect 800 37064 29200 37192
rect 880 36784 29120 37064
rect 800 36656 29200 36784
rect 880 36376 29120 36656
rect 800 36248 29200 36376
rect 880 35968 29120 36248
rect 800 35840 29200 35968
rect 880 35560 29120 35840
rect 800 35432 29200 35560
rect 880 35152 29120 35432
rect 800 35024 29200 35152
rect 880 34744 29120 35024
rect 800 34616 29200 34744
rect 880 34336 29120 34616
rect 800 34208 29200 34336
rect 880 33928 29120 34208
rect 800 33800 29200 33928
rect 880 33520 29120 33800
rect 800 33392 29200 33520
rect 880 33112 29120 33392
rect 800 32984 29200 33112
rect 880 32704 29120 32984
rect 800 32576 29200 32704
rect 880 32296 29120 32576
rect 800 32168 29200 32296
rect 880 31888 29120 32168
rect 800 31760 29200 31888
rect 880 31480 29120 31760
rect 800 31352 29200 31480
rect 880 31072 29120 31352
rect 800 30944 29200 31072
rect 880 30664 29120 30944
rect 800 30536 29200 30664
rect 880 30256 29120 30536
rect 800 30128 29200 30256
rect 880 29848 29120 30128
rect 800 29720 29200 29848
rect 880 29440 29120 29720
rect 800 29312 29200 29440
rect 880 29032 29120 29312
rect 800 28904 29200 29032
rect 880 28624 29120 28904
rect 800 28496 29200 28624
rect 880 28216 29120 28496
rect 800 28088 29200 28216
rect 880 27808 29120 28088
rect 800 27680 29200 27808
rect 880 27400 29120 27680
rect 800 27272 29200 27400
rect 880 26992 29120 27272
rect 800 26864 29200 26992
rect 880 26584 29120 26864
rect 800 26456 29200 26584
rect 880 26176 29120 26456
rect 800 26048 29200 26176
rect 880 25768 29120 26048
rect 800 25640 29200 25768
rect 880 25360 29120 25640
rect 800 25232 29200 25360
rect 880 24952 29120 25232
rect 800 24824 29200 24952
rect 880 24544 29120 24824
rect 800 24416 29200 24544
rect 880 24136 29120 24416
rect 800 24008 29200 24136
rect 880 23728 29120 24008
rect 800 23600 29200 23728
rect 880 23320 29120 23600
rect 800 23192 29200 23320
rect 880 22912 29120 23192
rect 800 22784 29200 22912
rect 880 22504 29120 22784
rect 800 22376 29200 22504
rect 880 22096 29120 22376
rect 800 21968 29200 22096
rect 880 21688 29120 21968
rect 800 21560 29200 21688
rect 880 21280 29120 21560
rect 800 21152 29200 21280
rect 880 20872 29120 21152
rect 800 20744 29200 20872
rect 880 20464 29120 20744
rect 800 20336 29200 20464
rect 880 20056 29120 20336
rect 800 19928 29200 20056
rect 880 19648 29120 19928
rect 800 19520 29200 19648
rect 880 19240 29120 19520
rect 800 19112 29200 19240
rect 880 18832 29120 19112
rect 800 18704 29200 18832
rect 880 18424 29120 18704
rect 800 18296 29200 18424
rect 880 18016 29120 18296
rect 800 17888 29200 18016
rect 880 17608 29120 17888
rect 800 17480 29200 17608
rect 880 17200 29120 17480
rect 800 17072 29200 17200
rect 880 16792 29120 17072
rect 800 16664 29200 16792
rect 880 16384 29120 16664
rect 800 16256 29200 16384
rect 880 15976 29120 16256
rect 800 15848 29200 15976
rect 880 15568 29120 15848
rect 800 15440 29200 15568
rect 880 15160 29120 15440
rect 800 15032 29200 15160
rect 880 14752 29120 15032
rect 800 14624 29200 14752
rect 880 14344 29120 14624
rect 800 14216 29200 14344
rect 880 13936 29120 14216
rect 800 13808 29200 13936
rect 880 13528 29120 13808
rect 800 13400 29200 13528
rect 880 13120 29120 13400
rect 800 12992 29200 13120
rect 880 12712 29120 12992
rect 800 12584 29200 12712
rect 880 12304 29120 12584
rect 800 12176 29200 12304
rect 880 11896 29120 12176
rect 800 11768 29200 11896
rect 880 11488 29120 11768
rect 800 11360 29200 11488
rect 880 11080 29120 11360
rect 800 10952 29200 11080
rect 880 10672 29120 10952
rect 800 10544 29200 10672
rect 880 10264 29120 10544
rect 800 10136 29200 10264
rect 880 9856 29120 10136
rect 800 9728 29200 9856
rect 880 9448 29120 9728
rect 800 9320 29200 9448
rect 880 9040 29120 9320
rect 800 8912 29200 9040
rect 880 8632 29120 8912
rect 800 8504 29200 8632
rect 880 8224 29120 8504
rect 800 8096 29200 8224
rect 880 7816 29120 8096
rect 800 7688 29200 7816
rect 880 7408 29120 7688
rect 800 7280 29200 7408
rect 880 7000 29120 7280
rect 800 6872 29200 7000
rect 880 6592 29120 6872
rect 800 6464 29200 6592
rect 880 6184 29120 6464
rect 800 6056 29200 6184
rect 880 5776 29120 6056
rect 800 5648 29200 5776
rect 880 5368 29120 5648
rect 800 5240 29200 5368
rect 880 4960 29120 5240
rect 800 4832 29200 4960
rect 880 4552 29120 4832
rect 800 4424 29200 4552
rect 880 4144 29120 4424
rect 800 4016 29200 4144
rect 880 3736 29120 4016
rect 800 3608 29200 3736
rect 880 3328 29120 3608
rect 800 3200 29200 3328
rect 880 2920 29120 3200
rect 800 2792 29200 2920
rect 880 2512 29120 2792
rect 800 2384 29200 2512
rect 880 2104 29120 2384
rect 800 1976 29200 2104
rect 880 1696 29120 1976
rect 800 1568 29200 1696
rect 880 1288 29120 1568
rect 800 1160 29200 1288
rect 880 880 29120 1160
rect 800 752 29200 880
rect 880 472 29120 752
rect 800 344 29200 472
rect 880 171 29120 344
<< metal4 >>
rect 5576 2128 5896 53360
rect 10208 2128 10528 53360
rect 14840 2128 15160 53360
rect 19472 2128 19792 53360
rect 24104 2128 24424 53360
<< labels >>
rlabel metal2 s 6090 -800 6146 800 8 io_adr_i[0]
port 1 nsew signal input
rlabel metal2 s 7470 -800 7526 800 8 io_adr_i[1]
port 2 nsew signal input
rlabel metal2 s 3330 -800 3386 800 8 io_cs_i
port 3 nsew signal input
rlabel metal2 s 8758 -800 8814 800 8 io_dat_i[0]
port 4 nsew signal input
rlabel metal2 s 22466 -800 22522 800 8 io_dat_i[10]
port 5 nsew signal input
rlabel metal2 s 23754 -800 23810 800 8 io_dat_i[11]
port 6 nsew signal input
rlabel metal2 s 25134 -800 25190 800 8 io_dat_i[12]
port 7 nsew signal input
rlabel metal2 s 26514 -800 26570 800 8 io_dat_i[13]
port 8 nsew signal input
rlabel metal2 s 27894 -800 27950 800 8 io_dat_i[14]
port 9 nsew signal input
rlabel metal2 s 29274 -800 29330 800 8 io_dat_i[15]
port 10 nsew signal input
rlabel metal2 s 10138 -800 10194 800 8 io_dat_i[1]
port 11 nsew signal input
rlabel metal2 s 11518 -800 11574 800 8 io_dat_i[2]
port 12 nsew signal input
rlabel metal2 s 12898 -800 12954 800 8 io_dat_i[3]
port 13 nsew signal input
rlabel metal2 s 14278 -800 14334 800 8 io_dat_i[4]
port 14 nsew signal input
rlabel metal2 s 15658 -800 15714 800 8 io_dat_i[5]
port 15 nsew signal input
rlabel metal2 s 16946 -800 17002 800 8 io_dat_i[6]
port 16 nsew signal input
rlabel metal2 s 18326 -800 18382 800 8 io_dat_i[7]
port 17 nsew signal input
rlabel metal2 s 19706 -800 19762 800 8 io_dat_i[8]
port 18 nsew signal input
rlabel metal2 s 21086 -800 21142 800 8 io_dat_i[9]
port 19 nsew signal input
rlabel metal2 s 846 55200 902 56800 6 io_dat_o[0]
port 20 nsew signal output
rlabel metal2 s 18418 55200 18474 56800 6 io_dat_o[10]
port 21 nsew signal output
rlabel metal2 s 20166 55200 20222 56800 6 io_dat_o[11]
port 22 nsew signal output
rlabel metal2 s 22006 55200 22062 56800 6 io_dat_o[12]
port 23 nsew signal output
rlabel metal2 s 23754 55200 23810 56800 6 io_dat_o[13]
port 24 nsew signal output
rlabel metal2 s 25502 55200 25558 56800 6 io_dat_o[14]
port 25 nsew signal output
rlabel metal2 s 27250 55200 27306 56800 6 io_dat_o[15]
port 26 nsew signal output
rlabel metal2 s 2594 55200 2650 56800 6 io_dat_o[1]
port 27 nsew signal output
rlabel metal2 s 4342 55200 4398 56800 6 io_dat_o[2]
port 28 nsew signal output
rlabel metal2 s 6090 55200 6146 56800 6 io_dat_o[3]
port 29 nsew signal output
rlabel metal2 s 7838 55200 7894 56800 6 io_dat_o[4]
port 30 nsew signal output
rlabel metal2 s 9586 55200 9642 56800 6 io_dat_o[5]
port 31 nsew signal output
rlabel metal2 s 11426 55200 11482 56800 6 io_dat_o[6]
port 32 nsew signal output
rlabel metal2 s 13174 55200 13230 56800 6 io_dat_o[7]
port 33 nsew signal output
rlabel metal2 s 14922 55200 14978 56800 6 io_dat_o[8]
port 34 nsew signal output
rlabel metal2 s 16670 55200 16726 56800 6 io_dat_o[9]
port 35 nsew signal output
rlabel metal3 s 29200 29520 30800 29640 6 io_eo[0]
port 36 nsew signal input
rlabel metal3 s 29200 33600 30800 33720 6 io_eo[10]
port 37 nsew signal input
rlabel metal3 s 29200 34008 30800 34128 6 io_eo[11]
port 38 nsew signal input
rlabel metal3 s 29200 34416 30800 34536 6 io_eo[12]
port 39 nsew signal input
rlabel metal3 s 29200 34824 30800 34944 6 io_eo[13]
port 40 nsew signal input
rlabel metal3 s 29200 35232 30800 35352 6 io_eo[14]
port 41 nsew signal input
rlabel metal3 s 29200 35640 30800 35760 6 io_eo[15]
port 42 nsew signal input
rlabel metal3 s 29200 36048 30800 36168 6 io_eo[16]
port 43 nsew signal input
rlabel metal3 s 29200 36456 30800 36576 6 io_eo[17]
port 44 nsew signal input
rlabel metal3 s 29200 36864 30800 36984 6 io_eo[18]
port 45 nsew signal input
rlabel metal3 s 29200 37272 30800 37392 6 io_eo[19]
port 46 nsew signal input
rlabel metal3 s 29200 29928 30800 30048 6 io_eo[1]
port 47 nsew signal input
rlabel metal3 s 29200 37680 30800 37800 6 io_eo[20]
port 48 nsew signal input
rlabel metal3 s 29200 38088 30800 38208 6 io_eo[21]
port 49 nsew signal input
rlabel metal3 s 29200 38496 30800 38616 6 io_eo[22]
port 50 nsew signal input
rlabel metal3 s 29200 38904 30800 39024 6 io_eo[23]
port 51 nsew signal input
rlabel metal3 s 29200 39312 30800 39432 6 io_eo[24]
port 52 nsew signal input
rlabel metal3 s 29200 39720 30800 39840 6 io_eo[25]
port 53 nsew signal input
rlabel metal3 s 29200 40128 30800 40248 6 io_eo[26]
port 54 nsew signal input
rlabel metal3 s 29200 40536 30800 40656 6 io_eo[27]
port 55 nsew signal input
rlabel metal3 s 29200 40944 30800 41064 6 io_eo[28]
port 56 nsew signal input
rlabel metal3 s 29200 41352 30800 41472 6 io_eo[29]
port 57 nsew signal input
rlabel metal3 s 29200 30336 30800 30456 6 io_eo[2]
port 58 nsew signal input
rlabel metal3 s 29200 41760 30800 41880 6 io_eo[30]
port 59 nsew signal input
rlabel metal3 s 29200 42168 30800 42288 6 io_eo[31]
port 60 nsew signal input
rlabel metal3 s 29200 42576 30800 42696 6 io_eo[32]
port 61 nsew signal input
rlabel metal3 s 29200 42984 30800 43104 6 io_eo[33]
port 62 nsew signal input
rlabel metal3 s 29200 43392 30800 43512 6 io_eo[34]
port 63 nsew signal input
rlabel metal3 s 29200 43800 30800 43920 6 io_eo[35]
port 64 nsew signal input
rlabel metal3 s 29200 44208 30800 44328 6 io_eo[36]
port 65 nsew signal input
rlabel metal3 s 29200 44616 30800 44736 6 io_eo[37]
port 66 nsew signal input
rlabel metal3 s 29200 45024 30800 45144 6 io_eo[38]
port 67 nsew signal input
rlabel metal3 s 29200 45432 30800 45552 6 io_eo[39]
port 68 nsew signal input
rlabel metal3 s 29200 30744 30800 30864 6 io_eo[3]
port 69 nsew signal input
rlabel metal3 s 29200 45840 30800 45960 6 io_eo[40]
port 70 nsew signal input
rlabel metal3 s 29200 46248 30800 46368 6 io_eo[41]
port 71 nsew signal input
rlabel metal3 s 29200 46656 30800 46776 6 io_eo[42]
port 72 nsew signal input
rlabel metal3 s 29200 47064 30800 47184 6 io_eo[43]
port 73 nsew signal input
rlabel metal3 s 29200 47472 30800 47592 6 io_eo[44]
port 74 nsew signal input
rlabel metal3 s 29200 47880 30800 48000 6 io_eo[45]
port 75 nsew signal input
rlabel metal3 s 29200 48288 30800 48408 6 io_eo[46]
port 76 nsew signal input
rlabel metal3 s 29200 48696 30800 48816 6 io_eo[47]
port 77 nsew signal input
rlabel metal3 s 29200 49104 30800 49224 6 io_eo[48]
port 78 nsew signal input
rlabel metal3 s 29200 49512 30800 49632 6 io_eo[49]
port 79 nsew signal input
rlabel metal3 s 29200 31152 30800 31272 6 io_eo[4]
port 80 nsew signal input
rlabel metal3 s 29200 49920 30800 50040 6 io_eo[50]
port 81 nsew signal input
rlabel metal3 s 29200 50328 30800 50448 6 io_eo[51]
port 82 nsew signal input
rlabel metal3 s 29200 50736 30800 50856 6 io_eo[52]
port 83 nsew signal input
rlabel metal3 s 29200 51144 30800 51264 6 io_eo[53]
port 84 nsew signal input
rlabel metal3 s 29200 51552 30800 51672 6 io_eo[54]
port 85 nsew signal input
rlabel metal3 s 29200 51960 30800 52080 6 io_eo[55]
port 86 nsew signal input
rlabel metal3 s 29200 52368 30800 52488 6 io_eo[56]
port 87 nsew signal input
rlabel metal3 s 29200 52776 30800 52896 6 io_eo[57]
port 88 nsew signal input
rlabel metal3 s 29200 53184 30800 53304 6 io_eo[58]
port 89 nsew signal input
rlabel metal3 s 29200 53592 30800 53712 6 io_eo[59]
port 90 nsew signal input
rlabel metal3 s 29200 31560 30800 31680 6 io_eo[5]
port 91 nsew signal input
rlabel metal3 s 29200 54000 30800 54120 6 io_eo[60]
port 92 nsew signal input
rlabel metal3 s 29200 54408 30800 54528 6 io_eo[61]
port 93 nsew signal input
rlabel metal3 s 29200 54816 30800 54936 6 io_eo[62]
port 94 nsew signal input
rlabel metal3 s 29200 55224 30800 55344 6 io_eo[63]
port 95 nsew signal input
rlabel metal3 s 29200 31968 30800 32088 6 io_eo[6]
port 96 nsew signal input
rlabel metal3 s 29200 32376 30800 32496 6 io_eo[7]
port 97 nsew signal input
rlabel metal3 s 29200 32784 30800 32904 6 io_eo[8]
port 98 nsew signal input
rlabel metal3 s 29200 33192 30800 33312 6 io_eo[9]
port 99 nsew signal input
rlabel metal3 s -800 144 800 264 4 io_i_0_ci
port 100 nsew signal input
rlabel metal3 s -800 3408 800 3528 4 io_i_0_in1[0]
port 101 nsew signal input
rlabel metal3 s -800 6672 800 6792 4 io_i_0_in1[1]
port 102 nsew signal input
rlabel metal3 s -800 9936 800 10056 4 io_i_0_in1[2]
port 103 nsew signal input
rlabel metal3 s -800 13200 800 13320 4 io_i_0_in1[3]
port 104 nsew signal input
rlabel metal3 s -800 16464 800 16584 4 io_i_0_in1[4]
port 105 nsew signal input
rlabel metal3 s -800 19728 800 19848 4 io_i_0_in1[5]
port 106 nsew signal input
rlabel metal3 s -800 22992 800 23112 4 io_i_0_in1[6]
port 107 nsew signal input
rlabel metal3 s -800 26256 800 26376 4 io_i_0_in1[7]
port 108 nsew signal input
rlabel metal3 s -800 552 800 672 4 io_i_1_ci
port 109 nsew signal input
rlabel metal3 s -800 3816 800 3936 4 io_i_1_in1[0]
port 110 nsew signal input
rlabel metal3 s -800 7080 800 7200 4 io_i_1_in1[1]
port 111 nsew signal input
rlabel metal3 s -800 10344 800 10464 4 io_i_1_in1[2]
port 112 nsew signal input
rlabel metal3 s -800 13608 800 13728 4 io_i_1_in1[3]
port 113 nsew signal input
rlabel metal3 s -800 16872 800 16992 4 io_i_1_in1[4]
port 114 nsew signal input
rlabel metal3 s -800 20136 800 20256 4 io_i_1_in1[5]
port 115 nsew signal input
rlabel metal3 s -800 23400 800 23520 4 io_i_1_in1[6]
port 116 nsew signal input
rlabel metal3 s -800 26664 800 26784 4 io_i_1_in1[7]
port 117 nsew signal input
rlabel metal3 s -800 960 800 1080 4 io_i_2_ci
port 118 nsew signal input
rlabel metal3 s -800 4224 800 4344 4 io_i_2_in1[0]
port 119 nsew signal input
rlabel metal3 s -800 7488 800 7608 4 io_i_2_in1[1]
port 120 nsew signal input
rlabel metal3 s -800 10752 800 10872 4 io_i_2_in1[2]
port 121 nsew signal input
rlabel metal3 s -800 14016 800 14136 4 io_i_2_in1[3]
port 122 nsew signal input
rlabel metal3 s -800 17280 800 17400 4 io_i_2_in1[4]
port 123 nsew signal input
rlabel metal3 s -800 20544 800 20664 4 io_i_2_in1[5]
port 124 nsew signal input
rlabel metal3 s -800 23808 800 23928 4 io_i_2_in1[6]
port 125 nsew signal input
rlabel metal3 s -800 27072 800 27192 4 io_i_2_in1[7]
port 126 nsew signal input
rlabel metal3 s -800 1368 800 1488 4 io_i_3_ci
port 127 nsew signal input
rlabel metal3 s -800 4632 800 4752 4 io_i_3_in1[0]
port 128 nsew signal input
rlabel metal3 s -800 7896 800 8016 4 io_i_3_in1[1]
port 129 nsew signal input
rlabel metal3 s -800 11160 800 11280 4 io_i_3_in1[2]
port 130 nsew signal input
rlabel metal3 s -800 14424 800 14544 4 io_i_3_in1[3]
port 131 nsew signal input
rlabel metal3 s -800 17688 800 17808 4 io_i_3_in1[4]
port 132 nsew signal input
rlabel metal3 s -800 20952 800 21072 4 io_i_3_in1[5]
port 133 nsew signal input
rlabel metal3 s -800 24216 800 24336 4 io_i_3_in1[6]
port 134 nsew signal input
rlabel metal3 s -800 27480 800 27600 4 io_i_3_in1[7]
port 135 nsew signal input
rlabel metal3 s -800 1776 800 1896 4 io_i_4_ci
port 136 nsew signal input
rlabel metal3 s -800 5040 800 5160 4 io_i_4_in1[0]
port 137 nsew signal input
rlabel metal3 s -800 8304 800 8424 4 io_i_4_in1[1]
port 138 nsew signal input
rlabel metal3 s -800 11568 800 11688 4 io_i_4_in1[2]
port 139 nsew signal input
rlabel metal3 s -800 14832 800 14952 4 io_i_4_in1[3]
port 140 nsew signal input
rlabel metal3 s -800 18096 800 18216 4 io_i_4_in1[4]
port 141 nsew signal input
rlabel metal3 s -800 21360 800 21480 4 io_i_4_in1[5]
port 142 nsew signal input
rlabel metal3 s -800 24624 800 24744 4 io_i_4_in1[6]
port 143 nsew signal input
rlabel metal3 s -800 27888 800 28008 4 io_i_4_in1[7]
port 144 nsew signal input
rlabel metal3 s -800 2184 800 2304 4 io_i_5_ci
port 145 nsew signal input
rlabel metal3 s -800 5448 800 5568 4 io_i_5_in1[0]
port 146 nsew signal input
rlabel metal3 s -800 8712 800 8832 4 io_i_5_in1[1]
port 147 nsew signal input
rlabel metal3 s -800 11976 800 12096 4 io_i_5_in1[2]
port 148 nsew signal input
rlabel metal3 s -800 15240 800 15360 4 io_i_5_in1[3]
port 149 nsew signal input
rlabel metal3 s -800 18504 800 18624 4 io_i_5_in1[4]
port 150 nsew signal input
rlabel metal3 s -800 21768 800 21888 4 io_i_5_in1[5]
port 151 nsew signal input
rlabel metal3 s -800 25032 800 25152 4 io_i_5_in1[6]
port 152 nsew signal input
rlabel metal3 s -800 28296 800 28416 4 io_i_5_in1[7]
port 153 nsew signal input
rlabel metal3 s -800 2592 800 2712 4 io_i_6_ci
port 154 nsew signal input
rlabel metal3 s -800 5856 800 5976 4 io_i_6_in1[0]
port 155 nsew signal input
rlabel metal3 s -800 9120 800 9240 4 io_i_6_in1[1]
port 156 nsew signal input
rlabel metal3 s -800 12384 800 12504 4 io_i_6_in1[2]
port 157 nsew signal input
rlabel metal3 s -800 15648 800 15768 4 io_i_6_in1[3]
port 158 nsew signal input
rlabel metal3 s -800 18912 800 19032 4 io_i_6_in1[4]
port 159 nsew signal input
rlabel metal3 s -800 22176 800 22296 4 io_i_6_in1[5]
port 160 nsew signal input
rlabel metal3 s -800 25440 800 25560 4 io_i_6_in1[6]
port 161 nsew signal input
rlabel metal3 s -800 28704 800 28824 4 io_i_6_in1[7]
port 162 nsew signal input
rlabel metal3 s -800 3000 800 3120 4 io_i_7_ci
port 163 nsew signal input
rlabel metal3 s -800 6264 800 6384 4 io_i_7_in1[0]
port 164 nsew signal input
rlabel metal3 s -800 9528 800 9648 4 io_i_7_in1[1]
port 165 nsew signal input
rlabel metal3 s -800 12792 800 12912 4 io_i_7_in1[2]
port 166 nsew signal input
rlabel metal3 s -800 16056 800 16176 4 io_i_7_in1[3]
port 167 nsew signal input
rlabel metal3 s -800 19320 800 19440 4 io_i_7_in1[4]
port 168 nsew signal input
rlabel metal3 s -800 22584 800 22704 4 io_i_7_in1[5]
port 169 nsew signal input
rlabel metal3 s -800 25848 800 25968 4 io_i_7_in1[6]
port 170 nsew signal input
rlabel metal3 s -800 29112 800 29232 4 io_i_7_in1[7]
port 171 nsew signal input
rlabel metal3 s 29200 144 30800 264 6 io_o_0_co
port 172 nsew signal output
rlabel metal3 s 29200 3408 30800 3528 6 io_o_0_out[0]
port 173 nsew signal output
rlabel metal3 s 29200 6672 30800 6792 6 io_o_0_out[1]
port 174 nsew signal output
rlabel metal3 s 29200 9936 30800 10056 6 io_o_0_out[2]
port 175 nsew signal output
rlabel metal3 s 29200 13200 30800 13320 6 io_o_0_out[3]
port 176 nsew signal output
rlabel metal3 s 29200 16464 30800 16584 6 io_o_0_out[4]
port 177 nsew signal output
rlabel metal3 s 29200 19728 30800 19848 6 io_o_0_out[5]
port 178 nsew signal output
rlabel metal3 s 29200 22992 30800 23112 6 io_o_0_out[6]
port 179 nsew signal output
rlabel metal3 s 29200 26256 30800 26376 6 io_o_0_out[7]
port 180 nsew signal output
rlabel metal3 s 29200 552 30800 672 6 io_o_1_co
port 181 nsew signal output
rlabel metal3 s 29200 3816 30800 3936 6 io_o_1_out[0]
port 182 nsew signal output
rlabel metal3 s 29200 7080 30800 7200 6 io_o_1_out[1]
port 183 nsew signal output
rlabel metal3 s 29200 10344 30800 10464 6 io_o_1_out[2]
port 184 nsew signal output
rlabel metal3 s 29200 13608 30800 13728 6 io_o_1_out[3]
port 185 nsew signal output
rlabel metal3 s 29200 16872 30800 16992 6 io_o_1_out[4]
port 186 nsew signal output
rlabel metal3 s 29200 20136 30800 20256 6 io_o_1_out[5]
port 187 nsew signal output
rlabel metal3 s 29200 23400 30800 23520 6 io_o_1_out[6]
port 188 nsew signal output
rlabel metal3 s 29200 26664 30800 26784 6 io_o_1_out[7]
port 189 nsew signal output
rlabel metal3 s 29200 960 30800 1080 6 io_o_2_co
port 190 nsew signal output
rlabel metal3 s 29200 4224 30800 4344 6 io_o_2_out[0]
port 191 nsew signal output
rlabel metal3 s 29200 7488 30800 7608 6 io_o_2_out[1]
port 192 nsew signal output
rlabel metal3 s 29200 10752 30800 10872 6 io_o_2_out[2]
port 193 nsew signal output
rlabel metal3 s 29200 14016 30800 14136 6 io_o_2_out[3]
port 194 nsew signal output
rlabel metal3 s 29200 17280 30800 17400 6 io_o_2_out[4]
port 195 nsew signal output
rlabel metal3 s 29200 20544 30800 20664 6 io_o_2_out[5]
port 196 nsew signal output
rlabel metal3 s 29200 23808 30800 23928 6 io_o_2_out[6]
port 197 nsew signal output
rlabel metal3 s 29200 27072 30800 27192 6 io_o_2_out[7]
port 198 nsew signal output
rlabel metal3 s 29200 1368 30800 1488 6 io_o_3_co
port 199 nsew signal output
rlabel metal3 s 29200 4632 30800 4752 6 io_o_3_out[0]
port 200 nsew signal output
rlabel metal3 s 29200 7896 30800 8016 6 io_o_3_out[1]
port 201 nsew signal output
rlabel metal3 s 29200 11160 30800 11280 6 io_o_3_out[2]
port 202 nsew signal output
rlabel metal3 s 29200 14424 30800 14544 6 io_o_3_out[3]
port 203 nsew signal output
rlabel metal3 s 29200 17688 30800 17808 6 io_o_3_out[4]
port 204 nsew signal output
rlabel metal3 s 29200 20952 30800 21072 6 io_o_3_out[5]
port 205 nsew signal output
rlabel metal3 s 29200 24216 30800 24336 6 io_o_3_out[6]
port 206 nsew signal output
rlabel metal3 s 29200 27480 30800 27600 6 io_o_3_out[7]
port 207 nsew signal output
rlabel metal3 s 29200 1776 30800 1896 6 io_o_4_co
port 208 nsew signal output
rlabel metal3 s 29200 5040 30800 5160 6 io_o_4_out[0]
port 209 nsew signal output
rlabel metal3 s 29200 8304 30800 8424 6 io_o_4_out[1]
port 210 nsew signal output
rlabel metal3 s 29200 11568 30800 11688 6 io_o_4_out[2]
port 211 nsew signal output
rlabel metal3 s 29200 14832 30800 14952 6 io_o_4_out[3]
port 212 nsew signal output
rlabel metal3 s 29200 18096 30800 18216 6 io_o_4_out[4]
port 213 nsew signal output
rlabel metal3 s 29200 21360 30800 21480 6 io_o_4_out[5]
port 214 nsew signal output
rlabel metal3 s 29200 24624 30800 24744 6 io_o_4_out[6]
port 215 nsew signal output
rlabel metal3 s 29200 27888 30800 28008 6 io_o_4_out[7]
port 216 nsew signal output
rlabel metal3 s 29200 2184 30800 2304 6 io_o_5_co
port 217 nsew signal output
rlabel metal3 s 29200 5448 30800 5568 6 io_o_5_out[0]
port 218 nsew signal output
rlabel metal3 s 29200 8712 30800 8832 6 io_o_5_out[1]
port 219 nsew signal output
rlabel metal3 s 29200 11976 30800 12096 6 io_o_5_out[2]
port 220 nsew signal output
rlabel metal3 s 29200 15240 30800 15360 6 io_o_5_out[3]
port 221 nsew signal output
rlabel metal3 s 29200 18504 30800 18624 6 io_o_5_out[4]
port 222 nsew signal output
rlabel metal3 s 29200 21768 30800 21888 6 io_o_5_out[5]
port 223 nsew signal output
rlabel metal3 s 29200 25032 30800 25152 6 io_o_5_out[6]
port 224 nsew signal output
rlabel metal3 s 29200 28296 30800 28416 6 io_o_5_out[7]
port 225 nsew signal output
rlabel metal3 s 29200 2592 30800 2712 6 io_o_6_co
port 226 nsew signal output
rlabel metal3 s 29200 5856 30800 5976 6 io_o_6_out[0]
port 227 nsew signal output
rlabel metal3 s 29200 9120 30800 9240 6 io_o_6_out[1]
port 228 nsew signal output
rlabel metal3 s 29200 12384 30800 12504 6 io_o_6_out[2]
port 229 nsew signal output
rlabel metal3 s 29200 15648 30800 15768 6 io_o_6_out[3]
port 230 nsew signal output
rlabel metal3 s 29200 18912 30800 19032 6 io_o_6_out[4]
port 231 nsew signal output
rlabel metal3 s 29200 22176 30800 22296 6 io_o_6_out[5]
port 232 nsew signal output
rlabel metal3 s 29200 25440 30800 25560 6 io_o_6_out[6]
port 233 nsew signal output
rlabel metal3 s 29200 28704 30800 28824 6 io_o_6_out[7]
port 234 nsew signal output
rlabel metal3 s 29200 3000 30800 3120 6 io_o_7_co
port 235 nsew signal output
rlabel metal3 s 29200 6264 30800 6384 6 io_o_7_out[0]
port 236 nsew signal output
rlabel metal3 s 29200 9528 30800 9648 6 io_o_7_out[1]
port 237 nsew signal output
rlabel metal3 s 29200 12792 30800 12912 6 io_o_7_out[2]
port 238 nsew signal output
rlabel metal3 s 29200 16056 30800 16176 6 io_o_7_out[3]
port 239 nsew signal output
rlabel metal3 s 29200 19320 30800 19440 6 io_o_7_out[4]
port 240 nsew signal output
rlabel metal3 s 29200 22584 30800 22704 6 io_o_7_out[5]
port 241 nsew signal output
rlabel metal3 s 29200 25848 30800 25968 6 io_o_7_out[6]
port 242 nsew signal output
rlabel metal3 s 29200 29112 30800 29232 6 io_o_7_out[7]
port 243 nsew signal output
rlabel metal2 s 662 -800 718 800 8 io_vci
port 244 nsew signal input
rlabel metal2 s 1950 -800 2006 800 8 io_vco
port 245 nsew signal output
rlabel metal2 s 28998 55200 29054 56800 6 io_vi
port 246 nsew signal input
rlabel metal2 s 4710 -800 4766 800 8 io_we_i
port 247 nsew signal input
rlabel metal3 s -800 29520 800 29640 4 io_wo[0]
port 248 nsew signal output
rlabel metal3 s -800 33600 800 33720 4 io_wo[10]
port 249 nsew signal output
rlabel metal3 s -800 34008 800 34128 4 io_wo[11]
port 250 nsew signal output
rlabel metal3 s -800 34416 800 34536 4 io_wo[12]
port 251 nsew signal output
rlabel metal3 s -800 34824 800 34944 4 io_wo[13]
port 252 nsew signal output
rlabel metal3 s -800 35232 800 35352 4 io_wo[14]
port 253 nsew signal output
rlabel metal3 s -800 35640 800 35760 4 io_wo[15]
port 254 nsew signal output
rlabel metal3 s -800 36048 800 36168 4 io_wo[16]
port 255 nsew signal output
rlabel metal3 s -800 36456 800 36576 4 io_wo[17]
port 256 nsew signal output
rlabel metal3 s -800 36864 800 36984 4 io_wo[18]
port 257 nsew signal output
rlabel metal3 s -800 37272 800 37392 4 io_wo[19]
port 258 nsew signal output
rlabel metal3 s -800 29928 800 30048 4 io_wo[1]
port 259 nsew signal output
rlabel metal3 s -800 37680 800 37800 4 io_wo[20]
port 260 nsew signal output
rlabel metal3 s -800 38088 800 38208 4 io_wo[21]
port 261 nsew signal output
rlabel metal3 s -800 38496 800 38616 4 io_wo[22]
port 262 nsew signal output
rlabel metal3 s -800 38904 800 39024 4 io_wo[23]
port 263 nsew signal output
rlabel metal3 s -800 39312 800 39432 4 io_wo[24]
port 264 nsew signal output
rlabel metal3 s -800 39720 800 39840 4 io_wo[25]
port 265 nsew signal output
rlabel metal3 s -800 40128 800 40248 4 io_wo[26]
port 266 nsew signal output
rlabel metal3 s -800 40536 800 40656 4 io_wo[27]
port 267 nsew signal output
rlabel metal3 s -800 40944 800 41064 4 io_wo[28]
port 268 nsew signal output
rlabel metal3 s -800 41352 800 41472 4 io_wo[29]
port 269 nsew signal output
rlabel metal3 s -800 30336 800 30456 4 io_wo[2]
port 270 nsew signal output
rlabel metal3 s -800 41760 800 41880 4 io_wo[30]
port 271 nsew signal output
rlabel metal3 s -800 42168 800 42288 4 io_wo[31]
port 272 nsew signal output
rlabel metal3 s -800 42576 800 42696 4 io_wo[32]
port 273 nsew signal output
rlabel metal3 s -800 42984 800 43104 4 io_wo[33]
port 274 nsew signal output
rlabel metal3 s -800 43392 800 43512 4 io_wo[34]
port 275 nsew signal output
rlabel metal3 s -800 43800 800 43920 4 io_wo[35]
port 276 nsew signal output
rlabel metal3 s -800 44208 800 44328 4 io_wo[36]
port 277 nsew signal output
rlabel metal3 s -800 44616 800 44736 4 io_wo[37]
port 278 nsew signal output
rlabel metal3 s -800 45024 800 45144 4 io_wo[38]
port 279 nsew signal output
rlabel metal3 s -800 45432 800 45552 4 io_wo[39]
port 280 nsew signal output
rlabel metal3 s -800 30744 800 30864 4 io_wo[3]
port 281 nsew signal output
rlabel metal3 s -800 45840 800 45960 4 io_wo[40]
port 282 nsew signal output
rlabel metal3 s -800 46248 800 46368 4 io_wo[41]
port 283 nsew signal output
rlabel metal3 s -800 46656 800 46776 4 io_wo[42]
port 284 nsew signal output
rlabel metal3 s -800 47064 800 47184 4 io_wo[43]
port 285 nsew signal output
rlabel metal3 s -800 47472 800 47592 4 io_wo[44]
port 286 nsew signal output
rlabel metal3 s -800 47880 800 48000 4 io_wo[45]
port 287 nsew signal output
rlabel metal3 s -800 48288 800 48408 4 io_wo[46]
port 288 nsew signal output
rlabel metal3 s -800 48696 800 48816 4 io_wo[47]
port 289 nsew signal output
rlabel metal3 s -800 49104 800 49224 4 io_wo[48]
port 290 nsew signal output
rlabel metal3 s -800 49512 800 49632 4 io_wo[49]
port 291 nsew signal output
rlabel metal3 s -800 31152 800 31272 4 io_wo[4]
port 292 nsew signal output
rlabel metal3 s -800 49920 800 50040 4 io_wo[50]
port 293 nsew signal output
rlabel metal3 s -800 50328 800 50448 4 io_wo[51]
port 294 nsew signal output
rlabel metal3 s -800 50736 800 50856 4 io_wo[52]
port 295 nsew signal output
rlabel metal3 s -800 51144 800 51264 4 io_wo[53]
port 296 nsew signal output
rlabel metal3 s -800 51552 800 51672 4 io_wo[54]
port 297 nsew signal output
rlabel metal3 s -800 51960 800 52080 4 io_wo[55]
port 298 nsew signal output
rlabel metal3 s -800 52368 800 52488 4 io_wo[56]
port 299 nsew signal output
rlabel metal3 s -800 52776 800 52896 4 io_wo[57]
port 300 nsew signal output
rlabel metal3 s -800 53184 800 53304 4 io_wo[58]
port 301 nsew signal output
rlabel metal3 s -800 53592 800 53712 4 io_wo[59]
port 302 nsew signal output
rlabel metal3 s -800 31560 800 31680 4 io_wo[5]
port 303 nsew signal output
rlabel metal3 s -800 54000 800 54120 4 io_wo[60]
port 304 nsew signal output
rlabel metal3 s -800 54408 800 54528 4 io_wo[61]
port 305 nsew signal output
rlabel metal3 s -800 54816 800 54936 4 io_wo[62]
port 306 nsew signal output
rlabel metal3 s -800 55224 800 55344 4 io_wo[63]
port 307 nsew signal output
rlabel metal3 s -800 31968 800 32088 4 io_wo[6]
port 308 nsew signal output
rlabel metal3 s -800 32376 800 32496 4 io_wo[7]
port 309 nsew signal output
rlabel metal3 s -800 32784 800 32904 4 io_wo[8]
port 310 nsew signal output
rlabel metal3 s -800 33192 800 33312 4 io_wo[9]
port 311 nsew signal output
rlabel metal3 s 29200 55632 30800 55752 6 wb_clk_i
port 312 nsew signal input
rlabel metal3 s -800 55632 800 55752 4 wb_rst_i
port 313 nsew signal input
rlabel metal4 s 24104 2128 24424 53360 6 vccd1
port 314 nsew power bidirectional
rlabel metal4 s 14840 2128 15160 53360 6 vccd1
port 315 nsew power bidirectional
rlabel metal4 s 5576 2128 5896 53360 6 vccd1
port 316 nsew power bidirectional
rlabel metal4 s 19472 2128 19792 53360 6 vssd1
port 317 nsew ground bidirectional
rlabel metal4 s 10208 2128 10528 53360 6 vssd1
port 318 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 30000 56000
string LEFview TRUE
string GDS_FILE /project/openlane/cic_block/runs/cic_block/results/magic/cic_block.gds
string GDS_END 4901764
string GDS_START 636668
<< end >>

