module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vccd1,
    vssd1,
    vccd2,
    vssd2,
    vdda1,
    vssa1,
    vdda2,
    vssa2,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vccd1;
 input vssd1;
 input vccd2;
 input vssd2;
 input vdda1;
 input vssa1;
 input vdda2;
 input vssa2;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 cic_block cb_0_0 (.io_cs_i(cb_0_0_io_cs_i),
    .io_i_0_ci(cb_0_0_io_i_0_ci),
    .io_o_0_co(cb_0_0_io_o_0_co),
    .io_o_1_co(cb_0_0_io_o_1_co),
    .io_o_2_co(cb_0_0_io_o_2_co),
    .io_o_3_co(cb_0_0_io_o_3_co),
    .io_o_4_co(cb_0_0_io_o_4_co),
    .io_o_5_co(cb_0_0_io_o_5_co),
    .io_o_6_co(cb_0_0_io_o_6_co),
    .io_o_7_co(cb_0_0_io_o_7_co),
    .io_vco(cb_0_0_io_vco),
    .io_vi(cb_0_0_io_vi),
    .io_we_i(cb_0_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_0_0_io_adr_i[1] ,
    \cb_0_0_io_adr_i[0] }),
    .io_dat_i({\cb_0_0_io_dat_i[15] ,
    \cb_0_0_io_dat_i[14] ,
    \cb_0_0_io_dat_i[13] ,
    \cb_0_0_io_dat_i[12] ,
    \cb_0_0_io_dat_i[11] ,
    \cb_0_0_io_dat_i[10] ,
    \cb_0_0_io_dat_i[9] ,
    \cb_0_0_io_dat_i[8] ,
    \cb_0_0_io_dat_i[7] ,
    \cb_0_0_io_dat_i[6] ,
    \cb_0_0_io_dat_i[5] ,
    \cb_0_0_io_dat_i[4] ,
    \cb_0_0_io_dat_i[3] ,
    \cb_0_0_io_dat_i[2] ,
    \cb_0_0_io_dat_i[1] ,
    \cb_0_0_io_dat_i[0] }),
    .io_dat_o({\cb_0_0_io_dat_o[15] ,
    \cb_0_0_io_dat_o[14] ,
    \cb_0_0_io_dat_o[13] ,
    \cb_0_0_io_dat_o[12] ,
    \cb_0_0_io_dat_o[11] ,
    \cb_0_0_io_dat_o[10] ,
    \cb_0_0_io_dat_o[9] ,
    \cb_0_0_io_dat_o[8] ,
    \cb_0_0_io_dat_o[7] ,
    \cb_0_0_io_dat_o[6] ,
    \cb_0_0_io_dat_o[5] ,
    \cb_0_0_io_dat_o[4] ,
    \cb_0_0_io_dat_o[3] ,
    \cb_0_0_io_dat_o[2] ,
    \cb_0_0_io_dat_o[1] ,
    \cb_0_0_io_dat_o[0] }),
    .io_eo({\cb_0_0_io_eo[63] ,
    \cb_0_0_io_eo[62] ,
    \cb_0_0_io_eo[61] ,
    \cb_0_0_io_eo[60] ,
    \cb_0_0_io_eo[59] ,
    \cb_0_0_io_eo[58] ,
    \cb_0_0_io_eo[57] ,
    \cb_0_0_io_eo[56] ,
    \cb_0_0_io_eo[55] ,
    \cb_0_0_io_eo[54] ,
    \cb_0_0_io_eo[53] ,
    \cb_0_0_io_eo[52] ,
    \cb_0_0_io_eo[51] ,
    \cb_0_0_io_eo[50] ,
    \cb_0_0_io_eo[49] ,
    \cb_0_0_io_eo[48] ,
    \cb_0_0_io_eo[47] ,
    \cb_0_0_io_eo[46] ,
    \cb_0_0_io_eo[45] ,
    \cb_0_0_io_eo[44] ,
    \cb_0_0_io_eo[43] ,
    \cb_0_0_io_eo[42] ,
    \cb_0_0_io_eo[41] ,
    \cb_0_0_io_eo[40] ,
    \cb_0_0_io_eo[39] ,
    \cb_0_0_io_eo[38] ,
    \cb_0_0_io_eo[37] ,
    \cb_0_0_io_eo[36] ,
    \cb_0_0_io_eo[35] ,
    \cb_0_0_io_eo[34] ,
    \cb_0_0_io_eo[33] ,
    \cb_0_0_io_eo[32] ,
    \cb_0_0_io_eo[31] ,
    \cb_0_0_io_eo[30] ,
    \cb_0_0_io_eo[29] ,
    \cb_0_0_io_eo[28] ,
    \cb_0_0_io_eo[27] ,
    \cb_0_0_io_eo[26] ,
    \cb_0_0_io_eo[25] ,
    \cb_0_0_io_eo[24] ,
    \cb_0_0_io_eo[23] ,
    \cb_0_0_io_eo[22] ,
    \cb_0_0_io_eo[21] ,
    \cb_0_0_io_eo[20] ,
    \cb_0_0_io_eo[19] ,
    \cb_0_0_io_eo[18] ,
    \cb_0_0_io_eo[17] ,
    \cb_0_0_io_eo[16] ,
    \cb_0_0_io_eo[15] ,
    \cb_0_0_io_eo[14] ,
    \cb_0_0_io_eo[13] ,
    \cb_0_0_io_eo[12] ,
    \cb_0_0_io_eo[11] ,
    \cb_0_0_io_eo[10] ,
    \cb_0_0_io_eo[9] ,
    \cb_0_0_io_eo[8] ,
    \cb_0_0_io_eo[7] ,
    \cb_0_0_io_eo[6] ,
    \cb_0_0_io_eo[5] ,
    \cb_0_0_io_eo[4] ,
    \cb_0_0_io_eo[3] ,
    \cb_0_0_io_eo[2] ,
    \cb_0_0_io_eo[1] ,
    \cb_0_0_io_eo[0] }),
    .io_i_0_in1({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8}),
    .io_i_1_in1({_NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16}),
    .io_i_2_in1({_NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24}),
    .io_i_3_in1({_NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32}),
    .io_i_4_in1({_NC33,
    _NC34,
    _NC35,
    _NC36,
    _NC37,
    _NC38,
    _NC39,
    _NC40}),
    .io_i_5_in1({_NC41,
    _NC42,
    _NC43,
    _NC44,
    _NC45,
    _NC46,
    _NC47,
    _NC48}),
    .io_i_6_in1({_NC49,
    _NC50,
    _NC51,
    _NC52,
    _NC53,
    _NC54,
    _NC55,
    _NC56}),
    .io_i_7_in1({_NC57,
    _NC58,
    _NC59,
    _NC60,
    _NC61,
    _NC62,
    _NC63,
    _NC64}),
    .io_o_0_out({\cb_0_0_io_o_0_out[7] ,
    \cb_0_0_io_o_0_out[6] ,
    \cb_0_0_io_o_0_out[5] ,
    \cb_0_0_io_o_0_out[4] ,
    \cb_0_0_io_o_0_out[3] ,
    \cb_0_0_io_o_0_out[2] ,
    \cb_0_0_io_o_0_out[1] ,
    \cb_0_0_io_o_0_out[0] }),
    .io_o_1_out({\cb_0_0_io_o_1_out[7] ,
    \cb_0_0_io_o_1_out[6] ,
    \cb_0_0_io_o_1_out[5] ,
    \cb_0_0_io_o_1_out[4] ,
    \cb_0_0_io_o_1_out[3] ,
    \cb_0_0_io_o_1_out[2] ,
    \cb_0_0_io_o_1_out[1] ,
    \cb_0_0_io_o_1_out[0] }),
    .io_o_2_out({\cb_0_0_io_o_2_out[7] ,
    \cb_0_0_io_o_2_out[6] ,
    \cb_0_0_io_o_2_out[5] ,
    \cb_0_0_io_o_2_out[4] ,
    \cb_0_0_io_o_2_out[3] ,
    \cb_0_0_io_o_2_out[2] ,
    \cb_0_0_io_o_2_out[1] ,
    \cb_0_0_io_o_2_out[0] }),
    .io_o_3_out({\cb_0_0_io_o_3_out[7] ,
    \cb_0_0_io_o_3_out[6] ,
    \cb_0_0_io_o_3_out[5] ,
    \cb_0_0_io_o_3_out[4] ,
    \cb_0_0_io_o_3_out[3] ,
    \cb_0_0_io_o_3_out[2] ,
    \cb_0_0_io_o_3_out[1] ,
    \cb_0_0_io_o_3_out[0] }),
    .io_o_4_out({\cb_0_0_io_o_4_out[7] ,
    \cb_0_0_io_o_4_out[6] ,
    \cb_0_0_io_o_4_out[5] ,
    \cb_0_0_io_o_4_out[4] ,
    \cb_0_0_io_o_4_out[3] ,
    \cb_0_0_io_o_4_out[2] ,
    \cb_0_0_io_o_4_out[1] ,
    \cb_0_0_io_o_4_out[0] }),
    .io_o_5_out({\cb_0_0_io_o_5_out[7] ,
    \cb_0_0_io_o_5_out[6] ,
    \cb_0_0_io_o_5_out[5] ,
    \cb_0_0_io_o_5_out[4] ,
    \cb_0_0_io_o_5_out[3] ,
    \cb_0_0_io_o_5_out[2] ,
    \cb_0_0_io_o_5_out[1] ,
    \cb_0_0_io_o_5_out[0] }),
    .io_o_6_out({\cb_0_0_io_o_6_out[7] ,
    \cb_0_0_io_o_6_out[6] ,
    \cb_0_0_io_o_6_out[5] ,
    \cb_0_0_io_o_6_out[4] ,
    \cb_0_0_io_o_6_out[3] ,
    \cb_0_0_io_o_6_out[2] ,
    \cb_0_0_io_o_6_out[1] ,
    \cb_0_0_io_o_6_out[0] }),
    .io_o_7_out({\cb_0_0_io_o_7_out[7] ,
    \cb_0_0_io_o_7_out[6] ,
    \cb_0_0_io_o_7_out[5] ,
    \cb_0_0_io_o_7_out[4] ,
    \cb_0_0_io_o_7_out[3] ,
    \cb_0_0_io_o_7_out[2] ,
    \cb_0_0_io_o_7_out[1] ,
    \cb_0_0_io_o_7_out[0] }),
    .io_wo({\cb_0_0_io_wo[63] ,
    \cb_0_0_io_wo[62] ,
    \cb_0_0_io_wo[61] ,
    \cb_0_0_io_wo[60] ,
    \cb_0_0_io_wo[59] ,
    \cb_0_0_io_wo[58] ,
    \cb_0_0_io_wo[57] ,
    \cb_0_0_io_wo[56] ,
    \cb_0_0_io_wo[55] ,
    \cb_0_0_io_wo[54] ,
    \cb_0_0_io_wo[53] ,
    \cb_0_0_io_wo[52] ,
    \cb_0_0_io_wo[51] ,
    \cb_0_0_io_wo[50] ,
    \cb_0_0_io_wo[49] ,
    \cb_0_0_io_wo[48] ,
    \cb_0_0_io_wo[47] ,
    \cb_0_0_io_wo[46] ,
    \cb_0_0_io_wo[45] ,
    \cb_0_0_io_wo[44] ,
    \cb_0_0_io_wo[43] ,
    \cb_0_0_io_wo[42] ,
    \cb_0_0_io_wo[41] ,
    \cb_0_0_io_wo[40] ,
    \cb_0_0_io_wo[39] ,
    \cb_0_0_io_wo[38] ,
    \cb_0_0_io_wo[37] ,
    \cb_0_0_io_wo[36] ,
    \cb_0_0_io_wo[35] ,
    \cb_0_0_io_wo[34] ,
    \cb_0_0_io_wo[33] ,
    \cb_0_0_io_wo[32] ,
    \cb_0_0_io_wo[31] ,
    \cb_0_0_io_wo[30] ,
    \cb_0_0_io_wo[29] ,
    \cb_0_0_io_wo[28] ,
    \cb_0_0_io_wo[27] ,
    \cb_0_0_io_wo[26] ,
    \cb_0_0_io_wo[25] ,
    \cb_0_0_io_wo[24] ,
    \cb_0_0_io_wo[23] ,
    \cb_0_0_io_wo[22] ,
    \cb_0_0_io_wo[21] ,
    \cb_0_0_io_wo[20] ,
    \cb_0_0_io_wo[19] ,
    \cb_0_0_io_wo[18] ,
    \cb_0_0_io_wo[17] ,
    \cb_0_0_io_wo[16] ,
    \cb_0_0_io_wo[15] ,
    \cb_0_0_io_wo[14] ,
    \cb_0_0_io_wo[13] ,
    \cb_0_0_io_wo[12] ,
    \cb_0_0_io_wo[11] ,
    \cb_0_0_io_wo[10] ,
    \cb_0_0_io_wo[9] ,
    \cb_0_0_io_wo[8] ,
    \cb_0_0_io_wo[7] ,
    \cb_0_0_io_wo[6] ,
    \cb_0_0_io_wo[5] ,
    \cb_0_0_io_wo[4] ,
    \cb_0_0_io_wo[3] ,
    \cb_0_0_io_wo[2] ,
    \cb_0_0_io_wo[1] ,
    \cb_0_0_io_wo[0] }));
 cic_block cb_0_1 (.io_cs_i(cb_0_1_io_cs_i),
    .io_i_0_ci(cb_0_0_io_o_0_co),
    .io_i_1_ci(cb_0_0_io_o_1_co),
    .io_i_2_ci(cb_0_0_io_o_2_co),
    .io_i_3_ci(cb_0_0_io_o_3_co),
    .io_i_4_ci(cb_0_0_io_o_4_co),
    .io_i_5_ci(cb_0_0_io_o_5_co),
    .io_i_6_ci(cb_0_0_io_o_6_co),
    .io_i_7_ci(cb_0_0_io_o_7_co),
    .io_o_0_co(cb_0_1_io_o_0_co),
    .io_o_1_co(cb_0_1_io_o_1_co),
    .io_o_2_co(cb_0_1_io_o_2_co),
    .io_o_3_co(cb_0_1_io_o_3_co),
    .io_o_4_co(cb_0_1_io_o_4_co),
    .io_o_5_co(cb_0_1_io_o_5_co),
    .io_o_6_co(cb_0_1_io_o_6_co),
    .io_o_7_co(cb_0_1_io_o_7_co),
    .io_vci(cb_0_0_io_vco),
    .io_vco(cb_0_1_io_vco),
    .io_vi(cb_0_1_io_vi),
    .io_we_i(cb_0_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_0_0_io_adr_i[1] ,
    \cb_0_0_io_adr_i[0] }),
    .io_dat_i({\cb_0_0_io_dat_i[15] ,
    \cb_0_0_io_dat_i[14] ,
    \cb_0_0_io_dat_i[13] ,
    \cb_0_0_io_dat_i[12] ,
    \cb_0_0_io_dat_i[11] ,
    \cb_0_0_io_dat_i[10] ,
    \cb_0_0_io_dat_i[9] ,
    \cb_0_0_io_dat_i[8] ,
    \cb_0_0_io_dat_i[7] ,
    \cb_0_0_io_dat_i[6] ,
    \cb_0_0_io_dat_i[5] ,
    \cb_0_0_io_dat_i[4] ,
    \cb_0_0_io_dat_i[3] ,
    \cb_0_0_io_dat_i[2] ,
    \cb_0_0_io_dat_i[1] ,
    \cb_0_0_io_dat_i[0] }),
    .io_dat_o({\cb_0_1_io_dat_o[15] ,
    \cb_0_1_io_dat_o[14] ,
    \cb_0_1_io_dat_o[13] ,
    \cb_0_1_io_dat_o[12] ,
    \cb_0_1_io_dat_o[11] ,
    \cb_0_1_io_dat_o[10] ,
    \cb_0_1_io_dat_o[9] ,
    \cb_0_1_io_dat_o[8] ,
    \cb_0_1_io_dat_o[7] ,
    \cb_0_1_io_dat_o[6] ,
    \cb_0_1_io_dat_o[5] ,
    \cb_0_1_io_dat_o[4] ,
    \cb_0_1_io_dat_o[3] ,
    \cb_0_1_io_dat_o[2] ,
    \cb_0_1_io_dat_o[1] ,
    \cb_0_1_io_dat_o[0] }),
    .io_eo({\cb_0_1_io_eo[63] ,
    \cb_0_1_io_eo[62] ,
    \cb_0_1_io_eo[61] ,
    \cb_0_1_io_eo[60] ,
    \cb_0_1_io_eo[59] ,
    \cb_0_1_io_eo[58] ,
    \cb_0_1_io_eo[57] ,
    \cb_0_1_io_eo[56] ,
    \cb_0_1_io_eo[55] ,
    \cb_0_1_io_eo[54] ,
    \cb_0_1_io_eo[53] ,
    \cb_0_1_io_eo[52] ,
    \cb_0_1_io_eo[51] ,
    \cb_0_1_io_eo[50] ,
    \cb_0_1_io_eo[49] ,
    \cb_0_1_io_eo[48] ,
    \cb_0_1_io_eo[47] ,
    \cb_0_1_io_eo[46] ,
    \cb_0_1_io_eo[45] ,
    \cb_0_1_io_eo[44] ,
    \cb_0_1_io_eo[43] ,
    \cb_0_1_io_eo[42] ,
    \cb_0_1_io_eo[41] ,
    \cb_0_1_io_eo[40] ,
    \cb_0_1_io_eo[39] ,
    \cb_0_1_io_eo[38] ,
    \cb_0_1_io_eo[37] ,
    \cb_0_1_io_eo[36] ,
    \cb_0_1_io_eo[35] ,
    \cb_0_1_io_eo[34] ,
    \cb_0_1_io_eo[33] ,
    \cb_0_1_io_eo[32] ,
    \cb_0_1_io_eo[31] ,
    \cb_0_1_io_eo[30] ,
    \cb_0_1_io_eo[29] ,
    \cb_0_1_io_eo[28] ,
    \cb_0_1_io_eo[27] ,
    \cb_0_1_io_eo[26] ,
    \cb_0_1_io_eo[25] ,
    \cb_0_1_io_eo[24] ,
    \cb_0_1_io_eo[23] ,
    \cb_0_1_io_eo[22] ,
    \cb_0_1_io_eo[21] ,
    \cb_0_1_io_eo[20] ,
    \cb_0_1_io_eo[19] ,
    \cb_0_1_io_eo[18] ,
    \cb_0_1_io_eo[17] ,
    \cb_0_1_io_eo[16] ,
    \cb_0_1_io_eo[15] ,
    \cb_0_1_io_eo[14] ,
    \cb_0_1_io_eo[13] ,
    \cb_0_1_io_eo[12] ,
    \cb_0_1_io_eo[11] ,
    \cb_0_1_io_eo[10] ,
    \cb_0_1_io_eo[9] ,
    \cb_0_1_io_eo[8] ,
    \cb_0_1_io_eo[7] ,
    \cb_0_1_io_eo[6] ,
    \cb_0_1_io_eo[5] ,
    \cb_0_1_io_eo[4] ,
    \cb_0_1_io_eo[3] ,
    \cb_0_1_io_eo[2] ,
    \cb_0_1_io_eo[1] ,
    \cb_0_1_io_eo[0] }),
    .io_i_0_in1({\cb_0_0_io_o_0_out[7] ,
    \cb_0_0_io_o_0_out[6] ,
    \cb_0_0_io_o_0_out[5] ,
    \cb_0_0_io_o_0_out[4] ,
    \cb_0_0_io_o_0_out[3] ,
    \cb_0_0_io_o_0_out[2] ,
    \cb_0_0_io_o_0_out[1] ,
    \cb_0_0_io_o_0_out[0] }),
    .io_i_1_in1({\cb_0_0_io_o_1_out[7] ,
    \cb_0_0_io_o_1_out[6] ,
    \cb_0_0_io_o_1_out[5] ,
    \cb_0_0_io_o_1_out[4] ,
    \cb_0_0_io_o_1_out[3] ,
    \cb_0_0_io_o_1_out[2] ,
    \cb_0_0_io_o_1_out[1] ,
    \cb_0_0_io_o_1_out[0] }),
    .io_i_2_in1({\cb_0_0_io_o_2_out[7] ,
    \cb_0_0_io_o_2_out[6] ,
    \cb_0_0_io_o_2_out[5] ,
    \cb_0_0_io_o_2_out[4] ,
    \cb_0_0_io_o_2_out[3] ,
    \cb_0_0_io_o_2_out[2] ,
    \cb_0_0_io_o_2_out[1] ,
    \cb_0_0_io_o_2_out[0] }),
    .io_i_3_in1({\cb_0_0_io_o_3_out[7] ,
    \cb_0_0_io_o_3_out[6] ,
    \cb_0_0_io_o_3_out[5] ,
    \cb_0_0_io_o_3_out[4] ,
    \cb_0_0_io_o_3_out[3] ,
    \cb_0_0_io_o_3_out[2] ,
    \cb_0_0_io_o_3_out[1] ,
    \cb_0_0_io_o_3_out[0] }),
    .io_i_4_in1({\cb_0_0_io_o_4_out[7] ,
    \cb_0_0_io_o_4_out[6] ,
    \cb_0_0_io_o_4_out[5] ,
    \cb_0_0_io_o_4_out[4] ,
    \cb_0_0_io_o_4_out[3] ,
    \cb_0_0_io_o_4_out[2] ,
    \cb_0_0_io_o_4_out[1] ,
    \cb_0_0_io_o_4_out[0] }),
    .io_i_5_in1({\cb_0_0_io_o_5_out[7] ,
    \cb_0_0_io_o_5_out[6] ,
    \cb_0_0_io_o_5_out[5] ,
    \cb_0_0_io_o_5_out[4] ,
    \cb_0_0_io_o_5_out[3] ,
    \cb_0_0_io_o_5_out[2] ,
    \cb_0_0_io_o_5_out[1] ,
    \cb_0_0_io_o_5_out[0] }),
    .io_i_6_in1({\cb_0_0_io_o_6_out[7] ,
    \cb_0_0_io_o_6_out[6] ,
    \cb_0_0_io_o_6_out[5] ,
    \cb_0_0_io_o_6_out[4] ,
    \cb_0_0_io_o_6_out[3] ,
    \cb_0_0_io_o_6_out[2] ,
    \cb_0_0_io_o_6_out[1] ,
    \cb_0_0_io_o_6_out[0] }),
    .io_i_7_in1({\cb_0_0_io_o_7_out[7] ,
    \cb_0_0_io_o_7_out[6] ,
    \cb_0_0_io_o_7_out[5] ,
    \cb_0_0_io_o_7_out[4] ,
    \cb_0_0_io_o_7_out[3] ,
    \cb_0_0_io_o_7_out[2] ,
    \cb_0_0_io_o_7_out[1] ,
    \cb_0_0_io_o_7_out[0] }),
    .io_o_0_out({\cb_0_1_io_o_0_out[7] ,
    \cb_0_1_io_o_0_out[6] ,
    \cb_0_1_io_o_0_out[5] ,
    \cb_0_1_io_o_0_out[4] ,
    \cb_0_1_io_o_0_out[3] ,
    \cb_0_1_io_o_0_out[2] ,
    \cb_0_1_io_o_0_out[1] ,
    \cb_0_1_io_o_0_out[0] }),
    .io_o_1_out({\cb_0_1_io_o_1_out[7] ,
    \cb_0_1_io_o_1_out[6] ,
    \cb_0_1_io_o_1_out[5] ,
    \cb_0_1_io_o_1_out[4] ,
    \cb_0_1_io_o_1_out[3] ,
    \cb_0_1_io_o_1_out[2] ,
    \cb_0_1_io_o_1_out[1] ,
    \cb_0_1_io_o_1_out[0] }),
    .io_o_2_out({\cb_0_1_io_o_2_out[7] ,
    \cb_0_1_io_o_2_out[6] ,
    \cb_0_1_io_o_2_out[5] ,
    \cb_0_1_io_o_2_out[4] ,
    \cb_0_1_io_o_2_out[3] ,
    \cb_0_1_io_o_2_out[2] ,
    \cb_0_1_io_o_2_out[1] ,
    \cb_0_1_io_o_2_out[0] }),
    .io_o_3_out({\cb_0_1_io_o_3_out[7] ,
    \cb_0_1_io_o_3_out[6] ,
    \cb_0_1_io_o_3_out[5] ,
    \cb_0_1_io_o_3_out[4] ,
    \cb_0_1_io_o_3_out[3] ,
    \cb_0_1_io_o_3_out[2] ,
    \cb_0_1_io_o_3_out[1] ,
    \cb_0_1_io_o_3_out[0] }),
    .io_o_4_out({\cb_0_1_io_o_4_out[7] ,
    \cb_0_1_io_o_4_out[6] ,
    \cb_0_1_io_o_4_out[5] ,
    \cb_0_1_io_o_4_out[4] ,
    \cb_0_1_io_o_4_out[3] ,
    \cb_0_1_io_o_4_out[2] ,
    \cb_0_1_io_o_4_out[1] ,
    \cb_0_1_io_o_4_out[0] }),
    .io_o_5_out({\cb_0_1_io_o_5_out[7] ,
    \cb_0_1_io_o_5_out[6] ,
    \cb_0_1_io_o_5_out[5] ,
    \cb_0_1_io_o_5_out[4] ,
    \cb_0_1_io_o_5_out[3] ,
    \cb_0_1_io_o_5_out[2] ,
    \cb_0_1_io_o_5_out[1] ,
    \cb_0_1_io_o_5_out[0] }),
    .io_o_6_out({\cb_0_1_io_o_6_out[7] ,
    \cb_0_1_io_o_6_out[6] ,
    \cb_0_1_io_o_6_out[5] ,
    \cb_0_1_io_o_6_out[4] ,
    \cb_0_1_io_o_6_out[3] ,
    \cb_0_1_io_o_6_out[2] ,
    \cb_0_1_io_o_6_out[1] ,
    \cb_0_1_io_o_6_out[0] }),
    .io_o_7_out({\cb_0_1_io_o_7_out[7] ,
    \cb_0_1_io_o_7_out[6] ,
    \cb_0_1_io_o_7_out[5] ,
    \cb_0_1_io_o_7_out[4] ,
    \cb_0_1_io_o_7_out[3] ,
    \cb_0_1_io_o_7_out[2] ,
    \cb_0_1_io_o_7_out[1] ,
    \cb_0_1_io_o_7_out[0] }),
    .io_wo({\cb_0_0_io_eo[63] ,
    \cb_0_0_io_eo[62] ,
    \cb_0_0_io_eo[61] ,
    \cb_0_0_io_eo[60] ,
    \cb_0_0_io_eo[59] ,
    \cb_0_0_io_eo[58] ,
    \cb_0_0_io_eo[57] ,
    \cb_0_0_io_eo[56] ,
    \cb_0_0_io_eo[55] ,
    \cb_0_0_io_eo[54] ,
    \cb_0_0_io_eo[53] ,
    \cb_0_0_io_eo[52] ,
    \cb_0_0_io_eo[51] ,
    \cb_0_0_io_eo[50] ,
    \cb_0_0_io_eo[49] ,
    \cb_0_0_io_eo[48] ,
    \cb_0_0_io_eo[47] ,
    \cb_0_0_io_eo[46] ,
    \cb_0_0_io_eo[45] ,
    \cb_0_0_io_eo[44] ,
    \cb_0_0_io_eo[43] ,
    \cb_0_0_io_eo[42] ,
    \cb_0_0_io_eo[41] ,
    \cb_0_0_io_eo[40] ,
    \cb_0_0_io_eo[39] ,
    \cb_0_0_io_eo[38] ,
    \cb_0_0_io_eo[37] ,
    \cb_0_0_io_eo[36] ,
    \cb_0_0_io_eo[35] ,
    \cb_0_0_io_eo[34] ,
    \cb_0_0_io_eo[33] ,
    \cb_0_0_io_eo[32] ,
    \cb_0_0_io_eo[31] ,
    \cb_0_0_io_eo[30] ,
    \cb_0_0_io_eo[29] ,
    \cb_0_0_io_eo[28] ,
    \cb_0_0_io_eo[27] ,
    \cb_0_0_io_eo[26] ,
    \cb_0_0_io_eo[25] ,
    \cb_0_0_io_eo[24] ,
    \cb_0_0_io_eo[23] ,
    \cb_0_0_io_eo[22] ,
    \cb_0_0_io_eo[21] ,
    \cb_0_0_io_eo[20] ,
    \cb_0_0_io_eo[19] ,
    \cb_0_0_io_eo[18] ,
    \cb_0_0_io_eo[17] ,
    \cb_0_0_io_eo[16] ,
    \cb_0_0_io_eo[15] ,
    \cb_0_0_io_eo[14] ,
    \cb_0_0_io_eo[13] ,
    \cb_0_0_io_eo[12] ,
    \cb_0_0_io_eo[11] ,
    \cb_0_0_io_eo[10] ,
    \cb_0_0_io_eo[9] ,
    \cb_0_0_io_eo[8] ,
    \cb_0_0_io_eo[7] ,
    \cb_0_0_io_eo[6] ,
    \cb_0_0_io_eo[5] ,
    \cb_0_0_io_eo[4] ,
    \cb_0_0_io_eo[3] ,
    \cb_0_0_io_eo[2] ,
    \cb_0_0_io_eo[1] ,
    \cb_0_0_io_eo[0] }));
 cic_block cb_0_10 (.io_cs_i(cb_0_10_io_cs_i),
    .io_i_0_ci(cb_0_10_io_i_0_ci),
    .io_i_1_ci(cb_0_10_io_i_1_ci),
    .io_i_2_ci(cb_0_10_io_i_2_ci),
    .io_i_3_ci(cb_0_10_io_i_3_ci),
    .io_i_4_ci(cb_0_10_io_i_4_ci),
    .io_i_5_ci(cb_0_10_io_i_5_ci),
    .io_i_6_ci(cb_0_10_io_i_6_ci),
    .io_i_7_ci(cb_0_10_io_i_7_ci),
    .io_o_0_co(cb_0_10_io_o_0_co),
    .io_o_1_co(cb_0_10_io_o_1_co),
    .io_o_2_co(cb_0_10_io_o_2_co),
    .io_o_3_co(cb_0_10_io_o_3_co),
    .io_o_4_co(cb_0_10_io_o_4_co),
    .io_o_5_co(cb_0_10_io_o_5_co),
    .io_o_6_co(cb_0_10_io_o_6_co),
    .io_o_7_co(cb_0_10_io_o_7_co),
    .io_vci(cb_0_10_io_vci),
    .io_vco(cb_0_10_io_vco),
    .io_vi(cb_0_10_io_vi),
    .io_we_i(cb_0_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_0_0_io_adr_i[1] ,
    \cb_0_0_io_adr_i[0] }),
    .io_dat_i({\cb_0_0_io_dat_i[15] ,
    \cb_0_0_io_dat_i[14] ,
    \cb_0_0_io_dat_i[13] ,
    \cb_0_0_io_dat_i[12] ,
    \cb_0_0_io_dat_i[11] ,
    \cb_0_0_io_dat_i[10] ,
    \cb_0_0_io_dat_i[9] ,
    \cb_0_0_io_dat_i[8] ,
    \cb_0_0_io_dat_i[7] ,
    \cb_0_0_io_dat_i[6] ,
    \cb_0_0_io_dat_i[5] ,
    \cb_0_0_io_dat_i[4] ,
    \cb_0_0_io_dat_i[3] ,
    \cb_0_0_io_dat_i[2] ,
    \cb_0_0_io_dat_i[1] ,
    \cb_0_0_io_dat_i[0] }),
    .io_dat_o({\cb_0_10_io_dat_o[15] ,
    \cb_0_10_io_dat_o[14] ,
    \cb_0_10_io_dat_o[13] ,
    \cb_0_10_io_dat_o[12] ,
    \cb_0_10_io_dat_o[11] ,
    \cb_0_10_io_dat_o[10] ,
    \cb_0_10_io_dat_o[9] ,
    \cb_0_10_io_dat_o[8] ,
    \cb_0_10_io_dat_o[7] ,
    \cb_0_10_io_dat_o[6] ,
    \cb_0_10_io_dat_o[5] ,
    \cb_0_10_io_dat_o[4] ,
    \cb_0_10_io_dat_o[3] ,
    \cb_0_10_io_dat_o[2] ,
    \cb_0_10_io_dat_o[1] ,
    \cb_0_10_io_dat_o[0] }),
    .io_eo({\_T_28[31] ,
    \_T_28[30] ,
    \_T_28[29] ,
    \_T_28[28] ,
    \_T_28[27] ,
    \_T_28[26] ,
    \_T_28[25] ,
    \_T_28[24] ,
    \_T_28[23] ,
    \_T_28[22] ,
    \_T_28[21] ,
    \_T_28[20] ,
    \_T_28[19] ,
    \_T_28[18] ,
    \_T_28[17] ,
    \_T_28[16] ,
    \_T_28[15] ,
    \_T_28[14] ,
    \_T_28[13] ,
    \_T_28[12] ,
    \_T_28[11] ,
    \_T_28[10] ,
    \_T_28[9] ,
    \_T_28[8] ,
    \_T_28[7] ,
    \_T_28[6] ,
    \_T_28[5] ,
    \_T_28[4] ,
    \_T_28[3] ,
    \_T_28[2] ,
    \_T_28[1] ,
    \_T_28[0] ,
    \_T_25[31] ,
    \_T_25[30] ,
    \_T_25[29] ,
    \_T_25[28] ,
    \_T_25[27] ,
    \_T_25[26] ,
    \_T_25[25] ,
    \_T_25[24] ,
    \_T_25[23] ,
    \_T_25[22] ,
    \_T_25[21] ,
    \_T_25[20] ,
    \_T_25[19] ,
    \_T_25[18] ,
    \_T_25[17] ,
    \_T_25[16] ,
    \_T_25[15] ,
    \_T_25[14] ,
    \_T_25[13] ,
    \_T_25[12] ,
    \_T_25[11] ,
    \_T_25[10] ,
    \_T_25[9] ,
    \_T_25[8] ,
    \_T_25[7] ,
    \_T_25[6] ,
    \_T_25[5] ,
    \_T_25[4] ,
    \_T_25[3] ,
    \_T_25[2] ,
    \_T_25[1] ,
    \_T_25[0] }),
    .io_i_0_in1({\cb_0_10_io_i_0_in1[7] ,
    \cb_0_10_io_i_0_in1[6] ,
    \cb_0_10_io_i_0_in1[5] ,
    \cb_0_10_io_i_0_in1[4] ,
    \cb_0_10_io_i_0_in1[3] ,
    \cb_0_10_io_i_0_in1[2] ,
    \cb_0_10_io_i_0_in1[1] ,
    \cb_0_10_io_i_0_in1[0] }),
    .io_i_1_in1({\cb_0_10_io_i_1_in1[7] ,
    \cb_0_10_io_i_1_in1[6] ,
    \cb_0_10_io_i_1_in1[5] ,
    \cb_0_10_io_i_1_in1[4] ,
    \cb_0_10_io_i_1_in1[3] ,
    \cb_0_10_io_i_1_in1[2] ,
    \cb_0_10_io_i_1_in1[1] ,
    \cb_0_10_io_i_1_in1[0] }),
    .io_i_2_in1({\cb_0_10_io_i_2_in1[7] ,
    \cb_0_10_io_i_2_in1[6] ,
    \cb_0_10_io_i_2_in1[5] ,
    \cb_0_10_io_i_2_in1[4] ,
    \cb_0_10_io_i_2_in1[3] ,
    \cb_0_10_io_i_2_in1[2] ,
    \cb_0_10_io_i_2_in1[1] ,
    \cb_0_10_io_i_2_in1[0] }),
    .io_i_3_in1({\cb_0_10_io_i_3_in1[7] ,
    \cb_0_10_io_i_3_in1[6] ,
    \cb_0_10_io_i_3_in1[5] ,
    \cb_0_10_io_i_3_in1[4] ,
    \cb_0_10_io_i_3_in1[3] ,
    \cb_0_10_io_i_3_in1[2] ,
    \cb_0_10_io_i_3_in1[1] ,
    \cb_0_10_io_i_3_in1[0] }),
    .io_i_4_in1({\cb_0_10_io_i_4_in1[7] ,
    \cb_0_10_io_i_4_in1[6] ,
    \cb_0_10_io_i_4_in1[5] ,
    \cb_0_10_io_i_4_in1[4] ,
    \cb_0_10_io_i_4_in1[3] ,
    \cb_0_10_io_i_4_in1[2] ,
    \cb_0_10_io_i_4_in1[1] ,
    \cb_0_10_io_i_4_in1[0] }),
    .io_i_5_in1({\cb_0_10_io_i_5_in1[7] ,
    \cb_0_10_io_i_5_in1[6] ,
    \cb_0_10_io_i_5_in1[5] ,
    \cb_0_10_io_i_5_in1[4] ,
    \cb_0_10_io_i_5_in1[3] ,
    \cb_0_10_io_i_5_in1[2] ,
    \cb_0_10_io_i_5_in1[1] ,
    \cb_0_10_io_i_5_in1[0] }),
    .io_i_6_in1({\cb_0_10_io_i_6_in1[7] ,
    \cb_0_10_io_i_6_in1[6] ,
    \cb_0_10_io_i_6_in1[5] ,
    \cb_0_10_io_i_6_in1[4] ,
    \cb_0_10_io_i_6_in1[3] ,
    \cb_0_10_io_i_6_in1[2] ,
    \cb_0_10_io_i_6_in1[1] ,
    \cb_0_10_io_i_6_in1[0] }),
    .io_i_7_in1({\cb_0_10_io_i_7_in1[7] ,
    \cb_0_10_io_i_7_in1[6] ,
    \cb_0_10_io_i_7_in1[5] ,
    \cb_0_10_io_i_7_in1[4] ,
    \cb_0_10_io_i_7_in1[3] ,
    \cb_0_10_io_i_7_in1[2] ,
    \cb_0_10_io_i_7_in1[1] ,
    \cb_0_10_io_i_7_in1[0] }),
    .io_o_0_out({\_T_25[7] ,
    \_T_25[6] ,
    \_T_25[5] ,
    \_T_25[4] ,
    \_T_25[3] ,
    \_T_25[2] ,
    \_T_25[1] ,
    \_T_25[0] }),
    .io_o_1_out({\_T_25[15] ,
    \_T_25[14] ,
    \_T_25[13] ,
    \_T_25[12] ,
    \_T_25[11] ,
    \_T_25[10] ,
    \_T_25[9] ,
    \_T_25[8] }),
    .io_o_2_out({\_T_25[23] ,
    \_T_25[22] ,
    \_T_25[21] ,
    \_T_25[20] ,
    \_T_25[19] ,
    \_T_25[18] ,
    \_T_25[17] ,
    \_T_25[16] }),
    .io_o_3_out({\_T_25[31] ,
    \_T_25[30] ,
    \_T_25[29] ,
    \_T_25[28] ,
    \_T_25[27] ,
    \_T_25[26] ,
    \_T_25[25] ,
    \_T_25[24] }),
    .io_o_4_out({\_T_28[7] ,
    \_T_28[6] ,
    \_T_28[5] ,
    \_T_28[4] ,
    \_T_28[3] ,
    \_T_28[2] ,
    \_T_28[1] ,
    \_T_28[0] }),
    .io_o_5_out({\_T_28[15] ,
    \_T_28[14] ,
    \_T_28[13] ,
    \_T_28[12] ,
    \_T_28[11] ,
    \_T_28[10] ,
    \_T_28[9] ,
    \_T_28[8] }),
    .io_o_6_out({\_T_28[23] ,
    \_T_28[22] ,
    \_T_28[21] ,
    \_T_28[20] ,
    \_T_28[19] ,
    \_T_28[18] ,
    \_T_28[17] ,
    \_T_28[16] }),
    .io_o_7_out({\_T_28[31] ,
    \_T_28[30] ,
    \_T_28[29] ,
    \_T_28[28] ,
    \_T_28[27] ,
    \_T_28[26] ,
    \_T_28[25] ,
    \_T_28[24] }),
    .io_wo({\cb_0_10_io_wo[63] ,
    \cb_0_10_io_wo[62] ,
    \cb_0_10_io_wo[61] ,
    \cb_0_10_io_wo[60] ,
    \cb_0_10_io_wo[59] ,
    \cb_0_10_io_wo[58] ,
    \cb_0_10_io_wo[57] ,
    \cb_0_10_io_wo[56] ,
    \cb_0_10_io_wo[55] ,
    \cb_0_10_io_wo[54] ,
    \cb_0_10_io_wo[53] ,
    \cb_0_10_io_wo[52] ,
    \cb_0_10_io_wo[51] ,
    \cb_0_10_io_wo[50] ,
    \cb_0_10_io_wo[49] ,
    \cb_0_10_io_wo[48] ,
    \cb_0_10_io_wo[47] ,
    \cb_0_10_io_wo[46] ,
    \cb_0_10_io_wo[45] ,
    \cb_0_10_io_wo[44] ,
    \cb_0_10_io_wo[43] ,
    \cb_0_10_io_wo[42] ,
    \cb_0_10_io_wo[41] ,
    \cb_0_10_io_wo[40] ,
    \cb_0_10_io_wo[39] ,
    \cb_0_10_io_wo[38] ,
    \cb_0_10_io_wo[37] ,
    \cb_0_10_io_wo[36] ,
    \cb_0_10_io_wo[35] ,
    \cb_0_10_io_wo[34] ,
    \cb_0_10_io_wo[33] ,
    \cb_0_10_io_wo[32] ,
    \cb_0_10_io_wo[31] ,
    \cb_0_10_io_wo[30] ,
    \cb_0_10_io_wo[29] ,
    \cb_0_10_io_wo[28] ,
    \cb_0_10_io_wo[27] ,
    \cb_0_10_io_wo[26] ,
    \cb_0_10_io_wo[25] ,
    \cb_0_10_io_wo[24] ,
    \cb_0_10_io_wo[23] ,
    \cb_0_10_io_wo[22] ,
    \cb_0_10_io_wo[21] ,
    \cb_0_10_io_wo[20] ,
    \cb_0_10_io_wo[19] ,
    \cb_0_10_io_wo[18] ,
    \cb_0_10_io_wo[17] ,
    \cb_0_10_io_wo[16] ,
    \cb_0_10_io_wo[15] ,
    \cb_0_10_io_wo[14] ,
    \cb_0_10_io_wo[13] ,
    \cb_0_10_io_wo[12] ,
    \cb_0_10_io_wo[11] ,
    \cb_0_10_io_wo[10] ,
    \cb_0_10_io_wo[9] ,
    \cb_0_10_io_wo[8] ,
    \cb_0_10_io_wo[7] ,
    \cb_0_10_io_wo[6] ,
    \cb_0_10_io_wo[5] ,
    \cb_0_10_io_wo[4] ,
    \cb_0_10_io_wo[3] ,
    \cb_0_10_io_wo[2] ,
    \cb_0_10_io_wo[1] ,
    \cb_0_10_io_wo[0] }));
 cic_block cb_0_2 (.io_cs_i(cb_0_2_io_cs_i),
    .io_i_0_ci(cb_0_1_io_o_0_co),
    .io_i_1_ci(cb_0_1_io_o_1_co),
    .io_i_2_ci(cb_0_1_io_o_2_co),
    .io_i_3_ci(cb_0_1_io_o_3_co),
    .io_i_4_ci(cb_0_1_io_o_4_co),
    .io_i_5_ci(cb_0_1_io_o_5_co),
    .io_i_6_ci(cb_0_1_io_o_6_co),
    .io_i_7_ci(cb_0_1_io_o_7_co),
    .io_o_0_co(cb_0_2_io_o_0_co),
    .io_o_1_co(cb_0_2_io_o_1_co),
    .io_o_2_co(cb_0_2_io_o_2_co),
    .io_o_3_co(cb_0_2_io_o_3_co),
    .io_o_4_co(cb_0_2_io_o_4_co),
    .io_o_5_co(cb_0_2_io_o_5_co),
    .io_o_6_co(cb_0_2_io_o_6_co),
    .io_o_7_co(cb_0_2_io_o_7_co),
    .io_vci(cb_0_1_io_vco),
    .io_vco(cb_0_2_io_vco),
    .io_vi(cb_0_2_io_vi),
    .io_we_i(cb_0_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_0_0_io_adr_i[1] ,
    \cb_0_0_io_adr_i[0] }),
    .io_dat_i({\cb_0_0_io_dat_i[15] ,
    \cb_0_0_io_dat_i[14] ,
    \cb_0_0_io_dat_i[13] ,
    \cb_0_0_io_dat_i[12] ,
    \cb_0_0_io_dat_i[11] ,
    \cb_0_0_io_dat_i[10] ,
    \cb_0_0_io_dat_i[9] ,
    \cb_0_0_io_dat_i[8] ,
    \cb_0_0_io_dat_i[7] ,
    \cb_0_0_io_dat_i[6] ,
    \cb_0_0_io_dat_i[5] ,
    \cb_0_0_io_dat_i[4] ,
    \cb_0_0_io_dat_i[3] ,
    \cb_0_0_io_dat_i[2] ,
    \cb_0_0_io_dat_i[1] ,
    \cb_0_0_io_dat_i[0] }),
    .io_dat_o({\cb_0_2_io_dat_o[15] ,
    \cb_0_2_io_dat_o[14] ,
    \cb_0_2_io_dat_o[13] ,
    \cb_0_2_io_dat_o[12] ,
    \cb_0_2_io_dat_o[11] ,
    \cb_0_2_io_dat_o[10] ,
    \cb_0_2_io_dat_o[9] ,
    \cb_0_2_io_dat_o[8] ,
    \cb_0_2_io_dat_o[7] ,
    \cb_0_2_io_dat_o[6] ,
    \cb_0_2_io_dat_o[5] ,
    \cb_0_2_io_dat_o[4] ,
    \cb_0_2_io_dat_o[3] ,
    \cb_0_2_io_dat_o[2] ,
    \cb_0_2_io_dat_o[1] ,
    \cb_0_2_io_dat_o[0] }),
    .io_eo({\cb_0_2_io_eo[63] ,
    \cb_0_2_io_eo[62] ,
    \cb_0_2_io_eo[61] ,
    \cb_0_2_io_eo[60] ,
    \cb_0_2_io_eo[59] ,
    \cb_0_2_io_eo[58] ,
    \cb_0_2_io_eo[57] ,
    \cb_0_2_io_eo[56] ,
    \cb_0_2_io_eo[55] ,
    \cb_0_2_io_eo[54] ,
    \cb_0_2_io_eo[53] ,
    \cb_0_2_io_eo[52] ,
    \cb_0_2_io_eo[51] ,
    \cb_0_2_io_eo[50] ,
    \cb_0_2_io_eo[49] ,
    \cb_0_2_io_eo[48] ,
    \cb_0_2_io_eo[47] ,
    \cb_0_2_io_eo[46] ,
    \cb_0_2_io_eo[45] ,
    \cb_0_2_io_eo[44] ,
    \cb_0_2_io_eo[43] ,
    \cb_0_2_io_eo[42] ,
    \cb_0_2_io_eo[41] ,
    \cb_0_2_io_eo[40] ,
    \cb_0_2_io_eo[39] ,
    \cb_0_2_io_eo[38] ,
    \cb_0_2_io_eo[37] ,
    \cb_0_2_io_eo[36] ,
    \cb_0_2_io_eo[35] ,
    \cb_0_2_io_eo[34] ,
    \cb_0_2_io_eo[33] ,
    \cb_0_2_io_eo[32] ,
    \cb_0_2_io_eo[31] ,
    \cb_0_2_io_eo[30] ,
    \cb_0_2_io_eo[29] ,
    \cb_0_2_io_eo[28] ,
    \cb_0_2_io_eo[27] ,
    \cb_0_2_io_eo[26] ,
    \cb_0_2_io_eo[25] ,
    \cb_0_2_io_eo[24] ,
    \cb_0_2_io_eo[23] ,
    \cb_0_2_io_eo[22] ,
    \cb_0_2_io_eo[21] ,
    \cb_0_2_io_eo[20] ,
    \cb_0_2_io_eo[19] ,
    \cb_0_2_io_eo[18] ,
    \cb_0_2_io_eo[17] ,
    \cb_0_2_io_eo[16] ,
    \cb_0_2_io_eo[15] ,
    \cb_0_2_io_eo[14] ,
    \cb_0_2_io_eo[13] ,
    \cb_0_2_io_eo[12] ,
    \cb_0_2_io_eo[11] ,
    \cb_0_2_io_eo[10] ,
    \cb_0_2_io_eo[9] ,
    \cb_0_2_io_eo[8] ,
    \cb_0_2_io_eo[7] ,
    \cb_0_2_io_eo[6] ,
    \cb_0_2_io_eo[5] ,
    \cb_0_2_io_eo[4] ,
    \cb_0_2_io_eo[3] ,
    \cb_0_2_io_eo[2] ,
    \cb_0_2_io_eo[1] ,
    \cb_0_2_io_eo[0] }),
    .io_i_0_in1({\cb_0_1_io_o_0_out[7] ,
    \cb_0_1_io_o_0_out[6] ,
    \cb_0_1_io_o_0_out[5] ,
    \cb_0_1_io_o_0_out[4] ,
    \cb_0_1_io_o_0_out[3] ,
    \cb_0_1_io_o_0_out[2] ,
    \cb_0_1_io_o_0_out[1] ,
    \cb_0_1_io_o_0_out[0] }),
    .io_i_1_in1({\cb_0_1_io_o_1_out[7] ,
    \cb_0_1_io_o_1_out[6] ,
    \cb_0_1_io_o_1_out[5] ,
    \cb_0_1_io_o_1_out[4] ,
    \cb_0_1_io_o_1_out[3] ,
    \cb_0_1_io_o_1_out[2] ,
    \cb_0_1_io_o_1_out[1] ,
    \cb_0_1_io_o_1_out[0] }),
    .io_i_2_in1({\cb_0_1_io_o_2_out[7] ,
    \cb_0_1_io_o_2_out[6] ,
    \cb_0_1_io_o_2_out[5] ,
    \cb_0_1_io_o_2_out[4] ,
    \cb_0_1_io_o_2_out[3] ,
    \cb_0_1_io_o_2_out[2] ,
    \cb_0_1_io_o_2_out[1] ,
    \cb_0_1_io_o_2_out[0] }),
    .io_i_3_in1({\cb_0_1_io_o_3_out[7] ,
    \cb_0_1_io_o_3_out[6] ,
    \cb_0_1_io_o_3_out[5] ,
    \cb_0_1_io_o_3_out[4] ,
    \cb_0_1_io_o_3_out[3] ,
    \cb_0_1_io_o_3_out[2] ,
    \cb_0_1_io_o_3_out[1] ,
    \cb_0_1_io_o_3_out[0] }),
    .io_i_4_in1({\cb_0_1_io_o_4_out[7] ,
    \cb_0_1_io_o_4_out[6] ,
    \cb_0_1_io_o_4_out[5] ,
    \cb_0_1_io_o_4_out[4] ,
    \cb_0_1_io_o_4_out[3] ,
    \cb_0_1_io_o_4_out[2] ,
    \cb_0_1_io_o_4_out[1] ,
    \cb_0_1_io_o_4_out[0] }),
    .io_i_5_in1({\cb_0_1_io_o_5_out[7] ,
    \cb_0_1_io_o_5_out[6] ,
    \cb_0_1_io_o_5_out[5] ,
    \cb_0_1_io_o_5_out[4] ,
    \cb_0_1_io_o_5_out[3] ,
    \cb_0_1_io_o_5_out[2] ,
    \cb_0_1_io_o_5_out[1] ,
    \cb_0_1_io_o_5_out[0] }),
    .io_i_6_in1({\cb_0_1_io_o_6_out[7] ,
    \cb_0_1_io_o_6_out[6] ,
    \cb_0_1_io_o_6_out[5] ,
    \cb_0_1_io_o_6_out[4] ,
    \cb_0_1_io_o_6_out[3] ,
    \cb_0_1_io_o_6_out[2] ,
    \cb_0_1_io_o_6_out[1] ,
    \cb_0_1_io_o_6_out[0] }),
    .io_i_7_in1({\cb_0_1_io_o_7_out[7] ,
    \cb_0_1_io_o_7_out[6] ,
    \cb_0_1_io_o_7_out[5] ,
    \cb_0_1_io_o_7_out[4] ,
    \cb_0_1_io_o_7_out[3] ,
    \cb_0_1_io_o_7_out[2] ,
    \cb_0_1_io_o_7_out[1] ,
    \cb_0_1_io_o_7_out[0] }),
    .io_o_0_out({\cb_0_2_io_o_0_out[7] ,
    \cb_0_2_io_o_0_out[6] ,
    \cb_0_2_io_o_0_out[5] ,
    \cb_0_2_io_o_0_out[4] ,
    \cb_0_2_io_o_0_out[3] ,
    \cb_0_2_io_o_0_out[2] ,
    \cb_0_2_io_o_0_out[1] ,
    \cb_0_2_io_o_0_out[0] }),
    .io_o_1_out({\cb_0_2_io_o_1_out[7] ,
    \cb_0_2_io_o_1_out[6] ,
    \cb_0_2_io_o_1_out[5] ,
    \cb_0_2_io_o_1_out[4] ,
    \cb_0_2_io_o_1_out[3] ,
    \cb_0_2_io_o_1_out[2] ,
    \cb_0_2_io_o_1_out[1] ,
    \cb_0_2_io_o_1_out[0] }),
    .io_o_2_out({\cb_0_2_io_o_2_out[7] ,
    \cb_0_2_io_o_2_out[6] ,
    \cb_0_2_io_o_2_out[5] ,
    \cb_0_2_io_o_2_out[4] ,
    \cb_0_2_io_o_2_out[3] ,
    \cb_0_2_io_o_2_out[2] ,
    \cb_0_2_io_o_2_out[1] ,
    \cb_0_2_io_o_2_out[0] }),
    .io_o_3_out({\cb_0_2_io_o_3_out[7] ,
    \cb_0_2_io_o_3_out[6] ,
    \cb_0_2_io_o_3_out[5] ,
    \cb_0_2_io_o_3_out[4] ,
    \cb_0_2_io_o_3_out[3] ,
    \cb_0_2_io_o_3_out[2] ,
    \cb_0_2_io_o_3_out[1] ,
    \cb_0_2_io_o_3_out[0] }),
    .io_o_4_out({\cb_0_2_io_o_4_out[7] ,
    \cb_0_2_io_o_4_out[6] ,
    \cb_0_2_io_o_4_out[5] ,
    \cb_0_2_io_o_4_out[4] ,
    \cb_0_2_io_o_4_out[3] ,
    \cb_0_2_io_o_4_out[2] ,
    \cb_0_2_io_o_4_out[1] ,
    \cb_0_2_io_o_4_out[0] }),
    .io_o_5_out({\cb_0_2_io_o_5_out[7] ,
    \cb_0_2_io_o_5_out[6] ,
    \cb_0_2_io_o_5_out[5] ,
    \cb_0_2_io_o_5_out[4] ,
    \cb_0_2_io_o_5_out[3] ,
    \cb_0_2_io_o_5_out[2] ,
    \cb_0_2_io_o_5_out[1] ,
    \cb_0_2_io_o_5_out[0] }),
    .io_o_6_out({\cb_0_2_io_o_6_out[7] ,
    \cb_0_2_io_o_6_out[6] ,
    \cb_0_2_io_o_6_out[5] ,
    \cb_0_2_io_o_6_out[4] ,
    \cb_0_2_io_o_6_out[3] ,
    \cb_0_2_io_o_6_out[2] ,
    \cb_0_2_io_o_6_out[1] ,
    \cb_0_2_io_o_6_out[0] }),
    .io_o_7_out({\cb_0_2_io_o_7_out[7] ,
    \cb_0_2_io_o_7_out[6] ,
    \cb_0_2_io_o_7_out[5] ,
    \cb_0_2_io_o_7_out[4] ,
    \cb_0_2_io_o_7_out[3] ,
    \cb_0_2_io_o_7_out[2] ,
    \cb_0_2_io_o_7_out[1] ,
    \cb_0_2_io_o_7_out[0] }),
    .io_wo({\cb_0_1_io_eo[63] ,
    \cb_0_1_io_eo[62] ,
    \cb_0_1_io_eo[61] ,
    \cb_0_1_io_eo[60] ,
    \cb_0_1_io_eo[59] ,
    \cb_0_1_io_eo[58] ,
    \cb_0_1_io_eo[57] ,
    \cb_0_1_io_eo[56] ,
    \cb_0_1_io_eo[55] ,
    \cb_0_1_io_eo[54] ,
    \cb_0_1_io_eo[53] ,
    \cb_0_1_io_eo[52] ,
    \cb_0_1_io_eo[51] ,
    \cb_0_1_io_eo[50] ,
    \cb_0_1_io_eo[49] ,
    \cb_0_1_io_eo[48] ,
    \cb_0_1_io_eo[47] ,
    \cb_0_1_io_eo[46] ,
    \cb_0_1_io_eo[45] ,
    \cb_0_1_io_eo[44] ,
    \cb_0_1_io_eo[43] ,
    \cb_0_1_io_eo[42] ,
    \cb_0_1_io_eo[41] ,
    \cb_0_1_io_eo[40] ,
    \cb_0_1_io_eo[39] ,
    \cb_0_1_io_eo[38] ,
    \cb_0_1_io_eo[37] ,
    \cb_0_1_io_eo[36] ,
    \cb_0_1_io_eo[35] ,
    \cb_0_1_io_eo[34] ,
    \cb_0_1_io_eo[33] ,
    \cb_0_1_io_eo[32] ,
    \cb_0_1_io_eo[31] ,
    \cb_0_1_io_eo[30] ,
    \cb_0_1_io_eo[29] ,
    \cb_0_1_io_eo[28] ,
    \cb_0_1_io_eo[27] ,
    \cb_0_1_io_eo[26] ,
    \cb_0_1_io_eo[25] ,
    \cb_0_1_io_eo[24] ,
    \cb_0_1_io_eo[23] ,
    \cb_0_1_io_eo[22] ,
    \cb_0_1_io_eo[21] ,
    \cb_0_1_io_eo[20] ,
    \cb_0_1_io_eo[19] ,
    \cb_0_1_io_eo[18] ,
    \cb_0_1_io_eo[17] ,
    \cb_0_1_io_eo[16] ,
    \cb_0_1_io_eo[15] ,
    \cb_0_1_io_eo[14] ,
    \cb_0_1_io_eo[13] ,
    \cb_0_1_io_eo[12] ,
    \cb_0_1_io_eo[11] ,
    \cb_0_1_io_eo[10] ,
    \cb_0_1_io_eo[9] ,
    \cb_0_1_io_eo[8] ,
    \cb_0_1_io_eo[7] ,
    \cb_0_1_io_eo[6] ,
    \cb_0_1_io_eo[5] ,
    \cb_0_1_io_eo[4] ,
    \cb_0_1_io_eo[3] ,
    \cb_0_1_io_eo[2] ,
    \cb_0_1_io_eo[1] ,
    \cb_0_1_io_eo[0] }));
 cic_block cb_0_3 (.io_cs_i(cb_0_3_io_cs_i),
    .io_i_0_ci(cb_0_2_io_o_0_co),
    .io_i_1_ci(cb_0_2_io_o_1_co),
    .io_i_2_ci(cb_0_2_io_o_2_co),
    .io_i_3_ci(cb_0_2_io_o_3_co),
    .io_i_4_ci(cb_0_2_io_o_4_co),
    .io_i_5_ci(cb_0_2_io_o_5_co),
    .io_i_6_ci(cb_0_2_io_o_6_co),
    .io_i_7_ci(cb_0_2_io_o_7_co),
    .io_o_0_co(cb_0_3_io_o_0_co),
    .io_o_1_co(cb_0_3_io_o_1_co),
    .io_o_2_co(cb_0_3_io_o_2_co),
    .io_o_3_co(cb_0_3_io_o_3_co),
    .io_o_4_co(cb_0_3_io_o_4_co),
    .io_o_5_co(cb_0_3_io_o_5_co),
    .io_o_6_co(cb_0_3_io_o_6_co),
    .io_o_7_co(cb_0_3_io_o_7_co),
    .io_vci(cb_0_2_io_vco),
    .io_vco(cb_0_3_io_vco),
    .io_vi(cb_0_3_io_vi),
    .io_we_i(cb_0_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_0_0_io_adr_i[1] ,
    \cb_0_0_io_adr_i[0] }),
    .io_dat_i({\cb_0_0_io_dat_i[15] ,
    \cb_0_0_io_dat_i[14] ,
    \cb_0_0_io_dat_i[13] ,
    \cb_0_0_io_dat_i[12] ,
    \cb_0_0_io_dat_i[11] ,
    \cb_0_0_io_dat_i[10] ,
    \cb_0_0_io_dat_i[9] ,
    \cb_0_0_io_dat_i[8] ,
    \cb_0_0_io_dat_i[7] ,
    \cb_0_0_io_dat_i[6] ,
    \cb_0_0_io_dat_i[5] ,
    \cb_0_0_io_dat_i[4] ,
    \cb_0_0_io_dat_i[3] ,
    \cb_0_0_io_dat_i[2] ,
    \cb_0_0_io_dat_i[1] ,
    \cb_0_0_io_dat_i[0] }),
    .io_dat_o({\cb_0_3_io_dat_o[15] ,
    \cb_0_3_io_dat_o[14] ,
    \cb_0_3_io_dat_o[13] ,
    \cb_0_3_io_dat_o[12] ,
    \cb_0_3_io_dat_o[11] ,
    \cb_0_3_io_dat_o[10] ,
    \cb_0_3_io_dat_o[9] ,
    \cb_0_3_io_dat_o[8] ,
    \cb_0_3_io_dat_o[7] ,
    \cb_0_3_io_dat_o[6] ,
    \cb_0_3_io_dat_o[5] ,
    \cb_0_3_io_dat_o[4] ,
    \cb_0_3_io_dat_o[3] ,
    \cb_0_3_io_dat_o[2] ,
    \cb_0_3_io_dat_o[1] ,
    \cb_0_3_io_dat_o[0] }),
    .io_eo({\cb_0_3_io_eo[63] ,
    \cb_0_3_io_eo[62] ,
    \cb_0_3_io_eo[61] ,
    \cb_0_3_io_eo[60] ,
    \cb_0_3_io_eo[59] ,
    \cb_0_3_io_eo[58] ,
    \cb_0_3_io_eo[57] ,
    \cb_0_3_io_eo[56] ,
    \cb_0_3_io_eo[55] ,
    \cb_0_3_io_eo[54] ,
    \cb_0_3_io_eo[53] ,
    \cb_0_3_io_eo[52] ,
    \cb_0_3_io_eo[51] ,
    \cb_0_3_io_eo[50] ,
    \cb_0_3_io_eo[49] ,
    \cb_0_3_io_eo[48] ,
    \cb_0_3_io_eo[47] ,
    \cb_0_3_io_eo[46] ,
    \cb_0_3_io_eo[45] ,
    \cb_0_3_io_eo[44] ,
    \cb_0_3_io_eo[43] ,
    \cb_0_3_io_eo[42] ,
    \cb_0_3_io_eo[41] ,
    \cb_0_3_io_eo[40] ,
    \cb_0_3_io_eo[39] ,
    \cb_0_3_io_eo[38] ,
    \cb_0_3_io_eo[37] ,
    \cb_0_3_io_eo[36] ,
    \cb_0_3_io_eo[35] ,
    \cb_0_3_io_eo[34] ,
    \cb_0_3_io_eo[33] ,
    \cb_0_3_io_eo[32] ,
    \cb_0_3_io_eo[31] ,
    \cb_0_3_io_eo[30] ,
    \cb_0_3_io_eo[29] ,
    \cb_0_3_io_eo[28] ,
    \cb_0_3_io_eo[27] ,
    \cb_0_3_io_eo[26] ,
    \cb_0_3_io_eo[25] ,
    \cb_0_3_io_eo[24] ,
    \cb_0_3_io_eo[23] ,
    \cb_0_3_io_eo[22] ,
    \cb_0_3_io_eo[21] ,
    \cb_0_3_io_eo[20] ,
    \cb_0_3_io_eo[19] ,
    \cb_0_3_io_eo[18] ,
    \cb_0_3_io_eo[17] ,
    \cb_0_3_io_eo[16] ,
    \cb_0_3_io_eo[15] ,
    \cb_0_3_io_eo[14] ,
    \cb_0_3_io_eo[13] ,
    \cb_0_3_io_eo[12] ,
    \cb_0_3_io_eo[11] ,
    \cb_0_3_io_eo[10] ,
    \cb_0_3_io_eo[9] ,
    \cb_0_3_io_eo[8] ,
    \cb_0_3_io_eo[7] ,
    \cb_0_3_io_eo[6] ,
    \cb_0_3_io_eo[5] ,
    \cb_0_3_io_eo[4] ,
    \cb_0_3_io_eo[3] ,
    \cb_0_3_io_eo[2] ,
    \cb_0_3_io_eo[1] ,
    \cb_0_3_io_eo[0] }),
    .io_i_0_in1({\cb_0_2_io_o_0_out[7] ,
    \cb_0_2_io_o_0_out[6] ,
    \cb_0_2_io_o_0_out[5] ,
    \cb_0_2_io_o_0_out[4] ,
    \cb_0_2_io_o_0_out[3] ,
    \cb_0_2_io_o_0_out[2] ,
    \cb_0_2_io_o_0_out[1] ,
    \cb_0_2_io_o_0_out[0] }),
    .io_i_1_in1({\cb_0_2_io_o_1_out[7] ,
    \cb_0_2_io_o_1_out[6] ,
    \cb_0_2_io_o_1_out[5] ,
    \cb_0_2_io_o_1_out[4] ,
    \cb_0_2_io_o_1_out[3] ,
    \cb_0_2_io_o_1_out[2] ,
    \cb_0_2_io_o_1_out[1] ,
    \cb_0_2_io_o_1_out[0] }),
    .io_i_2_in1({\cb_0_2_io_o_2_out[7] ,
    \cb_0_2_io_o_2_out[6] ,
    \cb_0_2_io_o_2_out[5] ,
    \cb_0_2_io_o_2_out[4] ,
    \cb_0_2_io_o_2_out[3] ,
    \cb_0_2_io_o_2_out[2] ,
    \cb_0_2_io_o_2_out[1] ,
    \cb_0_2_io_o_2_out[0] }),
    .io_i_3_in1({\cb_0_2_io_o_3_out[7] ,
    \cb_0_2_io_o_3_out[6] ,
    \cb_0_2_io_o_3_out[5] ,
    \cb_0_2_io_o_3_out[4] ,
    \cb_0_2_io_o_3_out[3] ,
    \cb_0_2_io_o_3_out[2] ,
    \cb_0_2_io_o_3_out[1] ,
    \cb_0_2_io_o_3_out[0] }),
    .io_i_4_in1({\cb_0_2_io_o_4_out[7] ,
    \cb_0_2_io_o_4_out[6] ,
    \cb_0_2_io_o_4_out[5] ,
    \cb_0_2_io_o_4_out[4] ,
    \cb_0_2_io_o_4_out[3] ,
    \cb_0_2_io_o_4_out[2] ,
    \cb_0_2_io_o_4_out[1] ,
    \cb_0_2_io_o_4_out[0] }),
    .io_i_5_in1({\cb_0_2_io_o_5_out[7] ,
    \cb_0_2_io_o_5_out[6] ,
    \cb_0_2_io_o_5_out[5] ,
    \cb_0_2_io_o_5_out[4] ,
    \cb_0_2_io_o_5_out[3] ,
    \cb_0_2_io_o_5_out[2] ,
    \cb_0_2_io_o_5_out[1] ,
    \cb_0_2_io_o_5_out[0] }),
    .io_i_6_in1({\cb_0_2_io_o_6_out[7] ,
    \cb_0_2_io_o_6_out[6] ,
    \cb_0_2_io_o_6_out[5] ,
    \cb_0_2_io_o_6_out[4] ,
    \cb_0_2_io_o_6_out[3] ,
    \cb_0_2_io_o_6_out[2] ,
    \cb_0_2_io_o_6_out[1] ,
    \cb_0_2_io_o_6_out[0] }),
    .io_i_7_in1({\cb_0_2_io_o_7_out[7] ,
    \cb_0_2_io_o_7_out[6] ,
    \cb_0_2_io_o_7_out[5] ,
    \cb_0_2_io_o_7_out[4] ,
    \cb_0_2_io_o_7_out[3] ,
    \cb_0_2_io_o_7_out[2] ,
    \cb_0_2_io_o_7_out[1] ,
    \cb_0_2_io_o_7_out[0] }),
    .io_o_0_out({\cb_0_3_io_o_0_out[7] ,
    \cb_0_3_io_o_0_out[6] ,
    \cb_0_3_io_o_0_out[5] ,
    \cb_0_3_io_o_0_out[4] ,
    \cb_0_3_io_o_0_out[3] ,
    \cb_0_3_io_o_0_out[2] ,
    \cb_0_3_io_o_0_out[1] ,
    \cb_0_3_io_o_0_out[0] }),
    .io_o_1_out({\cb_0_3_io_o_1_out[7] ,
    \cb_0_3_io_o_1_out[6] ,
    \cb_0_3_io_o_1_out[5] ,
    \cb_0_3_io_o_1_out[4] ,
    \cb_0_3_io_o_1_out[3] ,
    \cb_0_3_io_o_1_out[2] ,
    \cb_0_3_io_o_1_out[1] ,
    \cb_0_3_io_o_1_out[0] }),
    .io_o_2_out({\cb_0_3_io_o_2_out[7] ,
    \cb_0_3_io_o_2_out[6] ,
    \cb_0_3_io_o_2_out[5] ,
    \cb_0_3_io_o_2_out[4] ,
    \cb_0_3_io_o_2_out[3] ,
    \cb_0_3_io_o_2_out[2] ,
    \cb_0_3_io_o_2_out[1] ,
    \cb_0_3_io_o_2_out[0] }),
    .io_o_3_out({\cb_0_3_io_o_3_out[7] ,
    \cb_0_3_io_o_3_out[6] ,
    \cb_0_3_io_o_3_out[5] ,
    \cb_0_3_io_o_3_out[4] ,
    \cb_0_3_io_o_3_out[3] ,
    \cb_0_3_io_o_3_out[2] ,
    \cb_0_3_io_o_3_out[1] ,
    \cb_0_3_io_o_3_out[0] }),
    .io_o_4_out({\cb_0_3_io_o_4_out[7] ,
    \cb_0_3_io_o_4_out[6] ,
    \cb_0_3_io_o_4_out[5] ,
    \cb_0_3_io_o_4_out[4] ,
    \cb_0_3_io_o_4_out[3] ,
    \cb_0_3_io_o_4_out[2] ,
    \cb_0_3_io_o_4_out[1] ,
    \cb_0_3_io_o_4_out[0] }),
    .io_o_5_out({\cb_0_3_io_o_5_out[7] ,
    \cb_0_3_io_o_5_out[6] ,
    \cb_0_3_io_o_5_out[5] ,
    \cb_0_3_io_o_5_out[4] ,
    \cb_0_3_io_o_5_out[3] ,
    \cb_0_3_io_o_5_out[2] ,
    \cb_0_3_io_o_5_out[1] ,
    \cb_0_3_io_o_5_out[0] }),
    .io_o_6_out({\cb_0_3_io_o_6_out[7] ,
    \cb_0_3_io_o_6_out[6] ,
    \cb_0_3_io_o_6_out[5] ,
    \cb_0_3_io_o_6_out[4] ,
    \cb_0_3_io_o_6_out[3] ,
    \cb_0_3_io_o_6_out[2] ,
    \cb_0_3_io_o_6_out[1] ,
    \cb_0_3_io_o_6_out[0] }),
    .io_o_7_out({\cb_0_3_io_o_7_out[7] ,
    \cb_0_3_io_o_7_out[6] ,
    \cb_0_3_io_o_7_out[5] ,
    \cb_0_3_io_o_7_out[4] ,
    \cb_0_3_io_o_7_out[3] ,
    \cb_0_3_io_o_7_out[2] ,
    \cb_0_3_io_o_7_out[1] ,
    \cb_0_3_io_o_7_out[0] }),
    .io_wo({\cb_0_2_io_eo[63] ,
    \cb_0_2_io_eo[62] ,
    \cb_0_2_io_eo[61] ,
    \cb_0_2_io_eo[60] ,
    \cb_0_2_io_eo[59] ,
    \cb_0_2_io_eo[58] ,
    \cb_0_2_io_eo[57] ,
    \cb_0_2_io_eo[56] ,
    \cb_0_2_io_eo[55] ,
    \cb_0_2_io_eo[54] ,
    \cb_0_2_io_eo[53] ,
    \cb_0_2_io_eo[52] ,
    \cb_0_2_io_eo[51] ,
    \cb_0_2_io_eo[50] ,
    \cb_0_2_io_eo[49] ,
    \cb_0_2_io_eo[48] ,
    \cb_0_2_io_eo[47] ,
    \cb_0_2_io_eo[46] ,
    \cb_0_2_io_eo[45] ,
    \cb_0_2_io_eo[44] ,
    \cb_0_2_io_eo[43] ,
    \cb_0_2_io_eo[42] ,
    \cb_0_2_io_eo[41] ,
    \cb_0_2_io_eo[40] ,
    \cb_0_2_io_eo[39] ,
    \cb_0_2_io_eo[38] ,
    \cb_0_2_io_eo[37] ,
    \cb_0_2_io_eo[36] ,
    \cb_0_2_io_eo[35] ,
    \cb_0_2_io_eo[34] ,
    \cb_0_2_io_eo[33] ,
    \cb_0_2_io_eo[32] ,
    \cb_0_2_io_eo[31] ,
    \cb_0_2_io_eo[30] ,
    \cb_0_2_io_eo[29] ,
    \cb_0_2_io_eo[28] ,
    \cb_0_2_io_eo[27] ,
    \cb_0_2_io_eo[26] ,
    \cb_0_2_io_eo[25] ,
    \cb_0_2_io_eo[24] ,
    \cb_0_2_io_eo[23] ,
    \cb_0_2_io_eo[22] ,
    \cb_0_2_io_eo[21] ,
    \cb_0_2_io_eo[20] ,
    \cb_0_2_io_eo[19] ,
    \cb_0_2_io_eo[18] ,
    \cb_0_2_io_eo[17] ,
    \cb_0_2_io_eo[16] ,
    \cb_0_2_io_eo[15] ,
    \cb_0_2_io_eo[14] ,
    \cb_0_2_io_eo[13] ,
    \cb_0_2_io_eo[12] ,
    \cb_0_2_io_eo[11] ,
    \cb_0_2_io_eo[10] ,
    \cb_0_2_io_eo[9] ,
    \cb_0_2_io_eo[8] ,
    \cb_0_2_io_eo[7] ,
    \cb_0_2_io_eo[6] ,
    \cb_0_2_io_eo[5] ,
    \cb_0_2_io_eo[4] ,
    \cb_0_2_io_eo[3] ,
    \cb_0_2_io_eo[2] ,
    \cb_0_2_io_eo[1] ,
    \cb_0_2_io_eo[0] }));
 cic_block cb_0_4 (.io_cs_i(cb_0_4_io_cs_i),
    .io_i_0_ci(cb_0_3_io_o_0_co),
    .io_i_1_ci(cb_0_3_io_o_1_co),
    .io_i_2_ci(cb_0_3_io_o_2_co),
    .io_i_3_ci(cb_0_3_io_o_3_co),
    .io_i_4_ci(cb_0_3_io_o_4_co),
    .io_i_5_ci(cb_0_3_io_o_5_co),
    .io_i_6_ci(cb_0_3_io_o_6_co),
    .io_i_7_ci(cb_0_3_io_o_7_co),
    .io_o_0_co(cb_0_4_io_o_0_co),
    .io_o_1_co(cb_0_4_io_o_1_co),
    .io_o_2_co(cb_0_4_io_o_2_co),
    .io_o_3_co(cb_0_4_io_o_3_co),
    .io_o_4_co(cb_0_4_io_o_4_co),
    .io_o_5_co(cb_0_4_io_o_5_co),
    .io_o_6_co(cb_0_4_io_o_6_co),
    .io_o_7_co(cb_0_4_io_o_7_co),
    .io_vci(cb_0_3_io_vco),
    .io_vco(cb_0_4_io_vco),
    .io_vi(cb_0_4_io_vi),
    .io_we_i(cb_0_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_0_0_io_adr_i[1] ,
    \cb_0_0_io_adr_i[0] }),
    .io_dat_i({\cb_0_0_io_dat_i[15] ,
    \cb_0_0_io_dat_i[14] ,
    \cb_0_0_io_dat_i[13] ,
    \cb_0_0_io_dat_i[12] ,
    \cb_0_0_io_dat_i[11] ,
    \cb_0_0_io_dat_i[10] ,
    \cb_0_0_io_dat_i[9] ,
    \cb_0_0_io_dat_i[8] ,
    \cb_0_0_io_dat_i[7] ,
    \cb_0_0_io_dat_i[6] ,
    \cb_0_0_io_dat_i[5] ,
    \cb_0_0_io_dat_i[4] ,
    \cb_0_0_io_dat_i[3] ,
    \cb_0_0_io_dat_i[2] ,
    \cb_0_0_io_dat_i[1] ,
    \cb_0_0_io_dat_i[0] }),
    .io_dat_o({\cb_0_4_io_dat_o[15] ,
    \cb_0_4_io_dat_o[14] ,
    \cb_0_4_io_dat_o[13] ,
    \cb_0_4_io_dat_o[12] ,
    \cb_0_4_io_dat_o[11] ,
    \cb_0_4_io_dat_o[10] ,
    \cb_0_4_io_dat_o[9] ,
    \cb_0_4_io_dat_o[8] ,
    \cb_0_4_io_dat_o[7] ,
    \cb_0_4_io_dat_o[6] ,
    \cb_0_4_io_dat_o[5] ,
    \cb_0_4_io_dat_o[4] ,
    \cb_0_4_io_dat_o[3] ,
    \cb_0_4_io_dat_o[2] ,
    \cb_0_4_io_dat_o[1] ,
    \cb_0_4_io_dat_o[0] }),
    .io_eo({\cb_0_4_io_eo[63] ,
    \cb_0_4_io_eo[62] ,
    \cb_0_4_io_eo[61] ,
    \cb_0_4_io_eo[60] ,
    \cb_0_4_io_eo[59] ,
    \cb_0_4_io_eo[58] ,
    \cb_0_4_io_eo[57] ,
    \cb_0_4_io_eo[56] ,
    \cb_0_4_io_eo[55] ,
    \cb_0_4_io_eo[54] ,
    \cb_0_4_io_eo[53] ,
    \cb_0_4_io_eo[52] ,
    \cb_0_4_io_eo[51] ,
    \cb_0_4_io_eo[50] ,
    \cb_0_4_io_eo[49] ,
    \cb_0_4_io_eo[48] ,
    \cb_0_4_io_eo[47] ,
    \cb_0_4_io_eo[46] ,
    \cb_0_4_io_eo[45] ,
    \cb_0_4_io_eo[44] ,
    \cb_0_4_io_eo[43] ,
    \cb_0_4_io_eo[42] ,
    \cb_0_4_io_eo[41] ,
    \cb_0_4_io_eo[40] ,
    \cb_0_4_io_eo[39] ,
    \cb_0_4_io_eo[38] ,
    \cb_0_4_io_eo[37] ,
    \cb_0_4_io_eo[36] ,
    \cb_0_4_io_eo[35] ,
    \cb_0_4_io_eo[34] ,
    \cb_0_4_io_eo[33] ,
    \cb_0_4_io_eo[32] ,
    \cb_0_4_io_eo[31] ,
    \cb_0_4_io_eo[30] ,
    \cb_0_4_io_eo[29] ,
    \cb_0_4_io_eo[28] ,
    \cb_0_4_io_eo[27] ,
    \cb_0_4_io_eo[26] ,
    \cb_0_4_io_eo[25] ,
    \cb_0_4_io_eo[24] ,
    \cb_0_4_io_eo[23] ,
    \cb_0_4_io_eo[22] ,
    \cb_0_4_io_eo[21] ,
    \cb_0_4_io_eo[20] ,
    \cb_0_4_io_eo[19] ,
    \cb_0_4_io_eo[18] ,
    \cb_0_4_io_eo[17] ,
    \cb_0_4_io_eo[16] ,
    \cb_0_4_io_eo[15] ,
    \cb_0_4_io_eo[14] ,
    \cb_0_4_io_eo[13] ,
    \cb_0_4_io_eo[12] ,
    \cb_0_4_io_eo[11] ,
    \cb_0_4_io_eo[10] ,
    \cb_0_4_io_eo[9] ,
    \cb_0_4_io_eo[8] ,
    \cb_0_4_io_eo[7] ,
    \cb_0_4_io_eo[6] ,
    \cb_0_4_io_eo[5] ,
    \cb_0_4_io_eo[4] ,
    \cb_0_4_io_eo[3] ,
    \cb_0_4_io_eo[2] ,
    \cb_0_4_io_eo[1] ,
    \cb_0_4_io_eo[0] }),
    .io_i_0_in1({\cb_0_3_io_o_0_out[7] ,
    \cb_0_3_io_o_0_out[6] ,
    \cb_0_3_io_o_0_out[5] ,
    \cb_0_3_io_o_0_out[4] ,
    \cb_0_3_io_o_0_out[3] ,
    \cb_0_3_io_o_0_out[2] ,
    \cb_0_3_io_o_0_out[1] ,
    \cb_0_3_io_o_0_out[0] }),
    .io_i_1_in1({\cb_0_3_io_o_1_out[7] ,
    \cb_0_3_io_o_1_out[6] ,
    \cb_0_3_io_o_1_out[5] ,
    \cb_0_3_io_o_1_out[4] ,
    \cb_0_3_io_o_1_out[3] ,
    \cb_0_3_io_o_1_out[2] ,
    \cb_0_3_io_o_1_out[1] ,
    \cb_0_3_io_o_1_out[0] }),
    .io_i_2_in1({\cb_0_3_io_o_2_out[7] ,
    \cb_0_3_io_o_2_out[6] ,
    \cb_0_3_io_o_2_out[5] ,
    \cb_0_3_io_o_2_out[4] ,
    \cb_0_3_io_o_2_out[3] ,
    \cb_0_3_io_o_2_out[2] ,
    \cb_0_3_io_o_2_out[1] ,
    \cb_0_3_io_o_2_out[0] }),
    .io_i_3_in1({\cb_0_3_io_o_3_out[7] ,
    \cb_0_3_io_o_3_out[6] ,
    \cb_0_3_io_o_3_out[5] ,
    \cb_0_3_io_o_3_out[4] ,
    \cb_0_3_io_o_3_out[3] ,
    \cb_0_3_io_o_3_out[2] ,
    \cb_0_3_io_o_3_out[1] ,
    \cb_0_3_io_o_3_out[0] }),
    .io_i_4_in1({\cb_0_3_io_o_4_out[7] ,
    \cb_0_3_io_o_4_out[6] ,
    \cb_0_3_io_o_4_out[5] ,
    \cb_0_3_io_o_4_out[4] ,
    \cb_0_3_io_o_4_out[3] ,
    \cb_0_3_io_o_4_out[2] ,
    \cb_0_3_io_o_4_out[1] ,
    \cb_0_3_io_o_4_out[0] }),
    .io_i_5_in1({\cb_0_3_io_o_5_out[7] ,
    \cb_0_3_io_o_5_out[6] ,
    \cb_0_3_io_o_5_out[5] ,
    \cb_0_3_io_o_5_out[4] ,
    \cb_0_3_io_o_5_out[3] ,
    \cb_0_3_io_o_5_out[2] ,
    \cb_0_3_io_o_5_out[1] ,
    \cb_0_3_io_o_5_out[0] }),
    .io_i_6_in1({\cb_0_3_io_o_6_out[7] ,
    \cb_0_3_io_o_6_out[6] ,
    \cb_0_3_io_o_6_out[5] ,
    \cb_0_3_io_o_6_out[4] ,
    \cb_0_3_io_o_6_out[3] ,
    \cb_0_3_io_o_6_out[2] ,
    \cb_0_3_io_o_6_out[1] ,
    \cb_0_3_io_o_6_out[0] }),
    .io_i_7_in1({\cb_0_3_io_o_7_out[7] ,
    \cb_0_3_io_o_7_out[6] ,
    \cb_0_3_io_o_7_out[5] ,
    \cb_0_3_io_o_7_out[4] ,
    \cb_0_3_io_o_7_out[3] ,
    \cb_0_3_io_o_7_out[2] ,
    \cb_0_3_io_o_7_out[1] ,
    \cb_0_3_io_o_7_out[0] }),
    .io_o_0_out({\cb_0_4_io_o_0_out[7] ,
    \cb_0_4_io_o_0_out[6] ,
    \cb_0_4_io_o_0_out[5] ,
    \cb_0_4_io_o_0_out[4] ,
    \cb_0_4_io_o_0_out[3] ,
    \cb_0_4_io_o_0_out[2] ,
    \cb_0_4_io_o_0_out[1] ,
    \cb_0_4_io_o_0_out[0] }),
    .io_o_1_out({\cb_0_4_io_o_1_out[7] ,
    \cb_0_4_io_o_1_out[6] ,
    \cb_0_4_io_o_1_out[5] ,
    \cb_0_4_io_o_1_out[4] ,
    \cb_0_4_io_o_1_out[3] ,
    \cb_0_4_io_o_1_out[2] ,
    \cb_0_4_io_o_1_out[1] ,
    \cb_0_4_io_o_1_out[0] }),
    .io_o_2_out({\cb_0_4_io_o_2_out[7] ,
    \cb_0_4_io_o_2_out[6] ,
    \cb_0_4_io_o_2_out[5] ,
    \cb_0_4_io_o_2_out[4] ,
    \cb_0_4_io_o_2_out[3] ,
    \cb_0_4_io_o_2_out[2] ,
    \cb_0_4_io_o_2_out[1] ,
    \cb_0_4_io_o_2_out[0] }),
    .io_o_3_out({\cb_0_4_io_o_3_out[7] ,
    \cb_0_4_io_o_3_out[6] ,
    \cb_0_4_io_o_3_out[5] ,
    \cb_0_4_io_o_3_out[4] ,
    \cb_0_4_io_o_3_out[3] ,
    \cb_0_4_io_o_3_out[2] ,
    \cb_0_4_io_o_3_out[1] ,
    \cb_0_4_io_o_3_out[0] }),
    .io_o_4_out({\cb_0_4_io_o_4_out[7] ,
    \cb_0_4_io_o_4_out[6] ,
    \cb_0_4_io_o_4_out[5] ,
    \cb_0_4_io_o_4_out[4] ,
    \cb_0_4_io_o_4_out[3] ,
    \cb_0_4_io_o_4_out[2] ,
    \cb_0_4_io_o_4_out[1] ,
    \cb_0_4_io_o_4_out[0] }),
    .io_o_5_out({\cb_0_4_io_o_5_out[7] ,
    \cb_0_4_io_o_5_out[6] ,
    \cb_0_4_io_o_5_out[5] ,
    \cb_0_4_io_o_5_out[4] ,
    \cb_0_4_io_o_5_out[3] ,
    \cb_0_4_io_o_5_out[2] ,
    \cb_0_4_io_o_5_out[1] ,
    \cb_0_4_io_o_5_out[0] }),
    .io_o_6_out({\cb_0_4_io_o_6_out[7] ,
    \cb_0_4_io_o_6_out[6] ,
    \cb_0_4_io_o_6_out[5] ,
    \cb_0_4_io_o_6_out[4] ,
    \cb_0_4_io_o_6_out[3] ,
    \cb_0_4_io_o_6_out[2] ,
    \cb_0_4_io_o_6_out[1] ,
    \cb_0_4_io_o_6_out[0] }),
    .io_o_7_out({\cb_0_4_io_o_7_out[7] ,
    \cb_0_4_io_o_7_out[6] ,
    \cb_0_4_io_o_7_out[5] ,
    \cb_0_4_io_o_7_out[4] ,
    \cb_0_4_io_o_7_out[3] ,
    \cb_0_4_io_o_7_out[2] ,
    \cb_0_4_io_o_7_out[1] ,
    \cb_0_4_io_o_7_out[0] }),
    .io_wo({\cb_0_3_io_eo[63] ,
    \cb_0_3_io_eo[62] ,
    \cb_0_3_io_eo[61] ,
    \cb_0_3_io_eo[60] ,
    \cb_0_3_io_eo[59] ,
    \cb_0_3_io_eo[58] ,
    \cb_0_3_io_eo[57] ,
    \cb_0_3_io_eo[56] ,
    \cb_0_3_io_eo[55] ,
    \cb_0_3_io_eo[54] ,
    \cb_0_3_io_eo[53] ,
    \cb_0_3_io_eo[52] ,
    \cb_0_3_io_eo[51] ,
    \cb_0_3_io_eo[50] ,
    \cb_0_3_io_eo[49] ,
    \cb_0_3_io_eo[48] ,
    \cb_0_3_io_eo[47] ,
    \cb_0_3_io_eo[46] ,
    \cb_0_3_io_eo[45] ,
    \cb_0_3_io_eo[44] ,
    \cb_0_3_io_eo[43] ,
    \cb_0_3_io_eo[42] ,
    \cb_0_3_io_eo[41] ,
    \cb_0_3_io_eo[40] ,
    \cb_0_3_io_eo[39] ,
    \cb_0_3_io_eo[38] ,
    \cb_0_3_io_eo[37] ,
    \cb_0_3_io_eo[36] ,
    \cb_0_3_io_eo[35] ,
    \cb_0_3_io_eo[34] ,
    \cb_0_3_io_eo[33] ,
    \cb_0_3_io_eo[32] ,
    \cb_0_3_io_eo[31] ,
    \cb_0_3_io_eo[30] ,
    \cb_0_3_io_eo[29] ,
    \cb_0_3_io_eo[28] ,
    \cb_0_3_io_eo[27] ,
    \cb_0_3_io_eo[26] ,
    \cb_0_3_io_eo[25] ,
    \cb_0_3_io_eo[24] ,
    \cb_0_3_io_eo[23] ,
    \cb_0_3_io_eo[22] ,
    \cb_0_3_io_eo[21] ,
    \cb_0_3_io_eo[20] ,
    \cb_0_3_io_eo[19] ,
    \cb_0_3_io_eo[18] ,
    \cb_0_3_io_eo[17] ,
    \cb_0_3_io_eo[16] ,
    \cb_0_3_io_eo[15] ,
    \cb_0_3_io_eo[14] ,
    \cb_0_3_io_eo[13] ,
    \cb_0_3_io_eo[12] ,
    \cb_0_3_io_eo[11] ,
    \cb_0_3_io_eo[10] ,
    \cb_0_3_io_eo[9] ,
    \cb_0_3_io_eo[8] ,
    \cb_0_3_io_eo[7] ,
    \cb_0_3_io_eo[6] ,
    \cb_0_3_io_eo[5] ,
    \cb_0_3_io_eo[4] ,
    \cb_0_3_io_eo[3] ,
    \cb_0_3_io_eo[2] ,
    \cb_0_3_io_eo[1] ,
    \cb_0_3_io_eo[0] }));
 cic_block cb_0_5 (.io_cs_i(cb_0_5_io_cs_i),
    .io_i_0_ci(cb_0_4_io_o_0_co),
    .io_i_1_ci(cb_0_4_io_o_1_co),
    .io_i_2_ci(cb_0_4_io_o_2_co),
    .io_i_3_ci(cb_0_4_io_o_3_co),
    .io_i_4_ci(cb_0_4_io_o_4_co),
    .io_i_5_ci(cb_0_4_io_o_5_co),
    .io_i_6_ci(cb_0_4_io_o_6_co),
    .io_i_7_ci(cb_0_4_io_o_7_co),
    .io_o_0_co(cb_0_5_io_o_0_co),
    .io_o_1_co(cb_0_5_io_o_1_co),
    .io_o_2_co(cb_0_5_io_o_2_co),
    .io_o_3_co(cb_0_5_io_o_3_co),
    .io_o_4_co(cb_0_5_io_o_4_co),
    .io_o_5_co(cb_0_5_io_o_5_co),
    .io_o_6_co(cb_0_5_io_o_6_co),
    .io_o_7_co(cb_0_5_io_o_7_co),
    .io_vci(cb_0_4_io_vco),
    .io_vco(cb_0_5_io_vco),
    .io_vi(cb_0_5_io_vi),
    .io_we_i(cb_0_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_0_0_io_adr_i[1] ,
    \cb_0_0_io_adr_i[0] }),
    .io_dat_i({\cb_0_0_io_dat_i[15] ,
    \cb_0_0_io_dat_i[14] ,
    \cb_0_0_io_dat_i[13] ,
    \cb_0_0_io_dat_i[12] ,
    \cb_0_0_io_dat_i[11] ,
    \cb_0_0_io_dat_i[10] ,
    \cb_0_0_io_dat_i[9] ,
    \cb_0_0_io_dat_i[8] ,
    \cb_0_0_io_dat_i[7] ,
    \cb_0_0_io_dat_i[6] ,
    \cb_0_0_io_dat_i[5] ,
    \cb_0_0_io_dat_i[4] ,
    \cb_0_0_io_dat_i[3] ,
    \cb_0_0_io_dat_i[2] ,
    \cb_0_0_io_dat_i[1] ,
    \cb_0_0_io_dat_i[0] }),
    .io_dat_o({\cb_0_5_io_dat_o[15] ,
    \cb_0_5_io_dat_o[14] ,
    \cb_0_5_io_dat_o[13] ,
    \cb_0_5_io_dat_o[12] ,
    \cb_0_5_io_dat_o[11] ,
    \cb_0_5_io_dat_o[10] ,
    \cb_0_5_io_dat_o[9] ,
    \cb_0_5_io_dat_o[8] ,
    \cb_0_5_io_dat_o[7] ,
    \cb_0_5_io_dat_o[6] ,
    \cb_0_5_io_dat_o[5] ,
    \cb_0_5_io_dat_o[4] ,
    \cb_0_5_io_dat_o[3] ,
    \cb_0_5_io_dat_o[2] ,
    \cb_0_5_io_dat_o[1] ,
    \cb_0_5_io_dat_o[0] }),
    .io_eo({\cb_0_5_io_eo[63] ,
    \cb_0_5_io_eo[62] ,
    \cb_0_5_io_eo[61] ,
    \cb_0_5_io_eo[60] ,
    \cb_0_5_io_eo[59] ,
    \cb_0_5_io_eo[58] ,
    \cb_0_5_io_eo[57] ,
    \cb_0_5_io_eo[56] ,
    \cb_0_5_io_eo[55] ,
    \cb_0_5_io_eo[54] ,
    \cb_0_5_io_eo[53] ,
    \cb_0_5_io_eo[52] ,
    \cb_0_5_io_eo[51] ,
    \cb_0_5_io_eo[50] ,
    \cb_0_5_io_eo[49] ,
    \cb_0_5_io_eo[48] ,
    \cb_0_5_io_eo[47] ,
    \cb_0_5_io_eo[46] ,
    \cb_0_5_io_eo[45] ,
    \cb_0_5_io_eo[44] ,
    \cb_0_5_io_eo[43] ,
    \cb_0_5_io_eo[42] ,
    \cb_0_5_io_eo[41] ,
    \cb_0_5_io_eo[40] ,
    \cb_0_5_io_eo[39] ,
    \cb_0_5_io_eo[38] ,
    \cb_0_5_io_eo[37] ,
    \cb_0_5_io_eo[36] ,
    \cb_0_5_io_eo[35] ,
    \cb_0_5_io_eo[34] ,
    \cb_0_5_io_eo[33] ,
    \cb_0_5_io_eo[32] ,
    \cb_0_5_io_eo[31] ,
    \cb_0_5_io_eo[30] ,
    \cb_0_5_io_eo[29] ,
    \cb_0_5_io_eo[28] ,
    \cb_0_5_io_eo[27] ,
    \cb_0_5_io_eo[26] ,
    \cb_0_5_io_eo[25] ,
    \cb_0_5_io_eo[24] ,
    \cb_0_5_io_eo[23] ,
    \cb_0_5_io_eo[22] ,
    \cb_0_5_io_eo[21] ,
    \cb_0_5_io_eo[20] ,
    \cb_0_5_io_eo[19] ,
    \cb_0_5_io_eo[18] ,
    \cb_0_5_io_eo[17] ,
    \cb_0_5_io_eo[16] ,
    \cb_0_5_io_eo[15] ,
    \cb_0_5_io_eo[14] ,
    \cb_0_5_io_eo[13] ,
    \cb_0_5_io_eo[12] ,
    \cb_0_5_io_eo[11] ,
    \cb_0_5_io_eo[10] ,
    \cb_0_5_io_eo[9] ,
    \cb_0_5_io_eo[8] ,
    \cb_0_5_io_eo[7] ,
    \cb_0_5_io_eo[6] ,
    \cb_0_5_io_eo[5] ,
    \cb_0_5_io_eo[4] ,
    \cb_0_5_io_eo[3] ,
    \cb_0_5_io_eo[2] ,
    \cb_0_5_io_eo[1] ,
    \cb_0_5_io_eo[0] }),
    .io_i_0_in1({\cb_0_4_io_o_0_out[7] ,
    \cb_0_4_io_o_0_out[6] ,
    \cb_0_4_io_o_0_out[5] ,
    \cb_0_4_io_o_0_out[4] ,
    \cb_0_4_io_o_0_out[3] ,
    \cb_0_4_io_o_0_out[2] ,
    \cb_0_4_io_o_0_out[1] ,
    \cb_0_4_io_o_0_out[0] }),
    .io_i_1_in1({\cb_0_4_io_o_1_out[7] ,
    \cb_0_4_io_o_1_out[6] ,
    \cb_0_4_io_o_1_out[5] ,
    \cb_0_4_io_o_1_out[4] ,
    \cb_0_4_io_o_1_out[3] ,
    \cb_0_4_io_o_1_out[2] ,
    \cb_0_4_io_o_1_out[1] ,
    \cb_0_4_io_o_1_out[0] }),
    .io_i_2_in1({\cb_0_4_io_o_2_out[7] ,
    \cb_0_4_io_o_2_out[6] ,
    \cb_0_4_io_o_2_out[5] ,
    \cb_0_4_io_o_2_out[4] ,
    \cb_0_4_io_o_2_out[3] ,
    \cb_0_4_io_o_2_out[2] ,
    \cb_0_4_io_o_2_out[1] ,
    \cb_0_4_io_o_2_out[0] }),
    .io_i_3_in1({\cb_0_4_io_o_3_out[7] ,
    \cb_0_4_io_o_3_out[6] ,
    \cb_0_4_io_o_3_out[5] ,
    \cb_0_4_io_o_3_out[4] ,
    \cb_0_4_io_o_3_out[3] ,
    \cb_0_4_io_o_3_out[2] ,
    \cb_0_4_io_o_3_out[1] ,
    \cb_0_4_io_o_3_out[0] }),
    .io_i_4_in1({\cb_0_4_io_o_4_out[7] ,
    \cb_0_4_io_o_4_out[6] ,
    \cb_0_4_io_o_4_out[5] ,
    \cb_0_4_io_o_4_out[4] ,
    \cb_0_4_io_o_4_out[3] ,
    \cb_0_4_io_o_4_out[2] ,
    \cb_0_4_io_o_4_out[1] ,
    \cb_0_4_io_o_4_out[0] }),
    .io_i_5_in1({\cb_0_4_io_o_5_out[7] ,
    \cb_0_4_io_o_5_out[6] ,
    \cb_0_4_io_o_5_out[5] ,
    \cb_0_4_io_o_5_out[4] ,
    \cb_0_4_io_o_5_out[3] ,
    \cb_0_4_io_o_5_out[2] ,
    \cb_0_4_io_o_5_out[1] ,
    \cb_0_4_io_o_5_out[0] }),
    .io_i_6_in1({\cb_0_4_io_o_6_out[7] ,
    \cb_0_4_io_o_6_out[6] ,
    \cb_0_4_io_o_6_out[5] ,
    \cb_0_4_io_o_6_out[4] ,
    \cb_0_4_io_o_6_out[3] ,
    \cb_0_4_io_o_6_out[2] ,
    \cb_0_4_io_o_6_out[1] ,
    \cb_0_4_io_o_6_out[0] }),
    .io_i_7_in1({\cb_0_4_io_o_7_out[7] ,
    \cb_0_4_io_o_7_out[6] ,
    \cb_0_4_io_o_7_out[5] ,
    \cb_0_4_io_o_7_out[4] ,
    \cb_0_4_io_o_7_out[3] ,
    \cb_0_4_io_o_7_out[2] ,
    \cb_0_4_io_o_7_out[1] ,
    \cb_0_4_io_o_7_out[0] }),
    .io_o_0_out({\cb_0_5_io_o_0_out[7] ,
    \cb_0_5_io_o_0_out[6] ,
    \cb_0_5_io_o_0_out[5] ,
    \cb_0_5_io_o_0_out[4] ,
    \cb_0_5_io_o_0_out[3] ,
    \cb_0_5_io_o_0_out[2] ,
    \cb_0_5_io_o_0_out[1] ,
    \cb_0_5_io_o_0_out[0] }),
    .io_o_1_out({\cb_0_5_io_o_1_out[7] ,
    \cb_0_5_io_o_1_out[6] ,
    \cb_0_5_io_o_1_out[5] ,
    \cb_0_5_io_o_1_out[4] ,
    \cb_0_5_io_o_1_out[3] ,
    \cb_0_5_io_o_1_out[2] ,
    \cb_0_5_io_o_1_out[1] ,
    \cb_0_5_io_o_1_out[0] }),
    .io_o_2_out({\cb_0_5_io_o_2_out[7] ,
    \cb_0_5_io_o_2_out[6] ,
    \cb_0_5_io_o_2_out[5] ,
    \cb_0_5_io_o_2_out[4] ,
    \cb_0_5_io_o_2_out[3] ,
    \cb_0_5_io_o_2_out[2] ,
    \cb_0_5_io_o_2_out[1] ,
    \cb_0_5_io_o_2_out[0] }),
    .io_o_3_out({\cb_0_5_io_o_3_out[7] ,
    \cb_0_5_io_o_3_out[6] ,
    \cb_0_5_io_o_3_out[5] ,
    \cb_0_5_io_o_3_out[4] ,
    \cb_0_5_io_o_3_out[3] ,
    \cb_0_5_io_o_3_out[2] ,
    \cb_0_5_io_o_3_out[1] ,
    \cb_0_5_io_o_3_out[0] }),
    .io_o_4_out({\cb_0_5_io_o_4_out[7] ,
    \cb_0_5_io_o_4_out[6] ,
    \cb_0_5_io_o_4_out[5] ,
    \cb_0_5_io_o_4_out[4] ,
    \cb_0_5_io_o_4_out[3] ,
    \cb_0_5_io_o_4_out[2] ,
    \cb_0_5_io_o_4_out[1] ,
    \cb_0_5_io_o_4_out[0] }),
    .io_o_5_out({\cb_0_5_io_o_5_out[7] ,
    \cb_0_5_io_o_5_out[6] ,
    \cb_0_5_io_o_5_out[5] ,
    \cb_0_5_io_o_5_out[4] ,
    \cb_0_5_io_o_5_out[3] ,
    \cb_0_5_io_o_5_out[2] ,
    \cb_0_5_io_o_5_out[1] ,
    \cb_0_5_io_o_5_out[0] }),
    .io_o_6_out({\cb_0_5_io_o_6_out[7] ,
    \cb_0_5_io_o_6_out[6] ,
    \cb_0_5_io_o_6_out[5] ,
    \cb_0_5_io_o_6_out[4] ,
    \cb_0_5_io_o_6_out[3] ,
    \cb_0_5_io_o_6_out[2] ,
    \cb_0_5_io_o_6_out[1] ,
    \cb_0_5_io_o_6_out[0] }),
    .io_o_7_out({\cb_0_5_io_o_7_out[7] ,
    \cb_0_5_io_o_7_out[6] ,
    \cb_0_5_io_o_7_out[5] ,
    \cb_0_5_io_o_7_out[4] ,
    \cb_0_5_io_o_7_out[3] ,
    \cb_0_5_io_o_7_out[2] ,
    \cb_0_5_io_o_7_out[1] ,
    \cb_0_5_io_o_7_out[0] }),
    .io_wo({\cb_0_4_io_eo[63] ,
    \cb_0_4_io_eo[62] ,
    \cb_0_4_io_eo[61] ,
    \cb_0_4_io_eo[60] ,
    \cb_0_4_io_eo[59] ,
    \cb_0_4_io_eo[58] ,
    \cb_0_4_io_eo[57] ,
    \cb_0_4_io_eo[56] ,
    \cb_0_4_io_eo[55] ,
    \cb_0_4_io_eo[54] ,
    \cb_0_4_io_eo[53] ,
    \cb_0_4_io_eo[52] ,
    \cb_0_4_io_eo[51] ,
    \cb_0_4_io_eo[50] ,
    \cb_0_4_io_eo[49] ,
    \cb_0_4_io_eo[48] ,
    \cb_0_4_io_eo[47] ,
    \cb_0_4_io_eo[46] ,
    \cb_0_4_io_eo[45] ,
    \cb_0_4_io_eo[44] ,
    \cb_0_4_io_eo[43] ,
    \cb_0_4_io_eo[42] ,
    \cb_0_4_io_eo[41] ,
    \cb_0_4_io_eo[40] ,
    \cb_0_4_io_eo[39] ,
    \cb_0_4_io_eo[38] ,
    \cb_0_4_io_eo[37] ,
    \cb_0_4_io_eo[36] ,
    \cb_0_4_io_eo[35] ,
    \cb_0_4_io_eo[34] ,
    \cb_0_4_io_eo[33] ,
    \cb_0_4_io_eo[32] ,
    \cb_0_4_io_eo[31] ,
    \cb_0_4_io_eo[30] ,
    \cb_0_4_io_eo[29] ,
    \cb_0_4_io_eo[28] ,
    \cb_0_4_io_eo[27] ,
    \cb_0_4_io_eo[26] ,
    \cb_0_4_io_eo[25] ,
    \cb_0_4_io_eo[24] ,
    \cb_0_4_io_eo[23] ,
    \cb_0_4_io_eo[22] ,
    \cb_0_4_io_eo[21] ,
    \cb_0_4_io_eo[20] ,
    \cb_0_4_io_eo[19] ,
    \cb_0_4_io_eo[18] ,
    \cb_0_4_io_eo[17] ,
    \cb_0_4_io_eo[16] ,
    \cb_0_4_io_eo[15] ,
    \cb_0_4_io_eo[14] ,
    \cb_0_4_io_eo[13] ,
    \cb_0_4_io_eo[12] ,
    \cb_0_4_io_eo[11] ,
    \cb_0_4_io_eo[10] ,
    \cb_0_4_io_eo[9] ,
    \cb_0_4_io_eo[8] ,
    \cb_0_4_io_eo[7] ,
    \cb_0_4_io_eo[6] ,
    \cb_0_4_io_eo[5] ,
    \cb_0_4_io_eo[4] ,
    \cb_0_4_io_eo[3] ,
    \cb_0_4_io_eo[2] ,
    \cb_0_4_io_eo[1] ,
    \cb_0_4_io_eo[0] }));
 cic_block cb_0_6 (.io_cs_i(cb_0_6_io_cs_i),
    .io_i_0_ci(cb_0_5_io_o_0_co),
    .io_i_1_ci(cb_0_5_io_o_1_co),
    .io_i_2_ci(cb_0_5_io_o_2_co),
    .io_i_3_ci(cb_0_5_io_o_3_co),
    .io_i_4_ci(cb_0_5_io_o_4_co),
    .io_i_5_ci(cb_0_5_io_o_5_co),
    .io_i_6_ci(cb_0_5_io_o_6_co),
    .io_i_7_ci(cb_0_5_io_o_7_co),
    .io_o_0_co(cb_0_6_io_o_0_co),
    .io_o_1_co(cb_0_6_io_o_1_co),
    .io_o_2_co(cb_0_6_io_o_2_co),
    .io_o_3_co(cb_0_6_io_o_3_co),
    .io_o_4_co(cb_0_6_io_o_4_co),
    .io_o_5_co(cb_0_6_io_o_5_co),
    .io_o_6_co(cb_0_6_io_o_6_co),
    .io_o_7_co(cb_0_6_io_o_7_co),
    .io_vci(cb_0_5_io_vco),
    .io_vco(cb_0_6_io_vco),
    .io_vi(cb_0_6_io_vi),
    .io_we_i(cb_0_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_0_0_io_adr_i[1] ,
    \cb_0_0_io_adr_i[0] }),
    .io_dat_i({\cb_0_0_io_dat_i[15] ,
    \cb_0_0_io_dat_i[14] ,
    \cb_0_0_io_dat_i[13] ,
    \cb_0_0_io_dat_i[12] ,
    \cb_0_0_io_dat_i[11] ,
    \cb_0_0_io_dat_i[10] ,
    \cb_0_0_io_dat_i[9] ,
    \cb_0_0_io_dat_i[8] ,
    \cb_0_0_io_dat_i[7] ,
    \cb_0_0_io_dat_i[6] ,
    \cb_0_0_io_dat_i[5] ,
    \cb_0_0_io_dat_i[4] ,
    \cb_0_0_io_dat_i[3] ,
    \cb_0_0_io_dat_i[2] ,
    \cb_0_0_io_dat_i[1] ,
    \cb_0_0_io_dat_i[0] }),
    .io_dat_o({\cb_0_6_io_dat_o[15] ,
    \cb_0_6_io_dat_o[14] ,
    \cb_0_6_io_dat_o[13] ,
    \cb_0_6_io_dat_o[12] ,
    \cb_0_6_io_dat_o[11] ,
    \cb_0_6_io_dat_o[10] ,
    \cb_0_6_io_dat_o[9] ,
    \cb_0_6_io_dat_o[8] ,
    \cb_0_6_io_dat_o[7] ,
    \cb_0_6_io_dat_o[6] ,
    \cb_0_6_io_dat_o[5] ,
    \cb_0_6_io_dat_o[4] ,
    \cb_0_6_io_dat_o[3] ,
    \cb_0_6_io_dat_o[2] ,
    \cb_0_6_io_dat_o[1] ,
    \cb_0_6_io_dat_o[0] }),
    .io_eo({\cb_0_6_io_eo[63] ,
    \cb_0_6_io_eo[62] ,
    \cb_0_6_io_eo[61] ,
    \cb_0_6_io_eo[60] ,
    \cb_0_6_io_eo[59] ,
    \cb_0_6_io_eo[58] ,
    \cb_0_6_io_eo[57] ,
    \cb_0_6_io_eo[56] ,
    \cb_0_6_io_eo[55] ,
    \cb_0_6_io_eo[54] ,
    \cb_0_6_io_eo[53] ,
    \cb_0_6_io_eo[52] ,
    \cb_0_6_io_eo[51] ,
    \cb_0_6_io_eo[50] ,
    \cb_0_6_io_eo[49] ,
    \cb_0_6_io_eo[48] ,
    \cb_0_6_io_eo[47] ,
    \cb_0_6_io_eo[46] ,
    \cb_0_6_io_eo[45] ,
    \cb_0_6_io_eo[44] ,
    \cb_0_6_io_eo[43] ,
    \cb_0_6_io_eo[42] ,
    \cb_0_6_io_eo[41] ,
    \cb_0_6_io_eo[40] ,
    \cb_0_6_io_eo[39] ,
    \cb_0_6_io_eo[38] ,
    \cb_0_6_io_eo[37] ,
    \cb_0_6_io_eo[36] ,
    \cb_0_6_io_eo[35] ,
    \cb_0_6_io_eo[34] ,
    \cb_0_6_io_eo[33] ,
    \cb_0_6_io_eo[32] ,
    \cb_0_6_io_eo[31] ,
    \cb_0_6_io_eo[30] ,
    \cb_0_6_io_eo[29] ,
    \cb_0_6_io_eo[28] ,
    \cb_0_6_io_eo[27] ,
    \cb_0_6_io_eo[26] ,
    \cb_0_6_io_eo[25] ,
    \cb_0_6_io_eo[24] ,
    \cb_0_6_io_eo[23] ,
    \cb_0_6_io_eo[22] ,
    \cb_0_6_io_eo[21] ,
    \cb_0_6_io_eo[20] ,
    \cb_0_6_io_eo[19] ,
    \cb_0_6_io_eo[18] ,
    \cb_0_6_io_eo[17] ,
    \cb_0_6_io_eo[16] ,
    \cb_0_6_io_eo[15] ,
    \cb_0_6_io_eo[14] ,
    \cb_0_6_io_eo[13] ,
    \cb_0_6_io_eo[12] ,
    \cb_0_6_io_eo[11] ,
    \cb_0_6_io_eo[10] ,
    \cb_0_6_io_eo[9] ,
    \cb_0_6_io_eo[8] ,
    \cb_0_6_io_eo[7] ,
    \cb_0_6_io_eo[6] ,
    \cb_0_6_io_eo[5] ,
    \cb_0_6_io_eo[4] ,
    \cb_0_6_io_eo[3] ,
    \cb_0_6_io_eo[2] ,
    \cb_0_6_io_eo[1] ,
    \cb_0_6_io_eo[0] }),
    .io_i_0_in1({\cb_0_5_io_o_0_out[7] ,
    \cb_0_5_io_o_0_out[6] ,
    \cb_0_5_io_o_0_out[5] ,
    \cb_0_5_io_o_0_out[4] ,
    \cb_0_5_io_o_0_out[3] ,
    \cb_0_5_io_o_0_out[2] ,
    \cb_0_5_io_o_0_out[1] ,
    \cb_0_5_io_o_0_out[0] }),
    .io_i_1_in1({\cb_0_5_io_o_1_out[7] ,
    \cb_0_5_io_o_1_out[6] ,
    \cb_0_5_io_o_1_out[5] ,
    \cb_0_5_io_o_1_out[4] ,
    \cb_0_5_io_o_1_out[3] ,
    \cb_0_5_io_o_1_out[2] ,
    \cb_0_5_io_o_1_out[1] ,
    \cb_0_5_io_o_1_out[0] }),
    .io_i_2_in1({\cb_0_5_io_o_2_out[7] ,
    \cb_0_5_io_o_2_out[6] ,
    \cb_0_5_io_o_2_out[5] ,
    \cb_0_5_io_o_2_out[4] ,
    \cb_0_5_io_o_2_out[3] ,
    \cb_0_5_io_o_2_out[2] ,
    \cb_0_5_io_o_2_out[1] ,
    \cb_0_5_io_o_2_out[0] }),
    .io_i_3_in1({\cb_0_5_io_o_3_out[7] ,
    \cb_0_5_io_o_3_out[6] ,
    \cb_0_5_io_o_3_out[5] ,
    \cb_0_5_io_o_3_out[4] ,
    \cb_0_5_io_o_3_out[3] ,
    \cb_0_5_io_o_3_out[2] ,
    \cb_0_5_io_o_3_out[1] ,
    \cb_0_5_io_o_3_out[0] }),
    .io_i_4_in1({\cb_0_5_io_o_4_out[7] ,
    \cb_0_5_io_o_4_out[6] ,
    \cb_0_5_io_o_4_out[5] ,
    \cb_0_5_io_o_4_out[4] ,
    \cb_0_5_io_o_4_out[3] ,
    \cb_0_5_io_o_4_out[2] ,
    \cb_0_5_io_o_4_out[1] ,
    \cb_0_5_io_o_4_out[0] }),
    .io_i_5_in1({\cb_0_5_io_o_5_out[7] ,
    \cb_0_5_io_o_5_out[6] ,
    \cb_0_5_io_o_5_out[5] ,
    \cb_0_5_io_o_5_out[4] ,
    \cb_0_5_io_o_5_out[3] ,
    \cb_0_5_io_o_5_out[2] ,
    \cb_0_5_io_o_5_out[1] ,
    \cb_0_5_io_o_5_out[0] }),
    .io_i_6_in1({\cb_0_5_io_o_6_out[7] ,
    \cb_0_5_io_o_6_out[6] ,
    \cb_0_5_io_o_6_out[5] ,
    \cb_0_5_io_o_6_out[4] ,
    \cb_0_5_io_o_6_out[3] ,
    \cb_0_5_io_o_6_out[2] ,
    \cb_0_5_io_o_6_out[1] ,
    \cb_0_5_io_o_6_out[0] }),
    .io_i_7_in1({\cb_0_5_io_o_7_out[7] ,
    \cb_0_5_io_o_7_out[6] ,
    \cb_0_5_io_o_7_out[5] ,
    \cb_0_5_io_o_7_out[4] ,
    \cb_0_5_io_o_7_out[3] ,
    \cb_0_5_io_o_7_out[2] ,
    \cb_0_5_io_o_7_out[1] ,
    \cb_0_5_io_o_7_out[0] }),
    .io_o_0_out({\cb_0_6_io_o_0_out[7] ,
    \cb_0_6_io_o_0_out[6] ,
    \cb_0_6_io_o_0_out[5] ,
    \cb_0_6_io_o_0_out[4] ,
    \cb_0_6_io_o_0_out[3] ,
    \cb_0_6_io_o_0_out[2] ,
    \cb_0_6_io_o_0_out[1] ,
    \cb_0_6_io_o_0_out[0] }),
    .io_o_1_out({\cb_0_6_io_o_1_out[7] ,
    \cb_0_6_io_o_1_out[6] ,
    \cb_0_6_io_o_1_out[5] ,
    \cb_0_6_io_o_1_out[4] ,
    \cb_0_6_io_o_1_out[3] ,
    \cb_0_6_io_o_1_out[2] ,
    \cb_0_6_io_o_1_out[1] ,
    \cb_0_6_io_o_1_out[0] }),
    .io_o_2_out({\cb_0_6_io_o_2_out[7] ,
    \cb_0_6_io_o_2_out[6] ,
    \cb_0_6_io_o_2_out[5] ,
    \cb_0_6_io_o_2_out[4] ,
    \cb_0_6_io_o_2_out[3] ,
    \cb_0_6_io_o_2_out[2] ,
    \cb_0_6_io_o_2_out[1] ,
    \cb_0_6_io_o_2_out[0] }),
    .io_o_3_out({\cb_0_6_io_o_3_out[7] ,
    \cb_0_6_io_o_3_out[6] ,
    \cb_0_6_io_o_3_out[5] ,
    \cb_0_6_io_o_3_out[4] ,
    \cb_0_6_io_o_3_out[3] ,
    \cb_0_6_io_o_3_out[2] ,
    \cb_0_6_io_o_3_out[1] ,
    \cb_0_6_io_o_3_out[0] }),
    .io_o_4_out({\cb_0_6_io_o_4_out[7] ,
    \cb_0_6_io_o_4_out[6] ,
    \cb_0_6_io_o_4_out[5] ,
    \cb_0_6_io_o_4_out[4] ,
    \cb_0_6_io_o_4_out[3] ,
    \cb_0_6_io_o_4_out[2] ,
    \cb_0_6_io_o_4_out[1] ,
    \cb_0_6_io_o_4_out[0] }),
    .io_o_5_out({\cb_0_6_io_o_5_out[7] ,
    \cb_0_6_io_o_5_out[6] ,
    \cb_0_6_io_o_5_out[5] ,
    \cb_0_6_io_o_5_out[4] ,
    \cb_0_6_io_o_5_out[3] ,
    \cb_0_6_io_o_5_out[2] ,
    \cb_0_6_io_o_5_out[1] ,
    \cb_0_6_io_o_5_out[0] }),
    .io_o_6_out({\cb_0_6_io_o_6_out[7] ,
    \cb_0_6_io_o_6_out[6] ,
    \cb_0_6_io_o_6_out[5] ,
    \cb_0_6_io_o_6_out[4] ,
    \cb_0_6_io_o_6_out[3] ,
    \cb_0_6_io_o_6_out[2] ,
    \cb_0_6_io_o_6_out[1] ,
    \cb_0_6_io_o_6_out[0] }),
    .io_o_7_out({\cb_0_6_io_o_7_out[7] ,
    \cb_0_6_io_o_7_out[6] ,
    \cb_0_6_io_o_7_out[5] ,
    \cb_0_6_io_o_7_out[4] ,
    \cb_0_6_io_o_7_out[3] ,
    \cb_0_6_io_o_7_out[2] ,
    \cb_0_6_io_o_7_out[1] ,
    \cb_0_6_io_o_7_out[0] }),
    .io_wo({\cb_0_5_io_eo[63] ,
    \cb_0_5_io_eo[62] ,
    \cb_0_5_io_eo[61] ,
    \cb_0_5_io_eo[60] ,
    \cb_0_5_io_eo[59] ,
    \cb_0_5_io_eo[58] ,
    \cb_0_5_io_eo[57] ,
    \cb_0_5_io_eo[56] ,
    \cb_0_5_io_eo[55] ,
    \cb_0_5_io_eo[54] ,
    \cb_0_5_io_eo[53] ,
    \cb_0_5_io_eo[52] ,
    \cb_0_5_io_eo[51] ,
    \cb_0_5_io_eo[50] ,
    \cb_0_5_io_eo[49] ,
    \cb_0_5_io_eo[48] ,
    \cb_0_5_io_eo[47] ,
    \cb_0_5_io_eo[46] ,
    \cb_0_5_io_eo[45] ,
    \cb_0_5_io_eo[44] ,
    \cb_0_5_io_eo[43] ,
    \cb_0_5_io_eo[42] ,
    \cb_0_5_io_eo[41] ,
    \cb_0_5_io_eo[40] ,
    \cb_0_5_io_eo[39] ,
    \cb_0_5_io_eo[38] ,
    \cb_0_5_io_eo[37] ,
    \cb_0_5_io_eo[36] ,
    \cb_0_5_io_eo[35] ,
    \cb_0_5_io_eo[34] ,
    \cb_0_5_io_eo[33] ,
    \cb_0_5_io_eo[32] ,
    \cb_0_5_io_eo[31] ,
    \cb_0_5_io_eo[30] ,
    \cb_0_5_io_eo[29] ,
    \cb_0_5_io_eo[28] ,
    \cb_0_5_io_eo[27] ,
    \cb_0_5_io_eo[26] ,
    \cb_0_5_io_eo[25] ,
    \cb_0_5_io_eo[24] ,
    \cb_0_5_io_eo[23] ,
    \cb_0_5_io_eo[22] ,
    \cb_0_5_io_eo[21] ,
    \cb_0_5_io_eo[20] ,
    \cb_0_5_io_eo[19] ,
    \cb_0_5_io_eo[18] ,
    \cb_0_5_io_eo[17] ,
    \cb_0_5_io_eo[16] ,
    \cb_0_5_io_eo[15] ,
    \cb_0_5_io_eo[14] ,
    \cb_0_5_io_eo[13] ,
    \cb_0_5_io_eo[12] ,
    \cb_0_5_io_eo[11] ,
    \cb_0_5_io_eo[10] ,
    \cb_0_5_io_eo[9] ,
    \cb_0_5_io_eo[8] ,
    \cb_0_5_io_eo[7] ,
    \cb_0_5_io_eo[6] ,
    \cb_0_5_io_eo[5] ,
    \cb_0_5_io_eo[4] ,
    \cb_0_5_io_eo[3] ,
    \cb_0_5_io_eo[2] ,
    \cb_0_5_io_eo[1] ,
    \cb_0_5_io_eo[0] }));
 cic_block cb_0_7 (.io_cs_i(cb_0_7_io_cs_i),
    .io_i_0_ci(cb_0_6_io_o_0_co),
    .io_i_1_ci(cb_0_6_io_o_1_co),
    .io_i_2_ci(cb_0_6_io_o_2_co),
    .io_i_3_ci(cb_0_6_io_o_3_co),
    .io_i_4_ci(cb_0_6_io_o_4_co),
    .io_i_5_ci(cb_0_6_io_o_5_co),
    .io_i_6_ci(cb_0_6_io_o_6_co),
    .io_i_7_ci(cb_0_6_io_o_7_co),
    .io_o_0_co(cb_0_7_io_o_0_co),
    .io_o_1_co(cb_0_7_io_o_1_co),
    .io_o_2_co(cb_0_7_io_o_2_co),
    .io_o_3_co(cb_0_7_io_o_3_co),
    .io_o_4_co(cb_0_7_io_o_4_co),
    .io_o_5_co(cb_0_7_io_o_5_co),
    .io_o_6_co(cb_0_7_io_o_6_co),
    .io_o_7_co(cb_0_7_io_o_7_co),
    .io_vci(cb_0_6_io_vco),
    .io_vco(cb_0_7_io_vco),
    .io_vi(cb_0_7_io_vi),
    .io_we_i(cb_0_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_0_0_io_adr_i[1] ,
    \cb_0_0_io_adr_i[0] }),
    .io_dat_i({\cb_0_0_io_dat_i[15] ,
    \cb_0_0_io_dat_i[14] ,
    \cb_0_0_io_dat_i[13] ,
    \cb_0_0_io_dat_i[12] ,
    \cb_0_0_io_dat_i[11] ,
    \cb_0_0_io_dat_i[10] ,
    \cb_0_0_io_dat_i[9] ,
    \cb_0_0_io_dat_i[8] ,
    \cb_0_0_io_dat_i[7] ,
    \cb_0_0_io_dat_i[6] ,
    \cb_0_0_io_dat_i[5] ,
    \cb_0_0_io_dat_i[4] ,
    \cb_0_0_io_dat_i[3] ,
    \cb_0_0_io_dat_i[2] ,
    \cb_0_0_io_dat_i[1] ,
    \cb_0_0_io_dat_i[0] }),
    .io_dat_o({\cb_0_7_io_dat_o[15] ,
    \cb_0_7_io_dat_o[14] ,
    \cb_0_7_io_dat_o[13] ,
    \cb_0_7_io_dat_o[12] ,
    \cb_0_7_io_dat_o[11] ,
    \cb_0_7_io_dat_o[10] ,
    \cb_0_7_io_dat_o[9] ,
    \cb_0_7_io_dat_o[8] ,
    \cb_0_7_io_dat_o[7] ,
    \cb_0_7_io_dat_o[6] ,
    \cb_0_7_io_dat_o[5] ,
    \cb_0_7_io_dat_o[4] ,
    \cb_0_7_io_dat_o[3] ,
    \cb_0_7_io_dat_o[2] ,
    \cb_0_7_io_dat_o[1] ,
    \cb_0_7_io_dat_o[0] }),
    .io_eo({\cb_0_7_io_eo[63] ,
    \cb_0_7_io_eo[62] ,
    \cb_0_7_io_eo[61] ,
    \cb_0_7_io_eo[60] ,
    \cb_0_7_io_eo[59] ,
    \cb_0_7_io_eo[58] ,
    \cb_0_7_io_eo[57] ,
    \cb_0_7_io_eo[56] ,
    \cb_0_7_io_eo[55] ,
    \cb_0_7_io_eo[54] ,
    \cb_0_7_io_eo[53] ,
    \cb_0_7_io_eo[52] ,
    \cb_0_7_io_eo[51] ,
    \cb_0_7_io_eo[50] ,
    \cb_0_7_io_eo[49] ,
    \cb_0_7_io_eo[48] ,
    \cb_0_7_io_eo[47] ,
    \cb_0_7_io_eo[46] ,
    \cb_0_7_io_eo[45] ,
    \cb_0_7_io_eo[44] ,
    \cb_0_7_io_eo[43] ,
    \cb_0_7_io_eo[42] ,
    \cb_0_7_io_eo[41] ,
    \cb_0_7_io_eo[40] ,
    \cb_0_7_io_eo[39] ,
    \cb_0_7_io_eo[38] ,
    \cb_0_7_io_eo[37] ,
    \cb_0_7_io_eo[36] ,
    \cb_0_7_io_eo[35] ,
    \cb_0_7_io_eo[34] ,
    \cb_0_7_io_eo[33] ,
    \cb_0_7_io_eo[32] ,
    \cb_0_7_io_eo[31] ,
    \cb_0_7_io_eo[30] ,
    \cb_0_7_io_eo[29] ,
    \cb_0_7_io_eo[28] ,
    \cb_0_7_io_eo[27] ,
    \cb_0_7_io_eo[26] ,
    \cb_0_7_io_eo[25] ,
    \cb_0_7_io_eo[24] ,
    \cb_0_7_io_eo[23] ,
    \cb_0_7_io_eo[22] ,
    \cb_0_7_io_eo[21] ,
    \cb_0_7_io_eo[20] ,
    \cb_0_7_io_eo[19] ,
    \cb_0_7_io_eo[18] ,
    \cb_0_7_io_eo[17] ,
    \cb_0_7_io_eo[16] ,
    \cb_0_7_io_eo[15] ,
    \cb_0_7_io_eo[14] ,
    \cb_0_7_io_eo[13] ,
    \cb_0_7_io_eo[12] ,
    \cb_0_7_io_eo[11] ,
    \cb_0_7_io_eo[10] ,
    \cb_0_7_io_eo[9] ,
    \cb_0_7_io_eo[8] ,
    \cb_0_7_io_eo[7] ,
    \cb_0_7_io_eo[6] ,
    \cb_0_7_io_eo[5] ,
    \cb_0_7_io_eo[4] ,
    \cb_0_7_io_eo[3] ,
    \cb_0_7_io_eo[2] ,
    \cb_0_7_io_eo[1] ,
    \cb_0_7_io_eo[0] }),
    .io_i_0_in1({\cb_0_6_io_o_0_out[7] ,
    \cb_0_6_io_o_0_out[6] ,
    \cb_0_6_io_o_0_out[5] ,
    \cb_0_6_io_o_0_out[4] ,
    \cb_0_6_io_o_0_out[3] ,
    \cb_0_6_io_o_0_out[2] ,
    \cb_0_6_io_o_0_out[1] ,
    \cb_0_6_io_o_0_out[0] }),
    .io_i_1_in1({\cb_0_6_io_o_1_out[7] ,
    \cb_0_6_io_o_1_out[6] ,
    \cb_0_6_io_o_1_out[5] ,
    \cb_0_6_io_o_1_out[4] ,
    \cb_0_6_io_o_1_out[3] ,
    \cb_0_6_io_o_1_out[2] ,
    \cb_0_6_io_o_1_out[1] ,
    \cb_0_6_io_o_1_out[0] }),
    .io_i_2_in1({\cb_0_6_io_o_2_out[7] ,
    \cb_0_6_io_o_2_out[6] ,
    \cb_0_6_io_o_2_out[5] ,
    \cb_0_6_io_o_2_out[4] ,
    \cb_0_6_io_o_2_out[3] ,
    \cb_0_6_io_o_2_out[2] ,
    \cb_0_6_io_o_2_out[1] ,
    \cb_0_6_io_o_2_out[0] }),
    .io_i_3_in1({\cb_0_6_io_o_3_out[7] ,
    \cb_0_6_io_o_3_out[6] ,
    \cb_0_6_io_o_3_out[5] ,
    \cb_0_6_io_o_3_out[4] ,
    \cb_0_6_io_o_3_out[3] ,
    \cb_0_6_io_o_3_out[2] ,
    \cb_0_6_io_o_3_out[1] ,
    \cb_0_6_io_o_3_out[0] }),
    .io_i_4_in1({\cb_0_6_io_o_4_out[7] ,
    \cb_0_6_io_o_4_out[6] ,
    \cb_0_6_io_o_4_out[5] ,
    \cb_0_6_io_o_4_out[4] ,
    \cb_0_6_io_o_4_out[3] ,
    \cb_0_6_io_o_4_out[2] ,
    \cb_0_6_io_o_4_out[1] ,
    \cb_0_6_io_o_4_out[0] }),
    .io_i_5_in1({\cb_0_6_io_o_5_out[7] ,
    \cb_0_6_io_o_5_out[6] ,
    \cb_0_6_io_o_5_out[5] ,
    \cb_0_6_io_o_5_out[4] ,
    \cb_0_6_io_o_5_out[3] ,
    \cb_0_6_io_o_5_out[2] ,
    \cb_0_6_io_o_5_out[1] ,
    \cb_0_6_io_o_5_out[0] }),
    .io_i_6_in1({\cb_0_6_io_o_6_out[7] ,
    \cb_0_6_io_o_6_out[6] ,
    \cb_0_6_io_o_6_out[5] ,
    \cb_0_6_io_o_6_out[4] ,
    \cb_0_6_io_o_6_out[3] ,
    \cb_0_6_io_o_6_out[2] ,
    \cb_0_6_io_o_6_out[1] ,
    \cb_0_6_io_o_6_out[0] }),
    .io_i_7_in1({\cb_0_6_io_o_7_out[7] ,
    \cb_0_6_io_o_7_out[6] ,
    \cb_0_6_io_o_7_out[5] ,
    \cb_0_6_io_o_7_out[4] ,
    \cb_0_6_io_o_7_out[3] ,
    \cb_0_6_io_o_7_out[2] ,
    \cb_0_6_io_o_7_out[1] ,
    \cb_0_6_io_o_7_out[0] }),
    .io_o_0_out({\cb_0_7_io_o_0_out[7] ,
    \cb_0_7_io_o_0_out[6] ,
    \cb_0_7_io_o_0_out[5] ,
    \cb_0_7_io_o_0_out[4] ,
    \cb_0_7_io_o_0_out[3] ,
    \cb_0_7_io_o_0_out[2] ,
    \cb_0_7_io_o_0_out[1] ,
    \cb_0_7_io_o_0_out[0] }),
    .io_o_1_out({\cb_0_7_io_o_1_out[7] ,
    \cb_0_7_io_o_1_out[6] ,
    \cb_0_7_io_o_1_out[5] ,
    \cb_0_7_io_o_1_out[4] ,
    \cb_0_7_io_o_1_out[3] ,
    \cb_0_7_io_o_1_out[2] ,
    \cb_0_7_io_o_1_out[1] ,
    \cb_0_7_io_o_1_out[0] }),
    .io_o_2_out({\cb_0_7_io_o_2_out[7] ,
    \cb_0_7_io_o_2_out[6] ,
    \cb_0_7_io_o_2_out[5] ,
    \cb_0_7_io_o_2_out[4] ,
    \cb_0_7_io_o_2_out[3] ,
    \cb_0_7_io_o_2_out[2] ,
    \cb_0_7_io_o_2_out[1] ,
    \cb_0_7_io_o_2_out[0] }),
    .io_o_3_out({\cb_0_7_io_o_3_out[7] ,
    \cb_0_7_io_o_3_out[6] ,
    \cb_0_7_io_o_3_out[5] ,
    \cb_0_7_io_o_3_out[4] ,
    \cb_0_7_io_o_3_out[3] ,
    \cb_0_7_io_o_3_out[2] ,
    \cb_0_7_io_o_3_out[1] ,
    \cb_0_7_io_o_3_out[0] }),
    .io_o_4_out({\cb_0_7_io_o_4_out[7] ,
    \cb_0_7_io_o_4_out[6] ,
    \cb_0_7_io_o_4_out[5] ,
    \cb_0_7_io_o_4_out[4] ,
    \cb_0_7_io_o_4_out[3] ,
    \cb_0_7_io_o_4_out[2] ,
    \cb_0_7_io_o_4_out[1] ,
    \cb_0_7_io_o_4_out[0] }),
    .io_o_5_out({\cb_0_7_io_o_5_out[7] ,
    \cb_0_7_io_o_5_out[6] ,
    \cb_0_7_io_o_5_out[5] ,
    \cb_0_7_io_o_5_out[4] ,
    \cb_0_7_io_o_5_out[3] ,
    \cb_0_7_io_o_5_out[2] ,
    \cb_0_7_io_o_5_out[1] ,
    \cb_0_7_io_o_5_out[0] }),
    .io_o_6_out({\cb_0_7_io_o_6_out[7] ,
    \cb_0_7_io_o_6_out[6] ,
    \cb_0_7_io_o_6_out[5] ,
    \cb_0_7_io_o_6_out[4] ,
    \cb_0_7_io_o_6_out[3] ,
    \cb_0_7_io_o_6_out[2] ,
    \cb_0_7_io_o_6_out[1] ,
    \cb_0_7_io_o_6_out[0] }),
    .io_o_7_out({\cb_0_7_io_o_7_out[7] ,
    \cb_0_7_io_o_7_out[6] ,
    \cb_0_7_io_o_7_out[5] ,
    \cb_0_7_io_o_7_out[4] ,
    \cb_0_7_io_o_7_out[3] ,
    \cb_0_7_io_o_7_out[2] ,
    \cb_0_7_io_o_7_out[1] ,
    \cb_0_7_io_o_7_out[0] }),
    .io_wo({\cb_0_6_io_eo[63] ,
    \cb_0_6_io_eo[62] ,
    \cb_0_6_io_eo[61] ,
    \cb_0_6_io_eo[60] ,
    \cb_0_6_io_eo[59] ,
    \cb_0_6_io_eo[58] ,
    \cb_0_6_io_eo[57] ,
    \cb_0_6_io_eo[56] ,
    \cb_0_6_io_eo[55] ,
    \cb_0_6_io_eo[54] ,
    \cb_0_6_io_eo[53] ,
    \cb_0_6_io_eo[52] ,
    \cb_0_6_io_eo[51] ,
    \cb_0_6_io_eo[50] ,
    \cb_0_6_io_eo[49] ,
    \cb_0_6_io_eo[48] ,
    \cb_0_6_io_eo[47] ,
    \cb_0_6_io_eo[46] ,
    \cb_0_6_io_eo[45] ,
    \cb_0_6_io_eo[44] ,
    \cb_0_6_io_eo[43] ,
    \cb_0_6_io_eo[42] ,
    \cb_0_6_io_eo[41] ,
    \cb_0_6_io_eo[40] ,
    \cb_0_6_io_eo[39] ,
    \cb_0_6_io_eo[38] ,
    \cb_0_6_io_eo[37] ,
    \cb_0_6_io_eo[36] ,
    \cb_0_6_io_eo[35] ,
    \cb_0_6_io_eo[34] ,
    \cb_0_6_io_eo[33] ,
    \cb_0_6_io_eo[32] ,
    \cb_0_6_io_eo[31] ,
    \cb_0_6_io_eo[30] ,
    \cb_0_6_io_eo[29] ,
    \cb_0_6_io_eo[28] ,
    \cb_0_6_io_eo[27] ,
    \cb_0_6_io_eo[26] ,
    \cb_0_6_io_eo[25] ,
    \cb_0_6_io_eo[24] ,
    \cb_0_6_io_eo[23] ,
    \cb_0_6_io_eo[22] ,
    \cb_0_6_io_eo[21] ,
    \cb_0_6_io_eo[20] ,
    \cb_0_6_io_eo[19] ,
    \cb_0_6_io_eo[18] ,
    \cb_0_6_io_eo[17] ,
    \cb_0_6_io_eo[16] ,
    \cb_0_6_io_eo[15] ,
    \cb_0_6_io_eo[14] ,
    \cb_0_6_io_eo[13] ,
    \cb_0_6_io_eo[12] ,
    \cb_0_6_io_eo[11] ,
    \cb_0_6_io_eo[10] ,
    \cb_0_6_io_eo[9] ,
    \cb_0_6_io_eo[8] ,
    \cb_0_6_io_eo[7] ,
    \cb_0_6_io_eo[6] ,
    \cb_0_6_io_eo[5] ,
    \cb_0_6_io_eo[4] ,
    \cb_0_6_io_eo[3] ,
    \cb_0_6_io_eo[2] ,
    \cb_0_6_io_eo[1] ,
    \cb_0_6_io_eo[0] }));
 cic_block cb_0_8 (.io_cs_i(cb_0_8_io_cs_i),
    .io_i_0_ci(cb_0_7_io_o_0_co),
    .io_i_1_ci(cb_0_7_io_o_1_co),
    .io_i_2_ci(cb_0_7_io_o_2_co),
    .io_i_3_ci(cb_0_7_io_o_3_co),
    .io_i_4_ci(cb_0_7_io_o_4_co),
    .io_i_5_ci(cb_0_7_io_o_5_co),
    .io_i_6_ci(cb_0_7_io_o_6_co),
    .io_i_7_ci(cb_0_7_io_o_7_co),
    .io_o_0_co(cb_0_8_io_o_0_co),
    .io_o_1_co(cb_0_8_io_o_1_co),
    .io_o_2_co(cb_0_8_io_o_2_co),
    .io_o_3_co(cb_0_8_io_o_3_co),
    .io_o_4_co(cb_0_8_io_o_4_co),
    .io_o_5_co(cb_0_8_io_o_5_co),
    .io_o_6_co(cb_0_8_io_o_6_co),
    .io_o_7_co(cb_0_8_io_o_7_co),
    .io_vci(cb_0_7_io_vco),
    .io_vco(cb_0_8_io_vco),
    .io_vi(cb_0_8_io_vi),
    .io_we_i(cb_0_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_0_0_io_adr_i[1] ,
    \cb_0_0_io_adr_i[0] }),
    .io_dat_i({\cb_0_0_io_dat_i[15] ,
    \cb_0_0_io_dat_i[14] ,
    \cb_0_0_io_dat_i[13] ,
    \cb_0_0_io_dat_i[12] ,
    \cb_0_0_io_dat_i[11] ,
    \cb_0_0_io_dat_i[10] ,
    \cb_0_0_io_dat_i[9] ,
    \cb_0_0_io_dat_i[8] ,
    \cb_0_0_io_dat_i[7] ,
    \cb_0_0_io_dat_i[6] ,
    \cb_0_0_io_dat_i[5] ,
    \cb_0_0_io_dat_i[4] ,
    \cb_0_0_io_dat_i[3] ,
    \cb_0_0_io_dat_i[2] ,
    \cb_0_0_io_dat_i[1] ,
    \cb_0_0_io_dat_i[0] }),
    .io_dat_o({\cb_0_8_io_dat_o[15] ,
    \cb_0_8_io_dat_o[14] ,
    \cb_0_8_io_dat_o[13] ,
    \cb_0_8_io_dat_o[12] ,
    \cb_0_8_io_dat_o[11] ,
    \cb_0_8_io_dat_o[10] ,
    \cb_0_8_io_dat_o[9] ,
    \cb_0_8_io_dat_o[8] ,
    \cb_0_8_io_dat_o[7] ,
    \cb_0_8_io_dat_o[6] ,
    \cb_0_8_io_dat_o[5] ,
    \cb_0_8_io_dat_o[4] ,
    \cb_0_8_io_dat_o[3] ,
    \cb_0_8_io_dat_o[2] ,
    \cb_0_8_io_dat_o[1] ,
    \cb_0_8_io_dat_o[0] }),
    .io_eo({\cb_0_8_io_eo[63] ,
    \cb_0_8_io_eo[62] ,
    \cb_0_8_io_eo[61] ,
    \cb_0_8_io_eo[60] ,
    \cb_0_8_io_eo[59] ,
    \cb_0_8_io_eo[58] ,
    \cb_0_8_io_eo[57] ,
    \cb_0_8_io_eo[56] ,
    \cb_0_8_io_eo[55] ,
    \cb_0_8_io_eo[54] ,
    \cb_0_8_io_eo[53] ,
    \cb_0_8_io_eo[52] ,
    \cb_0_8_io_eo[51] ,
    \cb_0_8_io_eo[50] ,
    \cb_0_8_io_eo[49] ,
    \cb_0_8_io_eo[48] ,
    \cb_0_8_io_eo[47] ,
    \cb_0_8_io_eo[46] ,
    \cb_0_8_io_eo[45] ,
    \cb_0_8_io_eo[44] ,
    \cb_0_8_io_eo[43] ,
    \cb_0_8_io_eo[42] ,
    \cb_0_8_io_eo[41] ,
    \cb_0_8_io_eo[40] ,
    \cb_0_8_io_eo[39] ,
    \cb_0_8_io_eo[38] ,
    \cb_0_8_io_eo[37] ,
    \cb_0_8_io_eo[36] ,
    \cb_0_8_io_eo[35] ,
    \cb_0_8_io_eo[34] ,
    \cb_0_8_io_eo[33] ,
    \cb_0_8_io_eo[32] ,
    \cb_0_8_io_eo[31] ,
    \cb_0_8_io_eo[30] ,
    \cb_0_8_io_eo[29] ,
    \cb_0_8_io_eo[28] ,
    \cb_0_8_io_eo[27] ,
    \cb_0_8_io_eo[26] ,
    \cb_0_8_io_eo[25] ,
    \cb_0_8_io_eo[24] ,
    \cb_0_8_io_eo[23] ,
    \cb_0_8_io_eo[22] ,
    \cb_0_8_io_eo[21] ,
    \cb_0_8_io_eo[20] ,
    \cb_0_8_io_eo[19] ,
    \cb_0_8_io_eo[18] ,
    \cb_0_8_io_eo[17] ,
    \cb_0_8_io_eo[16] ,
    \cb_0_8_io_eo[15] ,
    \cb_0_8_io_eo[14] ,
    \cb_0_8_io_eo[13] ,
    \cb_0_8_io_eo[12] ,
    \cb_0_8_io_eo[11] ,
    \cb_0_8_io_eo[10] ,
    \cb_0_8_io_eo[9] ,
    \cb_0_8_io_eo[8] ,
    \cb_0_8_io_eo[7] ,
    \cb_0_8_io_eo[6] ,
    \cb_0_8_io_eo[5] ,
    \cb_0_8_io_eo[4] ,
    \cb_0_8_io_eo[3] ,
    \cb_0_8_io_eo[2] ,
    \cb_0_8_io_eo[1] ,
    \cb_0_8_io_eo[0] }),
    .io_i_0_in1({\cb_0_7_io_o_0_out[7] ,
    \cb_0_7_io_o_0_out[6] ,
    \cb_0_7_io_o_0_out[5] ,
    \cb_0_7_io_o_0_out[4] ,
    \cb_0_7_io_o_0_out[3] ,
    \cb_0_7_io_o_0_out[2] ,
    \cb_0_7_io_o_0_out[1] ,
    \cb_0_7_io_o_0_out[0] }),
    .io_i_1_in1({\cb_0_7_io_o_1_out[7] ,
    \cb_0_7_io_o_1_out[6] ,
    \cb_0_7_io_o_1_out[5] ,
    \cb_0_7_io_o_1_out[4] ,
    \cb_0_7_io_o_1_out[3] ,
    \cb_0_7_io_o_1_out[2] ,
    \cb_0_7_io_o_1_out[1] ,
    \cb_0_7_io_o_1_out[0] }),
    .io_i_2_in1({\cb_0_7_io_o_2_out[7] ,
    \cb_0_7_io_o_2_out[6] ,
    \cb_0_7_io_o_2_out[5] ,
    \cb_0_7_io_o_2_out[4] ,
    \cb_0_7_io_o_2_out[3] ,
    \cb_0_7_io_o_2_out[2] ,
    \cb_0_7_io_o_2_out[1] ,
    \cb_0_7_io_o_2_out[0] }),
    .io_i_3_in1({\cb_0_7_io_o_3_out[7] ,
    \cb_0_7_io_o_3_out[6] ,
    \cb_0_7_io_o_3_out[5] ,
    \cb_0_7_io_o_3_out[4] ,
    \cb_0_7_io_o_3_out[3] ,
    \cb_0_7_io_o_3_out[2] ,
    \cb_0_7_io_o_3_out[1] ,
    \cb_0_7_io_o_3_out[0] }),
    .io_i_4_in1({\cb_0_7_io_o_4_out[7] ,
    \cb_0_7_io_o_4_out[6] ,
    \cb_0_7_io_o_4_out[5] ,
    \cb_0_7_io_o_4_out[4] ,
    \cb_0_7_io_o_4_out[3] ,
    \cb_0_7_io_o_4_out[2] ,
    \cb_0_7_io_o_4_out[1] ,
    \cb_0_7_io_o_4_out[0] }),
    .io_i_5_in1({\cb_0_7_io_o_5_out[7] ,
    \cb_0_7_io_o_5_out[6] ,
    \cb_0_7_io_o_5_out[5] ,
    \cb_0_7_io_o_5_out[4] ,
    \cb_0_7_io_o_5_out[3] ,
    \cb_0_7_io_o_5_out[2] ,
    \cb_0_7_io_o_5_out[1] ,
    \cb_0_7_io_o_5_out[0] }),
    .io_i_6_in1({\cb_0_7_io_o_6_out[7] ,
    \cb_0_7_io_o_6_out[6] ,
    \cb_0_7_io_o_6_out[5] ,
    \cb_0_7_io_o_6_out[4] ,
    \cb_0_7_io_o_6_out[3] ,
    \cb_0_7_io_o_6_out[2] ,
    \cb_0_7_io_o_6_out[1] ,
    \cb_0_7_io_o_6_out[0] }),
    .io_i_7_in1({\cb_0_7_io_o_7_out[7] ,
    \cb_0_7_io_o_7_out[6] ,
    \cb_0_7_io_o_7_out[5] ,
    \cb_0_7_io_o_7_out[4] ,
    \cb_0_7_io_o_7_out[3] ,
    \cb_0_7_io_o_7_out[2] ,
    \cb_0_7_io_o_7_out[1] ,
    \cb_0_7_io_o_7_out[0] }),
    .io_o_0_out({\cb_0_8_io_o_0_out[7] ,
    \cb_0_8_io_o_0_out[6] ,
    \cb_0_8_io_o_0_out[5] ,
    \cb_0_8_io_o_0_out[4] ,
    \cb_0_8_io_o_0_out[3] ,
    \cb_0_8_io_o_0_out[2] ,
    \cb_0_8_io_o_0_out[1] ,
    \cb_0_8_io_o_0_out[0] }),
    .io_o_1_out({\cb_0_8_io_o_1_out[7] ,
    \cb_0_8_io_o_1_out[6] ,
    \cb_0_8_io_o_1_out[5] ,
    \cb_0_8_io_o_1_out[4] ,
    \cb_0_8_io_o_1_out[3] ,
    \cb_0_8_io_o_1_out[2] ,
    \cb_0_8_io_o_1_out[1] ,
    \cb_0_8_io_o_1_out[0] }),
    .io_o_2_out({\cb_0_8_io_o_2_out[7] ,
    \cb_0_8_io_o_2_out[6] ,
    \cb_0_8_io_o_2_out[5] ,
    \cb_0_8_io_o_2_out[4] ,
    \cb_0_8_io_o_2_out[3] ,
    \cb_0_8_io_o_2_out[2] ,
    \cb_0_8_io_o_2_out[1] ,
    \cb_0_8_io_o_2_out[0] }),
    .io_o_3_out({\cb_0_8_io_o_3_out[7] ,
    \cb_0_8_io_o_3_out[6] ,
    \cb_0_8_io_o_3_out[5] ,
    \cb_0_8_io_o_3_out[4] ,
    \cb_0_8_io_o_3_out[3] ,
    \cb_0_8_io_o_3_out[2] ,
    \cb_0_8_io_o_3_out[1] ,
    \cb_0_8_io_o_3_out[0] }),
    .io_o_4_out({\cb_0_8_io_o_4_out[7] ,
    \cb_0_8_io_o_4_out[6] ,
    \cb_0_8_io_o_4_out[5] ,
    \cb_0_8_io_o_4_out[4] ,
    \cb_0_8_io_o_4_out[3] ,
    \cb_0_8_io_o_4_out[2] ,
    \cb_0_8_io_o_4_out[1] ,
    \cb_0_8_io_o_4_out[0] }),
    .io_o_5_out({\cb_0_8_io_o_5_out[7] ,
    \cb_0_8_io_o_5_out[6] ,
    \cb_0_8_io_o_5_out[5] ,
    \cb_0_8_io_o_5_out[4] ,
    \cb_0_8_io_o_5_out[3] ,
    \cb_0_8_io_o_5_out[2] ,
    \cb_0_8_io_o_5_out[1] ,
    \cb_0_8_io_o_5_out[0] }),
    .io_o_6_out({\cb_0_8_io_o_6_out[7] ,
    \cb_0_8_io_o_6_out[6] ,
    \cb_0_8_io_o_6_out[5] ,
    \cb_0_8_io_o_6_out[4] ,
    \cb_0_8_io_o_6_out[3] ,
    \cb_0_8_io_o_6_out[2] ,
    \cb_0_8_io_o_6_out[1] ,
    \cb_0_8_io_o_6_out[0] }),
    .io_o_7_out({\cb_0_8_io_o_7_out[7] ,
    \cb_0_8_io_o_7_out[6] ,
    \cb_0_8_io_o_7_out[5] ,
    \cb_0_8_io_o_7_out[4] ,
    \cb_0_8_io_o_7_out[3] ,
    \cb_0_8_io_o_7_out[2] ,
    \cb_0_8_io_o_7_out[1] ,
    \cb_0_8_io_o_7_out[0] }),
    .io_wo({\cb_0_7_io_eo[63] ,
    \cb_0_7_io_eo[62] ,
    \cb_0_7_io_eo[61] ,
    \cb_0_7_io_eo[60] ,
    \cb_0_7_io_eo[59] ,
    \cb_0_7_io_eo[58] ,
    \cb_0_7_io_eo[57] ,
    \cb_0_7_io_eo[56] ,
    \cb_0_7_io_eo[55] ,
    \cb_0_7_io_eo[54] ,
    \cb_0_7_io_eo[53] ,
    \cb_0_7_io_eo[52] ,
    \cb_0_7_io_eo[51] ,
    \cb_0_7_io_eo[50] ,
    \cb_0_7_io_eo[49] ,
    \cb_0_7_io_eo[48] ,
    \cb_0_7_io_eo[47] ,
    \cb_0_7_io_eo[46] ,
    \cb_0_7_io_eo[45] ,
    \cb_0_7_io_eo[44] ,
    \cb_0_7_io_eo[43] ,
    \cb_0_7_io_eo[42] ,
    \cb_0_7_io_eo[41] ,
    \cb_0_7_io_eo[40] ,
    \cb_0_7_io_eo[39] ,
    \cb_0_7_io_eo[38] ,
    \cb_0_7_io_eo[37] ,
    \cb_0_7_io_eo[36] ,
    \cb_0_7_io_eo[35] ,
    \cb_0_7_io_eo[34] ,
    \cb_0_7_io_eo[33] ,
    \cb_0_7_io_eo[32] ,
    \cb_0_7_io_eo[31] ,
    \cb_0_7_io_eo[30] ,
    \cb_0_7_io_eo[29] ,
    \cb_0_7_io_eo[28] ,
    \cb_0_7_io_eo[27] ,
    \cb_0_7_io_eo[26] ,
    \cb_0_7_io_eo[25] ,
    \cb_0_7_io_eo[24] ,
    \cb_0_7_io_eo[23] ,
    \cb_0_7_io_eo[22] ,
    \cb_0_7_io_eo[21] ,
    \cb_0_7_io_eo[20] ,
    \cb_0_7_io_eo[19] ,
    \cb_0_7_io_eo[18] ,
    \cb_0_7_io_eo[17] ,
    \cb_0_7_io_eo[16] ,
    \cb_0_7_io_eo[15] ,
    \cb_0_7_io_eo[14] ,
    \cb_0_7_io_eo[13] ,
    \cb_0_7_io_eo[12] ,
    \cb_0_7_io_eo[11] ,
    \cb_0_7_io_eo[10] ,
    \cb_0_7_io_eo[9] ,
    \cb_0_7_io_eo[8] ,
    \cb_0_7_io_eo[7] ,
    \cb_0_7_io_eo[6] ,
    \cb_0_7_io_eo[5] ,
    \cb_0_7_io_eo[4] ,
    \cb_0_7_io_eo[3] ,
    \cb_0_7_io_eo[2] ,
    \cb_0_7_io_eo[1] ,
    \cb_0_7_io_eo[0] }));
 cic_block cb_0_9 (.io_cs_i(cb_0_9_io_cs_i),
    .io_i_0_ci(cb_0_8_io_o_0_co),
    .io_i_1_ci(cb_0_8_io_o_1_co),
    .io_i_2_ci(cb_0_8_io_o_2_co),
    .io_i_3_ci(cb_0_8_io_o_3_co),
    .io_i_4_ci(cb_0_8_io_o_4_co),
    .io_i_5_ci(cb_0_8_io_o_5_co),
    .io_i_6_ci(cb_0_8_io_o_6_co),
    .io_i_7_ci(cb_0_8_io_o_7_co),
    .io_o_0_co(cb_0_10_io_i_0_ci),
    .io_o_1_co(cb_0_10_io_i_1_ci),
    .io_o_2_co(cb_0_10_io_i_2_ci),
    .io_o_3_co(cb_0_10_io_i_3_ci),
    .io_o_4_co(cb_0_10_io_i_4_ci),
    .io_o_5_co(cb_0_10_io_i_5_ci),
    .io_o_6_co(cb_0_10_io_i_6_ci),
    .io_o_7_co(cb_0_10_io_i_7_ci),
    .io_vci(cb_0_8_io_vco),
    .io_vco(cb_0_10_io_vci),
    .io_vi(cb_0_9_io_vi),
    .io_we_i(cb_0_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_0_0_io_adr_i[1] ,
    \cb_0_0_io_adr_i[0] }),
    .io_dat_i({\cb_0_0_io_dat_i[15] ,
    \cb_0_0_io_dat_i[14] ,
    \cb_0_0_io_dat_i[13] ,
    \cb_0_0_io_dat_i[12] ,
    \cb_0_0_io_dat_i[11] ,
    \cb_0_0_io_dat_i[10] ,
    \cb_0_0_io_dat_i[9] ,
    \cb_0_0_io_dat_i[8] ,
    \cb_0_0_io_dat_i[7] ,
    \cb_0_0_io_dat_i[6] ,
    \cb_0_0_io_dat_i[5] ,
    \cb_0_0_io_dat_i[4] ,
    \cb_0_0_io_dat_i[3] ,
    \cb_0_0_io_dat_i[2] ,
    \cb_0_0_io_dat_i[1] ,
    \cb_0_0_io_dat_i[0] }),
    .io_dat_o({\cb_0_9_io_dat_o[15] ,
    \cb_0_9_io_dat_o[14] ,
    \cb_0_9_io_dat_o[13] ,
    \cb_0_9_io_dat_o[12] ,
    \cb_0_9_io_dat_o[11] ,
    \cb_0_9_io_dat_o[10] ,
    \cb_0_9_io_dat_o[9] ,
    \cb_0_9_io_dat_o[8] ,
    \cb_0_9_io_dat_o[7] ,
    \cb_0_9_io_dat_o[6] ,
    \cb_0_9_io_dat_o[5] ,
    \cb_0_9_io_dat_o[4] ,
    \cb_0_9_io_dat_o[3] ,
    \cb_0_9_io_dat_o[2] ,
    \cb_0_9_io_dat_o[1] ,
    \cb_0_9_io_dat_o[0] }),
    .io_eo({\cb_0_10_io_wo[63] ,
    \cb_0_10_io_wo[62] ,
    \cb_0_10_io_wo[61] ,
    \cb_0_10_io_wo[60] ,
    \cb_0_10_io_wo[59] ,
    \cb_0_10_io_wo[58] ,
    \cb_0_10_io_wo[57] ,
    \cb_0_10_io_wo[56] ,
    \cb_0_10_io_wo[55] ,
    \cb_0_10_io_wo[54] ,
    \cb_0_10_io_wo[53] ,
    \cb_0_10_io_wo[52] ,
    \cb_0_10_io_wo[51] ,
    \cb_0_10_io_wo[50] ,
    \cb_0_10_io_wo[49] ,
    \cb_0_10_io_wo[48] ,
    \cb_0_10_io_wo[47] ,
    \cb_0_10_io_wo[46] ,
    \cb_0_10_io_wo[45] ,
    \cb_0_10_io_wo[44] ,
    \cb_0_10_io_wo[43] ,
    \cb_0_10_io_wo[42] ,
    \cb_0_10_io_wo[41] ,
    \cb_0_10_io_wo[40] ,
    \cb_0_10_io_wo[39] ,
    \cb_0_10_io_wo[38] ,
    \cb_0_10_io_wo[37] ,
    \cb_0_10_io_wo[36] ,
    \cb_0_10_io_wo[35] ,
    \cb_0_10_io_wo[34] ,
    \cb_0_10_io_wo[33] ,
    \cb_0_10_io_wo[32] ,
    \cb_0_10_io_wo[31] ,
    \cb_0_10_io_wo[30] ,
    \cb_0_10_io_wo[29] ,
    \cb_0_10_io_wo[28] ,
    \cb_0_10_io_wo[27] ,
    \cb_0_10_io_wo[26] ,
    \cb_0_10_io_wo[25] ,
    \cb_0_10_io_wo[24] ,
    \cb_0_10_io_wo[23] ,
    \cb_0_10_io_wo[22] ,
    \cb_0_10_io_wo[21] ,
    \cb_0_10_io_wo[20] ,
    \cb_0_10_io_wo[19] ,
    \cb_0_10_io_wo[18] ,
    \cb_0_10_io_wo[17] ,
    \cb_0_10_io_wo[16] ,
    \cb_0_10_io_wo[15] ,
    \cb_0_10_io_wo[14] ,
    \cb_0_10_io_wo[13] ,
    \cb_0_10_io_wo[12] ,
    \cb_0_10_io_wo[11] ,
    \cb_0_10_io_wo[10] ,
    \cb_0_10_io_wo[9] ,
    \cb_0_10_io_wo[8] ,
    \cb_0_10_io_wo[7] ,
    \cb_0_10_io_wo[6] ,
    \cb_0_10_io_wo[5] ,
    \cb_0_10_io_wo[4] ,
    \cb_0_10_io_wo[3] ,
    \cb_0_10_io_wo[2] ,
    \cb_0_10_io_wo[1] ,
    \cb_0_10_io_wo[0] }),
    .io_i_0_in1({\cb_0_8_io_o_0_out[7] ,
    \cb_0_8_io_o_0_out[6] ,
    \cb_0_8_io_o_0_out[5] ,
    \cb_0_8_io_o_0_out[4] ,
    \cb_0_8_io_o_0_out[3] ,
    \cb_0_8_io_o_0_out[2] ,
    \cb_0_8_io_o_0_out[1] ,
    \cb_0_8_io_o_0_out[0] }),
    .io_i_1_in1({\cb_0_8_io_o_1_out[7] ,
    \cb_0_8_io_o_1_out[6] ,
    \cb_0_8_io_o_1_out[5] ,
    \cb_0_8_io_o_1_out[4] ,
    \cb_0_8_io_o_1_out[3] ,
    \cb_0_8_io_o_1_out[2] ,
    \cb_0_8_io_o_1_out[1] ,
    \cb_0_8_io_o_1_out[0] }),
    .io_i_2_in1({\cb_0_8_io_o_2_out[7] ,
    \cb_0_8_io_o_2_out[6] ,
    \cb_0_8_io_o_2_out[5] ,
    \cb_0_8_io_o_2_out[4] ,
    \cb_0_8_io_o_2_out[3] ,
    \cb_0_8_io_o_2_out[2] ,
    \cb_0_8_io_o_2_out[1] ,
    \cb_0_8_io_o_2_out[0] }),
    .io_i_3_in1({\cb_0_8_io_o_3_out[7] ,
    \cb_0_8_io_o_3_out[6] ,
    \cb_0_8_io_o_3_out[5] ,
    \cb_0_8_io_o_3_out[4] ,
    \cb_0_8_io_o_3_out[3] ,
    \cb_0_8_io_o_3_out[2] ,
    \cb_0_8_io_o_3_out[1] ,
    \cb_0_8_io_o_3_out[0] }),
    .io_i_4_in1({\cb_0_8_io_o_4_out[7] ,
    \cb_0_8_io_o_4_out[6] ,
    \cb_0_8_io_o_4_out[5] ,
    \cb_0_8_io_o_4_out[4] ,
    \cb_0_8_io_o_4_out[3] ,
    \cb_0_8_io_o_4_out[2] ,
    \cb_0_8_io_o_4_out[1] ,
    \cb_0_8_io_o_4_out[0] }),
    .io_i_5_in1({\cb_0_8_io_o_5_out[7] ,
    \cb_0_8_io_o_5_out[6] ,
    \cb_0_8_io_o_5_out[5] ,
    \cb_0_8_io_o_5_out[4] ,
    \cb_0_8_io_o_5_out[3] ,
    \cb_0_8_io_o_5_out[2] ,
    \cb_0_8_io_o_5_out[1] ,
    \cb_0_8_io_o_5_out[0] }),
    .io_i_6_in1({\cb_0_8_io_o_6_out[7] ,
    \cb_0_8_io_o_6_out[6] ,
    \cb_0_8_io_o_6_out[5] ,
    \cb_0_8_io_o_6_out[4] ,
    \cb_0_8_io_o_6_out[3] ,
    \cb_0_8_io_o_6_out[2] ,
    \cb_0_8_io_o_6_out[1] ,
    \cb_0_8_io_o_6_out[0] }),
    .io_i_7_in1({\cb_0_8_io_o_7_out[7] ,
    \cb_0_8_io_o_7_out[6] ,
    \cb_0_8_io_o_7_out[5] ,
    \cb_0_8_io_o_7_out[4] ,
    \cb_0_8_io_o_7_out[3] ,
    \cb_0_8_io_o_7_out[2] ,
    \cb_0_8_io_o_7_out[1] ,
    \cb_0_8_io_o_7_out[0] }),
    .io_o_0_out({\cb_0_10_io_i_0_in1[7] ,
    \cb_0_10_io_i_0_in1[6] ,
    \cb_0_10_io_i_0_in1[5] ,
    \cb_0_10_io_i_0_in1[4] ,
    \cb_0_10_io_i_0_in1[3] ,
    \cb_0_10_io_i_0_in1[2] ,
    \cb_0_10_io_i_0_in1[1] ,
    \cb_0_10_io_i_0_in1[0] }),
    .io_o_1_out({\cb_0_10_io_i_1_in1[7] ,
    \cb_0_10_io_i_1_in1[6] ,
    \cb_0_10_io_i_1_in1[5] ,
    \cb_0_10_io_i_1_in1[4] ,
    \cb_0_10_io_i_1_in1[3] ,
    \cb_0_10_io_i_1_in1[2] ,
    \cb_0_10_io_i_1_in1[1] ,
    \cb_0_10_io_i_1_in1[0] }),
    .io_o_2_out({\cb_0_10_io_i_2_in1[7] ,
    \cb_0_10_io_i_2_in1[6] ,
    \cb_0_10_io_i_2_in1[5] ,
    \cb_0_10_io_i_2_in1[4] ,
    \cb_0_10_io_i_2_in1[3] ,
    \cb_0_10_io_i_2_in1[2] ,
    \cb_0_10_io_i_2_in1[1] ,
    \cb_0_10_io_i_2_in1[0] }),
    .io_o_3_out({\cb_0_10_io_i_3_in1[7] ,
    \cb_0_10_io_i_3_in1[6] ,
    \cb_0_10_io_i_3_in1[5] ,
    \cb_0_10_io_i_3_in1[4] ,
    \cb_0_10_io_i_3_in1[3] ,
    \cb_0_10_io_i_3_in1[2] ,
    \cb_0_10_io_i_3_in1[1] ,
    \cb_0_10_io_i_3_in1[0] }),
    .io_o_4_out({\cb_0_10_io_i_4_in1[7] ,
    \cb_0_10_io_i_4_in1[6] ,
    \cb_0_10_io_i_4_in1[5] ,
    \cb_0_10_io_i_4_in1[4] ,
    \cb_0_10_io_i_4_in1[3] ,
    \cb_0_10_io_i_4_in1[2] ,
    \cb_0_10_io_i_4_in1[1] ,
    \cb_0_10_io_i_4_in1[0] }),
    .io_o_5_out({\cb_0_10_io_i_5_in1[7] ,
    \cb_0_10_io_i_5_in1[6] ,
    \cb_0_10_io_i_5_in1[5] ,
    \cb_0_10_io_i_5_in1[4] ,
    \cb_0_10_io_i_5_in1[3] ,
    \cb_0_10_io_i_5_in1[2] ,
    \cb_0_10_io_i_5_in1[1] ,
    \cb_0_10_io_i_5_in1[0] }),
    .io_o_6_out({\cb_0_10_io_i_6_in1[7] ,
    \cb_0_10_io_i_6_in1[6] ,
    \cb_0_10_io_i_6_in1[5] ,
    \cb_0_10_io_i_6_in1[4] ,
    \cb_0_10_io_i_6_in1[3] ,
    \cb_0_10_io_i_6_in1[2] ,
    \cb_0_10_io_i_6_in1[1] ,
    \cb_0_10_io_i_6_in1[0] }),
    .io_o_7_out({\cb_0_10_io_i_7_in1[7] ,
    \cb_0_10_io_i_7_in1[6] ,
    \cb_0_10_io_i_7_in1[5] ,
    \cb_0_10_io_i_7_in1[4] ,
    \cb_0_10_io_i_7_in1[3] ,
    \cb_0_10_io_i_7_in1[2] ,
    \cb_0_10_io_i_7_in1[1] ,
    \cb_0_10_io_i_7_in1[0] }),
    .io_wo({\cb_0_8_io_eo[63] ,
    \cb_0_8_io_eo[62] ,
    \cb_0_8_io_eo[61] ,
    \cb_0_8_io_eo[60] ,
    \cb_0_8_io_eo[59] ,
    \cb_0_8_io_eo[58] ,
    \cb_0_8_io_eo[57] ,
    \cb_0_8_io_eo[56] ,
    \cb_0_8_io_eo[55] ,
    \cb_0_8_io_eo[54] ,
    \cb_0_8_io_eo[53] ,
    \cb_0_8_io_eo[52] ,
    \cb_0_8_io_eo[51] ,
    \cb_0_8_io_eo[50] ,
    \cb_0_8_io_eo[49] ,
    \cb_0_8_io_eo[48] ,
    \cb_0_8_io_eo[47] ,
    \cb_0_8_io_eo[46] ,
    \cb_0_8_io_eo[45] ,
    \cb_0_8_io_eo[44] ,
    \cb_0_8_io_eo[43] ,
    \cb_0_8_io_eo[42] ,
    \cb_0_8_io_eo[41] ,
    \cb_0_8_io_eo[40] ,
    \cb_0_8_io_eo[39] ,
    \cb_0_8_io_eo[38] ,
    \cb_0_8_io_eo[37] ,
    \cb_0_8_io_eo[36] ,
    \cb_0_8_io_eo[35] ,
    \cb_0_8_io_eo[34] ,
    \cb_0_8_io_eo[33] ,
    \cb_0_8_io_eo[32] ,
    \cb_0_8_io_eo[31] ,
    \cb_0_8_io_eo[30] ,
    \cb_0_8_io_eo[29] ,
    \cb_0_8_io_eo[28] ,
    \cb_0_8_io_eo[27] ,
    \cb_0_8_io_eo[26] ,
    \cb_0_8_io_eo[25] ,
    \cb_0_8_io_eo[24] ,
    \cb_0_8_io_eo[23] ,
    \cb_0_8_io_eo[22] ,
    \cb_0_8_io_eo[21] ,
    \cb_0_8_io_eo[20] ,
    \cb_0_8_io_eo[19] ,
    \cb_0_8_io_eo[18] ,
    \cb_0_8_io_eo[17] ,
    \cb_0_8_io_eo[16] ,
    \cb_0_8_io_eo[15] ,
    \cb_0_8_io_eo[14] ,
    \cb_0_8_io_eo[13] ,
    \cb_0_8_io_eo[12] ,
    \cb_0_8_io_eo[11] ,
    \cb_0_8_io_eo[10] ,
    \cb_0_8_io_eo[9] ,
    \cb_0_8_io_eo[8] ,
    \cb_0_8_io_eo[7] ,
    \cb_0_8_io_eo[6] ,
    \cb_0_8_io_eo[5] ,
    \cb_0_8_io_eo[4] ,
    \cb_0_8_io_eo[3] ,
    \cb_0_8_io_eo[2] ,
    \cb_0_8_io_eo[1] ,
    \cb_0_8_io_eo[0] }));
 cic_block cb_1_0 (.io_cs_i(cb_1_0_io_cs_i),
    .io_i_0_ci(cb_1_0_io_i_0_ci),
    .io_o_0_co(cb_1_0_io_o_0_co),
    .io_o_1_co(cb_1_0_io_o_1_co),
    .io_o_2_co(cb_1_0_io_o_2_co),
    .io_o_3_co(cb_1_0_io_o_3_co),
    .io_o_4_co(cb_1_0_io_o_4_co),
    .io_o_5_co(cb_1_0_io_o_5_co),
    .io_o_6_co(cb_1_0_io_o_6_co),
    .io_o_7_co(cb_1_0_io_o_7_co),
    .io_vco(cb_1_0_io_vco),
    .io_vi(cb_1_0_io_vi),
    .io_we_i(cb_1_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_1_0_io_adr_i[1] ,
    \cb_1_0_io_adr_i[0] }),
    .io_dat_i({\cb_1_0_io_dat_i[15] ,
    \cb_1_0_io_dat_i[14] ,
    \cb_1_0_io_dat_i[13] ,
    \cb_1_0_io_dat_i[12] ,
    \cb_1_0_io_dat_i[11] ,
    \cb_1_0_io_dat_i[10] ,
    \cb_1_0_io_dat_i[9] ,
    \cb_1_0_io_dat_i[8] ,
    \cb_1_0_io_dat_i[7] ,
    \cb_1_0_io_dat_i[6] ,
    \cb_1_0_io_dat_i[5] ,
    \cb_1_0_io_dat_i[4] ,
    \cb_1_0_io_dat_i[3] ,
    \cb_1_0_io_dat_i[2] ,
    \cb_1_0_io_dat_i[1] ,
    \cb_1_0_io_dat_i[0] }),
    .io_dat_o({\cb_1_0_io_dat_o[15] ,
    \cb_1_0_io_dat_o[14] ,
    \cb_1_0_io_dat_o[13] ,
    \cb_1_0_io_dat_o[12] ,
    \cb_1_0_io_dat_o[11] ,
    \cb_1_0_io_dat_o[10] ,
    \cb_1_0_io_dat_o[9] ,
    \cb_1_0_io_dat_o[8] ,
    \cb_1_0_io_dat_o[7] ,
    \cb_1_0_io_dat_o[6] ,
    \cb_1_0_io_dat_o[5] ,
    \cb_1_0_io_dat_o[4] ,
    \cb_1_0_io_dat_o[3] ,
    \cb_1_0_io_dat_o[2] ,
    \cb_1_0_io_dat_o[1] ,
    \cb_1_0_io_dat_o[0] }),
    .io_eo({\cb_1_0_io_eo[63] ,
    \cb_1_0_io_eo[62] ,
    \cb_1_0_io_eo[61] ,
    \cb_1_0_io_eo[60] ,
    \cb_1_0_io_eo[59] ,
    \cb_1_0_io_eo[58] ,
    \cb_1_0_io_eo[57] ,
    \cb_1_0_io_eo[56] ,
    \cb_1_0_io_eo[55] ,
    \cb_1_0_io_eo[54] ,
    \cb_1_0_io_eo[53] ,
    \cb_1_0_io_eo[52] ,
    \cb_1_0_io_eo[51] ,
    \cb_1_0_io_eo[50] ,
    \cb_1_0_io_eo[49] ,
    \cb_1_0_io_eo[48] ,
    \cb_1_0_io_eo[47] ,
    \cb_1_0_io_eo[46] ,
    \cb_1_0_io_eo[45] ,
    \cb_1_0_io_eo[44] ,
    \cb_1_0_io_eo[43] ,
    \cb_1_0_io_eo[42] ,
    \cb_1_0_io_eo[41] ,
    \cb_1_0_io_eo[40] ,
    \cb_1_0_io_eo[39] ,
    \cb_1_0_io_eo[38] ,
    \cb_1_0_io_eo[37] ,
    \cb_1_0_io_eo[36] ,
    \cb_1_0_io_eo[35] ,
    \cb_1_0_io_eo[34] ,
    \cb_1_0_io_eo[33] ,
    \cb_1_0_io_eo[32] ,
    \cb_1_0_io_eo[31] ,
    \cb_1_0_io_eo[30] ,
    \cb_1_0_io_eo[29] ,
    \cb_1_0_io_eo[28] ,
    \cb_1_0_io_eo[27] ,
    \cb_1_0_io_eo[26] ,
    \cb_1_0_io_eo[25] ,
    \cb_1_0_io_eo[24] ,
    \cb_1_0_io_eo[23] ,
    \cb_1_0_io_eo[22] ,
    \cb_1_0_io_eo[21] ,
    \cb_1_0_io_eo[20] ,
    \cb_1_0_io_eo[19] ,
    \cb_1_0_io_eo[18] ,
    \cb_1_0_io_eo[17] ,
    \cb_1_0_io_eo[16] ,
    \cb_1_0_io_eo[15] ,
    \cb_1_0_io_eo[14] ,
    \cb_1_0_io_eo[13] ,
    \cb_1_0_io_eo[12] ,
    \cb_1_0_io_eo[11] ,
    \cb_1_0_io_eo[10] ,
    \cb_1_0_io_eo[9] ,
    \cb_1_0_io_eo[8] ,
    \cb_1_0_io_eo[7] ,
    \cb_1_0_io_eo[6] ,
    \cb_1_0_io_eo[5] ,
    \cb_1_0_io_eo[4] ,
    \cb_1_0_io_eo[3] ,
    \cb_1_0_io_eo[2] ,
    \cb_1_0_io_eo[1] ,
    \cb_1_0_io_eo[0] }),
    .io_i_0_in1({_NC65,
    _NC66,
    _NC67,
    _NC68,
    _NC69,
    _NC70,
    _NC71,
    _NC72}),
    .io_i_1_in1({_NC73,
    _NC74,
    _NC75,
    _NC76,
    _NC77,
    _NC78,
    _NC79,
    _NC80}),
    .io_i_2_in1({_NC81,
    _NC82,
    _NC83,
    _NC84,
    _NC85,
    _NC86,
    _NC87,
    _NC88}),
    .io_i_3_in1({_NC89,
    _NC90,
    _NC91,
    _NC92,
    _NC93,
    _NC94,
    _NC95,
    _NC96}),
    .io_i_4_in1({_NC97,
    _NC98,
    _NC99,
    _NC100,
    _NC101,
    _NC102,
    _NC103,
    _NC104}),
    .io_i_5_in1({_NC105,
    _NC106,
    _NC107,
    _NC108,
    _NC109,
    _NC110,
    _NC111,
    _NC112}),
    .io_i_6_in1({_NC113,
    _NC114,
    _NC115,
    _NC116,
    _NC117,
    _NC118,
    _NC119,
    _NC120}),
    .io_i_7_in1({_NC121,
    _NC122,
    _NC123,
    _NC124,
    _NC125,
    _NC126,
    _NC127,
    _NC128}),
    .io_o_0_out({\cb_1_0_io_o_0_out[7] ,
    \cb_1_0_io_o_0_out[6] ,
    \cb_1_0_io_o_0_out[5] ,
    \cb_1_0_io_o_0_out[4] ,
    \cb_1_0_io_o_0_out[3] ,
    \cb_1_0_io_o_0_out[2] ,
    \cb_1_0_io_o_0_out[1] ,
    \cb_1_0_io_o_0_out[0] }),
    .io_o_1_out({\cb_1_0_io_o_1_out[7] ,
    \cb_1_0_io_o_1_out[6] ,
    \cb_1_0_io_o_1_out[5] ,
    \cb_1_0_io_o_1_out[4] ,
    \cb_1_0_io_o_1_out[3] ,
    \cb_1_0_io_o_1_out[2] ,
    \cb_1_0_io_o_1_out[1] ,
    \cb_1_0_io_o_1_out[0] }),
    .io_o_2_out({\cb_1_0_io_o_2_out[7] ,
    \cb_1_0_io_o_2_out[6] ,
    \cb_1_0_io_o_2_out[5] ,
    \cb_1_0_io_o_2_out[4] ,
    \cb_1_0_io_o_2_out[3] ,
    \cb_1_0_io_o_2_out[2] ,
    \cb_1_0_io_o_2_out[1] ,
    \cb_1_0_io_o_2_out[0] }),
    .io_o_3_out({\cb_1_0_io_o_3_out[7] ,
    \cb_1_0_io_o_3_out[6] ,
    \cb_1_0_io_o_3_out[5] ,
    \cb_1_0_io_o_3_out[4] ,
    \cb_1_0_io_o_3_out[3] ,
    \cb_1_0_io_o_3_out[2] ,
    \cb_1_0_io_o_3_out[1] ,
    \cb_1_0_io_o_3_out[0] }),
    .io_o_4_out({\cb_1_0_io_o_4_out[7] ,
    \cb_1_0_io_o_4_out[6] ,
    \cb_1_0_io_o_4_out[5] ,
    \cb_1_0_io_o_4_out[4] ,
    \cb_1_0_io_o_4_out[3] ,
    \cb_1_0_io_o_4_out[2] ,
    \cb_1_0_io_o_4_out[1] ,
    \cb_1_0_io_o_4_out[0] }),
    .io_o_5_out({\cb_1_0_io_o_5_out[7] ,
    \cb_1_0_io_o_5_out[6] ,
    \cb_1_0_io_o_5_out[5] ,
    \cb_1_0_io_o_5_out[4] ,
    \cb_1_0_io_o_5_out[3] ,
    \cb_1_0_io_o_5_out[2] ,
    \cb_1_0_io_o_5_out[1] ,
    \cb_1_0_io_o_5_out[0] }),
    .io_o_6_out({\cb_1_0_io_o_6_out[7] ,
    \cb_1_0_io_o_6_out[6] ,
    \cb_1_0_io_o_6_out[5] ,
    \cb_1_0_io_o_6_out[4] ,
    \cb_1_0_io_o_6_out[3] ,
    \cb_1_0_io_o_6_out[2] ,
    \cb_1_0_io_o_6_out[1] ,
    \cb_1_0_io_o_6_out[0] }),
    .io_o_7_out({\cb_1_0_io_o_7_out[7] ,
    \cb_1_0_io_o_7_out[6] ,
    \cb_1_0_io_o_7_out[5] ,
    \cb_1_0_io_o_7_out[4] ,
    \cb_1_0_io_o_7_out[3] ,
    \cb_1_0_io_o_7_out[2] ,
    \cb_1_0_io_o_7_out[1] ,
    \cb_1_0_io_o_7_out[0] }),
    .io_wo({\cb_1_0_io_wo[63] ,
    \cb_1_0_io_wo[62] ,
    \cb_1_0_io_wo[61] ,
    \cb_1_0_io_wo[60] ,
    \cb_1_0_io_wo[59] ,
    \cb_1_0_io_wo[58] ,
    \cb_1_0_io_wo[57] ,
    \cb_1_0_io_wo[56] ,
    \cb_1_0_io_wo[55] ,
    \cb_1_0_io_wo[54] ,
    \cb_1_0_io_wo[53] ,
    \cb_1_0_io_wo[52] ,
    \cb_1_0_io_wo[51] ,
    \cb_1_0_io_wo[50] ,
    \cb_1_0_io_wo[49] ,
    \cb_1_0_io_wo[48] ,
    \cb_1_0_io_wo[47] ,
    \cb_1_0_io_wo[46] ,
    \cb_1_0_io_wo[45] ,
    \cb_1_0_io_wo[44] ,
    \cb_1_0_io_wo[43] ,
    \cb_1_0_io_wo[42] ,
    \cb_1_0_io_wo[41] ,
    \cb_1_0_io_wo[40] ,
    \cb_1_0_io_wo[39] ,
    \cb_1_0_io_wo[38] ,
    \cb_1_0_io_wo[37] ,
    \cb_1_0_io_wo[36] ,
    \cb_1_0_io_wo[35] ,
    \cb_1_0_io_wo[34] ,
    \cb_1_0_io_wo[33] ,
    \cb_1_0_io_wo[32] ,
    \cb_1_0_io_wo[31] ,
    \cb_1_0_io_wo[30] ,
    \cb_1_0_io_wo[29] ,
    \cb_1_0_io_wo[28] ,
    \cb_1_0_io_wo[27] ,
    \cb_1_0_io_wo[26] ,
    \cb_1_0_io_wo[25] ,
    \cb_1_0_io_wo[24] ,
    \cb_1_0_io_wo[23] ,
    \cb_1_0_io_wo[22] ,
    \cb_1_0_io_wo[21] ,
    \cb_1_0_io_wo[20] ,
    \cb_1_0_io_wo[19] ,
    \cb_1_0_io_wo[18] ,
    \cb_1_0_io_wo[17] ,
    \cb_1_0_io_wo[16] ,
    \cb_1_0_io_wo[15] ,
    \cb_1_0_io_wo[14] ,
    \cb_1_0_io_wo[13] ,
    \cb_1_0_io_wo[12] ,
    \cb_1_0_io_wo[11] ,
    \cb_1_0_io_wo[10] ,
    \cb_1_0_io_wo[9] ,
    \cb_1_0_io_wo[8] ,
    \cb_1_0_io_wo[7] ,
    \cb_1_0_io_wo[6] ,
    \cb_1_0_io_wo[5] ,
    \cb_1_0_io_wo[4] ,
    \cb_1_0_io_wo[3] ,
    \cb_1_0_io_wo[2] ,
    \cb_1_0_io_wo[1] ,
    \cb_1_0_io_wo[0] }));
 cic_block cb_1_1 (.io_cs_i(cb_1_1_io_cs_i),
    .io_i_0_ci(cb_1_0_io_o_0_co),
    .io_i_1_ci(cb_1_0_io_o_1_co),
    .io_i_2_ci(cb_1_0_io_o_2_co),
    .io_i_3_ci(cb_1_0_io_o_3_co),
    .io_i_4_ci(cb_1_0_io_o_4_co),
    .io_i_5_ci(cb_1_0_io_o_5_co),
    .io_i_6_ci(cb_1_0_io_o_6_co),
    .io_i_7_ci(cb_1_0_io_o_7_co),
    .io_o_0_co(cb_1_1_io_o_0_co),
    .io_o_1_co(cb_1_1_io_o_1_co),
    .io_o_2_co(cb_1_1_io_o_2_co),
    .io_o_3_co(cb_1_1_io_o_3_co),
    .io_o_4_co(cb_1_1_io_o_4_co),
    .io_o_5_co(cb_1_1_io_o_5_co),
    .io_o_6_co(cb_1_1_io_o_6_co),
    .io_o_7_co(cb_1_1_io_o_7_co),
    .io_vci(cb_1_0_io_vco),
    .io_vco(cb_1_1_io_vco),
    .io_vi(cb_1_1_io_vi),
    .io_we_i(cb_1_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_1_0_io_adr_i[1] ,
    \cb_1_0_io_adr_i[0] }),
    .io_dat_i({\cb_1_0_io_dat_i[15] ,
    \cb_1_0_io_dat_i[14] ,
    \cb_1_0_io_dat_i[13] ,
    \cb_1_0_io_dat_i[12] ,
    \cb_1_0_io_dat_i[11] ,
    \cb_1_0_io_dat_i[10] ,
    \cb_1_0_io_dat_i[9] ,
    \cb_1_0_io_dat_i[8] ,
    \cb_1_0_io_dat_i[7] ,
    \cb_1_0_io_dat_i[6] ,
    \cb_1_0_io_dat_i[5] ,
    \cb_1_0_io_dat_i[4] ,
    \cb_1_0_io_dat_i[3] ,
    \cb_1_0_io_dat_i[2] ,
    \cb_1_0_io_dat_i[1] ,
    \cb_1_0_io_dat_i[0] }),
    .io_dat_o({\cb_1_1_io_dat_o[15] ,
    \cb_1_1_io_dat_o[14] ,
    \cb_1_1_io_dat_o[13] ,
    \cb_1_1_io_dat_o[12] ,
    \cb_1_1_io_dat_o[11] ,
    \cb_1_1_io_dat_o[10] ,
    \cb_1_1_io_dat_o[9] ,
    \cb_1_1_io_dat_o[8] ,
    \cb_1_1_io_dat_o[7] ,
    \cb_1_1_io_dat_o[6] ,
    \cb_1_1_io_dat_o[5] ,
    \cb_1_1_io_dat_o[4] ,
    \cb_1_1_io_dat_o[3] ,
    \cb_1_1_io_dat_o[2] ,
    \cb_1_1_io_dat_o[1] ,
    \cb_1_1_io_dat_o[0] }),
    .io_eo({\cb_1_1_io_eo[63] ,
    \cb_1_1_io_eo[62] ,
    \cb_1_1_io_eo[61] ,
    \cb_1_1_io_eo[60] ,
    \cb_1_1_io_eo[59] ,
    \cb_1_1_io_eo[58] ,
    \cb_1_1_io_eo[57] ,
    \cb_1_1_io_eo[56] ,
    \cb_1_1_io_eo[55] ,
    \cb_1_1_io_eo[54] ,
    \cb_1_1_io_eo[53] ,
    \cb_1_1_io_eo[52] ,
    \cb_1_1_io_eo[51] ,
    \cb_1_1_io_eo[50] ,
    \cb_1_1_io_eo[49] ,
    \cb_1_1_io_eo[48] ,
    \cb_1_1_io_eo[47] ,
    \cb_1_1_io_eo[46] ,
    \cb_1_1_io_eo[45] ,
    \cb_1_1_io_eo[44] ,
    \cb_1_1_io_eo[43] ,
    \cb_1_1_io_eo[42] ,
    \cb_1_1_io_eo[41] ,
    \cb_1_1_io_eo[40] ,
    \cb_1_1_io_eo[39] ,
    \cb_1_1_io_eo[38] ,
    \cb_1_1_io_eo[37] ,
    \cb_1_1_io_eo[36] ,
    \cb_1_1_io_eo[35] ,
    \cb_1_1_io_eo[34] ,
    \cb_1_1_io_eo[33] ,
    \cb_1_1_io_eo[32] ,
    \cb_1_1_io_eo[31] ,
    \cb_1_1_io_eo[30] ,
    \cb_1_1_io_eo[29] ,
    \cb_1_1_io_eo[28] ,
    \cb_1_1_io_eo[27] ,
    \cb_1_1_io_eo[26] ,
    \cb_1_1_io_eo[25] ,
    \cb_1_1_io_eo[24] ,
    \cb_1_1_io_eo[23] ,
    \cb_1_1_io_eo[22] ,
    \cb_1_1_io_eo[21] ,
    \cb_1_1_io_eo[20] ,
    \cb_1_1_io_eo[19] ,
    \cb_1_1_io_eo[18] ,
    \cb_1_1_io_eo[17] ,
    \cb_1_1_io_eo[16] ,
    \cb_1_1_io_eo[15] ,
    \cb_1_1_io_eo[14] ,
    \cb_1_1_io_eo[13] ,
    \cb_1_1_io_eo[12] ,
    \cb_1_1_io_eo[11] ,
    \cb_1_1_io_eo[10] ,
    \cb_1_1_io_eo[9] ,
    \cb_1_1_io_eo[8] ,
    \cb_1_1_io_eo[7] ,
    \cb_1_1_io_eo[6] ,
    \cb_1_1_io_eo[5] ,
    \cb_1_1_io_eo[4] ,
    \cb_1_1_io_eo[3] ,
    \cb_1_1_io_eo[2] ,
    \cb_1_1_io_eo[1] ,
    \cb_1_1_io_eo[0] }),
    .io_i_0_in1({\cb_1_0_io_o_0_out[7] ,
    \cb_1_0_io_o_0_out[6] ,
    \cb_1_0_io_o_0_out[5] ,
    \cb_1_0_io_o_0_out[4] ,
    \cb_1_0_io_o_0_out[3] ,
    \cb_1_0_io_o_0_out[2] ,
    \cb_1_0_io_o_0_out[1] ,
    \cb_1_0_io_o_0_out[0] }),
    .io_i_1_in1({\cb_1_0_io_o_1_out[7] ,
    \cb_1_0_io_o_1_out[6] ,
    \cb_1_0_io_o_1_out[5] ,
    \cb_1_0_io_o_1_out[4] ,
    \cb_1_0_io_o_1_out[3] ,
    \cb_1_0_io_o_1_out[2] ,
    \cb_1_0_io_o_1_out[1] ,
    \cb_1_0_io_o_1_out[0] }),
    .io_i_2_in1({\cb_1_0_io_o_2_out[7] ,
    \cb_1_0_io_o_2_out[6] ,
    \cb_1_0_io_o_2_out[5] ,
    \cb_1_0_io_o_2_out[4] ,
    \cb_1_0_io_o_2_out[3] ,
    \cb_1_0_io_o_2_out[2] ,
    \cb_1_0_io_o_2_out[1] ,
    \cb_1_0_io_o_2_out[0] }),
    .io_i_3_in1({\cb_1_0_io_o_3_out[7] ,
    \cb_1_0_io_o_3_out[6] ,
    \cb_1_0_io_o_3_out[5] ,
    \cb_1_0_io_o_3_out[4] ,
    \cb_1_0_io_o_3_out[3] ,
    \cb_1_0_io_o_3_out[2] ,
    \cb_1_0_io_o_3_out[1] ,
    \cb_1_0_io_o_3_out[0] }),
    .io_i_4_in1({\cb_1_0_io_o_4_out[7] ,
    \cb_1_0_io_o_4_out[6] ,
    \cb_1_0_io_o_4_out[5] ,
    \cb_1_0_io_o_4_out[4] ,
    \cb_1_0_io_o_4_out[3] ,
    \cb_1_0_io_o_4_out[2] ,
    \cb_1_0_io_o_4_out[1] ,
    \cb_1_0_io_o_4_out[0] }),
    .io_i_5_in1({\cb_1_0_io_o_5_out[7] ,
    \cb_1_0_io_o_5_out[6] ,
    \cb_1_0_io_o_5_out[5] ,
    \cb_1_0_io_o_5_out[4] ,
    \cb_1_0_io_o_5_out[3] ,
    \cb_1_0_io_o_5_out[2] ,
    \cb_1_0_io_o_5_out[1] ,
    \cb_1_0_io_o_5_out[0] }),
    .io_i_6_in1({\cb_1_0_io_o_6_out[7] ,
    \cb_1_0_io_o_6_out[6] ,
    \cb_1_0_io_o_6_out[5] ,
    \cb_1_0_io_o_6_out[4] ,
    \cb_1_0_io_o_6_out[3] ,
    \cb_1_0_io_o_6_out[2] ,
    \cb_1_0_io_o_6_out[1] ,
    \cb_1_0_io_o_6_out[0] }),
    .io_i_7_in1({\cb_1_0_io_o_7_out[7] ,
    \cb_1_0_io_o_7_out[6] ,
    \cb_1_0_io_o_7_out[5] ,
    \cb_1_0_io_o_7_out[4] ,
    \cb_1_0_io_o_7_out[3] ,
    \cb_1_0_io_o_7_out[2] ,
    \cb_1_0_io_o_7_out[1] ,
    \cb_1_0_io_o_7_out[0] }),
    .io_o_0_out({\cb_1_1_io_o_0_out[7] ,
    \cb_1_1_io_o_0_out[6] ,
    \cb_1_1_io_o_0_out[5] ,
    \cb_1_1_io_o_0_out[4] ,
    \cb_1_1_io_o_0_out[3] ,
    \cb_1_1_io_o_0_out[2] ,
    \cb_1_1_io_o_0_out[1] ,
    \cb_1_1_io_o_0_out[0] }),
    .io_o_1_out({\cb_1_1_io_o_1_out[7] ,
    \cb_1_1_io_o_1_out[6] ,
    \cb_1_1_io_o_1_out[5] ,
    \cb_1_1_io_o_1_out[4] ,
    \cb_1_1_io_o_1_out[3] ,
    \cb_1_1_io_o_1_out[2] ,
    \cb_1_1_io_o_1_out[1] ,
    \cb_1_1_io_o_1_out[0] }),
    .io_o_2_out({\cb_1_1_io_o_2_out[7] ,
    \cb_1_1_io_o_2_out[6] ,
    \cb_1_1_io_o_2_out[5] ,
    \cb_1_1_io_o_2_out[4] ,
    \cb_1_1_io_o_2_out[3] ,
    \cb_1_1_io_o_2_out[2] ,
    \cb_1_1_io_o_2_out[1] ,
    \cb_1_1_io_o_2_out[0] }),
    .io_o_3_out({\cb_1_1_io_o_3_out[7] ,
    \cb_1_1_io_o_3_out[6] ,
    \cb_1_1_io_o_3_out[5] ,
    \cb_1_1_io_o_3_out[4] ,
    \cb_1_1_io_o_3_out[3] ,
    \cb_1_1_io_o_3_out[2] ,
    \cb_1_1_io_o_3_out[1] ,
    \cb_1_1_io_o_3_out[0] }),
    .io_o_4_out({\cb_1_1_io_o_4_out[7] ,
    \cb_1_1_io_o_4_out[6] ,
    \cb_1_1_io_o_4_out[5] ,
    \cb_1_1_io_o_4_out[4] ,
    \cb_1_1_io_o_4_out[3] ,
    \cb_1_1_io_o_4_out[2] ,
    \cb_1_1_io_o_4_out[1] ,
    \cb_1_1_io_o_4_out[0] }),
    .io_o_5_out({\cb_1_1_io_o_5_out[7] ,
    \cb_1_1_io_o_5_out[6] ,
    \cb_1_1_io_o_5_out[5] ,
    \cb_1_1_io_o_5_out[4] ,
    \cb_1_1_io_o_5_out[3] ,
    \cb_1_1_io_o_5_out[2] ,
    \cb_1_1_io_o_5_out[1] ,
    \cb_1_1_io_o_5_out[0] }),
    .io_o_6_out({\cb_1_1_io_o_6_out[7] ,
    \cb_1_1_io_o_6_out[6] ,
    \cb_1_1_io_o_6_out[5] ,
    \cb_1_1_io_o_6_out[4] ,
    \cb_1_1_io_o_6_out[3] ,
    \cb_1_1_io_o_6_out[2] ,
    \cb_1_1_io_o_6_out[1] ,
    \cb_1_1_io_o_6_out[0] }),
    .io_o_7_out({\cb_1_1_io_o_7_out[7] ,
    \cb_1_1_io_o_7_out[6] ,
    \cb_1_1_io_o_7_out[5] ,
    \cb_1_1_io_o_7_out[4] ,
    \cb_1_1_io_o_7_out[3] ,
    \cb_1_1_io_o_7_out[2] ,
    \cb_1_1_io_o_7_out[1] ,
    \cb_1_1_io_o_7_out[0] }),
    .io_wo({\cb_1_0_io_eo[63] ,
    \cb_1_0_io_eo[62] ,
    \cb_1_0_io_eo[61] ,
    \cb_1_0_io_eo[60] ,
    \cb_1_0_io_eo[59] ,
    \cb_1_0_io_eo[58] ,
    \cb_1_0_io_eo[57] ,
    \cb_1_0_io_eo[56] ,
    \cb_1_0_io_eo[55] ,
    \cb_1_0_io_eo[54] ,
    \cb_1_0_io_eo[53] ,
    \cb_1_0_io_eo[52] ,
    \cb_1_0_io_eo[51] ,
    \cb_1_0_io_eo[50] ,
    \cb_1_0_io_eo[49] ,
    \cb_1_0_io_eo[48] ,
    \cb_1_0_io_eo[47] ,
    \cb_1_0_io_eo[46] ,
    \cb_1_0_io_eo[45] ,
    \cb_1_0_io_eo[44] ,
    \cb_1_0_io_eo[43] ,
    \cb_1_0_io_eo[42] ,
    \cb_1_0_io_eo[41] ,
    \cb_1_0_io_eo[40] ,
    \cb_1_0_io_eo[39] ,
    \cb_1_0_io_eo[38] ,
    \cb_1_0_io_eo[37] ,
    \cb_1_0_io_eo[36] ,
    \cb_1_0_io_eo[35] ,
    \cb_1_0_io_eo[34] ,
    \cb_1_0_io_eo[33] ,
    \cb_1_0_io_eo[32] ,
    \cb_1_0_io_eo[31] ,
    \cb_1_0_io_eo[30] ,
    \cb_1_0_io_eo[29] ,
    \cb_1_0_io_eo[28] ,
    \cb_1_0_io_eo[27] ,
    \cb_1_0_io_eo[26] ,
    \cb_1_0_io_eo[25] ,
    \cb_1_0_io_eo[24] ,
    \cb_1_0_io_eo[23] ,
    \cb_1_0_io_eo[22] ,
    \cb_1_0_io_eo[21] ,
    \cb_1_0_io_eo[20] ,
    \cb_1_0_io_eo[19] ,
    \cb_1_0_io_eo[18] ,
    \cb_1_0_io_eo[17] ,
    \cb_1_0_io_eo[16] ,
    \cb_1_0_io_eo[15] ,
    \cb_1_0_io_eo[14] ,
    \cb_1_0_io_eo[13] ,
    \cb_1_0_io_eo[12] ,
    \cb_1_0_io_eo[11] ,
    \cb_1_0_io_eo[10] ,
    \cb_1_0_io_eo[9] ,
    \cb_1_0_io_eo[8] ,
    \cb_1_0_io_eo[7] ,
    \cb_1_0_io_eo[6] ,
    \cb_1_0_io_eo[5] ,
    \cb_1_0_io_eo[4] ,
    \cb_1_0_io_eo[3] ,
    \cb_1_0_io_eo[2] ,
    \cb_1_0_io_eo[1] ,
    \cb_1_0_io_eo[0] }));
 cic_block cb_1_10 (.io_cs_i(cb_1_10_io_cs_i),
    .io_i_0_ci(cb_1_10_io_i_0_ci),
    .io_i_1_ci(cb_1_10_io_i_1_ci),
    .io_i_2_ci(cb_1_10_io_i_2_ci),
    .io_i_3_ci(cb_1_10_io_i_3_ci),
    .io_i_4_ci(cb_1_10_io_i_4_ci),
    .io_i_5_ci(cb_1_10_io_i_5_ci),
    .io_i_6_ci(cb_1_10_io_i_6_ci),
    .io_i_7_ci(cb_1_10_io_i_7_ci),
    .io_o_0_co(cb_1_10_io_o_0_co),
    .io_o_1_co(cb_1_10_io_o_1_co),
    .io_o_2_co(cb_1_10_io_o_2_co),
    .io_o_3_co(cb_1_10_io_o_3_co),
    .io_o_4_co(cb_1_10_io_o_4_co),
    .io_o_5_co(cb_1_10_io_o_5_co),
    .io_o_6_co(cb_1_10_io_o_6_co),
    .io_o_7_co(cb_1_10_io_o_7_co),
    .io_vci(cb_1_10_io_vci),
    .io_vco(cb_1_10_io_vco),
    .io_vi(cb_1_10_io_vi),
    .io_we_i(cb_1_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_1_0_io_adr_i[1] ,
    \cb_1_0_io_adr_i[0] }),
    .io_dat_i({\cb_1_0_io_dat_i[15] ,
    \cb_1_0_io_dat_i[14] ,
    \cb_1_0_io_dat_i[13] ,
    \cb_1_0_io_dat_i[12] ,
    \cb_1_0_io_dat_i[11] ,
    \cb_1_0_io_dat_i[10] ,
    \cb_1_0_io_dat_i[9] ,
    \cb_1_0_io_dat_i[8] ,
    \cb_1_0_io_dat_i[7] ,
    \cb_1_0_io_dat_i[6] ,
    \cb_1_0_io_dat_i[5] ,
    \cb_1_0_io_dat_i[4] ,
    \cb_1_0_io_dat_i[3] ,
    \cb_1_0_io_dat_i[2] ,
    \cb_1_0_io_dat_i[1] ,
    \cb_1_0_io_dat_i[0] }),
    .io_dat_o({\cb_1_10_io_dat_o[15] ,
    \cb_1_10_io_dat_o[14] ,
    \cb_1_10_io_dat_o[13] ,
    \cb_1_10_io_dat_o[12] ,
    \cb_1_10_io_dat_o[11] ,
    \cb_1_10_io_dat_o[10] ,
    \cb_1_10_io_dat_o[9] ,
    \cb_1_10_io_dat_o[8] ,
    \cb_1_10_io_dat_o[7] ,
    \cb_1_10_io_dat_o[6] ,
    \cb_1_10_io_dat_o[5] ,
    \cb_1_10_io_dat_o[4] ,
    \cb_1_10_io_dat_o[3] ,
    \cb_1_10_io_dat_o[2] ,
    \cb_1_10_io_dat_o[1] ,
    \cb_1_10_io_dat_o[0] }),
    .io_eo({\_T_47[31] ,
    \_T_47[30] ,
    \_T_47[29] ,
    \_T_47[28] ,
    \_T_47[27] ,
    \_T_47[26] ,
    \_T_47[25] ,
    \_T_47[24] ,
    \_T_47[23] ,
    \_T_47[22] ,
    \_T_47[21] ,
    \_T_47[20] ,
    \_T_47[19] ,
    \_T_47[18] ,
    \_T_47[17] ,
    \_T_47[16] ,
    \_T_47[15] ,
    \_T_47[14] ,
    \_T_47[13] ,
    \_T_47[12] ,
    \_T_47[11] ,
    \_T_47[10] ,
    \_T_47[9] ,
    \_T_47[8] ,
    \_T_47[7] ,
    \_T_47[6] ,
    \_T_47[5] ,
    \_T_47[4] ,
    \_T_47[3] ,
    \_T_47[2] ,
    \_T_47[1] ,
    \_T_47[0] ,
    \_T_44[31] ,
    \_T_44[30] ,
    \_T_44[29] ,
    \_T_44[28] ,
    \_T_44[27] ,
    \_T_44[26] ,
    \_T_44[25] ,
    \_T_44[24] ,
    \_T_44[23] ,
    \_T_44[22] ,
    \_T_44[21] ,
    \_T_44[20] ,
    \_T_44[19] ,
    \_T_44[18] ,
    \_T_44[17] ,
    \_T_44[16] ,
    \_T_44[15] ,
    \_T_44[14] ,
    \_T_44[13] ,
    \_T_44[12] ,
    \_T_44[11] ,
    \_T_44[10] ,
    \_T_44[9] ,
    \_T_44[8] ,
    \_T_44[7] ,
    \_T_44[6] ,
    \_T_44[5] ,
    \_T_44[4] ,
    \_T_44[3] ,
    \_T_44[2] ,
    \_T_44[1] ,
    \_T_44[0] }),
    .io_i_0_in1({\cb_1_10_io_i_0_in1[7] ,
    \cb_1_10_io_i_0_in1[6] ,
    \cb_1_10_io_i_0_in1[5] ,
    \cb_1_10_io_i_0_in1[4] ,
    \cb_1_10_io_i_0_in1[3] ,
    \cb_1_10_io_i_0_in1[2] ,
    \cb_1_10_io_i_0_in1[1] ,
    \cb_1_10_io_i_0_in1[0] }),
    .io_i_1_in1({\cb_1_10_io_i_1_in1[7] ,
    \cb_1_10_io_i_1_in1[6] ,
    \cb_1_10_io_i_1_in1[5] ,
    \cb_1_10_io_i_1_in1[4] ,
    \cb_1_10_io_i_1_in1[3] ,
    \cb_1_10_io_i_1_in1[2] ,
    \cb_1_10_io_i_1_in1[1] ,
    \cb_1_10_io_i_1_in1[0] }),
    .io_i_2_in1({\cb_1_10_io_i_2_in1[7] ,
    \cb_1_10_io_i_2_in1[6] ,
    \cb_1_10_io_i_2_in1[5] ,
    \cb_1_10_io_i_2_in1[4] ,
    \cb_1_10_io_i_2_in1[3] ,
    \cb_1_10_io_i_2_in1[2] ,
    \cb_1_10_io_i_2_in1[1] ,
    \cb_1_10_io_i_2_in1[0] }),
    .io_i_3_in1({\cb_1_10_io_i_3_in1[7] ,
    \cb_1_10_io_i_3_in1[6] ,
    \cb_1_10_io_i_3_in1[5] ,
    \cb_1_10_io_i_3_in1[4] ,
    \cb_1_10_io_i_3_in1[3] ,
    \cb_1_10_io_i_3_in1[2] ,
    \cb_1_10_io_i_3_in1[1] ,
    \cb_1_10_io_i_3_in1[0] }),
    .io_i_4_in1({\cb_1_10_io_i_4_in1[7] ,
    \cb_1_10_io_i_4_in1[6] ,
    \cb_1_10_io_i_4_in1[5] ,
    \cb_1_10_io_i_4_in1[4] ,
    \cb_1_10_io_i_4_in1[3] ,
    \cb_1_10_io_i_4_in1[2] ,
    \cb_1_10_io_i_4_in1[1] ,
    \cb_1_10_io_i_4_in1[0] }),
    .io_i_5_in1({\cb_1_10_io_i_5_in1[7] ,
    \cb_1_10_io_i_5_in1[6] ,
    \cb_1_10_io_i_5_in1[5] ,
    \cb_1_10_io_i_5_in1[4] ,
    \cb_1_10_io_i_5_in1[3] ,
    \cb_1_10_io_i_5_in1[2] ,
    \cb_1_10_io_i_5_in1[1] ,
    \cb_1_10_io_i_5_in1[0] }),
    .io_i_6_in1({\cb_1_10_io_i_6_in1[7] ,
    \cb_1_10_io_i_6_in1[6] ,
    \cb_1_10_io_i_6_in1[5] ,
    \cb_1_10_io_i_6_in1[4] ,
    \cb_1_10_io_i_6_in1[3] ,
    \cb_1_10_io_i_6_in1[2] ,
    \cb_1_10_io_i_6_in1[1] ,
    \cb_1_10_io_i_6_in1[0] }),
    .io_i_7_in1({\cb_1_10_io_i_7_in1[7] ,
    \cb_1_10_io_i_7_in1[6] ,
    \cb_1_10_io_i_7_in1[5] ,
    \cb_1_10_io_i_7_in1[4] ,
    \cb_1_10_io_i_7_in1[3] ,
    \cb_1_10_io_i_7_in1[2] ,
    \cb_1_10_io_i_7_in1[1] ,
    \cb_1_10_io_i_7_in1[0] }),
    .io_o_0_out({\_T_44[7] ,
    \_T_44[6] ,
    \_T_44[5] ,
    \_T_44[4] ,
    \_T_44[3] ,
    \_T_44[2] ,
    \_T_44[1] ,
    \_T_44[0] }),
    .io_o_1_out({\_T_44[15] ,
    \_T_44[14] ,
    \_T_44[13] ,
    \_T_44[12] ,
    \_T_44[11] ,
    \_T_44[10] ,
    \_T_44[9] ,
    \_T_44[8] }),
    .io_o_2_out({\_T_44[23] ,
    \_T_44[22] ,
    \_T_44[21] ,
    \_T_44[20] ,
    \_T_44[19] ,
    \_T_44[18] ,
    \_T_44[17] ,
    \_T_44[16] }),
    .io_o_3_out({\_T_44[31] ,
    \_T_44[30] ,
    \_T_44[29] ,
    \_T_44[28] ,
    \_T_44[27] ,
    \_T_44[26] ,
    \_T_44[25] ,
    \_T_44[24] }),
    .io_o_4_out({\_T_47[7] ,
    \_T_47[6] ,
    \_T_47[5] ,
    \_T_47[4] ,
    \_T_47[3] ,
    \_T_47[2] ,
    \_T_47[1] ,
    \_T_47[0] }),
    .io_o_5_out({\_T_47[15] ,
    \_T_47[14] ,
    \_T_47[13] ,
    \_T_47[12] ,
    \_T_47[11] ,
    \_T_47[10] ,
    \_T_47[9] ,
    \_T_47[8] }),
    .io_o_6_out({\_T_47[23] ,
    \_T_47[22] ,
    \_T_47[21] ,
    \_T_47[20] ,
    \_T_47[19] ,
    \_T_47[18] ,
    \_T_47[17] ,
    \_T_47[16] }),
    .io_o_7_out({\_T_47[31] ,
    \_T_47[30] ,
    \_T_47[29] ,
    \_T_47[28] ,
    \_T_47[27] ,
    \_T_47[26] ,
    \_T_47[25] ,
    \_T_47[24] }),
    .io_wo({\cb_1_10_io_wo[63] ,
    \cb_1_10_io_wo[62] ,
    \cb_1_10_io_wo[61] ,
    \cb_1_10_io_wo[60] ,
    \cb_1_10_io_wo[59] ,
    \cb_1_10_io_wo[58] ,
    \cb_1_10_io_wo[57] ,
    \cb_1_10_io_wo[56] ,
    \cb_1_10_io_wo[55] ,
    \cb_1_10_io_wo[54] ,
    \cb_1_10_io_wo[53] ,
    \cb_1_10_io_wo[52] ,
    \cb_1_10_io_wo[51] ,
    \cb_1_10_io_wo[50] ,
    \cb_1_10_io_wo[49] ,
    \cb_1_10_io_wo[48] ,
    \cb_1_10_io_wo[47] ,
    \cb_1_10_io_wo[46] ,
    \cb_1_10_io_wo[45] ,
    \cb_1_10_io_wo[44] ,
    \cb_1_10_io_wo[43] ,
    \cb_1_10_io_wo[42] ,
    \cb_1_10_io_wo[41] ,
    \cb_1_10_io_wo[40] ,
    \cb_1_10_io_wo[39] ,
    \cb_1_10_io_wo[38] ,
    \cb_1_10_io_wo[37] ,
    \cb_1_10_io_wo[36] ,
    \cb_1_10_io_wo[35] ,
    \cb_1_10_io_wo[34] ,
    \cb_1_10_io_wo[33] ,
    \cb_1_10_io_wo[32] ,
    \cb_1_10_io_wo[31] ,
    \cb_1_10_io_wo[30] ,
    \cb_1_10_io_wo[29] ,
    \cb_1_10_io_wo[28] ,
    \cb_1_10_io_wo[27] ,
    \cb_1_10_io_wo[26] ,
    \cb_1_10_io_wo[25] ,
    \cb_1_10_io_wo[24] ,
    \cb_1_10_io_wo[23] ,
    \cb_1_10_io_wo[22] ,
    \cb_1_10_io_wo[21] ,
    \cb_1_10_io_wo[20] ,
    \cb_1_10_io_wo[19] ,
    \cb_1_10_io_wo[18] ,
    \cb_1_10_io_wo[17] ,
    \cb_1_10_io_wo[16] ,
    \cb_1_10_io_wo[15] ,
    \cb_1_10_io_wo[14] ,
    \cb_1_10_io_wo[13] ,
    \cb_1_10_io_wo[12] ,
    \cb_1_10_io_wo[11] ,
    \cb_1_10_io_wo[10] ,
    \cb_1_10_io_wo[9] ,
    \cb_1_10_io_wo[8] ,
    \cb_1_10_io_wo[7] ,
    \cb_1_10_io_wo[6] ,
    \cb_1_10_io_wo[5] ,
    \cb_1_10_io_wo[4] ,
    \cb_1_10_io_wo[3] ,
    \cb_1_10_io_wo[2] ,
    \cb_1_10_io_wo[1] ,
    \cb_1_10_io_wo[0] }));
 cic_block cb_1_2 (.io_cs_i(cb_1_2_io_cs_i),
    .io_i_0_ci(cb_1_1_io_o_0_co),
    .io_i_1_ci(cb_1_1_io_o_1_co),
    .io_i_2_ci(cb_1_1_io_o_2_co),
    .io_i_3_ci(cb_1_1_io_o_3_co),
    .io_i_4_ci(cb_1_1_io_o_4_co),
    .io_i_5_ci(cb_1_1_io_o_5_co),
    .io_i_6_ci(cb_1_1_io_o_6_co),
    .io_i_7_ci(cb_1_1_io_o_7_co),
    .io_o_0_co(cb_1_2_io_o_0_co),
    .io_o_1_co(cb_1_2_io_o_1_co),
    .io_o_2_co(cb_1_2_io_o_2_co),
    .io_o_3_co(cb_1_2_io_o_3_co),
    .io_o_4_co(cb_1_2_io_o_4_co),
    .io_o_5_co(cb_1_2_io_o_5_co),
    .io_o_6_co(cb_1_2_io_o_6_co),
    .io_o_7_co(cb_1_2_io_o_7_co),
    .io_vci(cb_1_1_io_vco),
    .io_vco(cb_1_2_io_vco),
    .io_vi(cb_1_2_io_vi),
    .io_we_i(cb_1_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_1_0_io_adr_i[1] ,
    \cb_1_0_io_adr_i[0] }),
    .io_dat_i({\cb_1_0_io_dat_i[15] ,
    \cb_1_0_io_dat_i[14] ,
    \cb_1_0_io_dat_i[13] ,
    \cb_1_0_io_dat_i[12] ,
    \cb_1_0_io_dat_i[11] ,
    \cb_1_0_io_dat_i[10] ,
    \cb_1_0_io_dat_i[9] ,
    \cb_1_0_io_dat_i[8] ,
    \cb_1_0_io_dat_i[7] ,
    \cb_1_0_io_dat_i[6] ,
    \cb_1_0_io_dat_i[5] ,
    \cb_1_0_io_dat_i[4] ,
    \cb_1_0_io_dat_i[3] ,
    \cb_1_0_io_dat_i[2] ,
    \cb_1_0_io_dat_i[1] ,
    \cb_1_0_io_dat_i[0] }),
    .io_dat_o({\cb_1_2_io_dat_o[15] ,
    \cb_1_2_io_dat_o[14] ,
    \cb_1_2_io_dat_o[13] ,
    \cb_1_2_io_dat_o[12] ,
    \cb_1_2_io_dat_o[11] ,
    \cb_1_2_io_dat_o[10] ,
    \cb_1_2_io_dat_o[9] ,
    \cb_1_2_io_dat_o[8] ,
    \cb_1_2_io_dat_o[7] ,
    \cb_1_2_io_dat_o[6] ,
    \cb_1_2_io_dat_o[5] ,
    \cb_1_2_io_dat_o[4] ,
    \cb_1_2_io_dat_o[3] ,
    \cb_1_2_io_dat_o[2] ,
    \cb_1_2_io_dat_o[1] ,
    \cb_1_2_io_dat_o[0] }),
    .io_eo({\cb_1_2_io_eo[63] ,
    \cb_1_2_io_eo[62] ,
    \cb_1_2_io_eo[61] ,
    \cb_1_2_io_eo[60] ,
    \cb_1_2_io_eo[59] ,
    \cb_1_2_io_eo[58] ,
    \cb_1_2_io_eo[57] ,
    \cb_1_2_io_eo[56] ,
    \cb_1_2_io_eo[55] ,
    \cb_1_2_io_eo[54] ,
    \cb_1_2_io_eo[53] ,
    \cb_1_2_io_eo[52] ,
    \cb_1_2_io_eo[51] ,
    \cb_1_2_io_eo[50] ,
    \cb_1_2_io_eo[49] ,
    \cb_1_2_io_eo[48] ,
    \cb_1_2_io_eo[47] ,
    \cb_1_2_io_eo[46] ,
    \cb_1_2_io_eo[45] ,
    \cb_1_2_io_eo[44] ,
    \cb_1_2_io_eo[43] ,
    \cb_1_2_io_eo[42] ,
    \cb_1_2_io_eo[41] ,
    \cb_1_2_io_eo[40] ,
    \cb_1_2_io_eo[39] ,
    \cb_1_2_io_eo[38] ,
    \cb_1_2_io_eo[37] ,
    \cb_1_2_io_eo[36] ,
    \cb_1_2_io_eo[35] ,
    \cb_1_2_io_eo[34] ,
    \cb_1_2_io_eo[33] ,
    \cb_1_2_io_eo[32] ,
    \cb_1_2_io_eo[31] ,
    \cb_1_2_io_eo[30] ,
    \cb_1_2_io_eo[29] ,
    \cb_1_2_io_eo[28] ,
    \cb_1_2_io_eo[27] ,
    \cb_1_2_io_eo[26] ,
    \cb_1_2_io_eo[25] ,
    \cb_1_2_io_eo[24] ,
    \cb_1_2_io_eo[23] ,
    \cb_1_2_io_eo[22] ,
    \cb_1_2_io_eo[21] ,
    \cb_1_2_io_eo[20] ,
    \cb_1_2_io_eo[19] ,
    \cb_1_2_io_eo[18] ,
    \cb_1_2_io_eo[17] ,
    \cb_1_2_io_eo[16] ,
    \cb_1_2_io_eo[15] ,
    \cb_1_2_io_eo[14] ,
    \cb_1_2_io_eo[13] ,
    \cb_1_2_io_eo[12] ,
    \cb_1_2_io_eo[11] ,
    \cb_1_2_io_eo[10] ,
    \cb_1_2_io_eo[9] ,
    \cb_1_2_io_eo[8] ,
    \cb_1_2_io_eo[7] ,
    \cb_1_2_io_eo[6] ,
    \cb_1_2_io_eo[5] ,
    \cb_1_2_io_eo[4] ,
    \cb_1_2_io_eo[3] ,
    \cb_1_2_io_eo[2] ,
    \cb_1_2_io_eo[1] ,
    \cb_1_2_io_eo[0] }),
    .io_i_0_in1({\cb_1_1_io_o_0_out[7] ,
    \cb_1_1_io_o_0_out[6] ,
    \cb_1_1_io_o_0_out[5] ,
    \cb_1_1_io_o_0_out[4] ,
    \cb_1_1_io_o_0_out[3] ,
    \cb_1_1_io_o_0_out[2] ,
    \cb_1_1_io_o_0_out[1] ,
    \cb_1_1_io_o_0_out[0] }),
    .io_i_1_in1({\cb_1_1_io_o_1_out[7] ,
    \cb_1_1_io_o_1_out[6] ,
    \cb_1_1_io_o_1_out[5] ,
    \cb_1_1_io_o_1_out[4] ,
    \cb_1_1_io_o_1_out[3] ,
    \cb_1_1_io_o_1_out[2] ,
    \cb_1_1_io_o_1_out[1] ,
    \cb_1_1_io_o_1_out[0] }),
    .io_i_2_in1({\cb_1_1_io_o_2_out[7] ,
    \cb_1_1_io_o_2_out[6] ,
    \cb_1_1_io_o_2_out[5] ,
    \cb_1_1_io_o_2_out[4] ,
    \cb_1_1_io_o_2_out[3] ,
    \cb_1_1_io_o_2_out[2] ,
    \cb_1_1_io_o_2_out[1] ,
    \cb_1_1_io_o_2_out[0] }),
    .io_i_3_in1({\cb_1_1_io_o_3_out[7] ,
    \cb_1_1_io_o_3_out[6] ,
    \cb_1_1_io_o_3_out[5] ,
    \cb_1_1_io_o_3_out[4] ,
    \cb_1_1_io_o_3_out[3] ,
    \cb_1_1_io_o_3_out[2] ,
    \cb_1_1_io_o_3_out[1] ,
    \cb_1_1_io_o_3_out[0] }),
    .io_i_4_in1({\cb_1_1_io_o_4_out[7] ,
    \cb_1_1_io_o_4_out[6] ,
    \cb_1_1_io_o_4_out[5] ,
    \cb_1_1_io_o_4_out[4] ,
    \cb_1_1_io_o_4_out[3] ,
    \cb_1_1_io_o_4_out[2] ,
    \cb_1_1_io_o_4_out[1] ,
    \cb_1_1_io_o_4_out[0] }),
    .io_i_5_in1({\cb_1_1_io_o_5_out[7] ,
    \cb_1_1_io_o_5_out[6] ,
    \cb_1_1_io_o_5_out[5] ,
    \cb_1_1_io_o_5_out[4] ,
    \cb_1_1_io_o_5_out[3] ,
    \cb_1_1_io_o_5_out[2] ,
    \cb_1_1_io_o_5_out[1] ,
    \cb_1_1_io_o_5_out[0] }),
    .io_i_6_in1({\cb_1_1_io_o_6_out[7] ,
    \cb_1_1_io_o_6_out[6] ,
    \cb_1_1_io_o_6_out[5] ,
    \cb_1_1_io_o_6_out[4] ,
    \cb_1_1_io_o_6_out[3] ,
    \cb_1_1_io_o_6_out[2] ,
    \cb_1_1_io_o_6_out[1] ,
    \cb_1_1_io_o_6_out[0] }),
    .io_i_7_in1({\cb_1_1_io_o_7_out[7] ,
    \cb_1_1_io_o_7_out[6] ,
    \cb_1_1_io_o_7_out[5] ,
    \cb_1_1_io_o_7_out[4] ,
    \cb_1_1_io_o_7_out[3] ,
    \cb_1_1_io_o_7_out[2] ,
    \cb_1_1_io_o_7_out[1] ,
    \cb_1_1_io_o_7_out[0] }),
    .io_o_0_out({\cb_1_2_io_o_0_out[7] ,
    \cb_1_2_io_o_0_out[6] ,
    \cb_1_2_io_o_0_out[5] ,
    \cb_1_2_io_o_0_out[4] ,
    \cb_1_2_io_o_0_out[3] ,
    \cb_1_2_io_o_0_out[2] ,
    \cb_1_2_io_o_0_out[1] ,
    \cb_1_2_io_o_0_out[0] }),
    .io_o_1_out({\cb_1_2_io_o_1_out[7] ,
    \cb_1_2_io_o_1_out[6] ,
    \cb_1_2_io_o_1_out[5] ,
    \cb_1_2_io_o_1_out[4] ,
    \cb_1_2_io_o_1_out[3] ,
    \cb_1_2_io_o_1_out[2] ,
    \cb_1_2_io_o_1_out[1] ,
    \cb_1_2_io_o_1_out[0] }),
    .io_o_2_out({\cb_1_2_io_o_2_out[7] ,
    \cb_1_2_io_o_2_out[6] ,
    \cb_1_2_io_o_2_out[5] ,
    \cb_1_2_io_o_2_out[4] ,
    \cb_1_2_io_o_2_out[3] ,
    \cb_1_2_io_o_2_out[2] ,
    \cb_1_2_io_o_2_out[1] ,
    \cb_1_2_io_o_2_out[0] }),
    .io_o_3_out({\cb_1_2_io_o_3_out[7] ,
    \cb_1_2_io_o_3_out[6] ,
    \cb_1_2_io_o_3_out[5] ,
    \cb_1_2_io_o_3_out[4] ,
    \cb_1_2_io_o_3_out[3] ,
    \cb_1_2_io_o_3_out[2] ,
    \cb_1_2_io_o_3_out[1] ,
    \cb_1_2_io_o_3_out[0] }),
    .io_o_4_out({\cb_1_2_io_o_4_out[7] ,
    \cb_1_2_io_o_4_out[6] ,
    \cb_1_2_io_o_4_out[5] ,
    \cb_1_2_io_o_4_out[4] ,
    \cb_1_2_io_o_4_out[3] ,
    \cb_1_2_io_o_4_out[2] ,
    \cb_1_2_io_o_4_out[1] ,
    \cb_1_2_io_o_4_out[0] }),
    .io_o_5_out({\cb_1_2_io_o_5_out[7] ,
    \cb_1_2_io_o_5_out[6] ,
    \cb_1_2_io_o_5_out[5] ,
    \cb_1_2_io_o_5_out[4] ,
    \cb_1_2_io_o_5_out[3] ,
    \cb_1_2_io_o_5_out[2] ,
    \cb_1_2_io_o_5_out[1] ,
    \cb_1_2_io_o_5_out[0] }),
    .io_o_6_out({\cb_1_2_io_o_6_out[7] ,
    \cb_1_2_io_o_6_out[6] ,
    \cb_1_2_io_o_6_out[5] ,
    \cb_1_2_io_o_6_out[4] ,
    \cb_1_2_io_o_6_out[3] ,
    \cb_1_2_io_o_6_out[2] ,
    \cb_1_2_io_o_6_out[1] ,
    \cb_1_2_io_o_6_out[0] }),
    .io_o_7_out({\cb_1_2_io_o_7_out[7] ,
    \cb_1_2_io_o_7_out[6] ,
    \cb_1_2_io_o_7_out[5] ,
    \cb_1_2_io_o_7_out[4] ,
    \cb_1_2_io_o_7_out[3] ,
    \cb_1_2_io_o_7_out[2] ,
    \cb_1_2_io_o_7_out[1] ,
    \cb_1_2_io_o_7_out[0] }),
    .io_wo({\cb_1_1_io_eo[63] ,
    \cb_1_1_io_eo[62] ,
    \cb_1_1_io_eo[61] ,
    \cb_1_1_io_eo[60] ,
    \cb_1_1_io_eo[59] ,
    \cb_1_1_io_eo[58] ,
    \cb_1_1_io_eo[57] ,
    \cb_1_1_io_eo[56] ,
    \cb_1_1_io_eo[55] ,
    \cb_1_1_io_eo[54] ,
    \cb_1_1_io_eo[53] ,
    \cb_1_1_io_eo[52] ,
    \cb_1_1_io_eo[51] ,
    \cb_1_1_io_eo[50] ,
    \cb_1_1_io_eo[49] ,
    \cb_1_1_io_eo[48] ,
    \cb_1_1_io_eo[47] ,
    \cb_1_1_io_eo[46] ,
    \cb_1_1_io_eo[45] ,
    \cb_1_1_io_eo[44] ,
    \cb_1_1_io_eo[43] ,
    \cb_1_1_io_eo[42] ,
    \cb_1_1_io_eo[41] ,
    \cb_1_1_io_eo[40] ,
    \cb_1_1_io_eo[39] ,
    \cb_1_1_io_eo[38] ,
    \cb_1_1_io_eo[37] ,
    \cb_1_1_io_eo[36] ,
    \cb_1_1_io_eo[35] ,
    \cb_1_1_io_eo[34] ,
    \cb_1_1_io_eo[33] ,
    \cb_1_1_io_eo[32] ,
    \cb_1_1_io_eo[31] ,
    \cb_1_1_io_eo[30] ,
    \cb_1_1_io_eo[29] ,
    \cb_1_1_io_eo[28] ,
    \cb_1_1_io_eo[27] ,
    \cb_1_1_io_eo[26] ,
    \cb_1_1_io_eo[25] ,
    \cb_1_1_io_eo[24] ,
    \cb_1_1_io_eo[23] ,
    \cb_1_1_io_eo[22] ,
    \cb_1_1_io_eo[21] ,
    \cb_1_1_io_eo[20] ,
    \cb_1_1_io_eo[19] ,
    \cb_1_1_io_eo[18] ,
    \cb_1_1_io_eo[17] ,
    \cb_1_1_io_eo[16] ,
    \cb_1_1_io_eo[15] ,
    \cb_1_1_io_eo[14] ,
    \cb_1_1_io_eo[13] ,
    \cb_1_1_io_eo[12] ,
    \cb_1_1_io_eo[11] ,
    \cb_1_1_io_eo[10] ,
    \cb_1_1_io_eo[9] ,
    \cb_1_1_io_eo[8] ,
    \cb_1_1_io_eo[7] ,
    \cb_1_1_io_eo[6] ,
    \cb_1_1_io_eo[5] ,
    \cb_1_1_io_eo[4] ,
    \cb_1_1_io_eo[3] ,
    \cb_1_1_io_eo[2] ,
    \cb_1_1_io_eo[1] ,
    \cb_1_1_io_eo[0] }));
 cic_block cb_1_3 (.io_cs_i(cb_1_3_io_cs_i),
    .io_i_0_ci(cb_1_2_io_o_0_co),
    .io_i_1_ci(cb_1_2_io_o_1_co),
    .io_i_2_ci(cb_1_2_io_o_2_co),
    .io_i_3_ci(cb_1_2_io_o_3_co),
    .io_i_4_ci(cb_1_2_io_o_4_co),
    .io_i_5_ci(cb_1_2_io_o_5_co),
    .io_i_6_ci(cb_1_2_io_o_6_co),
    .io_i_7_ci(cb_1_2_io_o_7_co),
    .io_o_0_co(cb_1_3_io_o_0_co),
    .io_o_1_co(cb_1_3_io_o_1_co),
    .io_o_2_co(cb_1_3_io_o_2_co),
    .io_o_3_co(cb_1_3_io_o_3_co),
    .io_o_4_co(cb_1_3_io_o_4_co),
    .io_o_5_co(cb_1_3_io_o_5_co),
    .io_o_6_co(cb_1_3_io_o_6_co),
    .io_o_7_co(cb_1_3_io_o_7_co),
    .io_vci(cb_1_2_io_vco),
    .io_vco(cb_1_3_io_vco),
    .io_vi(cb_1_3_io_vi),
    .io_we_i(cb_1_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_1_0_io_adr_i[1] ,
    \cb_1_0_io_adr_i[0] }),
    .io_dat_i({\cb_1_0_io_dat_i[15] ,
    \cb_1_0_io_dat_i[14] ,
    \cb_1_0_io_dat_i[13] ,
    \cb_1_0_io_dat_i[12] ,
    \cb_1_0_io_dat_i[11] ,
    \cb_1_0_io_dat_i[10] ,
    \cb_1_0_io_dat_i[9] ,
    \cb_1_0_io_dat_i[8] ,
    \cb_1_0_io_dat_i[7] ,
    \cb_1_0_io_dat_i[6] ,
    \cb_1_0_io_dat_i[5] ,
    \cb_1_0_io_dat_i[4] ,
    \cb_1_0_io_dat_i[3] ,
    \cb_1_0_io_dat_i[2] ,
    \cb_1_0_io_dat_i[1] ,
    \cb_1_0_io_dat_i[0] }),
    .io_dat_o({\cb_1_3_io_dat_o[15] ,
    \cb_1_3_io_dat_o[14] ,
    \cb_1_3_io_dat_o[13] ,
    \cb_1_3_io_dat_o[12] ,
    \cb_1_3_io_dat_o[11] ,
    \cb_1_3_io_dat_o[10] ,
    \cb_1_3_io_dat_o[9] ,
    \cb_1_3_io_dat_o[8] ,
    \cb_1_3_io_dat_o[7] ,
    \cb_1_3_io_dat_o[6] ,
    \cb_1_3_io_dat_o[5] ,
    \cb_1_3_io_dat_o[4] ,
    \cb_1_3_io_dat_o[3] ,
    \cb_1_3_io_dat_o[2] ,
    \cb_1_3_io_dat_o[1] ,
    \cb_1_3_io_dat_o[0] }),
    .io_eo({\cb_1_3_io_eo[63] ,
    \cb_1_3_io_eo[62] ,
    \cb_1_3_io_eo[61] ,
    \cb_1_3_io_eo[60] ,
    \cb_1_3_io_eo[59] ,
    \cb_1_3_io_eo[58] ,
    \cb_1_3_io_eo[57] ,
    \cb_1_3_io_eo[56] ,
    \cb_1_3_io_eo[55] ,
    \cb_1_3_io_eo[54] ,
    \cb_1_3_io_eo[53] ,
    \cb_1_3_io_eo[52] ,
    \cb_1_3_io_eo[51] ,
    \cb_1_3_io_eo[50] ,
    \cb_1_3_io_eo[49] ,
    \cb_1_3_io_eo[48] ,
    \cb_1_3_io_eo[47] ,
    \cb_1_3_io_eo[46] ,
    \cb_1_3_io_eo[45] ,
    \cb_1_3_io_eo[44] ,
    \cb_1_3_io_eo[43] ,
    \cb_1_3_io_eo[42] ,
    \cb_1_3_io_eo[41] ,
    \cb_1_3_io_eo[40] ,
    \cb_1_3_io_eo[39] ,
    \cb_1_3_io_eo[38] ,
    \cb_1_3_io_eo[37] ,
    \cb_1_3_io_eo[36] ,
    \cb_1_3_io_eo[35] ,
    \cb_1_3_io_eo[34] ,
    \cb_1_3_io_eo[33] ,
    \cb_1_3_io_eo[32] ,
    \cb_1_3_io_eo[31] ,
    \cb_1_3_io_eo[30] ,
    \cb_1_3_io_eo[29] ,
    \cb_1_3_io_eo[28] ,
    \cb_1_3_io_eo[27] ,
    \cb_1_3_io_eo[26] ,
    \cb_1_3_io_eo[25] ,
    \cb_1_3_io_eo[24] ,
    \cb_1_3_io_eo[23] ,
    \cb_1_3_io_eo[22] ,
    \cb_1_3_io_eo[21] ,
    \cb_1_3_io_eo[20] ,
    \cb_1_3_io_eo[19] ,
    \cb_1_3_io_eo[18] ,
    \cb_1_3_io_eo[17] ,
    \cb_1_3_io_eo[16] ,
    \cb_1_3_io_eo[15] ,
    \cb_1_3_io_eo[14] ,
    \cb_1_3_io_eo[13] ,
    \cb_1_3_io_eo[12] ,
    \cb_1_3_io_eo[11] ,
    \cb_1_3_io_eo[10] ,
    \cb_1_3_io_eo[9] ,
    \cb_1_3_io_eo[8] ,
    \cb_1_3_io_eo[7] ,
    \cb_1_3_io_eo[6] ,
    \cb_1_3_io_eo[5] ,
    \cb_1_3_io_eo[4] ,
    \cb_1_3_io_eo[3] ,
    \cb_1_3_io_eo[2] ,
    \cb_1_3_io_eo[1] ,
    \cb_1_3_io_eo[0] }),
    .io_i_0_in1({\cb_1_2_io_o_0_out[7] ,
    \cb_1_2_io_o_0_out[6] ,
    \cb_1_2_io_o_0_out[5] ,
    \cb_1_2_io_o_0_out[4] ,
    \cb_1_2_io_o_0_out[3] ,
    \cb_1_2_io_o_0_out[2] ,
    \cb_1_2_io_o_0_out[1] ,
    \cb_1_2_io_o_0_out[0] }),
    .io_i_1_in1({\cb_1_2_io_o_1_out[7] ,
    \cb_1_2_io_o_1_out[6] ,
    \cb_1_2_io_o_1_out[5] ,
    \cb_1_2_io_o_1_out[4] ,
    \cb_1_2_io_o_1_out[3] ,
    \cb_1_2_io_o_1_out[2] ,
    \cb_1_2_io_o_1_out[1] ,
    \cb_1_2_io_o_1_out[0] }),
    .io_i_2_in1({\cb_1_2_io_o_2_out[7] ,
    \cb_1_2_io_o_2_out[6] ,
    \cb_1_2_io_o_2_out[5] ,
    \cb_1_2_io_o_2_out[4] ,
    \cb_1_2_io_o_2_out[3] ,
    \cb_1_2_io_o_2_out[2] ,
    \cb_1_2_io_o_2_out[1] ,
    \cb_1_2_io_o_2_out[0] }),
    .io_i_3_in1({\cb_1_2_io_o_3_out[7] ,
    \cb_1_2_io_o_3_out[6] ,
    \cb_1_2_io_o_3_out[5] ,
    \cb_1_2_io_o_3_out[4] ,
    \cb_1_2_io_o_3_out[3] ,
    \cb_1_2_io_o_3_out[2] ,
    \cb_1_2_io_o_3_out[1] ,
    \cb_1_2_io_o_3_out[0] }),
    .io_i_4_in1({\cb_1_2_io_o_4_out[7] ,
    \cb_1_2_io_o_4_out[6] ,
    \cb_1_2_io_o_4_out[5] ,
    \cb_1_2_io_o_4_out[4] ,
    \cb_1_2_io_o_4_out[3] ,
    \cb_1_2_io_o_4_out[2] ,
    \cb_1_2_io_o_4_out[1] ,
    \cb_1_2_io_o_4_out[0] }),
    .io_i_5_in1({\cb_1_2_io_o_5_out[7] ,
    \cb_1_2_io_o_5_out[6] ,
    \cb_1_2_io_o_5_out[5] ,
    \cb_1_2_io_o_5_out[4] ,
    \cb_1_2_io_o_5_out[3] ,
    \cb_1_2_io_o_5_out[2] ,
    \cb_1_2_io_o_5_out[1] ,
    \cb_1_2_io_o_5_out[0] }),
    .io_i_6_in1({\cb_1_2_io_o_6_out[7] ,
    \cb_1_2_io_o_6_out[6] ,
    \cb_1_2_io_o_6_out[5] ,
    \cb_1_2_io_o_6_out[4] ,
    \cb_1_2_io_o_6_out[3] ,
    \cb_1_2_io_o_6_out[2] ,
    \cb_1_2_io_o_6_out[1] ,
    \cb_1_2_io_o_6_out[0] }),
    .io_i_7_in1({\cb_1_2_io_o_7_out[7] ,
    \cb_1_2_io_o_7_out[6] ,
    \cb_1_2_io_o_7_out[5] ,
    \cb_1_2_io_o_7_out[4] ,
    \cb_1_2_io_o_7_out[3] ,
    \cb_1_2_io_o_7_out[2] ,
    \cb_1_2_io_o_7_out[1] ,
    \cb_1_2_io_o_7_out[0] }),
    .io_o_0_out({\cb_1_3_io_o_0_out[7] ,
    \cb_1_3_io_o_0_out[6] ,
    \cb_1_3_io_o_0_out[5] ,
    \cb_1_3_io_o_0_out[4] ,
    \cb_1_3_io_o_0_out[3] ,
    \cb_1_3_io_o_0_out[2] ,
    \cb_1_3_io_o_0_out[1] ,
    \cb_1_3_io_o_0_out[0] }),
    .io_o_1_out({\cb_1_3_io_o_1_out[7] ,
    \cb_1_3_io_o_1_out[6] ,
    \cb_1_3_io_o_1_out[5] ,
    \cb_1_3_io_o_1_out[4] ,
    \cb_1_3_io_o_1_out[3] ,
    \cb_1_3_io_o_1_out[2] ,
    \cb_1_3_io_o_1_out[1] ,
    \cb_1_3_io_o_1_out[0] }),
    .io_o_2_out({\cb_1_3_io_o_2_out[7] ,
    \cb_1_3_io_o_2_out[6] ,
    \cb_1_3_io_o_2_out[5] ,
    \cb_1_3_io_o_2_out[4] ,
    \cb_1_3_io_o_2_out[3] ,
    \cb_1_3_io_o_2_out[2] ,
    \cb_1_3_io_o_2_out[1] ,
    \cb_1_3_io_o_2_out[0] }),
    .io_o_3_out({\cb_1_3_io_o_3_out[7] ,
    \cb_1_3_io_o_3_out[6] ,
    \cb_1_3_io_o_3_out[5] ,
    \cb_1_3_io_o_3_out[4] ,
    \cb_1_3_io_o_3_out[3] ,
    \cb_1_3_io_o_3_out[2] ,
    \cb_1_3_io_o_3_out[1] ,
    \cb_1_3_io_o_3_out[0] }),
    .io_o_4_out({\cb_1_3_io_o_4_out[7] ,
    \cb_1_3_io_o_4_out[6] ,
    \cb_1_3_io_o_4_out[5] ,
    \cb_1_3_io_o_4_out[4] ,
    \cb_1_3_io_o_4_out[3] ,
    \cb_1_3_io_o_4_out[2] ,
    \cb_1_3_io_o_4_out[1] ,
    \cb_1_3_io_o_4_out[0] }),
    .io_o_5_out({\cb_1_3_io_o_5_out[7] ,
    \cb_1_3_io_o_5_out[6] ,
    \cb_1_3_io_o_5_out[5] ,
    \cb_1_3_io_o_5_out[4] ,
    \cb_1_3_io_o_5_out[3] ,
    \cb_1_3_io_o_5_out[2] ,
    \cb_1_3_io_o_5_out[1] ,
    \cb_1_3_io_o_5_out[0] }),
    .io_o_6_out({\cb_1_3_io_o_6_out[7] ,
    \cb_1_3_io_o_6_out[6] ,
    \cb_1_3_io_o_6_out[5] ,
    \cb_1_3_io_o_6_out[4] ,
    \cb_1_3_io_o_6_out[3] ,
    \cb_1_3_io_o_6_out[2] ,
    \cb_1_3_io_o_6_out[1] ,
    \cb_1_3_io_o_6_out[0] }),
    .io_o_7_out({\cb_1_3_io_o_7_out[7] ,
    \cb_1_3_io_o_7_out[6] ,
    \cb_1_3_io_o_7_out[5] ,
    \cb_1_3_io_o_7_out[4] ,
    \cb_1_3_io_o_7_out[3] ,
    \cb_1_3_io_o_7_out[2] ,
    \cb_1_3_io_o_7_out[1] ,
    \cb_1_3_io_o_7_out[0] }),
    .io_wo({\cb_1_2_io_eo[63] ,
    \cb_1_2_io_eo[62] ,
    \cb_1_2_io_eo[61] ,
    \cb_1_2_io_eo[60] ,
    \cb_1_2_io_eo[59] ,
    \cb_1_2_io_eo[58] ,
    \cb_1_2_io_eo[57] ,
    \cb_1_2_io_eo[56] ,
    \cb_1_2_io_eo[55] ,
    \cb_1_2_io_eo[54] ,
    \cb_1_2_io_eo[53] ,
    \cb_1_2_io_eo[52] ,
    \cb_1_2_io_eo[51] ,
    \cb_1_2_io_eo[50] ,
    \cb_1_2_io_eo[49] ,
    \cb_1_2_io_eo[48] ,
    \cb_1_2_io_eo[47] ,
    \cb_1_2_io_eo[46] ,
    \cb_1_2_io_eo[45] ,
    \cb_1_2_io_eo[44] ,
    \cb_1_2_io_eo[43] ,
    \cb_1_2_io_eo[42] ,
    \cb_1_2_io_eo[41] ,
    \cb_1_2_io_eo[40] ,
    \cb_1_2_io_eo[39] ,
    \cb_1_2_io_eo[38] ,
    \cb_1_2_io_eo[37] ,
    \cb_1_2_io_eo[36] ,
    \cb_1_2_io_eo[35] ,
    \cb_1_2_io_eo[34] ,
    \cb_1_2_io_eo[33] ,
    \cb_1_2_io_eo[32] ,
    \cb_1_2_io_eo[31] ,
    \cb_1_2_io_eo[30] ,
    \cb_1_2_io_eo[29] ,
    \cb_1_2_io_eo[28] ,
    \cb_1_2_io_eo[27] ,
    \cb_1_2_io_eo[26] ,
    \cb_1_2_io_eo[25] ,
    \cb_1_2_io_eo[24] ,
    \cb_1_2_io_eo[23] ,
    \cb_1_2_io_eo[22] ,
    \cb_1_2_io_eo[21] ,
    \cb_1_2_io_eo[20] ,
    \cb_1_2_io_eo[19] ,
    \cb_1_2_io_eo[18] ,
    \cb_1_2_io_eo[17] ,
    \cb_1_2_io_eo[16] ,
    \cb_1_2_io_eo[15] ,
    \cb_1_2_io_eo[14] ,
    \cb_1_2_io_eo[13] ,
    \cb_1_2_io_eo[12] ,
    \cb_1_2_io_eo[11] ,
    \cb_1_2_io_eo[10] ,
    \cb_1_2_io_eo[9] ,
    \cb_1_2_io_eo[8] ,
    \cb_1_2_io_eo[7] ,
    \cb_1_2_io_eo[6] ,
    \cb_1_2_io_eo[5] ,
    \cb_1_2_io_eo[4] ,
    \cb_1_2_io_eo[3] ,
    \cb_1_2_io_eo[2] ,
    \cb_1_2_io_eo[1] ,
    \cb_1_2_io_eo[0] }));
 cic_block cb_1_4 (.io_cs_i(cb_1_4_io_cs_i),
    .io_i_0_ci(cb_1_3_io_o_0_co),
    .io_i_1_ci(cb_1_3_io_o_1_co),
    .io_i_2_ci(cb_1_3_io_o_2_co),
    .io_i_3_ci(cb_1_3_io_o_3_co),
    .io_i_4_ci(cb_1_3_io_o_4_co),
    .io_i_5_ci(cb_1_3_io_o_5_co),
    .io_i_6_ci(cb_1_3_io_o_6_co),
    .io_i_7_ci(cb_1_3_io_o_7_co),
    .io_o_0_co(cb_1_4_io_o_0_co),
    .io_o_1_co(cb_1_4_io_o_1_co),
    .io_o_2_co(cb_1_4_io_o_2_co),
    .io_o_3_co(cb_1_4_io_o_3_co),
    .io_o_4_co(cb_1_4_io_o_4_co),
    .io_o_5_co(cb_1_4_io_o_5_co),
    .io_o_6_co(cb_1_4_io_o_6_co),
    .io_o_7_co(cb_1_4_io_o_7_co),
    .io_vci(cb_1_3_io_vco),
    .io_vco(cb_1_4_io_vco),
    .io_vi(cb_1_4_io_vi),
    .io_we_i(cb_1_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_1_0_io_adr_i[1] ,
    \cb_1_0_io_adr_i[0] }),
    .io_dat_i({\cb_1_0_io_dat_i[15] ,
    \cb_1_0_io_dat_i[14] ,
    \cb_1_0_io_dat_i[13] ,
    \cb_1_0_io_dat_i[12] ,
    \cb_1_0_io_dat_i[11] ,
    \cb_1_0_io_dat_i[10] ,
    \cb_1_0_io_dat_i[9] ,
    \cb_1_0_io_dat_i[8] ,
    \cb_1_0_io_dat_i[7] ,
    \cb_1_0_io_dat_i[6] ,
    \cb_1_0_io_dat_i[5] ,
    \cb_1_0_io_dat_i[4] ,
    \cb_1_0_io_dat_i[3] ,
    \cb_1_0_io_dat_i[2] ,
    \cb_1_0_io_dat_i[1] ,
    \cb_1_0_io_dat_i[0] }),
    .io_dat_o({\cb_1_4_io_dat_o[15] ,
    \cb_1_4_io_dat_o[14] ,
    \cb_1_4_io_dat_o[13] ,
    \cb_1_4_io_dat_o[12] ,
    \cb_1_4_io_dat_o[11] ,
    \cb_1_4_io_dat_o[10] ,
    \cb_1_4_io_dat_o[9] ,
    \cb_1_4_io_dat_o[8] ,
    \cb_1_4_io_dat_o[7] ,
    \cb_1_4_io_dat_o[6] ,
    \cb_1_4_io_dat_o[5] ,
    \cb_1_4_io_dat_o[4] ,
    \cb_1_4_io_dat_o[3] ,
    \cb_1_4_io_dat_o[2] ,
    \cb_1_4_io_dat_o[1] ,
    \cb_1_4_io_dat_o[0] }),
    .io_eo({\cb_1_4_io_eo[63] ,
    \cb_1_4_io_eo[62] ,
    \cb_1_4_io_eo[61] ,
    \cb_1_4_io_eo[60] ,
    \cb_1_4_io_eo[59] ,
    \cb_1_4_io_eo[58] ,
    \cb_1_4_io_eo[57] ,
    \cb_1_4_io_eo[56] ,
    \cb_1_4_io_eo[55] ,
    \cb_1_4_io_eo[54] ,
    \cb_1_4_io_eo[53] ,
    \cb_1_4_io_eo[52] ,
    \cb_1_4_io_eo[51] ,
    \cb_1_4_io_eo[50] ,
    \cb_1_4_io_eo[49] ,
    \cb_1_4_io_eo[48] ,
    \cb_1_4_io_eo[47] ,
    \cb_1_4_io_eo[46] ,
    \cb_1_4_io_eo[45] ,
    \cb_1_4_io_eo[44] ,
    \cb_1_4_io_eo[43] ,
    \cb_1_4_io_eo[42] ,
    \cb_1_4_io_eo[41] ,
    \cb_1_4_io_eo[40] ,
    \cb_1_4_io_eo[39] ,
    \cb_1_4_io_eo[38] ,
    \cb_1_4_io_eo[37] ,
    \cb_1_4_io_eo[36] ,
    \cb_1_4_io_eo[35] ,
    \cb_1_4_io_eo[34] ,
    \cb_1_4_io_eo[33] ,
    \cb_1_4_io_eo[32] ,
    \cb_1_4_io_eo[31] ,
    \cb_1_4_io_eo[30] ,
    \cb_1_4_io_eo[29] ,
    \cb_1_4_io_eo[28] ,
    \cb_1_4_io_eo[27] ,
    \cb_1_4_io_eo[26] ,
    \cb_1_4_io_eo[25] ,
    \cb_1_4_io_eo[24] ,
    \cb_1_4_io_eo[23] ,
    \cb_1_4_io_eo[22] ,
    \cb_1_4_io_eo[21] ,
    \cb_1_4_io_eo[20] ,
    \cb_1_4_io_eo[19] ,
    \cb_1_4_io_eo[18] ,
    \cb_1_4_io_eo[17] ,
    \cb_1_4_io_eo[16] ,
    \cb_1_4_io_eo[15] ,
    \cb_1_4_io_eo[14] ,
    \cb_1_4_io_eo[13] ,
    \cb_1_4_io_eo[12] ,
    \cb_1_4_io_eo[11] ,
    \cb_1_4_io_eo[10] ,
    \cb_1_4_io_eo[9] ,
    \cb_1_4_io_eo[8] ,
    \cb_1_4_io_eo[7] ,
    \cb_1_4_io_eo[6] ,
    \cb_1_4_io_eo[5] ,
    \cb_1_4_io_eo[4] ,
    \cb_1_4_io_eo[3] ,
    \cb_1_4_io_eo[2] ,
    \cb_1_4_io_eo[1] ,
    \cb_1_4_io_eo[0] }),
    .io_i_0_in1({\cb_1_3_io_o_0_out[7] ,
    \cb_1_3_io_o_0_out[6] ,
    \cb_1_3_io_o_0_out[5] ,
    \cb_1_3_io_o_0_out[4] ,
    \cb_1_3_io_o_0_out[3] ,
    \cb_1_3_io_o_0_out[2] ,
    \cb_1_3_io_o_0_out[1] ,
    \cb_1_3_io_o_0_out[0] }),
    .io_i_1_in1({\cb_1_3_io_o_1_out[7] ,
    \cb_1_3_io_o_1_out[6] ,
    \cb_1_3_io_o_1_out[5] ,
    \cb_1_3_io_o_1_out[4] ,
    \cb_1_3_io_o_1_out[3] ,
    \cb_1_3_io_o_1_out[2] ,
    \cb_1_3_io_o_1_out[1] ,
    \cb_1_3_io_o_1_out[0] }),
    .io_i_2_in1({\cb_1_3_io_o_2_out[7] ,
    \cb_1_3_io_o_2_out[6] ,
    \cb_1_3_io_o_2_out[5] ,
    \cb_1_3_io_o_2_out[4] ,
    \cb_1_3_io_o_2_out[3] ,
    \cb_1_3_io_o_2_out[2] ,
    \cb_1_3_io_o_2_out[1] ,
    \cb_1_3_io_o_2_out[0] }),
    .io_i_3_in1({\cb_1_3_io_o_3_out[7] ,
    \cb_1_3_io_o_3_out[6] ,
    \cb_1_3_io_o_3_out[5] ,
    \cb_1_3_io_o_3_out[4] ,
    \cb_1_3_io_o_3_out[3] ,
    \cb_1_3_io_o_3_out[2] ,
    \cb_1_3_io_o_3_out[1] ,
    \cb_1_3_io_o_3_out[0] }),
    .io_i_4_in1({\cb_1_3_io_o_4_out[7] ,
    \cb_1_3_io_o_4_out[6] ,
    \cb_1_3_io_o_4_out[5] ,
    \cb_1_3_io_o_4_out[4] ,
    \cb_1_3_io_o_4_out[3] ,
    \cb_1_3_io_o_4_out[2] ,
    \cb_1_3_io_o_4_out[1] ,
    \cb_1_3_io_o_4_out[0] }),
    .io_i_5_in1({\cb_1_3_io_o_5_out[7] ,
    \cb_1_3_io_o_5_out[6] ,
    \cb_1_3_io_o_5_out[5] ,
    \cb_1_3_io_o_5_out[4] ,
    \cb_1_3_io_o_5_out[3] ,
    \cb_1_3_io_o_5_out[2] ,
    \cb_1_3_io_o_5_out[1] ,
    \cb_1_3_io_o_5_out[0] }),
    .io_i_6_in1({\cb_1_3_io_o_6_out[7] ,
    \cb_1_3_io_o_6_out[6] ,
    \cb_1_3_io_o_6_out[5] ,
    \cb_1_3_io_o_6_out[4] ,
    \cb_1_3_io_o_6_out[3] ,
    \cb_1_3_io_o_6_out[2] ,
    \cb_1_3_io_o_6_out[1] ,
    \cb_1_3_io_o_6_out[0] }),
    .io_i_7_in1({\cb_1_3_io_o_7_out[7] ,
    \cb_1_3_io_o_7_out[6] ,
    \cb_1_3_io_o_7_out[5] ,
    \cb_1_3_io_o_7_out[4] ,
    \cb_1_3_io_o_7_out[3] ,
    \cb_1_3_io_o_7_out[2] ,
    \cb_1_3_io_o_7_out[1] ,
    \cb_1_3_io_o_7_out[0] }),
    .io_o_0_out({\cb_1_4_io_o_0_out[7] ,
    \cb_1_4_io_o_0_out[6] ,
    \cb_1_4_io_o_0_out[5] ,
    \cb_1_4_io_o_0_out[4] ,
    \cb_1_4_io_o_0_out[3] ,
    \cb_1_4_io_o_0_out[2] ,
    \cb_1_4_io_o_0_out[1] ,
    \cb_1_4_io_o_0_out[0] }),
    .io_o_1_out({\cb_1_4_io_o_1_out[7] ,
    \cb_1_4_io_o_1_out[6] ,
    \cb_1_4_io_o_1_out[5] ,
    \cb_1_4_io_o_1_out[4] ,
    \cb_1_4_io_o_1_out[3] ,
    \cb_1_4_io_o_1_out[2] ,
    \cb_1_4_io_o_1_out[1] ,
    \cb_1_4_io_o_1_out[0] }),
    .io_o_2_out({\cb_1_4_io_o_2_out[7] ,
    \cb_1_4_io_o_2_out[6] ,
    \cb_1_4_io_o_2_out[5] ,
    \cb_1_4_io_o_2_out[4] ,
    \cb_1_4_io_o_2_out[3] ,
    \cb_1_4_io_o_2_out[2] ,
    \cb_1_4_io_o_2_out[1] ,
    \cb_1_4_io_o_2_out[0] }),
    .io_o_3_out({\cb_1_4_io_o_3_out[7] ,
    \cb_1_4_io_o_3_out[6] ,
    \cb_1_4_io_o_3_out[5] ,
    \cb_1_4_io_o_3_out[4] ,
    \cb_1_4_io_o_3_out[3] ,
    \cb_1_4_io_o_3_out[2] ,
    \cb_1_4_io_o_3_out[1] ,
    \cb_1_4_io_o_3_out[0] }),
    .io_o_4_out({\cb_1_4_io_o_4_out[7] ,
    \cb_1_4_io_o_4_out[6] ,
    \cb_1_4_io_o_4_out[5] ,
    \cb_1_4_io_o_4_out[4] ,
    \cb_1_4_io_o_4_out[3] ,
    \cb_1_4_io_o_4_out[2] ,
    \cb_1_4_io_o_4_out[1] ,
    \cb_1_4_io_o_4_out[0] }),
    .io_o_5_out({\cb_1_4_io_o_5_out[7] ,
    \cb_1_4_io_o_5_out[6] ,
    \cb_1_4_io_o_5_out[5] ,
    \cb_1_4_io_o_5_out[4] ,
    \cb_1_4_io_o_5_out[3] ,
    \cb_1_4_io_o_5_out[2] ,
    \cb_1_4_io_o_5_out[1] ,
    \cb_1_4_io_o_5_out[0] }),
    .io_o_6_out({\cb_1_4_io_o_6_out[7] ,
    \cb_1_4_io_o_6_out[6] ,
    \cb_1_4_io_o_6_out[5] ,
    \cb_1_4_io_o_6_out[4] ,
    \cb_1_4_io_o_6_out[3] ,
    \cb_1_4_io_o_6_out[2] ,
    \cb_1_4_io_o_6_out[1] ,
    \cb_1_4_io_o_6_out[0] }),
    .io_o_7_out({\cb_1_4_io_o_7_out[7] ,
    \cb_1_4_io_o_7_out[6] ,
    \cb_1_4_io_o_7_out[5] ,
    \cb_1_4_io_o_7_out[4] ,
    \cb_1_4_io_o_7_out[3] ,
    \cb_1_4_io_o_7_out[2] ,
    \cb_1_4_io_o_7_out[1] ,
    \cb_1_4_io_o_7_out[0] }),
    .io_wo({\cb_1_3_io_eo[63] ,
    \cb_1_3_io_eo[62] ,
    \cb_1_3_io_eo[61] ,
    \cb_1_3_io_eo[60] ,
    \cb_1_3_io_eo[59] ,
    \cb_1_3_io_eo[58] ,
    \cb_1_3_io_eo[57] ,
    \cb_1_3_io_eo[56] ,
    \cb_1_3_io_eo[55] ,
    \cb_1_3_io_eo[54] ,
    \cb_1_3_io_eo[53] ,
    \cb_1_3_io_eo[52] ,
    \cb_1_3_io_eo[51] ,
    \cb_1_3_io_eo[50] ,
    \cb_1_3_io_eo[49] ,
    \cb_1_3_io_eo[48] ,
    \cb_1_3_io_eo[47] ,
    \cb_1_3_io_eo[46] ,
    \cb_1_3_io_eo[45] ,
    \cb_1_3_io_eo[44] ,
    \cb_1_3_io_eo[43] ,
    \cb_1_3_io_eo[42] ,
    \cb_1_3_io_eo[41] ,
    \cb_1_3_io_eo[40] ,
    \cb_1_3_io_eo[39] ,
    \cb_1_3_io_eo[38] ,
    \cb_1_3_io_eo[37] ,
    \cb_1_3_io_eo[36] ,
    \cb_1_3_io_eo[35] ,
    \cb_1_3_io_eo[34] ,
    \cb_1_3_io_eo[33] ,
    \cb_1_3_io_eo[32] ,
    \cb_1_3_io_eo[31] ,
    \cb_1_3_io_eo[30] ,
    \cb_1_3_io_eo[29] ,
    \cb_1_3_io_eo[28] ,
    \cb_1_3_io_eo[27] ,
    \cb_1_3_io_eo[26] ,
    \cb_1_3_io_eo[25] ,
    \cb_1_3_io_eo[24] ,
    \cb_1_3_io_eo[23] ,
    \cb_1_3_io_eo[22] ,
    \cb_1_3_io_eo[21] ,
    \cb_1_3_io_eo[20] ,
    \cb_1_3_io_eo[19] ,
    \cb_1_3_io_eo[18] ,
    \cb_1_3_io_eo[17] ,
    \cb_1_3_io_eo[16] ,
    \cb_1_3_io_eo[15] ,
    \cb_1_3_io_eo[14] ,
    \cb_1_3_io_eo[13] ,
    \cb_1_3_io_eo[12] ,
    \cb_1_3_io_eo[11] ,
    \cb_1_3_io_eo[10] ,
    \cb_1_3_io_eo[9] ,
    \cb_1_3_io_eo[8] ,
    \cb_1_3_io_eo[7] ,
    \cb_1_3_io_eo[6] ,
    \cb_1_3_io_eo[5] ,
    \cb_1_3_io_eo[4] ,
    \cb_1_3_io_eo[3] ,
    \cb_1_3_io_eo[2] ,
    \cb_1_3_io_eo[1] ,
    \cb_1_3_io_eo[0] }));
 cic_block cb_1_5 (.io_cs_i(cb_1_5_io_cs_i),
    .io_i_0_ci(cb_1_4_io_o_0_co),
    .io_i_1_ci(cb_1_4_io_o_1_co),
    .io_i_2_ci(cb_1_4_io_o_2_co),
    .io_i_3_ci(cb_1_4_io_o_3_co),
    .io_i_4_ci(cb_1_4_io_o_4_co),
    .io_i_5_ci(cb_1_4_io_o_5_co),
    .io_i_6_ci(cb_1_4_io_o_6_co),
    .io_i_7_ci(cb_1_4_io_o_7_co),
    .io_o_0_co(cb_1_5_io_o_0_co),
    .io_o_1_co(cb_1_5_io_o_1_co),
    .io_o_2_co(cb_1_5_io_o_2_co),
    .io_o_3_co(cb_1_5_io_o_3_co),
    .io_o_4_co(cb_1_5_io_o_4_co),
    .io_o_5_co(cb_1_5_io_o_5_co),
    .io_o_6_co(cb_1_5_io_o_6_co),
    .io_o_7_co(cb_1_5_io_o_7_co),
    .io_vci(cb_1_4_io_vco),
    .io_vco(cb_1_5_io_vco),
    .io_vi(cb_1_5_io_vi),
    .io_we_i(cb_1_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_1_0_io_adr_i[1] ,
    \cb_1_0_io_adr_i[0] }),
    .io_dat_i({\cb_1_0_io_dat_i[15] ,
    \cb_1_0_io_dat_i[14] ,
    \cb_1_0_io_dat_i[13] ,
    \cb_1_0_io_dat_i[12] ,
    \cb_1_0_io_dat_i[11] ,
    \cb_1_0_io_dat_i[10] ,
    \cb_1_0_io_dat_i[9] ,
    \cb_1_0_io_dat_i[8] ,
    \cb_1_0_io_dat_i[7] ,
    \cb_1_0_io_dat_i[6] ,
    \cb_1_0_io_dat_i[5] ,
    \cb_1_0_io_dat_i[4] ,
    \cb_1_0_io_dat_i[3] ,
    \cb_1_0_io_dat_i[2] ,
    \cb_1_0_io_dat_i[1] ,
    \cb_1_0_io_dat_i[0] }),
    .io_dat_o({\cb_1_5_io_dat_o[15] ,
    \cb_1_5_io_dat_o[14] ,
    \cb_1_5_io_dat_o[13] ,
    \cb_1_5_io_dat_o[12] ,
    \cb_1_5_io_dat_o[11] ,
    \cb_1_5_io_dat_o[10] ,
    \cb_1_5_io_dat_o[9] ,
    \cb_1_5_io_dat_o[8] ,
    \cb_1_5_io_dat_o[7] ,
    \cb_1_5_io_dat_o[6] ,
    \cb_1_5_io_dat_o[5] ,
    \cb_1_5_io_dat_o[4] ,
    \cb_1_5_io_dat_o[3] ,
    \cb_1_5_io_dat_o[2] ,
    \cb_1_5_io_dat_o[1] ,
    \cb_1_5_io_dat_o[0] }),
    .io_eo({\cb_1_5_io_eo[63] ,
    \cb_1_5_io_eo[62] ,
    \cb_1_5_io_eo[61] ,
    \cb_1_5_io_eo[60] ,
    \cb_1_5_io_eo[59] ,
    \cb_1_5_io_eo[58] ,
    \cb_1_5_io_eo[57] ,
    \cb_1_5_io_eo[56] ,
    \cb_1_5_io_eo[55] ,
    \cb_1_5_io_eo[54] ,
    \cb_1_5_io_eo[53] ,
    \cb_1_5_io_eo[52] ,
    \cb_1_5_io_eo[51] ,
    \cb_1_5_io_eo[50] ,
    \cb_1_5_io_eo[49] ,
    \cb_1_5_io_eo[48] ,
    \cb_1_5_io_eo[47] ,
    \cb_1_5_io_eo[46] ,
    \cb_1_5_io_eo[45] ,
    \cb_1_5_io_eo[44] ,
    \cb_1_5_io_eo[43] ,
    \cb_1_5_io_eo[42] ,
    \cb_1_5_io_eo[41] ,
    \cb_1_5_io_eo[40] ,
    \cb_1_5_io_eo[39] ,
    \cb_1_5_io_eo[38] ,
    \cb_1_5_io_eo[37] ,
    \cb_1_5_io_eo[36] ,
    \cb_1_5_io_eo[35] ,
    \cb_1_5_io_eo[34] ,
    \cb_1_5_io_eo[33] ,
    \cb_1_5_io_eo[32] ,
    \cb_1_5_io_eo[31] ,
    \cb_1_5_io_eo[30] ,
    \cb_1_5_io_eo[29] ,
    \cb_1_5_io_eo[28] ,
    \cb_1_5_io_eo[27] ,
    \cb_1_5_io_eo[26] ,
    \cb_1_5_io_eo[25] ,
    \cb_1_5_io_eo[24] ,
    \cb_1_5_io_eo[23] ,
    \cb_1_5_io_eo[22] ,
    \cb_1_5_io_eo[21] ,
    \cb_1_5_io_eo[20] ,
    \cb_1_5_io_eo[19] ,
    \cb_1_5_io_eo[18] ,
    \cb_1_5_io_eo[17] ,
    \cb_1_5_io_eo[16] ,
    \cb_1_5_io_eo[15] ,
    \cb_1_5_io_eo[14] ,
    \cb_1_5_io_eo[13] ,
    \cb_1_5_io_eo[12] ,
    \cb_1_5_io_eo[11] ,
    \cb_1_5_io_eo[10] ,
    \cb_1_5_io_eo[9] ,
    \cb_1_5_io_eo[8] ,
    \cb_1_5_io_eo[7] ,
    \cb_1_5_io_eo[6] ,
    \cb_1_5_io_eo[5] ,
    \cb_1_5_io_eo[4] ,
    \cb_1_5_io_eo[3] ,
    \cb_1_5_io_eo[2] ,
    \cb_1_5_io_eo[1] ,
    \cb_1_5_io_eo[0] }),
    .io_i_0_in1({\cb_1_4_io_o_0_out[7] ,
    \cb_1_4_io_o_0_out[6] ,
    \cb_1_4_io_o_0_out[5] ,
    \cb_1_4_io_o_0_out[4] ,
    \cb_1_4_io_o_0_out[3] ,
    \cb_1_4_io_o_0_out[2] ,
    \cb_1_4_io_o_0_out[1] ,
    \cb_1_4_io_o_0_out[0] }),
    .io_i_1_in1({\cb_1_4_io_o_1_out[7] ,
    \cb_1_4_io_o_1_out[6] ,
    \cb_1_4_io_o_1_out[5] ,
    \cb_1_4_io_o_1_out[4] ,
    \cb_1_4_io_o_1_out[3] ,
    \cb_1_4_io_o_1_out[2] ,
    \cb_1_4_io_o_1_out[1] ,
    \cb_1_4_io_o_1_out[0] }),
    .io_i_2_in1({\cb_1_4_io_o_2_out[7] ,
    \cb_1_4_io_o_2_out[6] ,
    \cb_1_4_io_o_2_out[5] ,
    \cb_1_4_io_o_2_out[4] ,
    \cb_1_4_io_o_2_out[3] ,
    \cb_1_4_io_o_2_out[2] ,
    \cb_1_4_io_o_2_out[1] ,
    \cb_1_4_io_o_2_out[0] }),
    .io_i_3_in1({\cb_1_4_io_o_3_out[7] ,
    \cb_1_4_io_o_3_out[6] ,
    \cb_1_4_io_o_3_out[5] ,
    \cb_1_4_io_o_3_out[4] ,
    \cb_1_4_io_o_3_out[3] ,
    \cb_1_4_io_o_3_out[2] ,
    \cb_1_4_io_o_3_out[1] ,
    \cb_1_4_io_o_3_out[0] }),
    .io_i_4_in1({\cb_1_4_io_o_4_out[7] ,
    \cb_1_4_io_o_4_out[6] ,
    \cb_1_4_io_o_4_out[5] ,
    \cb_1_4_io_o_4_out[4] ,
    \cb_1_4_io_o_4_out[3] ,
    \cb_1_4_io_o_4_out[2] ,
    \cb_1_4_io_o_4_out[1] ,
    \cb_1_4_io_o_4_out[0] }),
    .io_i_5_in1({\cb_1_4_io_o_5_out[7] ,
    \cb_1_4_io_o_5_out[6] ,
    \cb_1_4_io_o_5_out[5] ,
    \cb_1_4_io_o_5_out[4] ,
    \cb_1_4_io_o_5_out[3] ,
    \cb_1_4_io_o_5_out[2] ,
    \cb_1_4_io_o_5_out[1] ,
    \cb_1_4_io_o_5_out[0] }),
    .io_i_6_in1({\cb_1_4_io_o_6_out[7] ,
    \cb_1_4_io_o_6_out[6] ,
    \cb_1_4_io_o_6_out[5] ,
    \cb_1_4_io_o_6_out[4] ,
    \cb_1_4_io_o_6_out[3] ,
    \cb_1_4_io_o_6_out[2] ,
    \cb_1_4_io_o_6_out[1] ,
    \cb_1_4_io_o_6_out[0] }),
    .io_i_7_in1({\cb_1_4_io_o_7_out[7] ,
    \cb_1_4_io_o_7_out[6] ,
    \cb_1_4_io_o_7_out[5] ,
    \cb_1_4_io_o_7_out[4] ,
    \cb_1_4_io_o_7_out[3] ,
    \cb_1_4_io_o_7_out[2] ,
    \cb_1_4_io_o_7_out[1] ,
    \cb_1_4_io_o_7_out[0] }),
    .io_o_0_out({\cb_1_5_io_o_0_out[7] ,
    \cb_1_5_io_o_0_out[6] ,
    \cb_1_5_io_o_0_out[5] ,
    \cb_1_5_io_o_0_out[4] ,
    \cb_1_5_io_o_0_out[3] ,
    \cb_1_5_io_o_0_out[2] ,
    \cb_1_5_io_o_0_out[1] ,
    \cb_1_5_io_o_0_out[0] }),
    .io_o_1_out({\cb_1_5_io_o_1_out[7] ,
    \cb_1_5_io_o_1_out[6] ,
    \cb_1_5_io_o_1_out[5] ,
    \cb_1_5_io_o_1_out[4] ,
    \cb_1_5_io_o_1_out[3] ,
    \cb_1_5_io_o_1_out[2] ,
    \cb_1_5_io_o_1_out[1] ,
    \cb_1_5_io_o_1_out[0] }),
    .io_o_2_out({\cb_1_5_io_o_2_out[7] ,
    \cb_1_5_io_o_2_out[6] ,
    \cb_1_5_io_o_2_out[5] ,
    \cb_1_5_io_o_2_out[4] ,
    \cb_1_5_io_o_2_out[3] ,
    \cb_1_5_io_o_2_out[2] ,
    \cb_1_5_io_o_2_out[1] ,
    \cb_1_5_io_o_2_out[0] }),
    .io_o_3_out({\cb_1_5_io_o_3_out[7] ,
    \cb_1_5_io_o_3_out[6] ,
    \cb_1_5_io_o_3_out[5] ,
    \cb_1_5_io_o_3_out[4] ,
    \cb_1_5_io_o_3_out[3] ,
    \cb_1_5_io_o_3_out[2] ,
    \cb_1_5_io_o_3_out[1] ,
    \cb_1_5_io_o_3_out[0] }),
    .io_o_4_out({\cb_1_5_io_o_4_out[7] ,
    \cb_1_5_io_o_4_out[6] ,
    \cb_1_5_io_o_4_out[5] ,
    \cb_1_5_io_o_4_out[4] ,
    \cb_1_5_io_o_4_out[3] ,
    \cb_1_5_io_o_4_out[2] ,
    \cb_1_5_io_o_4_out[1] ,
    \cb_1_5_io_o_4_out[0] }),
    .io_o_5_out({\cb_1_5_io_o_5_out[7] ,
    \cb_1_5_io_o_5_out[6] ,
    \cb_1_5_io_o_5_out[5] ,
    \cb_1_5_io_o_5_out[4] ,
    \cb_1_5_io_o_5_out[3] ,
    \cb_1_5_io_o_5_out[2] ,
    \cb_1_5_io_o_5_out[1] ,
    \cb_1_5_io_o_5_out[0] }),
    .io_o_6_out({\cb_1_5_io_o_6_out[7] ,
    \cb_1_5_io_o_6_out[6] ,
    \cb_1_5_io_o_6_out[5] ,
    \cb_1_5_io_o_6_out[4] ,
    \cb_1_5_io_o_6_out[3] ,
    \cb_1_5_io_o_6_out[2] ,
    \cb_1_5_io_o_6_out[1] ,
    \cb_1_5_io_o_6_out[0] }),
    .io_o_7_out({\cb_1_5_io_o_7_out[7] ,
    \cb_1_5_io_o_7_out[6] ,
    \cb_1_5_io_o_7_out[5] ,
    \cb_1_5_io_o_7_out[4] ,
    \cb_1_5_io_o_7_out[3] ,
    \cb_1_5_io_o_7_out[2] ,
    \cb_1_5_io_o_7_out[1] ,
    \cb_1_5_io_o_7_out[0] }),
    .io_wo({\cb_1_4_io_eo[63] ,
    \cb_1_4_io_eo[62] ,
    \cb_1_4_io_eo[61] ,
    \cb_1_4_io_eo[60] ,
    \cb_1_4_io_eo[59] ,
    \cb_1_4_io_eo[58] ,
    \cb_1_4_io_eo[57] ,
    \cb_1_4_io_eo[56] ,
    \cb_1_4_io_eo[55] ,
    \cb_1_4_io_eo[54] ,
    \cb_1_4_io_eo[53] ,
    \cb_1_4_io_eo[52] ,
    \cb_1_4_io_eo[51] ,
    \cb_1_4_io_eo[50] ,
    \cb_1_4_io_eo[49] ,
    \cb_1_4_io_eo[48] ,
    \cb_1_4_io_eo[47] ,
    \cb_1_4_io_eo[46] ,
    \cb_1_4_io_eo[45] ,
    \cb_1_4_io_eo[44] ,
    \cb_1_4_io_eo[43] ,
    \cb_1_4_io_eo[42] ,
    \cb_1_4_io_eo[41] ,
    \cb_1_4_io_eo[40] ,
    \cb_1_4_io_eo[39] ,
    \cb_1_4_io_eo[38] ,
    \cb_1_4_io_eo[37] ,
    \cb_1_4_io_eo[36] ,
    \cb_1_4_io_eo[35] ,
    \cb_1_4_io_eo[34] ,
    \cb_1_4_io_eo[33] ,
    \cb_1_4_io_eo[32] ,
    \cb_1_4_io_eo[31] ,
    \cb_1_4_io_eo[30] ,
    \cb_1_4_io_eo[29] ,
    \cb_1_4_io_eo[28] ,
    \cb_1_4_io_eo[27] ,
    \cb_1_4_io_eo[26] ,
    \cb_1_4_io_eo[25] ,
    \cb_1_4_io_eo[24] ,
    \cb_1_4_io_eo[23] ,
    \cb_1_4_io_eo[22] ,
    \cb_1_4_io_eo[21] ,
    \cb_1_4_io_eo[20] ,
    \cb_1_4_io_eo[19] ,
    \cb_1_4_io_eo[18] ,
    \cb_1_4_io_eo[17] ,
    \cb_1_4_io_eo[16] ,
    \cb_1_4_io_eo[15] ,
    \cb_1_4_io_eo[14] ,
    \cb_1_4_io_eo[13] ,
    \cb_1_4_io_eo[12] ,
    \cb_1_4_io_eo[11] ,
    \cb_1_4_io_eo[10] ,
    \cb_1_4_io_eo[9] ,
    \cb_1_4_io_eo[8] ,
    \cb_1_4_io_eo[7] ,
    \cb_1_4_io_eo[6] ,
    \cb_1_4_io_eo[5] ,
    \cb_1_4_io_eo[4] ,
    \cb_1_4_io_eo[3] ,
    \cb_1_4_io_eo[2] ,
    \cb_1_4_io_eo[1] ,
    \cb_1_4_io_eo[0] }));
 cic_block cb_1_6 (.io_cs_i(cb_1_6_io_cs_i),
    .io_i_0_ci(cb_1_5_io_o_0_co),
    .io_i_1_ci(cb_1_5_io_o_1_co),
    .io_i_2_ci(cb_1_5_io_o_2_co),
    .io_i_3_ci(cb_1_5_io_o_3_co),
    .io_i_4_ci(cb_1_5_io_o_4_co),
    .io_i_5_ci(cb_1_5_io_o_5_co),
    .io_i_6_ci(cb_1_5_io_o_6_co),
    .io_i_7_ci(cb_1_5_io_o_7_co),
    .io_o_0_co(cb_1_6_io_o_0_co),
    .io_o_1_co(cb_1_6_io_o_1_co),
    .io_o_2_co(cb_1_6_io_o_2_co),
    .io_o_3_co(cb_1_6_io_o_3_co),
    .io_o_4_co(cb_1_6_io_o_4_co),
    .io_o_5_co(cb_1_6_io_o_5_co),
    .io_o_6_co(cb_1_6_io_o_6_co),
    .io_o_7_co(cb_1_6_io_o_7_co),
    .io_vci(cb_1_5_io_vco),
    .io_vco(cb_1_6_io_vco),
    .io_vi(cb_1_6_io_vi),
    .io_we_i(cb_1_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_1_0_io_adr_i[1] ,
    \cb_1_0_io_adr_i[0] }),
    .io_dat_i({\cb_1_0_io_dat_i[15] ,
    \cb_1_0_io_dat_i[14] ,
    \cb_1_0_io_dat_i[13] ,
    \cb_1_0_io_dat_i[12] ,
    \cb_1_0_io_dat_i[11] ,
    \cb_1_0_io_dat_i[10] ,
    \cb_1_0_io_dat_i[9] ,
    \cb_1_0_io_dat_i[8] ,
    \cb_1_0_io_dat_i[7] ,
    \cb_1_0_io_dat_i[6] ,
    \cb_1_0_io_dat_i[5] ,
    \cb_1_0_io_dat_i[4] ,
    \cb_1_0_io_dat_i[3] ,
    \cb_1_0_io_dat_i[2] ,
    \cb_1_0_io_dat_i[1] ,
    \cb_1_0_io_dat_i[0] }),
    .io_dat_o({\cb_1_6_io_dat_o[15] ,
    \cb_1_6_io_dat_o[14] ,
    \cb_1_6_io_dat_o[13] ,
    \cb_1_6_io_dat_o[12] ,
    \cb_1_6_io_dat_o[11] ,
    \cb_1_6_io_dat_o[10] ,
    \cb_1_6_io_dat_o[9] ,
    \cb_1_6_io_dat_o[8] ,
    \cb_1_6_io_dat_o[7] ,
    \cb_1_6_io_dat_o[6] ,
    \cb_1_6_io_dat_o[5] ,
    \cb_1_6_io_dat_o[4] ,
    \cb_1_6_io_dat_o[3] ,
    \cb_1_6_io_dat_o[2] ,
    \cb_1_6_io_dat_o[1] ,
    \cb_1_6_io_dat_o[0] }),
    .io_eo({\cb_1_6_io_eo[63] ,
    \cb_1_6_io_eo[62] ,
    \cb_1_6_io_eo[61] ,
    \cb_1_6_io_eo[60] ,
    \cb_1_6_io_eo[59] ,
    \cb_1_6_io_eo[58] ,
    \cb_1_6_io_eo[57] ,
    \cb_1_6_io_eo[56] ,
    \cb_1_6_io_eo[55] ,
    \cb_1_6_io_eo[54] ,
    \cb_1_6_io_eo[53] ,
    \cb_1_6_io_eo[52] ,
    \cb_1_6_io_eo[51] ,
    \cb_1_6_io_eo[50] ,
    \cb_1_6_io_eo[49] ,
    \cb_1_6_io_eo[48] ,
    \cb_1_6_io_eo[47] ,
    \cb_1_6_io_eo[46] ,
    \cb_1_6_io_eo[45] ,
    \cb_1_6_io_eo[44] ,
    \cb_1_6_io_eo[43] ,
    \cb_1_6_io_eo[42] ,
    \cb_1_6_io_eo[41] ,
    \cb_1_6_io_eo[40] ,
    \cb_1_6_io_eo[39] ,
    \cb_1_6_io_eo[38] ,
    \cb_1_6_io_eo[37] ,
    \cb_1_6_io_eo[36] ,
    \cb_1_6_io_eo[35] ,
    \cb_1_6_io_eo[34] ,
    \cb_1_6_io_eo[33] ,
    \cb_1_6_io_eo[32] ,
    \cb_1_6_io_eo[31] ,
    \cb_1_6_io_eo[30] ,
    \cb_1_6_io_eo[29] ,
    \cb_1_6_io_eo[28] ,
    \cb_1_6_io_eo[27] ,
    \cb_1_6_io_eo[26] ,
    \cb_1_6_io_eo[25] ,
    \cb_1_6_io_eo[24] ,
    \cb_1_6_io_eo[23] ,
    \cb_1_6_io_eo[22] ,
    \cb_1_6_io_eo[21] ,
    \cb_1_6_io_eo[20] ,
    \cb_1_6_io_eo[19] ,
    \cb_1_6_io_eo[18] ,
    \cb_1_6_io_eo[17] ,
    \cb_1_6_io_eo[16] ,
    \cb_1_6_io_eo[15] ,
    \cb_1_6_io_eo[14] ,
    \cb_1_6_io_eo[13] ,
    \cb_1_6_io_eo[12] ,
    \cb_1_6_io_eo[11] ,
    \cb_1_6_io_eo[10] ,
    \cb_1_6_io_eo[9] ,
    \cb_1_6_io_eo[8] ,
    \cb_1_6_io_eo[7] ,
    \cb_1_6_io_eo[6] ,
    \cb_1_6_io_eo[5] ,
    \cb_1_6_io_eo[4] ,
    \cb_1_6_io_eo[3] ,
    \cb_1_6_io_eo[2] ,
    \cb_1_6_io_eo[1] ,
    \cb_1_6_io_eo[0] }),
    .io_i_0_in1({\cb_1_5_io_o_0_out[7] ,
    \cb_1_5_io_o_0_out[6] ,
    \cb_1_5_io_o_0_out[5] ,
    \cb_1_5_io_o_0_out[4] ,
    \cb_1_5_io_o_0_out[3] ,
    \cb_1_5_io_o_0_out[2] ,
    \cb_1_5_io_o_0_out[1] ,
    \cb_1_5_io_o_0_out[0] }),
    .io_i_1_in1({\cb_1_5_io_o_1_out[7] ,
    \cb_1_5_io_o_1_out[6] ,
    \cb_1_5_io_o_1_out[5] ,
    \cb_1_5_io_o_1_out[4] ,
    \cb_1_5_io_o_1_out[3] ,
    \cb_1_5_io_o_1_out[2] ,
    \cb_1_5_io_o_1_out[1] ,
    \cb_1_5_io_o_1_out[0] }),
    .io_i_2_in1({\cb_1_5_io_o_2_out[7] ,
    \cb_1_5_io_o_2_out[6] ,
    \cb_1_5_io_o_2_out[5] ,
    \cb_1_5_io_o_2_out[4] ,
    \cb_1_5_io_o_2_out[3] ,
    \cb_1_5_io_o_2_out[2] ,
    \cb_1_5_io_o_2_out[1] ,
    \cb_1_5_io_o_2_out[0] }),
    .io_i_3_in1({\cb_1_5_io_o_3_out[7] ,
    \cb_1_5_io_o_3_out[6] ,
    \cb_1_5_io_o_3_out[5] ,
    \cb_1_5_io_o_3_out[4] ,
    \cb_1_5_io_o_3_out[3] ,
    \cb_1_5_io_o_3_out[2] ,
    \cb_1_5_io_o_3_out[1] ,
    \cb_1_5_io_o_3_out[0] }),
    .io_i_4_in1({\cb_1_5_io_o_4_out[7] ,
    \cb_1_5_io_o_4_out[6] ,
    \cb_1_5_io_o_4_out[5] ,
    \cb_1_5_io_o_4_out[4] ,
    \cb_1_5_io_o_4_out[3] ,
    \cb_1_5_io_o_4_out[2] ,
    \cb_1_5_io_o_4_out[1] ,
    \cb_1_5_io_o_4_out[0] }),
    .io_i_5_in1({\cb_1_5_io_o_5_out[7] ,
    \cb_1_5_io_o_5_out[6] ,
    \cb_1_5_io_o_5_out[5] ,
    \cb_1_5_io_o_5_out[4] ,
    \cb_1_5_io_o_5_out[3] ,
    \cb_1_5_io_o_5_out[2] ,
    \cb_1_5_io_o_5_out[1] ,
    \cb_1_5_io_o_5_out[0] }),
    .io_i_6_in1({\cb_1_5_io_o_6_out[7] ,
    \cb_1_5_io_o_6_out[6] ,
    \cb_1_5_io_o_6_out[5] ,
    \cb_1_5_io_o_6_out[4] ,
    \cb_1_5_io_o_6_out[3] ,
    \cb_1_5_io_o_6_out[2] ,
    \cb_1_5_io_o_6_out[1] ,
    \cb_1_5_io_o_6_out[0] }),
    .io_i_7_in1({\cb_1_5_io_o_7_out[7] ,
    \cb_1_5_io_o_7_out[6] ,
    \cb_1_5_io_o_7_out[5] ,
    \cb_1_5_io_o_7_out[4] ,
    \cb_1_5_io_o_7_out[3] ,
    \cb_1_5_io_o_7_out[2] ,
    \cb_1_5_io_o_7_out[1] ,
    \cb_1_5_io_o_7_out[0] }),
    .io_o_0_out({\cb_1_6_io_o_0_out[7] ,
    \cb_1_6_io_o_0_out[6] ,
    \cb_1_6_io_o_0_out[5] ,
    \cb_1_6_io_o_0_out[4] ,
    \cb_1_6_io_o_0_out[3] ,
    \cb_1_6_io_o_0_out[2] ,
    \cb_1_6_io_o_0_out[1] ,
    \cb_1_6_io_o_0_out[0] }),
    .io_o_1_out({\cb_1_6_io_o_1_out[7] ,
    \cb_1_6_io_o_1_out[6] ,
    \cb_1_6_io_o_1_out[5] ,
    \cb_1_6_io_o_1_out[4] ,
    \cb_1_6_io_o_1_out[3] ,
    \cb_1_6_io_o_1_out[2] ,
    \cb_1_6_io_o_1_out[1] ,
    \cb_1_6_io_o_1_out[0] }),
    .io_o_2_out({\cb_1_6_io_o_2_out[7] ,
    \cb_1_6_io_o_2_out[6] ,
    \cb_1_6_io_o_2_out[5] ,
    \cb_1_6_io_o_2_out[4] ,
    \cb_1_6_io_o_2_out[3] ,
    \cb_1_6_io_o_2_out[2] ,
    \cb_1_6_io_o_2_out[1] ,
    \cb_1_6_io_o_2_out[0] }),
    .io_o_3_out({\cb_1_6_io_o_3_out[7] ,
    \cb_1_6_io_o_3_out[6] ,
    \cb_1_6_io_o_3_out[5] ,
    \cb_1_6_io_o_3_out[4] ,
    \cb_1_6_io_o_3_out[3] ,
    \cb_1_6_io_o_3_out[2] ,
    \cb_1_6_io_o_3_out[1] ,
    \cb_1_6_io_o_3_out[0] }),
    .io_o_4_out({\cb_1_6_io_o_4_out[7] ,
    \cb_1_6_io_o_4_out[6] ,
    \cb_1_6_io_o_4_out[5] ,
    \cb_1_6_io_o_4_out[4] ,
    \cb_1_6_io_o_4_out[3] ,
    \cb_1_6_io_o_4_out[2] ,
    \cb_1_6_io_o_4_out[1] ,
    \cb_1_6_io_o_4_out[0] }),
    .io_o_5_out({\cb_1_6_io_o_5_out[7] ,
    \cb_1_6_io_o_5_out[6] ,
    \cb_1_6_io_o_5_out[5] ,
    \cb_1_6_io_o_5_out[4] ,
    \cb_1_6_io_o_5_out[3] ,
    \cb_1_6_io_o_5_out[2] ,
    \cb_1_6_io_o_5_out[1] ,
    \cb_1_6_io_o_5_out[0] }),
    .io_o_6_out({\cb_1_6_io_o_6_out[7] ,
    \cb_1_6_io_o_6_out[6] ,
    \cb_1_6_io_o_6_out[5] ,
    \cb_1_6_io_o_6_out[4] ,
    \cb_1_6_io_o_6_out[3] ,
    \cb_1_6_io_o_6_out[2] ,
    \cb_1_6_io_o_6_out[1] ,
    \cb_1_6_io_o_6_out[0] }),
    .io_o_7_out({\cb_1_6_io_o_7_out[7] ,
    \cb_1_6_io_o_7_out[6] ,
    \cb_1_6_io_o_7_out[5] ,
    \cb_1_6_io_o_7_out[4] ,
    \cb_1_6_io_o_7_out[3] ,
    \cb_1_6_io_o_7_out[2] ,
    \cb_1_6_io_o_7_out[1] ,
    \cb_1_6_io_o_7_out[0] }),
    .io_wo({\cb_1_5_io_eo[63] ,
    \cb_1_5_io_eo[62] ,
    \cb_1_5_io_eo[61] ,
    \cb_1_5_io_eo[60] ,
    \cb_1_5_io_eo[59] ,
    \cb_1_5_io_eo[58] ,
    \cb_1_5_io_eo[57] ,
    \cb_1_5_io_eo[56] ,
    \cb_1_5_io_eo[55] ,
    \cb_1_5_io_eo[54] ,
    \cb_1_5_io_eo[53] ,
    \cb_1_5_io_eo[52] ,
    \cb_1_5_io_eo[51] ,
    \cb_1_5_io_eo[50] ,
    \cb_1_5_io_eo[49] ,
    \cb_1_5_io_eo[48] ,
    \cb_1_5_io_eo[47] ,
    \cb_1_5_io_eo[46] ,
    \cb_1_5_io_eo[45] ,
    \cb_1_5_io_eo[44] ,
    \cb_1_5_io_eo[43] ,
    \cb_1_5_io_eo[42] ,
    \cb_1_5_io_eo[41] ,
    \cb_1_5_io_eo[40] ,
    \cb_1_5_io_eo[39] ,
    \cb_1_5_io_eo[38] ,
    \cb_1_5_io_eo[37] ,
    \cb_1_5_io_eo[36] ,
    \cb_1_5_io_eo[35] ,
    \cb_1_5_io_eo[34] ,
    \cb_1_5_io_eo[33] ,
    \cb_1_5_io_eo[32] ,
    \cb_1_5_io_eo[31] ,
    \cb_1_5_io_eo[30] ,
    \cb_1_5_io_eo[29] ,
    \cb_1_5_io_eo[28] ,
    \cb_1_5_io_eo[27] ,
    \cb_1_5_io_eo[26] ,
    \cb_1_5_io_eo[25] ,
    \cb_1_5_io_eo[24] ,
    \cb_1_5_io_eo[23] ,
    \cb_1_5_io_eo[22] ,
    \cb_1_5_io_eo[21] ,
    \cb_1_5_io_eo[20] ,
    \cb_1_5_io_eo[19] ,
    \cb_1_5_io_eo[18] ,
    \cb_1_5_io_eo[17] ,
    \cb_1_5_io_eo[16] ,
    \cb_1_5_io_eo[15] ,
    \cb_1_5_io_eo[14] ,
    \cb_1_5_io_eo[13] ,
    \cb_1_5_io_eo[12] ,
    \cb_1_5_io_eo[11] ,
    \cb_1_5_io_eo[10] ,
    \cb_1_5_io_eo[9] ,
    \cb_1_5_io_eo[8] ,
    \cb_1_5_io_eo[7] ,
    \cb_1_5_io_eo[6] ,
    \cb_1_5_io_eo[5] ,
    \cb_1_5_io_eo[4] ,
    \cb_1_5_io_eo[3] ,
    \cb_1_5_io_eo[2] ,
    \cb_1_5_io_eo[1] ,
    \cb_1_5_io_eo[0] }));
 cic_block cb_1_7 (.io_cs_i(cb_1_7_io_cs_i),
    .io_i_0_ci(cb_1_6_io_o_0_co),
    .io_i_1_ci(cb_1_6_io_o_1_co),
    .io_i_2_ci(cb_1_6_io_o_2_co),
    .io_i_3_ci(cb_1_6_io_o_3_co),
    .io_i_4_ci(cb_1_6_io_o_4_co),
    .io_i_5_ci(cb_1_6_io_o_5_co),
    .io_i_6_ci(cb_1_6_io_o_6_co),
    .io_i_7_ci(cb_1_6_io_o_7_co),
    .io_o_0_co(cb_1_7_io_o_0_co),
    .io_o_1_co(cb_1_7_io_o_1_co),
    .io_o_2_co(cb_1_7_io_o_2_co),
    .io_o_3_co(cb_1_7_io_o_3_co),
    .io_o_4_co(cb_1_7_io_o_4_co),
    .io_o_5_co(cb_1_7_io_o_5_co),
    .io_o_6_co(cb_1_7_io_o_6_co),
    .io_o_7_co(cb_1_7_io_o_7_co),
    .io_vci(cb_1_6_io_vco),
    .io_vco(cb_1_7_io_vco),
    .io_vi(cb_1_7_io_vi),
    .io_we_i(cb_1_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_1_0_io_adr_i[1] ,
    \cb_1_0_io_adr_i[0] }),
    .io_dat_i({\cb_1_0_io_dat_i[15] ,
    \cb_1_0_io_dat_i[14] ,
    \cb_1_0_io_dat_i[13] ,
    \cb_1_0_io_dat_i[12] ,
    \cb_1_0_io_dat_i[11] ,
    \cb_1_0_io_dat_i[10] ,
    \cb_1_0_io_dat_i[9] ,
    \cb_1_0_io_dat_i[8] ,
    \cb_1_0_io_dat_i[7] ,
    \cb_1_0_io_dat_i[6] ,
    \cb_1_0_io_dat_i[5] ,
    \cb_1_0_io_dat_i[4] ,
    \cb_1_0_io_dat_i[3] ,
    \cb_1_0_io_dat_i[2] ,
    \cb_1_0_io_dat_i[1] ,
    \cb_1_0_io_dat_i[0] }),
    .io_dat_o({\cb_1_7_io_dat_o[15] ,
    \cb_1_7_io_dat_o[14] ,
    \cb_1_7_io_dat_o[13] ,
    \cb_1_7_io_dat_o[12] ,
    \cb_1_7_io_dat_o[11] ,
    \cb_1_7_io_dat_o[10] ,
    \cb_1_7_io_dat_o[9] ,
    \cb_1_7_io_dat_o[8] ,
    \cb_1_7_io_dat_o[7] ,
    \cb_1_7_io_dat_o[6] ,
    \cb_1_7_io_dat_o[5] ,
    \cb_1_7_io_dat_o[4] ,
    \cb_1_7_io_dat_o[3] ,
    \cb_1_7_io_dat_o[2] ,
    \cb_1_7_io_dat_o[1] ,
    \cb_1_7_io_dat_o[0] }),
    .io_eo({\cb_1_7_io_eo[63] ,
    \cb_1_7_io_eo[62] ,
    \cb_1_7_io_eo[61] ,
    \cb_1_7_io_eo[60] ,
    \cb_1_7_io_eo[59] ,
    \cb_1_7_io_eo[58] ,
    \cb_1_7_io_eo[57] ,
    \cb_1_7_io_eo[56] ,
    \cb_1_7_io_eo[55] ,
    \cb_1_7_io_eo[54] ,
    \cb_1_7_io_eo[53] ,
    \cb_1_7_io_eo[52] ,
    \cb_1_7_io_eo[51] ,
    \cb_1_7_io_eo[50] ,
    \cb_1_7_io_eo[49] ,
    \cb_1_7_io_eo[48] ,
    \cb_1_7_io_eo[47] ,
    \cb_1_7_io_eo[46] ,
    \cb_1_7_io_eo[45] ,
    \cb_1_7_io_eo[44] ,
    \cb_1_7_io_eo[43] ,
    \cb_1_7_io_eo[42] ,
    \cb_1_7_io_eo[41] ,
    \cb_1_7_io_eo[40] ,
    \cb_1_7_io_eo[39] ,
    \cb_1_7_io_eo[38] ,
    \cb_1_7_io_eo[37] ,
    \cb_1_7_io_eo[36] ,
    \cb_1_7_io_eo[35] ,
    \cb_1_7_io_eo[34] ,
    \cb_1_7_io_eo[33] ,
    \cb_1_7_io_eo[32] ,
    \cb_1_7_io_eo[31] ,
    \cb_1_7_io_eo[30] ,
    \cb_1_7_io_eo[29] ,
    \cb_1_7_io_eo[28] ,
    \cb_1_7_io_eo[27] ,
    \cb_1_7_io_eo[26] ,
    \cb_1_7_io_eo[25] ,
    \cb_1_7_io_eo[24] ,
    \cb_1_7_io_eo[23] ,
    \cb_1_7_io_eo[22] ,
    \cb_1_7_io_eo[21] ,
    \cb_1_7_io_eo[20] ,
    \cb_1_7_io_eo[19] ,
    \cb_1_7_io_eo[18] ,
    \cb_1_7_io_eo[17] ,
    \cb_1_7_io_eo[16] ,
    \cb_1_7_io_eo[15] ,
    \cb_1_7_io_eo[14] ,
    \cb_1_7_io_eo[13] ,
    \cb_1_7_io_eo[12] ,
    \cb_1_7_io_eo[11] ,
    \cb_1_7_io_eo[10] ,
    \cb_1_7_io_eo[9] ,
    \cb_1_7_io_eo[8] ,
    \cb_1_7_io_eo[7] ,
    \cb_1_7_io_eo[6] ,
    \cb_1_7_io_eo[5] ,
    \cb_1_7_io_eo[4] ,
    \cb_1_7_io_eo[3] ,
    \cb_1_7_io_eo[2] ,
    \cb_1_7_io_eo[1] ,
    \cb_1_7_io_eo[0] }),
    .io_i_0_in1({\cb_1_6_io_o_0_out[7] ,
    \cb_1_6_io_o_0_out[6] ,
    \cb_1_6_io_o_0_out[5] ,
    \cb_1_6_io_o_0_out[4] ,
    \cb_1_6_io_o_0_out[3] ,
    \cb_1_6_io_o_0_out[2] ,
    \cb_1_6_io_o_0_out[1] ,
    \cb_1_6_io_o_0_out[0] }),
    .io_i_1_in1({\cb_1_6_io_o_1_out[7] ,
    \cb_1_6_io_o_1_out[6] ,
    \cb_1_6_io_o_1_out[5] ,
    \cb_1_6_io_o_1_out[4] ,
    \cb_1_6_io_o_1_out[3] ,
    \cb_1_6_io_o_1_out[2] ,
    \cb_1_6_io_o_1_out[1] ,
    \cb_1_6_io_o_1_out[0] }),
    .io_i_2_in1({\cb_1_6_io_o_2_out[7] ,
    \cb_1_6_io_o_2_out[6] ,
    \cb_1_6_io_o_2_out[5] ,
    \cb_1_6_io_o_2_out[4] ,
    \cb_1_6_io_o_2_out[3] ,
    \cb_1_6_io_o_2_out[2] ,
    \cb_1_6_io_o_2_out[1] ,
    \cb_1_6_io_o_2_out[0] }),
    .io_i_3_in1({\cb_1_6_io_o_3_out[7] ,
    \cb_1_6_io_o_3_out[6] ,
    \cb_1_6_io_o_3_out[5] ,
    \cb_1_6_io_o_3_out[4] ,
    \cb_1_6_io_o_3_out[3] ,
    \cb_1_6_io_o_3_out[2] ,
    \cb_1_6_io_o_3_out[1] ,
    \cb_1_6_io_o_3_out[0] }),
    .io_i_4_in1({\cb_1_6_io_o_4_out[7] ,
    \cb_1_6_io_o_4_out[6] ,
    \cb_1_6_io_o_4_out[5] ,
    \cb_1_6_io_o_4_out[4] ,
    \cb_1_6_io_o_4_out[3] ,
    \cb_1_6_io_o_4_out[2] ,
    \cb_1_6_io_o_4_out[1] ,
    \cb_1_6_io_o_4_out[0] }),
    .io_i_5_in1({\cb_1_6_io_o_5_out[7] ,
    \cb_1_6_io_o_5_out[6] ,
    \cb_1_6_io_o_5_out[5] ,
    \cb_1_6_io_o_5_out[4] ,
    \cb_1_6_io_o_5_out[3] ,
    \cb_1_6_io_o_5_out[2] ,
    \cb_1_6_io_o_5_out[1] ,
    \cb_1_6_io_o_5_out[0] }),
    .io_i_6_in1({\cb_1_6_io_o_6_out[7] ,
    \cb_1_6_io_o_6_out[6] ,
    \cb_1_6_io_o_6_out[5] ,
    \cb_1_6_io_o_6_out[4] ,
    \cb_1_6_io_o_6_out[3] ,
    \cb_1_6_io_o_6_out[2] ,
    \cb_1_6_io_o_6_out[1] ,
    \cb_1_6_io_o_6_out[0] }),
    .io_i_7_in1({\cb_1_6_io_o_7_out[7] ,
    \cb_1_6_io_o_7_out[6] ,
    \cb_1_6_io_o_7_out[5] ,
    \cb_1_6_io_o_7_out[4] ,
    \cb_1_6_io_o_7_out[3] ,
    \cb_1_6_io_o_7_out[2] ,
    \cb_1_6_io_o_7_out[1] ,
    \cb_1_6_io_o_7_out[0] }),
    .io_o_0_out({\cb_1_7_io_o_0_out[7] ,
    \cb_1_7_io_o_0_out[6] ,
    \cb_1_7_io_o_0_out[5] ,
    \cb_1_7_io_o_0_out[4] ,
    \cb_1_7_io_o_0_out[3] ,
    \cb_1_7_io_o_0_out[2] ,
    \cb_1_7_io_o_0_out[1] ,
    \cb_1_7_io_o_0_out[0] }),
    .io_o_1_out({\cb_1_7_io_o_1_out[7] ,
    \cb_1_7_io_o_1_out[6] ,
    \cb_1_7_io_o_1_out[5] ,
    \cb_1_7_io_o_1_out[4] ,
    \cb_1_7_io_o_1_out[3] ,
    \cb_1_7_io_o_1_out[2] ,
    \cb_1_7_io_o_1_out[1] ,
    \cb_1_7_io_o_1_out[0] }),
    .io_o_2_out({\cb_1_7_io_o_2_out[7] ,
    \cb_1_7_io_o_2_out[6] ,
    \cb_1_7_io_o_2_out[5] ,
    \cb_1_7_io_o_2_out[4] ,
    \cb_1_7_io_o_2_out[3] ,
    \cb_1_7_io_o_2_out[2] ,
    \cb_1_7_io_o_2_out[1] ,
    \cb_1_7_io_o_2_out[0] }),
    .io_o_3_out({\cb_1_7_io_o_3_out[7] ,
    \cb_1_7_io_o_3_out[6] ,
    \cb_1_7_io_o_3_out[5] ,
    \cb_1_7_io_o_3_out[4] ,
    \cb_1_7_io_o_3_out[3] ,
    \cb_1_7_io_o_3_out[2] ,
    \cb_1_7_io_o_3_out[1] ,
    \cb_1_7_io_o_3_out[0] }),
    .io_o_4_out({\cb_1_7_io_o_4_out[7] ,
    \cb_1_7_io_o_4_out[6] ,
    \cb_1_7_io_o_4_out[5] ,
    \cb_1_7_io_o_4_out[4] ,
    \cb_1_7_io_o_4_out[3] ,
    \cb_1_7_io_o_4_out[2] ,
    \cb_1_7_io_o_4_out[1] ,
    \cb_1_7_io_o_4_out[0] }),
    .io_o_5_out({\cb_1_7_io_o_5_out[7] ,
    \cb_1_7_io_o_5_out[6] ,
    \cb_1_7_io_o_5_out[5] ,
    \cb_1_7_io_o_5_out[4] ,
    \cb_1_7_io_o_5_out[3] ,
    \cb_1_7_io_o_5_out[2] ,
    \cb_1_7_io_o_5_out[1] ,
    \cb_1_7_io_o_5_out[0] }),
    .io_o_6_out({\cb_1_7_io_o_6_out[7] ,
    \cb_1_7_io_o_6_out[6] ,
    \cb_1_7_io_o_6_out[5] ,
    \cb_1_7_io_o_6_out[4] ,
    \cb_1_7_io_o_6_out[3] ,
    \cb_1_7_io_o_6_out[2] ,
    \cb_1_7_io_o_6_out[1] ,
    \cb_1_7_io_o_6_out[0] }),
    .io_o_7_out({\cb_1_7_io_o_7_out[7] ,
    \cb_1_7_io_o_7_out[6] ,
    \cb_1_7_io_o_7_out[5] ,
    \cb_1_7_io_o_7_out[4] ,
    \cb_1_7_io_o_7_out[3] ,
    \cb_1_7_io_o_7_out[2] ,
    \cb_1_7_io_o_7_out[1] ,
    \cb_1_7_io_o_7_out[0] }),
    .io_wo({\cb_1_6_io_eo[63] ,
    \cb_1_6_io_eo[62] ,
    \cb_1_6_io_eo[61] ,
    \cb_1_6_io_eo[60] ,
    \cb_1_6_io_eo[59] ,
    \cb_1_6_io_eo[58] ,
    \cb_1_6_io_eo[57] ,
    \cb_1_6_io_eo[56] ,
    \cb_1_6_io_eo[55] ,
    \cb_1_6_io_eo[54] ,
    \cb_1_6_io_eo[53] ,
    \cb_1_6_io_eo[52] ,
    \cb_1_6_io_eo[51] ,
    \cb_1_6_io_eo[50] ,
    \cb_1_6_io_eo[49] ,
    \cb_1_6_io_eo[48] ,
    \cb_1_6_io_eo[47] ,
    \cb_1_6_io_eo[46] ,
    \cb_1_6_io_eo[45] ,
    \cb_1_6_io_eo[44] ,
    \cb_1_6_io_eo[43] ,
    \cb_1_6_io_eo[42] ,
    \cb_1_6_io_eo[41] ,
    \cb_1_6_io_eo[40] ,
    \cb_1_6_io_eo[39] ,
    \cb_1_6_io_eo[38] ,
    \cb_1_6_io_eo[37] ,
    \cb_1_6_io_eo[36] ,
    \cb_1_6_io_eo[35] ,
    \cb_1_6_io_eo[34] ,
    \cb_1_6_io_eo[33] ,
    \cb_1_6_io_eo[32] ,
    \cb_1_6_io_eo[31] ,
    \cb_1_6_io_eo[30] ,
    \cb_1_6_io_eo[29] ,
    \cb_1_6_io_eo[28] ,
    \cb_1_6_io_eo[27] ,
    \cb_1_6_io_eo[26] ,
    \cb_1_6_io_eo[25] ,
    \cb_1_6_io_eo[24] ,
    \cb_1_6_io_eo[23] ,
    \cb_1_6_io_eo[22] ,
    \cb_1_6_io_eo[21] ,
    \cb_1_6_io_eo[20] ,
    \cb_1_6_io_eo[19] ,
    \cb_1_6_io_eo[18] ,
    \cb_1_6_io_eo[17] ,
    \cb_1_6_io_eo[16] ,
    \cb_1_6_io_eo[15] ,
    \cb_1_6_io_eo[14] ,
    \cb_1_6_io_eo[13] ,
    \cb_1_6_io_eo[12] ,
    \cb_1_6_io_eo[11] ,
    \cb_1_6_io_eo[10] ,
    \cb_1_6_io_eo[9] ,
    \cb_1_6_io_eo[8] ,
    \cb_1_6_io_eo[7] ,
    \cb_1_6_io_eo[6] ,
    \cb_1_6_io_eo[5] ,
    \cb_1_6_io_eo[4] ,
    \cb_1_6_io_eo[3] ,
    \cb_1_6_io_eo[2] ,
    \cb_1_6_io_eo[1] ,
    \cb_1_6_io_eo[0] }));
 cic_block cb_1_8 (.io_cs_i(cb_1_8_io_cs_i),
    .io_i_0_ci(cb_1_7_io_o_0_co),
    .io_i_1_ci(cb_1_7_io_o_1_co),
    .io_i_2_ci(cb_1_7_io_o_2_co),
    .io_i_3_ci(cb_1_7_io_o_3_co),
    .io_i_4_ci(cb_1_7_io_o_4_co),
    .io_i_5_ci(cb_1_7_io_o_5_co),
    .io_i_6_ci(cb_1_7_io_o_6_co),
    .io_i_7_ci(cb_1_7_io_o_7_co),
    .io_o_0_co(cb_1_8_io_o_0_co),
    .io_o_1_co(cb_1_8_io_o_1_co),
    .io_o_2_co(cb_1_8_io_o_2_co),
    .io_o_3_co(cb_1_8_io_o_3_co),
    .io_o_4_co(cb_1_8_io_o_4_co),
    .io_o_5_co(cb_1_8_io_o_5_co),
    .io_o_6_co(cb_1_8_io_o_6_co),
    .io_o_7_co(cb_1_8_io_o_7_co),
    .io_vci(cb_1_7_io_vco),
    .io_vco(cb_1_8_io_vco),
    .io_vi(cb_1_8_io_vi),
    .io_we_i(cb_1_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_1_0_io_adr_i[1] ,
    \cb_1_0_io_adr_i[0] }),
    .io_dat_i({\cb_1_0_io_dat_i[15] ,
    \cb_1_0_io_dat_i[14] ,
    \cb_1_0_io_dat_i[13] ,
    \cb_1_0_io_dat_i[12] ,
    \cb_1_0_io_dat_i[11] ,
    \cb_1_0_io_dat_i[10] ,
    \cb_1_0_io_dat_i[9] ,
    \cb_1_0_io_dat_i[8] ,
    \cb_1_0_io_dat_i[7] ,
    \cb_1_0_io_dat_i[6] ,
    \cb_1_0_io_dat_i[5] ,
    \cb_1_0_io_dat_i[4] ,
    \cb_1_0_io_dat_i[3] ,
    \cb_1_0_io_dat_i[2] ,
    \cb_1_0_io_dat_i[1] ,
    \cb_1_0_io_dat_i[0] }),
    .io_dat_o({\cb_1_8_io_dat_o[15] ,
    \cb_1_8_io_dat_o[14] ,
    \cb_1_8_io_dat_o[13] ,
    \cb_1_8_io_dat_o[12] ,
    \cb_1_8_io_dat_o[11] ,
    \cb_1_8_io_dat_o[10] ,
    \cb_1_8_io_dat_o[9] ,
    \cb_1_8_io_dat_o[8] ,
    \cb_1_8_io_dat_o[7] ,
    \cb_1_8_io_dat_o[6] ,
    \cb_1_8_io_dat_o[5] ,
    \cb_1_8_io_dat_o[4] ,
    \cb_1_8_io_dat_o[3] ,
    \cb_1_8_io_dat_o[2] ,
    \cb_1_8_io_dat_o[1] ,
    \cb_1_8_io_dat_o[0] }),
    .io_eo({\cb_1_8_io_eo[63] ,
    \cb_1_8_io_eo[62] ,
    \cb_1_8_io_eo[61] ,
    \cb_1_8_io_eo[60] ,
    \cb_1_8_io_eo[59] ,
    \cb_1_8_io_eo[58] ,
    \cb_1_8_io_eo[57] ,
    \cb_1_8_io_eo[56] ,
    \cb_1_8_io_eo[55] ,
    \cb_1_8_io_eo[54] ,
    \cb_1_8_io_eo[53] ,
    \cb_1_8_io_eo[52] ,
    \cb_1_8_io_eo[51] ,
    \cb_1_8_io_eo[50] ,
    \cb_1_8_io_eo[49] ,
    \cb_1_8_io_eo[48] ,
    \cb_1_8_io_eo[47] ,
    \cb_1_8_io_eo[46] ,
    \cb_1_8_io_eo[45] ,
    \cb_1_8_io_eo[44] ,
    \cb_1_8_io_eo[43] ,
    \cb_1_8_io_eo[42] ,
    \cb_1_8_io_eo[41] ,
    \cb_1_8_io_eo[40] ,
    \cb_1_8_io_eo[39] ,
    \cb_1_8_io_eo[38] ,
    \cb_1_8_io_eo[37] ,
    \cb_1_8_io_eo[36] ,
    \cb_1_8_io_eo[35] ,
    \cb_1_8_io_eo[34] ,
    \cb_1_8_io_eo[33] ,
    \cb_1_8_io_eo[32] ,
    \cb_1_8_io_eo[31] ,
    \cb_1_8_io_eo[30] ,
    \cb_1_8_io_eo[29] ,
    \cb_1_8_io_eo[28] ,
    \cb_1_8_io_eo[27] ,
    \cb_1_8_io_eo[26] ,
    \cb_1_8_io_eo[25] ,
    \cb_1_8_io_eo[24] ,
    \cb_1_8_io_eo[23] ,
    \cb_1_8_io_eo[22] ,
    \cb_1_8_io_eo[21] ,
    \cb_1_8_io_eo[20] ,
    \cb_1_8_io_eo[19] ,
    \cb_1_8_io_eo[18] ,
    \cb_1_8_io_eo[17] ,
    \cb_1_8_io_eo[16] ,
    \cb_1_8_io_eo[15] ,
    \cb_1_8_io_eo[14] ,
    \cb_1_8_io_eo[13] ,
    \cb_1_8_io_eo[12] ,
    \cb_1_8_io_eo[11] ,
    \cb_1_8_io_eo[10] ,
    \cb_1_8_io_eo[9] ,
    \cb_1_8_io_eo[8] ,
    \cb_1_8_io_eo[7] ,
    \cb_1_8_io_eo[6] ,
    \cb_1_8_io_eo[5] ,
    \cb_1_8_io_eo[4] ,
    \cb_1_8_io_eo[3] ,
    \cb_1_8_io_eo[2] ,
    \cb_1_8_io_eo[1] ,
    \cb_1_8_io_eo[0] }),
    .io_i_0_in1({\cb_1_7_io_o_0_out[7] ,
    \cb_1_7_io_o_0_out[6] ,
    \cb_1_7_io_o_0_out[5] ,
    \cb_1_7_io_o_0_out[4] ,
    \cb_1_7_io_o_0_out[3] ,
    \cb_1_7_io_o_0_out[2] ,
    \cb_1_7_io_o_0_out[1] ,
    \cb_1_7_io_o_0_out[0] }),
    .io_i_1_in1({\cb_1_7_io_o_1_out[7] ,
    \cb_1_7_io_o_1_out[6] ,
    \cb_1_7_io_o_1_out[5] ,
    \cb_1_7_io_o_1_out[4] ,
    \cb_1_7_io_o_1_out[3] ,
    \cb_1_7_io_o_1_out[2] ,
    \cb_1_7_io_o_1_out[1] ,
    \cb_1_7_io_o_1_out[0] }),
    .io_i_2_in1({\cb_1_7_io_o_2_out[7] ,
    \cb_1_7_io_o_2_out[6] ,
    \cb_1_7_io_o_2_out[5] ,
    \cb_1_7_io_o_2_out[4] ,
    \cb_1_7_io_o_2_out[3] ,
    \cb_1_7_io_o_2_out[2] ,
    \cb_1_7_io_o_2_out[1] ,
    \cb_1_7_io_o_2_out[0] }),
    .io_i_3_in1({\cb_1_7_io_o_3_out[7] ,
    \cb_1_7_io_o_3_out[6] ,
    \cb_1_7_io_o_3_out[5] ,
    \cb_1_7_io_o_3_out[4] ,
    \cb_1_7_io_o_3_out[3] ,
    \cb_1_7_io_o_3_out[2] ,
    \cb_1_7_io_o_3_out[1] ,
    \cb_1_7_io_o_3_out[0] }),
    .io_i_4_in1({\cb_1_7_io_o_4_out[7] ,
    \cb_1_7_io_o_4_out[6] ,
    \cb_1_7_io_o_4_out[5] ,
    \cb_1_7_io_o_4_out[4] ,
    \cb_1_7_io_o_4_out[3] ,
    \cb_1_7_io_o_4_out[2] ,
    \cb_1_7_io_o_4_out[1] ,
    \cb_1_7_io_o_4_out[0] }),
    .io_i_5_in1({\cb_1_7_io_o_5_out[7] ,
    \cb_1_7_io_o_5_out[6] ,
    \cb_1_7_io_o_5_out[5] ,
    \cb_1_7_io_o_5_out[4] ,
    \cb_1_7_io_o_5_out[3] ,
    \cb_1_7_io_o_5_out[2] ,
    \cb_1_7_io_o_5_out[1] ,
    \cb_1_7_io_o_5_out[0] }),
    .io_i_6_in1({\cb_1_7_io_o_6_out[7] ,
    \cb_1_7_io_o_6_out[6] ,
    \cb_1_7_io_o_6_out[5] ,
    \cb_1_7_io_o_6_out[4] ,
    \cb_1_7_io_o_6_out[3] ,
    \cb_1_7_io_o_6_out[2] ,
    \cb_1_7_io_o_6_out[1] ,
    \cb_1_7_io_o_6_out[0] }),
    .io_i_7_in1({\cb_1_7_io_o_7_out[7] ,
    \cb_1_7_io_o_7_out[6] ,
    \cb_1_7_io_o_7_out[5] ,
    \cb_1_7_io_o_7_out[4] ,
    \cb_1_7_io_o_7_out[3] ,
    \cb_1_7_io_o_7_out[2] ,
    \cb_1_7_io_o_7_out[1] ,
    \cb_1_7_io_o_7_out[0] }),
    .io_o_0_out({\cb_1_8_io_o_0_out[7] ,
    \cb_1_8_io_o_0_out[6] ,
    \cb_1_8_io_o_0_out[5] ,
    \cb_1_8_io_o_0_out[4] ,
    \cb_1_8_io_o_0_out[3] ,
    \cb_1_8_io_o_0_out[2] ,
    \cb_1_8_io_o_0_out[1] ,
    \cb_1_8_io_o_0_out[0] }),
    .io_o_1_out({\cb_1_8_io_o_1_out[7] ,
    \cb_1_8_io_o_1_out[6] ,
    \cb_1_8_io_o_1_out[5] ,
    \cb_1_8_io_o_1_out[4] ,
    \cb_1_8_io_o_1_out[3] ,
    \cb_1_8_io_o_1_out[2] ,
    \cb_1_8_io_o_1_out[1] ,
    \cb_1_8_io_o_1_out[0] }),
    .io_o_2_out({\cb_1_8_io_o_2_out[7] ,
    \cb_1_8_io_o_2_out[6] ,
    \cb_1_8_io_o_2_out[5] ,
    \cb_1_8_io_o_2_out[4] ,
    \cb_1_8_io_o_2_out[3] ,
    \cb_1_8_io_o_2_out[2] ,
    \cb_1_8_io_o_2_out[1] ,
    \cb_1_8_io_o_2_out[0] }),
    .io_o_3_out({\cb_1_8_io_o_3_out[7] ,
    \cb_1_8_io_o_3_out[6] ,
    \cb_1_8_io_o_3_out[5] ,
    \cb_1_8_io_o_3_out[4] ,
    \cb_1_8_io_o_3_out[3] ,
    \cb_1_8_io_o_3_out[2] ,
    \cb_1_8_io_o_3_out[1] ,
    \cb_1_8_io_o_3_out[0] }),
    .io_o_4_out({\cb_1_8_io_o_4_out[7] ,
    \cb_1_8_io_o_4_out[6] ,
    \cb_1_8_io_o_4_out[5] ,
    \cb_1_8_io_o_4_out[4] ,
    \cb_1_8_io_o_4_out[3] ,
    \cb_1_8_io_o_4_out[2] ,
    \cb_1_8_io_o_4_out[1] ,
    \cb_1_8_io_o_4_out[0] }),
    .io_o_5_out({\cb_1_8_io_o_5_out[7] ,
    \cb_1_8_io_o_5_out[6] ,
    \cb_1_8_io_o_5_out[5] ,
    \cb_1_8_io_o_5_out[4] ,
    \cb_1_8_io_o_5_out[3] ,
    \cb_1_8_io_o_5_out[2] ,
    \cb_1_8_io_o_5_out[1] ,
    \cb_1_8_io_o_5_out[0] }),
    .io_o_6_out({\cb_1_8_io_o_6_out[7] ,
    \cb_1_8_io_o_6_out[6] ,
    \cb_1_8_io_o_6_out[5] ,
    \cb_1_8_io_o_6_out[4] ,
    \cb_1_8_io_o_6_out[3] ,
    \cb_1_8_io_o_6_out[2] ,
    \cb_1_8_io_o_6_out[1] ,
    \cb_1_8_io_o_6_out[0] }),
    .io_o_7_out({\cb_1_8_io_o_7_out[7] ,
    \cb_1_8_io_o_7_out[6] ,
    \cb_1_8_io_o_7_out[5] ,
    \cb_1_8_io_o_7_out[4] ,
    \cb_1_8_io_o_7_out[3] ,
    \cb_1_8_io_o_7_out[2] ,
    \cb_1_8_io_o_7_out[1] ,
    \cb_1_8_io_o_7_out[0] }),
    .io_wo({\cb_1_7_io_eo[63] ,
    \cb_1_7_io_eo[62] ,
    \cb_1_7_io_eo[61] ,
    \cb_1_7_io_eo[60] ,
    \cb_1_7_io_eo[59] ,
    \cb_1_7_io_eo[58] ,
    \cb_1_7_io_eo[57] ,
    \cb_1_7_io_eo[56] ,
    \cb_1_7_io_eo[55] ,
    \cb_1_7_io_eo[54] ,
    \cb_1_7_io_eo[53] ,
    \cb_1_7_io_eo[52] ,
    \cb_1_7_io_eo[51] ,
    \cb_1_7_io_eo[50] ,
    \cb_1_7_io_eo[49] ,
    \cb_1_7_io_eo[48] ,
    \cb_1_7_io_eo[47] ,
    \cb_1_7_io_eo[46] ,
    \cb_1_7_io_eo[45] ,
    \cb_1_7_io_eo[44] ,
    \cb_1_7_io_eo[43] ,
    \cb_1_7_io_eo[42] ,
    \cb_1_7_io_eo[41] ,
    \cb_1_7_io_eo[40] ,
    \cb_1_7_io_eo[39] ,
    \cb_1_7_io_eo[38] ,
    \cb_1_7_io_eo[37] ,
    \cb_1_7_io_eo[36] ,
    \cb_1_7_io_eo[35] ,
    \cb_1_7_io_eo[34] ,
    \cb_1_7_io_eo[33] ,
    \cb_1_7_io_eo[32] ,
    \cb_1_7_io_eo[31] ,
    \cb_1_7_io_eo[30] ,
    \cb_1_7_io_eo[29] ,
    \cb_1_7_io_eo[28] ,
    \cb_1_7_io_eo[27] ,
    \cb_1_7_io_eo[26] ,
    \cb_1_7_io_eo[25] ,
    \cb_1_7_io_eo[24] ,
    \cb_1_7_io_eo[23] ,
    \cb_1_7_io_eo[22] ,
    \cb_1_7_io_eo[21] ,
    \cb_1_7_io_eo[20] ,
    \cb_1_7_io_eo[19] ,
    \cb_1_7_io_eo[18] ,
    \cb_1_7_io_eo[17] ,
    \cb_1_7_io_eo[16] ,
    \cb_1_7_io_eo[15] ,
    \cb_1_7_io_eo[14] ,
    \cb_1_7_io_eo[13] ,
    \cb_1_7_io_eo[12] ,
    \cb_1_7_io_eo[11] ,
    \cb_1_7_io_eo[10] ,
    \cb_1_7_io_eo[9] ,
    \cb_1_7_io_eo[8] ,
    \cb_1_7_io_eo[7] ,
    \cb_1_7_io_eo[6] ,
    \cb_1_7_io_eo[5] ,
    \cb_1_7_io_eo[4] ,
    \cb_1_7_io_eo[3] ,
    \cb_1_7_io_eo[2] ,
    \cb_1_7_io_eo[1] ,
    \cb_1_7_io_eo[0] }));
 cic_block cb_1_9 (.io_cs_i(cb_1_9_io_cs_i),
    .io_i_0_ci(cb_1_8_io_o_0_co),
    .io_i_1_ci(cb_1_8_io_o_1_co),
    .io_i_2_ci(cb_1_8_io_o_2_co),
    .io_i_3_ci(cb_1_8_io_o_3_co),
    .io_i_4_ci(cb_1_8_io_o_4_co),
    .io_i_5_ci(cb_1_8_io_o_5_co),
    .io_i_6_ci(cb_1_8_io_o_6_co),
    .io_i_7_ci(cb_1_8_io_o_7_co),
    .io_o_0_co(cb_1_10_io_i_0_ci),
    .io_o_1_co(cb_1_10_io_i_1_ci),
    .io_o_2_co(cb_1_10_io_i_2_ci),
    .io_o_3_co(cb_1_10_io_i_3_ci),
    .io_o_4_co(cb_1_10_io_i_4_ci),
    .io_o_5_co(cb_1_10_io_i_5_ci),
    .io_o_6_co(cb_1_10_io_i_6_ci),
    .io_o_7_co(cb_1_10_io_i_7_ci),
    .io_vci(cb_1_8_io_vco),
    .io_vco(cb_1_10_io_vci),
    .io_vi(cb_1_9_io_vi),
    .io_we_i(cb_1_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_1_0_io_adr_i[1] ,
    \cb_1_0_io_adr_i[0] }),
    .io_dat_i({\cb_1_0_io_dat_i[15] ,
    \cb_1_0_io_dat_i[14] ,
    \cb_1_0_io_dat_i[13] ,
    \cb_1_0_io_dat_i[12] ,
    \cb_1_0_io_dat_i[11] ,
    \cb_1_0_io_dat_i[10] ,
    \cb_1_0_io_dat_i[9] ,
    \cb_1_0_io_dat_i[8] ,
    \cb_1_0_io_dat_i[7] ,
    \cb_1_0_io_dat_i[6] ,
    \cb_1_0_io_dat_i[5] ,
    \cb_1_0_io_dat_i[4] ,
    \cb_1_0_io_dat_i[3] ,
    \cb_1_0_io_dat_i[2] ,
    \cb_1_0_io_dat_i[1] ,
    \cb_1_0_io_dat_i[0] }),
    .io_dat_o({\cb_1_9_io_dat_o[15] ,
    \cb_1_9_io_dat_o[14] ,
    \cb_1_9_io_dat_o[13] ,
    \cb_1_9_io_dat_o[12] ,
    \cb_1_9_io_dat_o[11] ,
    \cb_1_9_io_dat_o[10] ,
    \cb_1_9_io_dat_o[9] ,
    \cb_1_9_io_dat_o[8] ,
    \cb_1_9_io_dat_o[7] ,
    \cb_1_9_io_dat_o[6] ,
    \cb_1_9_io_dat_o[5] ,
    \cb_1_9_io_dat_o[4] ,
    \cb_1_9_io_dat_o[3] ,
    \cb_1_9_io_dat_o[2] ,
    \cb_1_9_io_dat_o[1] ,
    \cb_1_9_io_dat_o[0] }),
    .io_eo({\cb_1_10_io_wo[63] ,
    \cb_1_10_io_wo[62] ,
    \cb_1_10_io_wo[61] ,
    \cb_1_10_io_wo[60] ,
    \cb_1_10_io_wo[59] ,
    \cb_1_10_io_wo[58] ,
    \cb_1_10_io_wo[57] ,
    \cb_1_10_io_wo[56] ,
    \cb_1_10_io_wo[55] ,
    \cb_1_10_io_wo[54] ,
    \cb_1_10_io_wo[53] ,
    \cb_1_10_io_wo[52] ,
    \cb_1_10_io_wo[51] ,
    \cb_1_10_io_wo[50] ,
    \cb_1_10_io_wo[49] ,
    \cb_1_10_io_wo[48] ,
    \cb_1_10_io_wo[47] ,
    \cb_1_10_io_wo[46] ,
    \cb_1_10_io_wo[45] ,
    \cb_1_10_io_wo[44] ,
    \cb_1_10_io_wo[43] ,
    \cb_1_10_io_wo[42] ,
    \cb_1_10_io_wo[41] ,
    \cb_1_10_io_wo[40] ,
    \cb_1_10_io_wo[39] ,
    \cb_1_10_io_wo[38] ,
    \cb_1_10_io_wo[37] ,
    \cb_1_10_io_wo[36] ,
    \cb_1_10_io_wo[35] ,
    \cb_1_10_io_wo[34] ,
    \cb_1_10_io_wo[33] ,
    \cb_1_10_io_wo[32] ,
    \cb_1_10_io_wo[31] ,
    \cb_1_10_io_wo[30] ,
    \cb_1_10_io_wo[29] ,
    \cb_1_10_io_wo[28] ,
    \cb_1_10_io_wo[27] ,
    \cb_1_10_io_wo[26] ,
    \cb_1_10_io_wo[25] ,
    \cb_1_10_io_wo[24] ,
    \cb_1_10_io_wo[23] ,
    \cb_1_10_io_wo[22] ,
    \cb_1_10_io_wo[21] ,
    \cb_1_10_io_wo[20] ,
    \cb_1_10_io_wo[19] ,
    \cb_1_10_io_wo[18] ,
    \cb_1_10_io_wo[17] ,
    \cb_1_10_io_wo[16] ,
    \cb_1_10_io_wo[15] ,
    \cb_1_10_io_wo[14] ,
    \cb_1_10_io_wo[13] ,
    \cb_1_10_io_wo[12] ,
    \cb_1_10_io_wo[11] ,
    \cb_1_10_io_wo[10] ,
    \cb_1_10_io_wo[9] ,
    \cb_1_10_io_wo[8] ,
    \cb_1_10_io_wo[7] ,
    \cb_1_10_io_wo[6] ,
    \cb_1_10_io_wo[5] ,
    \cb_1_10_io_wo[4] ,
    \cb_1_10_io_wo[3] ,
    \cb_1_10_io_wo[2] ,
    \cb_1_10_io_wo[1] ,
    \cb_1_10_io_wo[0] }),
    .io_i_0_in1({\cb_1_8_io_o_0_out[7] ,
    \cb_1_8_io_o_0_out[6] ,
    \cb_1_8_io_o_0_out[5] ,
    \cb_1_8_io_o_0_out[4] ,
    \cb_1_8_io_o_0_out[3] ,
    \cb_1_8_io_o_0_out[2] ,
    \cb_1_8_io_o_0_out[1] ,
    \cb_1_8_io_o_0_out[0] }),
    .io_i_1_in1({\cb_1_8_io_o_1_out[7] ,
    \cb_1_8_io_o_1_out[6] ,
    \cb_1_8_io_o_1_out[5] ,
    \cb_1_8_io_o_1_out[4] ,
    \cb_1_8_io_o_1_out[3] ,
    \cb_1_8_io_o_1_out[2] ,
    \cb_1_8_io_o_1_out[1] ,
    \cb_1_8_io_o_1_out[0] }),
    .io_i_2_in1({\cb_1_8_io_o_2_out[7] ,
    \cb_1_8_io_o_2_out[6] ,
    \cb_1_8_io_o_2_out[5] ,
    \cb_1_8_io_o_2_out[4] ,
    \cb_1_8_io_o_2_out[3] ,
    \cb_1_8_io_o_2_out[2] ,
    \cb_1_8_io_o_2_out[1] ,
    \cb_1_8_io_o_2_out[0] }),
    .io_i_3_in1({\cb_1_8_io_o_3_out[7] ,
    \cb_1_8_io_o_3_out[6] ,
    \cb_1_8_io_o_3_out[5] ,
    \cb_1_8_io_o_3_out[4] ,
    \cb_1_8_io_o_3_out[3] ,
    \cb_1_8_io_o_3_out[2] ,
    \cb_1_8_io_o_3_out[1] ,
    \cb_1_8_io_o_3_out[0] }),
    .io_i_4_in1({\cb_1_8_io_o_4_out[7] ,
    \cb_1_8_io_o_4_out[6] ,
    \cb_1_8_io_o_4_out[5] ,
    \cb_1_8_io_o_4_out[4] ,
    \cb_1_8_io_o_4_out[3] ,
    \cb_1_8_io_o_4_out[2] ,
    \cb_1_8_io_o_4_out[1] ,
    \cb_1_8_io_o_4_out[0] }),
    .io_i_5_in1({\cb_1_8_io_o_5_out[7] ,
    \cb_1_8_io_o_5_out[6] ,
    \cb_1_8_io_o_5_out[5] ,
    \cb_1_8_io_o_5_out[4] ,
    \cb_1_8_io_o_5_out[3] ,
    \cb_1_8_io_o_5_out[2] ,
    \cb_1_8_io_o_5_out[1] ,
    \cb_1_8_io_o_5_out[0] }),
    .io_i_6_in1({\cb_1_8_io_o_6_out[7] ,
    \cb_1_8_io_o_6_out[6] ,
    \cb_1_8_io_o_6_out[5] ,
    \cb_1_8_io_o_6_out[4] ,
    \cb_1_8_io_o_6_out[3] ,
    \cb_1_8_io_o_6_out[2] ,
    \cb_1_8_io_o_6_out[1] ,
    \cb_1_8_io_o_6_out[0] }),
    .io_i_7_in1({\cb_1_8_io_o_7_out[7] ,
    \cb_1_8_io_o_7_out[6] ,
    \cb_1_8_io_o_7_out[5] ,
    \cb_1_8_io_o_7_out[4] ,
    \cb_1_8_io_o_7_out[3] ,
    \cb_1_8_io_o_7_out[2] ,
    \cb_1_8_io_o_7_out[1] ,
    \cb_1_8_io_o_7_out[0] }),
    .io_o_0_out({\cb_1_10_io_i_0_in1[7] ,
    \cb_1_10_io_i_0_in1[6] ,
    \cb_1_10_io_i_0_in1[5] ,
    \cb_1_10_io_i_0_in1[4] ,
    \cb_1_10_io_i_0_in1[3] ,
    \cb_1_10_io_i_0_in1[2] ,
    \cb_1_10_io_i_0_in1[1] ,
    \cb_1_10_io_i_0_in1[0] }),
    .io_o_1_out({\cb_1_10_io_i_1_in1[7] ,
    \cb_1_10_io_i_1_in1[6] ,
    \cb_1_10_io_i_1_in1[5] ,
    \cb_1_10_io_i_1_in1[4] ,
    \cb_1_10_io_i_1_in1[3] ,
    \cb_1_10_io_i_1_in1[2] ,
    \cb_1_10_io_i_1_in1[1] ,
    \cb_1_10_io_i_1_in1[0] }),
    .io_o_2_out({\cb_1_10_io_i_2_in1[7] ,
    \cb_1_10_io_i_2_in1[6] ,
    \cb_1_10_io_i_2_in1[5] ,
    \cb_1_10_io_i_2_in1[4] ,
    \cb_1_10_io_i_2_in1[3] ,
    \cb_1_10_io_i_2_in1[2] ,
    \cb_1_10_io_i_2_in1[1] ,
    \cb_1_10_io_i_2_in1[0] }),
    .io_o_3_out({\cb_1_10_io_i_3_in1[7] ,
    \cb_1_10_io_i_3_in1[6] ,
    \cb_1_10_io_i_3_in1[5] ,
    \cb_1_10_io_i_3_in1[4] ,
    \cb_1_10_io_i_3_in1[3] ,
    \cb_1_10_io_i_3_in1[2] ,
    \cb_1_10_io_i_3_in1[1] ,
    \cb_1_10_io_i_3_in1[0] }),
    .io_o_4_out({\cb_1_10_io_i_4_in1[7] ,
    \cb_1_10_io_i_4_in1[6] ,
    \cb_1_10_io_i_4_in1[5] ,
    \cb_1_10_io_i_4_in1[4] ,
    \cb_1_10_io_i_4_in1[3] ,
    \cb_1_10_io_i_4_in1[2] ,
    \cb_1_10_io_i_4_in1[1] ,
    \cb_1_10_io_i_4_in1[0] }),
    .io_o_5_out({\cb_1_10_io_i_5_in1[7] ,
    \cb_1_10_io_i_5_in1[6] ,
    \cb_1_10_io_i_5_in1[5] ,
    \cb_1_10_io_i_5_in1[4] ,
    \cb_1_10_io_i_5_in1[3] ,
    \cb_1_10_io_i_5_in1[2] ,
    \cb_1_10_io_i_5_in1[1] ,
    \cb_1_10_io_i_5_in1[0] }),
    .io_o_6_out({\cb_1_10_io_i_6_in1[7] ,
    \cb_1_10_io_i_6_in1[6] ,
    \cb_1_10_io_i_6_in1[5] ,
    \cb_1_10_io_i_6_in1[4] ,
    \cb_1_10_io_i_6_in1[3] ,
    \cb_1_10_io_i_6_in1[2] ,
    \cb_1_10_io_i_6_in1[1] ,
    \cb_1_10_io_i_6_in1[0] }),
    .io_o_7_out({\cb_1_10_io_i_7_in1[7] ,
    \cb_1_10_io_i_7_in1[6] ,
    \cb_1_10_io_i_7_in1[5] ,
    \cb_1_10_io_i_7_in1[4] ,
    \cb_1_10_io_i_7_in1[3] ,
    \cb_1_10_io_i_7_in1[2] ,
    \cb_1_10_io_i_7_in1[1] ,
    \cb_1_10_io_i_7_in1[0] }),
    .io_wo({\cb_1_8_io_eo[63] ,
    \cb_1_8_io_eo[62] ,
    \cb_1_8_io_eo[61] ,
    \cb_1_8_io_eo[60] ,
    \cb_1_8_io_eo[59] ,
    \cb_1_8_io_eo[58] ,
    \cb_1_8_io_eo[57] ,
    \cb_1_8_io_eo[56] ,
    \cb_1_8_io_eo[55] ,
    \cb_1_8_io_eo[54] ,
    \cb_1_8_io_eo[53] ,
    \cb_1_8_io_eo[52] ,
    \cb_1_8_io_eo[51] ,
    \cb_1_8_io_eo[50] ,
    \cb_1_8_io_eo[49] ,
    \cb_1_8_io_eo[48] ,
    \cb_1_8_io_eo[47] ,
    \cb_1_8_io_eo[46] ,
    \cb_1_8_io_eo[45] ,
    \cb_1_8_io_eo[44] ,
    \cb_1_8_io_eo[43] ,
    \cb_1_8_io_eo[42] ,
    \cb_1_8_io_eo[41] ,
    \cb_1_8_io_eo[40] ,
    \cb_1_8_io_eo[39] ,
    \cb_1_8_io_eo[38] ,
    \cb_1_8_io_eo[37] ,
    \cb_1_8_io_eo[36] ,
    \cb_1_8_io_eo[35] ,
    \cb_1_8_io_eo[34] ,
    \cb_1_8_io_eo[33] ,
    \cb_1_8_io_eo[32] ,
    \cb_1_8_io_eo[31] ,
    \cb_1_8_io_eo[30] ,
    \cb_1_8_io_eo[29] ,
    \cb_1_8_io_eo[28] ,
    \cb_1_8_io_eo[27] ,
    \cb_1_8_io_eo[26] ,
    \cb_1_8_io_eo[25] ,
    \cb_1_8_io_eo[24] ,
    \cb_1_8_io_eo[23] ,
    \cb_1_8_io_eo[22] ,
    \cb_1_8_io_eo[21] ,
    \cb_1_8_io_eo[20] ,
    \cb_1_8_io_eo[19] ,
    \cb_1_8_io_eo[18] ,
    \cb_1_8_io_eo[17] ,
    \cb_1_8_io_eo[16] ,
    \cb_1_8_io_eo[15] ,
    \cb_1_8_io_eo[14] ,
    \cb_1_8_io_eo[13] ,
    \cb_1_8_io_eo[12] ,
    \cb_1_8_io_eo[11] ,
    \cb_1_8_io_eo[10] ,
    \cb_1_8_io_eo[9] ,
    \cb_1_8_io_eo[8] ,
    \cb_1_8_io_eo[7] ,
    \cb_1_8_io_eo[6] ,
    \cb_1_8_io_eo[5] ,
    \cb_1_8_io_eo[4] ,
    \cb_1_8_io_eo[3] ,
    \cb_1_8_io_eo[2] ,
    \cb_1_8_io_eo[1] ,
    \cb_1_8_io_eo[0] }));
 cic_block cb_2_0 (.io_cs_i(cb_2_0_io_cs_i),
    .io_i_0_ci(cb_2_0_io_i_0_ci),
    .io_o_0_co(cb_2_0_io_o_0_co),
    .io_o_1_co(cb_2_0_io_o_1_co),
    .io_o_2_co(cb_2_0_io_o_2_co),
    .io_o_3_co(cb_2_0_io_o_3_co),
    .io_o_4_co(cb_2_0_io_o_4_co),
    .io_o_5_co(cb_2_0_io_o_5_co),
    .io_o_6_co(cb_2_0_io_o_6_co),
    .io_o_7_co(cb_2_0_io_o_7_co),
    .io_vco(cb_2_0_io_vco),
    .io_vi(cb_2_0_io_vi),
    .io_we_i(cb_2_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_2_0_io_adr_i[1] ,
    \cb_2_0_io_adr_i[0] }),
    .io_dat_i({\cb_2_0_io_dat_i[15] ,
    \cb_2_0_io_dat_i[14] ,
    \cb_2_0_io_dat_i[13] ,
    \cb_2_0_io_dat_i[12] ,
    \cb_2_0_io_dat_i[11] ,
    \cb_2_0_io_dat_i[10] ,
    \cb_2_0_io_dat_i[9] ,
    \cb_2_0_io_dat_i[8] ,
    \cb_2_0_io_dat_i[7] ,
    \cb_2_0_io_dat_i[6] ,
    \cb_2_0_io_dat_i[5] ,
    \cb_2_0_io_dat_i[4] ,
    \cb_2_0_io_dat_i[3] ,
    \cb_2_0_io_dat_i[2] ,
    \cb_2_0_io_dat_i[1] ,
    \cb_2_0_io_dat_i[0] }),
    .io_dat_o({\cb_2_0_io_dat_o[15] ,
    \cb_2_0_io_dat_o[14] ,
    \cb_2_0_io_dat_o[13] ,
    \cb_2_0_io_dat_o[12] ,
    \cb_2_0_io_dat_o[11] ,
    \cb_2_0_io_dat_o[10] ,
    \cb_2_0_io_dat_o[9] ,
    \cb_2_0_io_dat_o[8] ,
    \cb_2_0_io_dat_o[7] ,
    \cb_2_0_io_dat_o[6] ,
    \cb_2_0_io_dat_o[5] ,
    \cb_2_0_io_dat_o[4] ,
    \cb_2_0_io_dat_o[3] ,
    \cb_2_0_io_dat_o[2] ,
    \cb_2_0_io_dat_o[1] ,
    \cb_2_0_io_dat_o[0] }),
    .io_eo({\cb_2_0_io_eo[63] ,
    \cb_2_0_io_eo[62] ,
    \cb_2_0_io_eo[61] ,
    \cb_2_0_io_eo[60] ,
    \cb_2_0_io_eo[59] ,
    \cb_2_0_io_eo[58] ,
    \cb_2_0_io_eo[57] ,
    \cb_2_0_io_eo[56] ,
    \cb_2_0_io_eo[55] ,
    \cb_2_0_io_eo[54] ,
    \cb_2_0_io_eo[53] ,
    \cb_2_0_io_eo[52] ,
    \cb_2_0_io_eo[51] ,
    \cb_2_0_io_eo[50] ,
    \cb_2_0_io_eo[49] ,
    \cb_2_0_io_eo[48] ,
    \cb_2_0_io_eo[47] ,
    \cb_2_0_io_eo[46] ,
    \cb_2_0_io_eo[45] ,
    \cb_2_0_io_eo[44] ,
    \cb_2_0_io_eo[43] ,
    \cb_2_0_io_eo[42] ,
    \cb_2_0_io_eo[41] ,
    \cb_2_0_io_eo[40] ,
    \cb_2_0_io_eo[39] ,
    \cb_2_0_io_eo[38] ,
    \cb_2_0_io_eo[37] ,
    \cb_2_0_io_eo[36] ,
    \cb_2_0_io_eo[35] ,
    \cb_2_0_io_eo[34] ,
    \cb_2_0_io_eo[33] ,
    \cb_2_0_io_eo[32] ,
    \cb_2_0_io_eo[31] ,
    \cb_2_0_io_eo[30] ,
    \cb_2_0_io_eo[29] ,
    \cb_2_0_io_eo[28] ,
    \cb_2_0_io_eo[27] ,
    \cb_2_0_io_eo[26] ,
    \cb_2_0_io_eo[25] ,
    \cb_2_0_io_eo[24] ,
    \cb_2_0_io_eo[23] ,
    \cb_2_0_io_eo[22] ,
    \cb_2_0_io_eo[21] ,
    \cb_2_0_io_eo[20] ,
    \cb_2_0_io_eo[19] ,
    \cb_2_0_io_eo[18] ,
    \cb_2_0_io_eo[17] ,
    \cb_2_0_io_eo[16] ,
    \cb_2_0_io_eo[15] ,
    \cb_2_0_io_eo[14] ,
    \cb_2_0_io_eo[13] ,
    \cb_2_0_io_eo[12] ,
    \cb_2_0_io_eo[11] ,
    \cb_2_0_io_eo[10] ,
    \cb_2_0_io_eo[9] ,
    \cb_2_0_io_eo[8] ,
    \cb_2_0_io_eo[7] ,
    \cb_2_0_io_eo[6] ,
    \cb_2_0_io_eo[5] ,
    \cb_2_0_io_eo[4] ,
    \cb_2_0_io_eo[3] ,
    \cb_2_0_io_eo[2] ,
    \cb_2_0_io_eo[1] ,
    \cb_2_0_io_eo[0] }),
    .io_i_0_in1({_NC129,
    _NC130,
    _NC131,
    _NC132,
    _NC133,
    _NC134,
    _NC135,
    _NC136}),
    .io_i_1_in1({_NC137,
    _NC138,
    _NC139,
    _NC140,
    _NC141,
    _NC142,
    _NC143,
    _NC144}),
    .io_i_2_in1({_NC145,
    _NC146,
    _NC147,
    _NC148,
    _NC149,
    _NC150,
    _NC151,
    _NC152}),
    .io_i_3_in1({_NC153,
    _NC154,
    _NC155,
    _NC156,
    _NC157,
    _NC158,
    _NC159,
    _NC160}),
    .io_i_4_in1({_NC161,
    _NC162,
    _NC163,
    _NC164,
    _NC165,
    _NC166,
    _NC167,
    _NC168}),
    .io_i_5_in1({_NC169,
    _NC170,
    _NC171,
    _NC172,
    _NC173,
    _NC174,
    _NC175,
    _NC176}),
    .io_i_6_in1({_NC177,
    _NC178,
    _NC179,
    _NC180,
    _NC181,
    _NC182,
    _NC183,
    _NC184}),
    .io_i_7_in1({_NC185,
    _NC186,
    _NC187,
    _NC188,
    _NC189,
    _NC190,
    _NC191,
    _NC192}),
    .io_o_0_out({\cb_2_0_io_o_0_out[7] ,
    \cb_2_0_io_o_0_out[6] ,
    \cb_2_0_io_o_0_out[5] ,
    \cb_2_0_io_o_0_out[4] ,
    \cb_2_0_io_o_0_out[3] ,
    \cb_2_0_io_o_0_out[2] ,
    \cb_2_0_io_o_0_out[1] ,
    \cb_2_0_io_o_0_out[0] }),
    .io_o_1_out({\cb_2_0_io_o_1_out[7] ,
    \cb_2_0_io_o_1_out[6] ,
    \cb_2_0_io_o_1_out[5] ,
    \cb_2_0_io_o_1_out[4] ,
    \cb_2_0_io_o_1_out[3] ,
    \cb_2_0_io_o_1_out[2] ,
    \cb_2_0_io_o_1_out[1] ,
    \cb_2_0_io_o_1_out[0] }),
    .io_o_2_out({\cb_2_0_io_o_2_out[7] ,
    \cb_2_0_io_o_2_out[6] ,
    \cb_2_0_io_o_2_out[5] ,
    \cb_2_0_io_o_2_out[4] ,
    \cb_2_0_io_o_2_out[3] ,
    \cb_2_0_io_o_2_out[2] ,
    \cb_2_0_io_o_2_out[1] ,
    \cb_2_0_io_o_2_out[0] }),
    .io_o_3_out({\cb_2_0_io_o_3_out[7] ,
    \cb_2_0_io_o_3_out[6] ,
    \cb_2_0_io_o_3_out[5] ,
    \cb_2_0_io_o_3_out[4] ,
    \cb_2_0_io_o_3_out[3] ,
    \cb_2_0_io_o_3_out[2] ,
    \cb_2_0_io_o_3_out[1] ,
    \cb_2_0_io_o_3_out[0] }),
    .io_o_4_out({\cb_2_0_io_o_4_out[7] ,
    \cb_2_0_io_o_4_out[6] ,
    \cb_2_0_io_o_4_out[5] ,
    \cb_2_0_io_o_4_out[4] ,
    \cb_2_0_io_o_4_out[3] ,
    \cb_2_0_io_o_4_out[2] ,
    \cb_2_0_io_o_4_out[1] ,
    \cb_2_0_io_o_4_out[0] }),
    .io_o_5_out({\cb_2_0_io_o_5_out[7] ,
    \cb_2_0_io_o_5_out[6] ,
    \cb_2_0_io_o_5_out[5] ,
    \cb_2_0_io_o_5_out[4] ,
    \cb_2_0_io_o_5_out[3] ,
    \cb_2_0_io_o_5_out[2] ,
    \cb_2_0_io_o_5_out[1] ,
    \cb_2_0_io_o_5_out[0] }),
    .io_o_6_out({\cb_2_0_io_o_6_out[7] ,
    \cb_2_0_io_o_6_out[6] ,
    \cb_2_0_io_o_6_out[5] ,
    \cb_2_0_io_o_6_out[4] ,
    \cb_2_0_io_o_6_out[3] ,
    \cb_2_0_io_o_6_out[2] ,
    \cb_2_0_io_o_6_out[1] ,
    \cb_2_0_io_o_6_out[0] }),
    .io_o_7_out({\cb_2_0_io_o_7_out[7] ,
    \cb_2_0_io_o_7_out[6] ,
    \cb_2_0_io_o_7_out[5] ,
    \cb_2_0_io_o_7_out[4] ,
    \cb_2_0_io_o_7_out[3] ,
    \cb_2_0_io_o_7_out[2] ,
    \cb_2_0_io_o_7_out[1] ,
    \cb_2_0_io_o_7_out[0] }),
    .io_wo({\cb_2_0_io_wo[63] ,
    \cb_2_0_io_wo[62] ,
    \cb_2_0_io_wo[61] ,
    \cb_2_0_io_wo[60] ,
    \cb_2_0_io_wo[59] ,
    \cb_2_0_io_wo[58] ,
    \cb_2_0_io_wo[57] ,
    \cb_2_0_io_wo[56] ,
    \cb_2_0_io_wo[55] ,
    \cb_2_0_io_wo[54] ,
    \cb_2_0_io_wo[53] ,
    \cb_2_0_io_wo[52] ,
    \cb_2_0_io_wo[51] ,
    \cb_2_0_io_wo[50] ,
    \cb_2_0_io_wo[49] ,
    \cb_2_0_io_wo[48] ,
    \cb_2_0_io_wo[47] ,
    \cb_2_0_io_wo[46] ,
    \cb_2_0_io_wo[45] ,
    \cb_2_0_io_wo[44] ,
    \cb_2_0_io_wo[43] ,
    \cb_2_0_io_wo[42] ,
    \cb_2_0_io_wo[41] ,
    \cb_2_0_io_wo[40] ,
    \cb_2_0_io_wo[39] ,
    \cb_2_0_io_wo[38] ,
    \cb_2_0_io_wo[37] ,
    \cb_2_0_io_wo[36] ,
    \cb_2_0_io_wo[35] ,
    \cb_2_0_io_wo[34] ,
    \cb_2_0_io_wo[33] ,
    \cb_2_0_io_wo[32] ,
    \cb_2_0_io_wo[31] ,
    \cb_2_0_io_wo[30] ,
    \cb_2_0_io_wo[29] ,
    \cb_2_0_io_wo[28] ,
    \cb_2_0_io_wo[27] ,
    \cb_2_0_io_wo[26] ,
    \cb_2_0_io_wo[25] ,
    \cb_2_0_io_wo[24] ,
    \cb_2_0_io_wo[23] ,
    \cb_2_0_io_wo[22] ,
    \cb_2_0_io_wo[21] ,
    \cb_2_0_io_wo[20] ,
    \cb_2_0_io_wo[19] ,
    \cb_2_0_io_wo[18] ,
    \cb_2_0_io_wo[17] ,
    \cb_2_0_io_wo[16] ,
    \cb_2_0_io_wo[15] ,
    \cb_2_0_io_wo[14] ,
    \cb_2_0_io_wo[13] ,
    \cb_2_0_io_wo[12] ,
    \cb_2_0_io_wo[11] ,
    \cb_2_0_io_wo[10] ,
    \cb_2_0_io_wo[9] ,
    \cb_2_0_io_wo[8] ,
    \cb_2_0_io_wo[7] ,
    \cb_2_0_io_wo[6] ,
    \cb_2_0_io_wo[5] ,
    \cb_2_0_io_wo[4] ,
    \cb_2_0_io_wo[3] ,
    \cb_2_0_io_wo[2] ,
    \cb_2_0_io_wo[1] ,
    \cb_2_0_io_wo[0] }));
 cic_block cb_2_1 (.io_cs_i(cb_2_1_io_cs_i),
    .io_i_0_ci(cb_2_0_io_o_0_co),
    .io_i_1_ci(cb_2_0_io_o_1_co),
    .io_i_2_ci(cb_2_0_io_o_2_co),
    .io_i_3_ci(cb_2_0_io_o_3_co),
    .io_i_4_ci(cb_2_0_io_o_4_co),
    .io_i_5_ci(cb_2_0_io_o_5_co),
    .io_i_6_ci(cb_2_0_io_o_6_co),
    .io_i_7_ci(cb_2_0_io_o_7_co),
    .io_o_0_co(cb_2_1_io_o_0_co),
    .io_o_1_co(cb_2_1_io_o_1_co),
    .io_o_2_co(cb_2_1_io_o_2_co),
    .io_o_3_co(cb_2_1_io_o_3_co),
    .io_o_4_co(cb_2_1_io_o_4_co),
    .io_o_5_co(cb_2_1_io_o_5_co),
    .io_o_6_co(cb_2_1_io_o_6_co),
    .io_o_7_co(cb_2_1_io_o_7_co),
    .io_vci(cb_2_0_io_vco),
    .io_vco(cb_2_1_io_vco),
    .io_vi(cb_2_1_io_vi),
    .io_we_i(cb_2_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_2_0_io_adr_i[1] ,
    \cb_2_0_io_adr_i[0] }),
    .io_dat_i({\cb_2_0_io_dat_i[15] ,
    \cb_2_0_io_dat_i[14] ,
    \cb_2_0_io_dat_i[13] ,
    \cb_2_0_io_dat_i[12] ,
    \cb_2_0_io_dat_i[11] ,
    \cb_2_0_io_dat_i[10] ,
    \cb_2_0_io_dat_i[9] ,
    \cb_2_0_io_dat_i[8] ,
    \cb_2_0_io_dat_i[7] ,
    \cb_2_0_io_dat_i[6] ,
    \cb_2_0_io_dat_i[5] ,
    \cb_2_0_io_dat_i[4] ,
    \cb_2_0_io_dat_i[3] ,
    \cb_2_0_io_dat_i[2] ,
    \cb_2_0_io_dat_i[1] ,
    \cb_2_0_io_dat_i[0] }),
    .io_dat_o({\cb_2_1_io_dat_o[15] ,
    \cb_2_1_io_dat_o[14] ,
    \cb_2_1_io_dat_o[13] ,
    \cb_2_1_io_dat_o[12] ,
    \cb_2_1_io_dat_o[11] ,
    \cb_2_1_io_dat_o[10] ,
    \cb_2_1_io_dat_o[9] ,
    \cb_2_1_io_dat_o[8] ,
    \cb_2_1_io_dat_o[7] ,
    \cb_2_1_io_dat_o[6] ,
    \cb_2_1_io_dat_o[5] ,
    \cb_2_1_io_dat_o[4] ,
    \cb_2_1_io_dat_o[3] ,
    \cb_2_1_io_dat_o[2] ,
    \cb_2_1_io_dat_o[1] ,
    \cb_2_1_io_dat_o[0] }),
    .io_eo({\cb_2_1_io_eo[63] ,
    \cb_2_1_io_eo[62] ,
    \cb_2_1_io_eo[61] ,
    \cb_2_1_io_eo[60] ,
    \cb_2_1_io_eo[59] ,
    \cb_2_1_io_eo[58] ,
    \cb_2_1_io_eo[57] ,
    \cb_2_1_io_eo[56] ,
    \cb_2_1_io_eo[55] ,
    \cb_2_1_io_eo[54] ,
    \cb_2_1_io_eo[53] ,
    \cb_2_1_io_eo[52] ,
    \cb_2_1_io_eo[51] ,
    \cb_2_1_io_eo[50] ,
    \cb_2_1_io_eo[49] ,
    \cb_2_1_io_eo[48] ,
    \cb_2_1_io_eo[47] ,
    \cb_2_1_io_eo[46] ,
    \cb_2_1_io_eo[45] ,
    \cb_2_1_io_eo[44] ,
    \cb_2_1_io_eo[43] ,
    \cb_2_1_io_eo[42] ,
    \cb_2_1_io_eo[41] ,
    \cb_2_1_io_eo[40] ,
    \cb_2_1_io_eo[39] ,
    \cb_2_1_io_eo[38] ,
    \cb_2_1_io_eo[37] ,
    \cb_2_1_io_eo[36] ,
    \cb_2_1_io_eo[35] ,
    \cb_2_1_io_eo[34] ,
    \cb_2_1_io_eo[33] ,
    \cb_2_1_io_eo[32] ,
    \cb_2_1_io_eo[31] ,
    \cb_2_1_io_eo[30] ,
    \cb_2_1_io_eo[29] ,
    \cb_2_1_io_eo[28] ,
    \cb_2_1_io_eo[27] ,
    \cb_2_1_io_eo[26] ,
    \cb_2_1_io_eo[25] ,
    \cb_2_1_io_eo[24] ,
    \cb_2_1_io_eo[23] ,
    \cb_2_1_io_eo[22] ,
    \cb_2_1_io_eo[21] ,
    \cb_2_1_io_eo[20] ,
    \cb_2_1_io_eo[19] ,
    \cb_2_1_io_eo[18] ,
    \cb_2_1_io_eo[17] ,
    \cb_2_1_io_eo[16] ,
    \cb_2_1_io_eo[15] ,
    \cb_2_1_io_eo[14] ,
    \cb_2_1_io_eo[13] ,
    \cb_2_1_io_eo[12] ,
    \cb_2_1_io_eo[11] ,
    \cb_2_1_io_eo[10] ,
    \cb_2_1_io_eo[9] ,
    \cb_2_1_io_eo[8] ,
    \cb_2_1_io_eo[7] ,
    \cb_2_1_io_eo[6] ,
    \cb_2_1_io_eo[5] ,
    \cb_2_1_io_eo[4] ,
    \cb_2_1_io_eo[3] ,
    \cb_2_1_io_eo[2] ,
    \cb_2_1_io_eo[1] ,
    \cb_2_1_io_eo[0] }),
    .io_i_0_in1({\cb_2_0_io_o_0_out[7] ,
    \cb_2_0_io_o_0_out[6] ,
    \cb_2_0_io_o_0_out[5] ,
    \cb_2_0_io_o_0_out[4] ,
    \cb_2_0_io_o_0_out[3] ,
    \cb_2_0_io_o_0_out[2] ,
    \cb_2_0_io_o_0_out[1] ,
    \cb_2_0_io_o_0_out[0] }),
    .io_i_1_in1({\cb_2_0_io_o_1_out[7] ,
    \cb_2_0_io_o_1_out[6] ,
    \cb_2_0_io_o_1_out[5] ,
    \cb_2_0_io_o_1_out[4] ,
    \cb_2_0_io_o_1_out[3] ,
    \cb_2_0_io_o_1_out[2] ,
    \cb_2_0_io_o_1_out[1] ,
    \cb_2_0_io_o_1_out[0] }),
    .io_i_2_in1({\cb_2_0_io_o_2_out[7] ,
    \cb_2_0_io_o_2_out[6] ,
    \cb_2_0_io_o_2_out[5] ,
    \cb_2_0_io_o_2_out[4] ,
    \cb_2_0_io_o_2_out[3] ,
    \cb_2_0_io_o_2_out[2] ,
    \cb_2_0_io_o_2_out[1] ,
    \cb_2_0_io_o_2_out[0] }),
    .io_i_3_in1({\cb_2_0_io_o_3_out[7] ,
    \cb_2_0_io_o_3_out[6] ,
    \cb_2_0_io_o_3_out[5] ,
    \cb_2_0_io_o_3_out[4] ,
    \cb_2_0_io_o_3_out[3] ,
    \cb_2_0_io_o_3_out[2] ,
    \cb_2_0_io_o_3_out[1] ,
    \cb_2_0_io_o_3_out[0] }),
    .io_i_4_in1({\cb_2_0_io_o_4_out[7] ,
    \cb_2_0_io_o_4_out[6] ,
    \cb_2_0_io_o_4_out[5] ,
    \cb_2_0_io_o_4_out[4] ,
    \cb_2_0_io_o_4_out[3] ,
    \cb_2_0_io_o_4_out[2] ,
    \cb_2_0_io_o_4_out[1] ,
    \cb_2_0_io_o_4_out[0] }),
    .io_i_5_in1({\cb_2_0_io_o_5_out[7] ,
    \cb_2_0_io_o_5_out[6] ,
    \cb_2_0_io_o_5_out[5] ,
    \cb_2_0_io_o_5_out[4] ,
    \cb_2_0_io_o_5_out[3] ,
    \cb_2_0_io_o_5_out[2] ,
    \cb_2_0_io_o_5_out[1] ,
    \cb_2_0_io_o_5_out[0] }),
    .io_i_6_in1({\cb_2_0_io_o_6_out[7] ,
    \cb_2_0_io_o_6_out[6] ,
    \cb_2_0_io_o_6_out[5] ,
    \cb_2_0_io_o_6_out[4] ,
    \cb_2_0_io_o_6_out[3] ,
    \cb_2_0_io_o_6_out[2] ,
    \cb_2_0_io_o_6_out[1] ,
    \cb_2_0_io_o_6_out[0] }),
    .io_i_7_in1({\cb_2_0_io_o_7_out[7] ,
    \cb_2_0_io_o_7_out[6] ,
    \cb_2_0_io_o_7_out[5] ,
    \cb_2_0_io_o_7_out[4] ,
    \cb_2_0_io_o_7_out[3] ,
    \cb_2_0_io_o_7_out[2] ,
    \cb_2_0_io_o_7_out[1] ,
    \cb_2_0_io_o_7_out[0] }),
    .io_o_0_out({\cb_2_1_io_o_0_out[7] ,
    \cb_2_1_io_o_0_out[6] ,
    \cb_2_1_io_o_0_out[5] ,
    \cb_2_1_io_o_0_out[4] ,
    \cb_2_1_io_o_0_out[3] ,
    \cb_2_1_io_o_0_out[2] ,
    \cb_2_1_io_o_0_out[1] ,
    \cb_2_1_io_o_0_out[0] }),
    .io_o_1_out({\cb_2_1_io_o_1_out[7] ,
    \cb_2_1_io_o_1_out[6] ,
    \cb_2_1_io_o_1_out[5] ,
    \cb_2_1_io_o_1_out[4] ,
    \cb_2_1_io_o_1_out[3] ,
    \cb_2_1_io_o_1_out[2] ,
    \cb_2_1_io_o_1_out[1] ,
    \cb_2_1_io_o_1_out[0] }),
    .io_o_2_out({\cb_2_1_io_o_2_out[7] ,
    \cb_2_1_io_o_2_out[6] ,
    \cb_2_1_io_o_2_out[5] ,
    \cb_2_1_io_o_2_out[4] ,
    \cb_2_1_io_o_2_out[3] ,
    \cb_2_1_io_o_2_out[2] ,
    \cb_2_1_io_o_2_out[1] ,
    \cb_2_1_io_o_2_out[0] }),
    .io_o_3_out({\cb_2_1_io_o_3_out[7] ,
    \cb_2_1_io_o_3_out[6] ,
    \cb_2_1_io_o_3_out[5] ,
    \cb_2_1_io_o_3_out[4] ,
    \cb_2_1_io_o_3_out[3] ,
    \cb_2_1_io_o_3_out[2] ,
    \cb_2_1_io_o_3_out[1] ,
    \cb_2_1_io_o_3_out[0] }),
    .io_o_4_out({\cb_2_1_io_o_4_out[7] ,
    \cb_2_1_io_o_4_out[6] ,
    \cb_2_1_io_o_4_out[5] ,
    \cb_2_1_io_o_4_out[4] ,
    \cb_2_1_io_o_4_out[3] ,
    \cb_2_1_io_o_4_out[2] ,
    \cb_2_1_io_o_4_out[1] ,
    \cb_2_1_io_o_4_out[0] }),
    .io_o_5_out({\cb_2_1_io_o_5_out[7] ,
    \cb_2_1_io_o_5_out[6] ,
    \cb_2_1_io_o_5_out[5] ,
    \cb_2_1_io_o_5_out[4] ,
    \cb_2_1_io_o_5_out[3] ,
    \cb_2_1_io_o_5_out[2] ,
    \cb_2_1_io_o_5_out[1] ,
    \cb_2_1_io_o_5_out[0] }),
    .io_o_6_out({\cb_2_1_io_o_6_out[7] ,
    \cb_2_1_io_o_6_out[6] ,
    \cb_2_1_io_o_6_out[5] ,
    \cb_2_1_io_o_6_out[4] ,
    \cb_2_1_io_o_6_out[3] ,
    \cb_2_1_io_o_6_out[2] ,
    \cb_2_1_io_o_6_out[1] ,
    \cb_2_1_io_o_6_out[0] }),
    .io_o_7_out({\cb_2_1_io_o_7_out[7] ,
    \cb_2_1_io_o_7_out[6] ,
    \cb_2_1_io_o_7_out[5] ,
    \cb_2_1_io_o_7_out[4] ,
    \cb_2_1_io_o_7_out[3] ,
    \cb_2_1_io_o_7_out[2] ,
    \cb_2_1_io_o_7_out[1] ,
    \cb_2_1_io_o_7_out[0] }),
    .io_wo({\cb_2_0_io_eo[63] ,
    \cb_2_0_io_eo[62] ,
    \cb_2_0_io_eo[61] ,
    \cb_2_0_io_eo[60] ,
    \cb_2_0_io_eo[59] ,
    \cb_2_0_io_eo[58] ,
    \cb_2_0_io_eo[57] ,
    \cb_2_0_io_eo[56] ,
    \cb_2_0_io_eo[55] ,
    \cb_2_0_io_eo[54] ,
    \cb_2_0_io_eo[53] ,
    \cb_2_0_io_eo[52] ,
    \cb_2_0_io_eo[51] ,
    \cb_2_0_io_eo[50] ,
    \cb_2_0_io_eo[49] ,
    \cb_2_0_io_eo[48] ,
    \cb_2_0_io_eo[47] ,
    \cb_2_0_io_eo[46] ,
    \cb_2_0_io_eo[45] ,
    \cb_2_0_io_eo[44] ,
    \cb_2_0_io_eo[43] ,
    \cb_2_0_io_eo[42] ,
    \cb_2_0_io_eo[41] ,
    \cb_2_0_io_eo[40] ,
    \cb_2_0_io_eo[39] ,
    \cb_2_0_io_eo[38] ,
    \cb_2_0_io_eo[37] ,
    \cb_2_0_io_eo[36] ,
    \cb_2_0_io_eo[35] ,
    \cb_2_0_io_eo[34] ,
    \cb_2_0_io_eo[33] ,
    \cb_2_0_io_eo[32] ,
    \cb_2_0_io_eo[31] ,
    \cb_2_0_io_eo[30] ,
    \cb_2_0_io_eo[29] ,
    \cb_2_0_io_eo[28] ,
    \cb_2_0_io_eo[27] ,
    \cb_2_0_io_eo[26] ,
    \cb_2_0_io_eo[25] ,
    \cb_2_0_io_eo[24] ,
    \cb_2_0_io_eo[23] ,
    \cb_2_0_io_eo[22] ,
    \cb_2_0_io_eo[21] ,
    \cb_2_0_io_eo[20] ,
    \cb_2_0_io_eo[19] ,
    \cb_2_0_io_eo[18] ,
    \cb_2_0_io_eo[17] ,
    \cb_2_0_io_eo[16] ,
    \cb_2_0_io_eo[15] ,
    \cb_2_0_io_eo[14] ,
    \cb_2_0_io_eo[13] ,
    \cb_2_0_io_eo[12] ,
    \cb_2_0_io_eo[11] ,
    \cb_2_0_io_eo[10] ,
    \cb_2_0_io_eo[9] ,
    \cb_2_0_io_eo[8] ,
    \cb_2_0_io_eo[7] ,
    \cb_2_0_io_eo[6] ,
    \cb_2_0_io_eo[5] ,
    \cb_2_0_io_eo[4] ,
    \cb_2_0_io_eo[3] ,
    \cb_2_0_io_eo[2] ,
    \cb_2_0_io_eo[1] ,
    \cb_2_0_io_eo[0] }));
 cic_block cb_2_10 (.io_cs_i(cb_2_10_io_cs_i),
    .io_i_0_ci(cb_2_10_io_i_0_ci),
    .io_i_1_ci(cb_2_10_io_i_1_ci),
    .io_i_2_ci(cb_2_10_io_i_2_ci),
    .io_i_3_ci(cb_2_10_io_i_3_ci),
    .io_i_4_ci(cb_2_10_io_i_4_ci),
    .io_i_5_ci(cb_2_10_io_i_5_ci),
    .io_i_6_ci(cb_2_10_io_i_6_ci),
    .io_i_7_ci(cb_2_10_io_i_7_ci),
    .io_o_0_co(cb_2_10_io_o_0_co),
    .io_o_1_co(cb_2_10_io_o_1_co),
    .io_o_2_co(cb_2_10_io_o_2_co),
    .io_o_3_co(cb_2_10_io_o_3_co),
    .io_o_4_co(cb_2_10_io_o_4_co),
    .io_o_5_co(cb_2_10_io_o_5_co),
    .io_o_6_co(cb_2_10_io_o_6_co),
    .io_o_7_co(cb_2_10_io_o_7_co),
    .io_vci(cb_2_10_io_vci),
    .io_vco(cb_2_10_io_vco),
    .io_vi(cb_2_10_io_vi),
    .io_we_i(cb_2_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_2_0_io_adr_i[1] ,
    \cb_2_0_io_adr_i[0] }),
    .io_dat_i({\cb_2_0_io_dat_i[15] ,
    \cb_2_0_io_dat_i[14] ,
    \cb_2_0_io_dat_i[13] ,
    \cb_2_0_io_dat_i[12] ,
    \cb_2_0_io_dat_i[11] ,
    \cb_2_0_io_dat_i[10] ,
    \cb_2_0_io_dat_i[9] ,
    \cb_2_0_io_dat_i[8] ,
    \cb_2_0_io_dat_i[7] ,
    \cb_2_0_io_dat_i[6] ,
    \cb_2_0_io_dat_i[5] ,
    \cb_2_0_io_dat_i[4] ,
    \cb_2_0_io_dat_i[3] ,
    \cb_2_0_io_dat_i[2] ,
    \cb_2_0_io_dat_i[1] ,
    \cb_2_0_io_dat_i[0] }),
    .io_dat_o({\cb_2_10_io_dat_o[15] ,
    \cb_2_10_io_dat_o[14] ,
    \cb_2_10_io_dat_o[13] ,
    \cb_2_10_io_dat_o[12] ,
    \cb_2_10_io_dat_o[11] ,
    \cb_2_10_io_dat_o[10] ,
    \cb_2_10_io_dat_o[9] ,
    \cb_2_10_io_dat_o[8] ,
    \cb_2_10_io_dat_o[7] ,
    \cb_2_10_io_dat_o[6] ,
    \cb_2_10_io_dat_o[5] ,
    \cb_2_10_io_dat_o[4] ,
    \cb_2_10_io_dat_o[3] ,
    \cb_2_10_io_dat_o[2] ,
    \cb_2_10_io_dat_o[1] ,
    \cb_2_10_io_dat_o[0] }),
    .io_eo({\_T_66[31] ,
    \_T_66[30] ,
    \_T_66[29] ,
    \_T_66[28] ,
    \_T_66[27] ,
    \_T_66[26] ,
    \_T_66[25] ,
    \_T_66[24] ,
    \_T_66[23] ,
    \_T_66[22] ,
    \_T_66[21] ,
    \_T_66[20] ,
    \_T_66[19] ,
    \_T_66[18] ,
    \_T_66[17] ,
    \_T_66[16] ,
    \_T_66[15] ,
    \_T_66[14] ,
    \_T_66[13] ,
    \_T_66[12] ,
    \_T_66[11] ,
    \_T_66[10] ,
    \_T_66[9] ,
    \_T_66[8] ,
    \_T_66[7] ,
    \_T_66[6] ,
    \_T_66[5] ,
    \_T_66[4] ,
    \_T_66[3] ,
    \_T_66[2] ,
    \_T_66[1] ,
    \_T_66[0] ,
    \_T_63[31] ,
    \_T_63[30] ,
    \_T_63[29] ,
    \_T_63[28] ,
    \_T_63[27] ,
    \_T_63[26] ,
    \_T_63[25] ,
    \_T_63[24] ,
    \_T_63[23] ,
    \_T_63[22] ,
    \_T_63[21] ,
    \_T_63[20] ,
    \_T_63[19] ,
    \_T_63[18] ,
    \_T_63[17] ,
    \_T_63[16] ,
    \_T_63[15] ,
    \_T_63[14] ,
    \_T_63[13] ,
    \_T_63[12] ,
    \_T_63[11] ,
    \_T_63[10] ,
    \_T_63[9] ,
    \_T_63[8] ,
    \_T_63[7] ,
    \_T_63[6] ,
    \_T_63[5] ,
    \_T_63[4] ,
    \_T_63[3] ,
    \_T_63[2] ,
    \_T_63[1] ,
    \_T_63[0] }),
    .io_i_0_in1({\cb_2_10_io_i_0_in1[7] ,
    \cb_2_10_io_i_0_in1[6] ,
    \cb_2_10_io_i_0_in1[5] ,
    \cb_2_10_io_i_0_in1[4] ,
    \cb_2_10_io_i_0_in1[3] ,
    \cb_2_10_io_i_0_in1[2] ,
    \cb_2_10_io_i_0_in1[1] ,
    \cb_2_10_io_i_0_in1[0] }),
    .io_i_1_in1({\cb_2_10_io_i_1_in1[7] ,
    \cb_2_10_io_i_1_in1[6] ,
    \cb_2_10_io_i_1_in1[5] ,
    \cb_2_10_io_i_1_in1[4] ,
    \cb_2_10_io_i_1_in1[3] ,
    \cb_2_10_io_i_1_in1[2] ,
    \cb_2_10_io_i_1_in1[1] ,
    \cb_2_10_io_i_1_in1[0] }),
    .io_i_2_in1({\cb_2_10_io_i_2_in1[7] ,
    \cb_2_10_io_i_2_in1[6] ,
    \cb_2_10_io_i_2_in1[5] ,
    \cb_2_10_io_i_2_in1[4] ,
    \cb_2_10_io_i_2_in1[3] ,
    \cb_2_10_io_i_2_in1[2] ,
    \cb_2_10_io_i_2_in1[1] ,
    \cb_2_10_io_i_2_in1[0] }),
    .io_i_3_in1({\cb_2_10_io_i_3_in1[7] ,
    \cb_2_10_io_i_3_in1[6] ,
    \cb_2_10_io_i_3_in1[5] ,
    \cb_2_10_io_i_3_in1[4] ,
    \cb_2_10_io_i_3_in1[3] ,
    \cb_2_10_io_i_3_in1[2] ,
    \cb_2_10_io_i_3_in1[1] ,
    \cb_2_10_io_i_3_in1[0] }),
    .io_i_4_in1({\cb_2_10_io_i_4_in1[7] ,
    \cb_2_10_io_i_4_in1[6] ,
    \cb_2_10_io_i_4_in1[5] ,
    \cb_2_10_io_i_4_in1[4] ,
    \cb_2_10_io_i_4_in1[3] ,
    \cb_2_10_io_i_4_in1[2] ,
    \cb_2_10_io_i_4_in1[1] ,
    \cb_2_10_io_i_4_in1[0] }),
    .io_i_5_in1({\cb_2_10_io_i_5_in1[7] ,
    \cb_2_10_io_i_5_in1[6] ,
    \cb_2_10_io_i_5_in1[5] ,
    \cb_2_10_io_i_5_in1[4] ,
    \cb_2_10_io_i_5_in1[3] ,
    \cb_2_10_io_i_5_in1[2] ,
    \cb_2_10_io_i_5_in1[1] ,
    \cb_2_10_io_i_5_in1[0] }),
    .io_i_6_in1({\cb_2_10_io_i_6_in1[7] ,
    \cb_2_10_io_i_6_in1[6] ,
    \cb_2_10_io_i_6_in1[5] ,
    \cb_2_10_io_i_6_in1[4] ,
    \cb_2_10_io_i_6_in1[3] ,
    \cb_2_10_io_i_6_in1[2] ,
    \cb_2_10_io_i_6_in1[1] ,
    \cb_2_10_io_i_6_in1[0] }),
    .io_i_7_in1({\cb_2_10_io_i_7_in1[7] ,
    \cb_2_10_io_i_7_in1[6] ,
    \cb_2_10_io_i_7_in1[5] ,
    \cb_2_10_io_i_7_in1[4] ,
    \cb_2_10_io_i_7_in1[3] ,
    \cb_2_10_io_i_7_in1[2] ,
    \cb_2_10_io_i_7_in1[1] ,
    \cb_2_10_io_i_7_in1[0] }),
    .io_o_0_out({\_T_63[7] ,
    \_T_63[6] ,
    \_T_63[5] ,
    \_T_63[4] ,
    \_T_63[3] ,
    \_T_63[2] ,
    \_T_63[1] ,
    \_T_63[0] }),
    .io_o_1_out({\_T_63[15] ,
    \_T_63[14] ,
    \_T_63[13] ,
    \_T_63[12] ,
    \_T_63[11] ,
    \_T_63[10] ,
    \_T_63[9] ,
    \_T_63[8] }),
    .io_o_2_out({\_T_63[23] ,
    \_T_63[22] ,
    \_T_63[21] ,
    \_T_63[20] ,
    \_T_63[19] ,
    \_T_63[18] ,
    \_T_63[17] ,
    \_T_63[16] }),
    .io_o_3_out({\_T_63[31] ,
    \_T_63[30] ,
    \_T_63[29] ,
    \_T_63[28] ,
    \_T_63[27] ,
    \_T_63[26] ,
    \_T_63[25] ,
    \_T_63[24] }),
    .io_o_4_out({\_T_66[7] ,
    \_T_66[6] ,
    \_T_66[5] ,
    \_T_66[4] ,
    \_T_66[3] ,
    \_T_66[2] ,
    \_T_66[1] ,
    \_T_66[0] }),
    .io_o_5_out({\_T_66[15] ,
    \_T_66[14] ,
    \_T_66[13] ,
    \_T_66[12] ,
    \_T_66[11] ,
    \_T_66[10] ,
    \_T_66[9] ,
    \_T_66[8] }),
    .io_o_6_out({\_T_66[23] ,
    \_T_66[22] ,
    \_T_66[21] ,
    \_T_66[20] ,
    \_T_66[19] ,
    \_T_66[18] ,
    \_T_66[17] ,
    \_T_66[16] }),
    .io_o_7_out({\_T_66[31] ,
    \_T_66[30] ,
    \_T_66[29] ,
    \_T_66[28] ,
    \_T_66[27] ,
    \_T_66[26] ,
    \_T_66[25] ,
    \_T_66[24] }),
    .io_wo({\cb_2_10_io_wo[63] ,
    \cb_2_10_io_wo[62] ,
    \cb_2_10_io_wo[61] ,
    \cb_2_10_io_wo[60] ,
    \cb_2_10_io_wo[59] ,
    \cb_2_10_io_wo[58] ,
    \cb_2_10_io_wo[57] ,
    \cb_2_10_io_wo[56] ,
    \cb_2_10_io_wo[55] ,
    \cb_2_10_io_wo[54] ,
    \cb_2_10_io_wo[53] ,
    \cb_2_10_io_wo[52] ,
    \cb_2_10_io_wo[51] ,
    \cb_2_10_io_wo[50] ,
    \cb_2_10_io_wo[49] ,
    \cb_2_10_io_wo[48] ,
    \cb_2_10_io_wo[47] ,
    \cb_2_10_io_wo[46] ,
    \cb_2_10_io_wo[45] ,
    \cb_2_10_io_wo[44] ,
    \cb_2_10_io_wo[43] ,
    \cb_2_10_io_wo[42] ,
    \cb_2_10_io_wo[41] ,
    \cb_2_10_io_wo[40] ,
    \cb_2_10_io_wo[39] ,
    \cb_2_10_io_wo[38] ,
    \cb_2_10_io_wo[37] ,
    \cb_2_10_io_wo[36] ,
    \cb_2_10_io_wo[35] ,
    \cb_2_10_io_wo[34] ,
    \cb_2_10_io_wo[33] ,
    \cb_2_10_io_wo[32] ,
    \cb_2_10_io_wo[31] ,
    \cb_2_10_io_wo[30] ,
    \cb_2_10_io_wo[29] ,
    \cb_2_10_io_wo[28] ,
    \cb_2_10_io_wo[27] ,
    \cb_2_10_io_wo[26] ,
    \cb_2_10_io_wo[25] ,
    \cb_2_10_io_wo[24] ,
    \cb_2_10_io_wo[23] ,
    \cb_2_10_io_wo[22] ,
    \cb_2_10_io_wo[21] ,
    \cb_2_10_io_wo[20] ,
    \cb_2_10_io_wo[19] ,
    \cb_2_10_io_wo[18] ,
    \cb_2_10_io_wo[17] ,
    \cb_2_10_io_wo[16] ,
    \cb_2_10_io_wo[15] ,
    \cb_2_10_io_wo[14] ,
    \cb_2_10_io_wo[13] ,
    \cb_2_10_io_wo[12] ,
    \cb_2_10_io_wo[11] ,
    \cb_2_10_io_wo[10] ,
    \cb_2_10_io_wo[9] ,
    \cb_2_10_io_wo[8] ,
    \cb_2_10_io_wo[7] ,
    \cb_2_10_io_wo[6] ,
    \cb_2_10_io_wo[5] ,
    \cb_2_10_io_wo[4] ,
    \cb_2_10_io_wo[3] ,
    \cb_2_10_io_wo[2] ,
    \cb_2_10_io_wo[1] ,
    \cb_2_10_io_wo[0] }));
 cic_block cb_2_2 (.io_cs_i(cb_2_2_io_cs_i),
    .io_i_0_ci(cb_2_1_io_o_0_co),
    .io_i_1_ci(cb_2_1_io_o_1_co),
    .io_i_2_ci(cb_2_1_io_o_2_co),
    .io_i_3_ci(cb_2_1_io_o_3_co),
    .io_i_4_ci(cb_2_1_io_o_4_co),
    .io_i_5_ci(cb_2_1_io_o_5_co),
    .io_i_6_ci(cb_2_1_io_o_6_co),
    .io_i_7_ci(cb_2_1_io_o_7_co),
    .io_o_0_co(cb_2_2_io_o_0_co),
    .io_o_1_co(cb_2_2_io_o_1_co),
    .io_o_2_co(cb_2_2_io_o_2_co),
    .io_o_3_co(cb_2_2_io_o_3_co),
    .io_o_4_co(cb_2_2_io_o_4_co),
    .io_o_5_co(cb_2_2_io_o_5_co),
    .io_o_6_co(cb_2_2_io_o_6_co),
    .io_o_7_co(cb_2_2_io_o_7_co),
    .io_vci(cb_2_1_io_vco),
    .io_vco(cb_2_2_io_vco),
    .io_vi(cb_2_2_io_vi),
    .io_we_i(cb_2_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_2_0_io_adr_i[1] ,
    \cb_2_0_io_adr_i[0] }),
    .io_dat_i({\cb_2_0_io_dat_i[15] ,
    \cb_2_0_io_dat_i[14] ,
    \cb_2_0_io_dat_i[13] ,
    \cb_2_0_io_dat_i[12] ,
    \cb_2_0_io_dat_i[11] ,
    \cb_2_0_io_dat_i[10] ,
    \cb_2_0_io_dat_i[9] ,
    \cb_2_0_io_dat_i[8] ,
    \cb_2_0_io_dat_i[7] ,
    \cb_2_0_io_dat_i[6] ,
    \cb_2_0_io_dat_i[5] ,
    \cb_2_0_io_dat_i[4] ,
    \cb_2_0_io_dat_i[3] ,
    \cb_2_0_io_dat_i[2] ,
    \cb_2_0_io_dat_i[1] ,
    \cb_2_0_io_dat_i[0] }),
    .io_dat_o({\cb_2_2_io_dat_o[15] ,
    \cb_2_2_io_dat_o[14] ,
    \cb_2_2_io_dat_o[13] ,
    \cb_2_2_io_dat_o[12] ,
    \cb_2_2_io_dat_o[11] ,
    \cb_2_2_io_dat_o[10] ,
    \cb_2_2_io_dat_o[9] ,
    \cb_2_2_io_dat_o[8] ,
    \cb_2_2_io_dat_o[7] ,
    \cb_2_2_io_dat_o[6] ,
    \cb_2_2_io_dat_o[5] ,
    \cb_2_2_io_dat_o[4] ,
    \cb_2_2_io_dat_o[3] ,
    \cb_2_2_io_dat_o[2] ,
    \cb_2_2_io_dat_o[1] ,
    \cb_2_2_io_dat_o[0] }),
    .io_eo({\cb_2_2_io_eo[63] ,
    \cb_2_2_io_eo[62] ,
    \cb_2_2_io_eo[61] ,
    \cb_2_2_io_eo[60] ,
    \cb_2_2_io_eo[59] ,
    \cb_2_2_io_eo[58] ,
    \cb_2_2_io_eo[57] ,
    \cb_2_2_io_eo[56] ,
    \cb_2_2_io_eo[55] ,
    \cb_2_2_io_eo[54] ,
    \cb_2_2_io_eo[53] ,
    \cb_2_2_io_eo[52] ,
    \cb_2_2_io_eo[51] ,
    \cb_2_2_io_eo[50] ,
    \cb_2_2_io_eo[49] ,
    \cb_2_2_io_eo[48] ,
    \cb_2_2_io_eo[47] ,
    \cb_2_2_io_eo[46] ,
    \cb_2_2_io_eo[45] ,
    \cb_2_2_io_eo[44] ,
    \cb_2_2_io_eo[43] ,
    \cb_2_2_io_eo[42] ,
    \cb_2_2_io_eo[41] ,
    \cb_2_2_io_eo[40] ,
    \cb_2_2_io_eo[39] ,
    \cb_2_2_io_eo[38] ,
    \cb_2_2_io_eo[37] ,
    \cb_2_2_io_eo[36] ,
    \cb_2_2_io_eo[35] ,
    \cb_2_2_io_eo[34] ,
    \cb_2_2_io_eo[33] ,
    \cb_2_2_io_eo[32] ,
    \cb_2_2_io_eo[31] ,
    \cb_2_2_io_eo[30] ,
    \cb_2_2_io_eo[29] ,
    \cb_2_2_io_eo[28] ,
    \cb_2_2_io_eo[27] ,
    \cb_2_2_io_eo[26] ,
    \cb_2_2_io_eo[25] ,
    \cb_2_2_io_eo[24] ,
    \cb_2_2_io_eo[23] ,
    \cb_2_2_io_eo[22] ,
    \cb_2_2_io_eo[21] ,
    \cb_2_2_io_eo[20] ,
    \cb_2_2_io_eo[19] ,
    \cb_2_2_io_eo[18] ,
    \cb_2_2_io_eo[17] ,
    \cb_2_2_io_eo[16] ,
    \cb_2_2_io_eo[15] ,
    \cb_2_2_io_eo[14] ,
    \cb_2_2_io_eo[13] ,
    \cb_2_2_io_eo[12] ,
    \cb_2_2_io_eo[11] ,
    \cb_2_2_io_eo[10] ,
    \cb_2_2_io_eo[9] ,
    \cb_2_2_io_eo[8] ,
    \cb_2_2_io_eo[7] ,
    \cb_2_2_io_eo[6] ,
    \cb_2_2_io_eo[5] ,
    \cb_2_2_io_eo[4] ,
    \cb_2_2_io_eo[3] ,
    \cb_2_2_io_eo[2] ,
    \cb_2_2_io_eo[1] ,
    \cb_2_2_io_eo[0] }),
    .io_i_0_in1({\cb_2_1_io_o_0_out[7] ,
    \cb_2_1_io_o_0_out[6] ,
    \cb_2_1_io_o_0_out[5] ,
    \cb_2_1_io_o_0_out[4] ,
    \cb_2_1_io_o_0_out[3] ,
    \cb_2_1_io_o_0_out[2] ,
    \cb_2_1_io_o_0_out[1] ,
    \cb_2_1_io_o_0_out[0] }),
    .io_i_1_in1({\cb_2_1_io_o_1_out[7] ,
    \cb_2_1_io_o_1_out[6] ,
    \cb_2_1_io_o_1_out[5] ,
    \cb_2_1_io_o_1_out[4] ,
    \cb_2_1_io_o_1_out[3] ,
    \cb_2_1_io_o_1_out[2] ,
    \cb_2_1_io_o_1_out[1] ,
    \cb_2_1_io_o_1_out[0] }),
    .io_i_2_in1({\cb_2_1_io_o_2_out[7] ,
    \cb_2_1_io_o_2_out[6] ,
    \cb_2_1_io_o_2_out[5] ,
    \cb_2_1_io_o_2_out[4] ,
    \cb_2_1_io_o_2_out[3] ,
    \cb_2_1_io_o_2_out[2] ,
    \cb_2_1_io_o_2_out[1] ,
    \cb_2_1_io_o_2_out[0] }),
    .io_i_3_in1({\cb_2_1_io_o_3_out[7] ,
    \cb_2_1_io_o_3_out[6] ,
    \cb_2_1_io_o_3_out[5] ,
    \cb_2_1_io_o_3_out[4] ,
    \cb_2_1_io_o_3_out[3] ,
    \cb_2_1_io_o_3_out[2] ,
    \cb_2_1_io_o_3_out[1] ,
    \cb_2_1_io_o_3_out[0] }),
    .io_i_4_in1({\cb_2_1_io_o_4_out[7] ,
    \cb_2_1_io_o_4_out[6] ,
    \cb_2_1_io_o_4_out[5] ,
    \cb_2_1_io_o_4_out[4] ,
    \cb_2_1_io_o_4_out[3] ,
    \cb_2_1_io_o_4_out[2] ,
    \cb_2_1_io_o_4_out[1] ,
    \cb_2_1_io_o_4_out[0] }),
    .io_i_5_in1({\cb_2_1_io_o_5_out[7] ,
    \cb_2_1_io_o_5_out[6] ,
    \cb_2_1_io_o_5_out[5] ,
    \cb_2_1_io_o_5_out[4] ,
    \cb_2_1_io_o_5_out[3] ,
    \cb_2_1_io_o_5_out[2] ,
    \cb_2_1_io_o_5_out[1] ,
    \cb_2_1_io_o_5_out[0] }),
    .io_i_6_in1({\cb_2_1_io_o_6_out[7] ,
    \cb_2_1_io_o_6_out[6] ,
    \cb_2_1_io_o_6_out[5] ,
    \cb_2_1_io_o_6_out[4] ,
    \cb_2_1_io_o_6_out[3] ,
    \cb_2_1_io_o_6_out[2] ,
    \cb_2_1_io_o_6_out[1] ,
    \cb_2_1_io_o_6_out[0] }),
    .io_i_7_in1({\cb_2_1_io_o_7_out[7] ,
    \cb_2_1_io_o_7_out[6] ,
    \cb_2_1_io_o_7_out[5] ,
    \cb_2_1_io_o_7_out[4] ,
    \cb_2_1_io_o_7_out[3] ,
    \cb_2_1_io_o_7_out[2] ,
    \cb_2_1_io_o_7_out[1] ,
    \cb_2_1_io_o_7_out[0] }),
    .io_o_0_out({\cb_2_2_io_o_0_out[7] ,
    \cb_2_2_io_o_0_out[6] ,
    \cb_2_2_io_o_0_out[5] ,
    \cb_2_2_io_o_0_out[4] ,
    \cb_2_2_io_o_0_out[3] ,
    \cb_2_2_io_o_0_out[2] ,
    \cb_2_2_io_o_0_out[1] ,
    \cb_2_2_io_o_0_out[0] }),
    .io_o_1_out({\cb_2_2_io_o_1_out[7] ,
    \cb_2_2_io_o_1_out[6] ,
    \cb_2_2_io_o_1_out[5] ,
    \cb_2_2_io_o_1_out[4] ,
    \cb_2_2_io_o_1_out[3] ,
    \cb_2_2_io_o_1_out[2] ,
    \cb_2_2_io_o_1_out[1] ,
    \cb_2_2_io_o_1_out[0] }),
    .io_o_2_out({\cb_2_2_io_o_2_out[7] ,
    \cb_2_2_io_o_2_out[6] ,
    \cb_2_2_io_o_2_out[5] ,
    \cb_2_2_io_o_2_out[4] ,
    \cb_2_2_io_o_2_out[3] ,
    \cb_2_2_io_o_2_out[2] ,
    \cb_2_2_io_o_2_out[1] ,
    \cb_2_2_io_o_2_out[0] }),
    .io_o_3_out({\cb_2_2_io_o_3_out[7] ,
    \cb_2_2_io_o_3_out[6] ,
    \cb_2_2_io_o_3_out[5] ,
    \cb_2_2_io_o_3_out[4] ,
    \cb_2_2_io_o_3_out[3] ,
    \cb_2_2_io_o_3_out[2] ,
    \cb_2_2_io_o_3_out[1] ,
    \cb_2_2_io_o_3_out[0] }),
    .io_o_4_out({\cb_2_2_io_o_4_out[7] ,
    \cb_2_2_io_o_4_out[6] ,
    \cb_2_2_io_o_4_out[5] ,
    \cb_2_2_io_o_4_out[4] ,
    \cb_2_2_io_o_4_out[3] ,
    \cb_2_2_io_o_4_out[2] ,
    \cb_2_2_io_o_4_out[1] ,
    \cb_2_2_io_o_4_out[0] }),
    .io_o_5_out({\cb_2_2_io_o_5_out[7] ,
    \cb_2_2_io_o_5_out[6] ,
    \cb_2_2_io_o_5_out[5] ,
    \cb_2_2_io_o_5_out[4] ,
    \cb_2_2_io_o_5_out[3] ,
    \cb_2_2_io_o_5_out[2] ,
    \cb_2_2_io_o_5_out[1] ,
    \cb_2_2_io_o_5_out[0] }),
    .io_o_6_out({\cb_2_2_io_o_6_out[7] ,
    \cb_2_2_io_o_6_out[6] ,
    \cb_2_2_io_o_6_out[5] ,
    \cb_2_2_io_o_6_out[4] ,
    \cb_2_2_io_o_6_out[3] ,
    \cb_2_2_io_o_6_out[2] ,
    \cb_2_2_io_o_6_out[1] ,
    \cb_2_2_io_o_6_out[0] }),
    .io_o_7_out({\cb_2_2_io_o_7_out[7] ,
    \cb_2_2_io_o_7_out[6] ,
    \cb_2_2_io_o_7_out[5] ,
    \cb_2_2_io_o_7_out[4] ,
    \cb_2_2_io_o_7_out[3] ,
    \cb_2_2_io_o_7_out[2] ,
    \cb_2_2_io_o_7_out[1] ,
    \cb_2_2_io_o_7_out[0] }),
    .io_wo({\cb_2_1_io_eo[63] ,
    \cb_2_1_io_eo[62] ,
    \cb_2_1_io_eo[61] ,
    \cb_2_1_io_eo[60] ,
    \cb_2_1_io_eo[59] ,
    \cb_2_1_io_eo[58] ,
    \cb_2_1_io_eo[57] ,
    \cb_2_1_io_eo[56] ,
    \cb_2_1_io_eo[55] ,
    \cb_2_1_io_eo[54] ,
    \cb_2_1_io_eo[53] ,
    \cb_2_1_io_eo[52] ,
    \cb_2_1_io_eo[51] ,
    \cb_2_1_io_eo[50] ,
    \cb_2_1_io_eo[49] ,
    \cb_2_1_io_eo[48] ,
    \cb_2_1_io_eo[47] ,
    \cb_2_1_io_eo[46] ,
    \cb_2_1_io_eo[45] ,
    \cb_2_1_io_eo[44] ,
    \cb_2_1_io_eo[43] ,
    \cb_2_1_io_eo[42] ,
    \cb_2_1_io_eo[41] ,
    \cb_2_1_io_eo[40] ,
    \cb_2_1_io_eo[39] ,
    \cb_2_1_io_eo[38] ,
    \cb_2_1_io_eo[37] ,
    \cb_2_1_io_eo[36] ,
    \cb_2_1_io_eo[35] ,
    \cb_2_1_io_eo[34] ,
    \cb_2_1_io_eo[33] ,
    \cb_2_1_io_eo[32] ,
    \cb_2_1_io_eo[31] ,
    \cb_2_1_io_eo[30] ,
    \cb_2_1_io_eo[29] ,
    \cb_2_1_io_eo[28] ,
    \cb_2_1_io_eo[27] ,
    \cb_2_1_io_eo[26] ,
    \cb_2_1_io_eo[25] ,
    \cb_2_1_io_eo[24] ,
    \cb_2_1_io_eo[23] ,
    \cb_2_1_io_eo[22] ,
    \cb_2_1_io_eo[21] ,
    \cb_2_1_io_eo[20] ,
    \cb_2_1_io_eo[19] ,
    \cb_2_1_io_eo[18] ,
    \cb_2_1_io_eo[17] ,
    \cb_2_1_io_eo[16] ,
    \cb_2_1_io_eo[15] ,
    \cb_2_1_io_eo[14] ,
    \cb_2_1_io_eo[13] ,
    \cb_2_1_io_eo[12] ,
    \cb_2_1_io_eo[11] ,
    \cb_2_1_io_eo[10] ,
    \cb_2_1_io_eo[9] ,
    \cb_2_1_io_eo[8] ,
    \cb_2_1_io_eo[7] ,
    \cb_2_1_io_eo[6] ,
    \cb_2_1_io_eo[5] ,
    \cb_2_1_io_eo[4] ,
    \cb_2_1_io_eo[3] ,
    \cb_2_1_io_eo[2] ,
    \cb_2_1_io_eo[1] ,
    \cb_2_1_io_eo[0] }));
 cic_block cb_2_3 (.io_cs_i(cb_2_3_io_cs_i),
    .io_i_0_ci(cb_2_2_io_o_0_co),
    .io_i_1_ci(cb_2_2_io_o_1_co),
    .io_i_2_ci(cb_2_2_io_o_2_co),
    .io_i_3_ci(cb_2_2_io_o_3_co),
    .io_i_4_ci(cb_2_2_io_o_4_co),
    .io_i_5_ci(cb_2_2_io_o_5_co),
    .io_i_6_ci(cb_2_2_io_o_6_co),
    .io_i_7_ci(cb_2_2_io_o_7_co),
    .io_o_0_co(cb_2_3_io_o_0_co),
    .io_o_1_co(cb_2_3_io_o_1_co),
    .io_o_2_co(cb_2_3_io_o_2_co),
    .io_o_3_co(cb_2_3_io_o_3_co),
    .io_o_4_co(cb_2_3_io_o_4_co),
    .io_o_5_co(cb_2_3_io_o_5_co),
    .io_o_6_co(cb_2_3_io_o_6_co),
    .io_o_7_co(cb_2_3_io_o_7_co),
    .io_vci(cb_2_2_io_vco),
    .io_vco(cb_2_3_io_vco),
    .io_vi(cb_2_3_io_vi),
    .io_we_i(cb_2_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_2_0_io_adr_i[1] ,
    \cb_2_0_io_adr_i[0] }),
    .io_dat_i({\cb_2_0_io_dat_i[15] ,
    \cb_2_0_io_dat_i[14] ,
    \cb_2_0_io_dat_i[13] ,
    \cb_2_0_io_dat_i[12] ,
    \cb_2_0_io_dat_i[11] ,
    \cb_2_0_io_dat_i[10] ,
    \cb_2_0_io_dat_i[9] ,
    \cb_2_0_io_dat_i[8] ,
    \cb_2_0_io_dat_i[7] ,
    \cb_2_0_io_dat_i[6] ,
    \cb_2_0_io_dat_i[5] ,
    \cb_2_0_io_dat_i[4] ,
    \cb_2_0_io_dat_i[3] ,
    \cb_2_0_io_dat_i[2] ,
    \cb_2_0_io_dat_i[1] ,
    \cb_2_0_io_dat_i[0] }),
    .io_dat_o({\cb_2_3_io_dat_o[15] ,
    \cb_2_3_io_dat_o[14] ,
    \cb_2_3_io_dat_o[13] ,
    \cb_2_3_io_dat_o[12] ,
    \cb_2_3_io_dat_o[11] ,
    \cb_2_3_io_dat_o[10] ,
    \cb_2_3_io_dat_o[9] ,
    \cb_2_3_io_dat_o[8] ,
    \cb_2_3_io_dat_o[7] ,
    \cb_2_3_io_dat_o[6] ,
    \cb_2_3_io_dat_o[5] ,
    \cb_2_3_io_dat_o[4] ,
    \cb_2_3_io_dat_o[3] ,
    \cb_2_3_io_dat_o[2] ,
    \cb_2_3_io_dat_o[1] ,
    \cb_2_3_io_dat_o[0] }),
    .io_eo({\cb_2_3_io_eo[63] ,
    \cb_2_3_io_eo[62] ,
    \cb_2_3_io_eo[61] ,
    \cb_2_3_io_eo[60] ,
    \cb_2_3_io_eo[59] ,
    \cb_2_3_io_eo[58] ,
    \cb_2_3_io_eo[57] ,
    \cb_2_3_io_eo[56] ,
    \cb_2_3_io_eo[55] ,
    \cb_2_3_io_eo[54] ,
    \cb_2_3_io_eo[53] ,
    \cb_2_3_io_eo[52] ,
    \cb_2_3_io_eo[51] ,
    \cb_2_3_io_eo[50] ,
    \cb_2_3_io_eo[49] ,
    \cb_2_3_io_eo[48] ,
    \cb_2_3_io_eo[47] ,
    \cb_2_3_io_eo[46] ,
    \cb_2_3_io_eo[45] ,
    \cb_2_3_io_eo[44] ,
    \cb_2_3_io_eo[43] ,
    \cb_2_3_io_eo[42] ,
    \cb_2_3_io_eo[41] ,
    \cb_2_3_io_eo[40] ,
    \cb_2_3_io_eo[39] ,
    \cb_2_3_io_eo[38] ,
    \cb_2_3_io_eo[37] ,
    \cb_2_3_io_eo[36] ,
    \cb_2_3_io_eo[35] ,
    \cb_2_3_io_eo[34] ,
    \cb_2_3_io_eo[33] ,
    \cb_2_3_io_eo[32] ,
    \cb_2_3_io_eo[31] ,
    \cb_2_3_io_eo[30] ,
    \cb_2_3_io_eo[29] ,
    \cb_2_3_io_eo[28] ,
    \cb_2_3_io_eo[27] ,
    \cb_2_3_io_eo[26] ,
    \cb_2_3_io_eo[25] ,
    \cb_2_3_io_eo[24] ,
    \cb_2_3_io_eo[23] ,
    \cb_2_3_io_eo[22] ,
    \cb_2_3_io_eo[21] ,
    \cb_2_3_io_eo[20] ,
    \cb_2_3_io_eo[19] ,
    \cb_2_3_io_eo[18] ,
    \cb_2_3_io_eo[17] ,
    \cb_2_3_io_eo[16] ,
    \cb_2_3_io_eo[15] ,
    \cb_2_3_io_eo[14] ,
    \cb_2_3_io_eo[13] ,
    \cb_2_3_io_eo[12] ,
    \cb_2_3_io_eo[11] ,
    \cb_2_3_io_eo[10] ,
    \cb_2_3_io_eo[9] ,
    \cb_2_3_io_eo[8] ,
    \cb_2_3_io_eo[7] ,
    \cb_2_3_io_eo[6] ,
    \cb_2_3_io_eo[5] ,
    \cb_2_3_io_eo[4] ,
    \cb_2_3_io_eo[3] ,
    \cb_2_3_io_eo[2] ,
    \cb_2_3_io_eo[1] ,
    \cb_2_3_io_eo[0] }),
    .io_i_0_in1({\cb_2_2_io_o_0_out[7] ,
    \cb_2_2_io_o_0_out[6] ,
    \cb_2_2_io_o_0_out[5] ,
    \cb_2_2_io_o_0_out[4] ,
    \cb_2_2_io_o_0_out[3] ,
    \cb_2_2_io_o_0_out[2] ,
    \cb_2_2_io_o_0_out[1] ,
    \cb_2_2_io_o_0_out[0] }),
    .io_i_1_in1({\cb_2_2_io_o_1_out[7] ,
    \cb_2_2_io_o_1_out[6] ,
    \cb_2_2_io_o_1_out[5] ,
    \cb_2_2_io_o_1_out[4] ,
    \cb_2_2_io_o_1_out[3] ,
    \cb_2_2_io_o_1_out[2] ,
    \cb_2_2_io_o_1_out[1] ,
    \cb_2_2_io_o_1_out[0] }),
    .io_i_2_in1({\cb_2_2_io_o_2_out[7] ,
    \cb_2_2_io_o_2_out[6] ,
    \cb_2_2_io_o_2_out[5] ,
    \cb_2_2_io_o_2_out[4] ,
    \cb_2_2_io_o_2_out[3] ,
    \cb_2_2_io_o_2_out[2] ,
    \cb_2_2_io_o_2_out[1] ,
    \cb_2_2_io_o_2_out[0] }),
    .io_i_3_in1({\cb_2_2_io_o_3_out[7] ,
    \cb_2_2_io_o_3_out[6] ,
    \cb_2_2_io_o_3_out[5] ,
    \cb_2_2_io_o_3_out[4] ,
    \cb_2_2_io_o_3_out[3] ,
    \cb_2_2_io_o_3_out[2] ,
    \cb_2_2_io_o_3_out[1] ,
    \cb_2_2_io_o_3_out[0] }),
    .io_i_4_in1({\cb_2_2_io_o_4_out[7] ,
    \cb_2_2_io_o_4_out[6] ,
    \cb_2_2_io_o_4_out[5] ,
    \cb_2_2_io_o_4_out[4] ,
    \cb_2_2_io_o_4_out[3] ,
    \cb_2_2_io_o_4_out[2] ,
    \cb_2_2_io_o_4_out[1] ,
    \cb_2_2_io_o_4_out[0] }),
    .io_i_5_in1({\cb_2_2_io_o_5_out[7] ,
    \cb_2_2_io_o_5_out[6] ,
    \cb_2_2_io_o_5_out[5] ,
    \cb_2_2_io_o_5_out[4] ,
    \cb_2_2_io_o_5_out[3] ,
    \cb_2_2_io_o_5_out[2] ,
    \cb_2_2_io_o_5_out[1] ,
    \cb_2_2_io_o_5_out[0] }),
    .io_i_6_in1({\cb_2_2_io_o_6_out[7] ,
    \cb_2_2_io_o_6_out[6] ,
    \cb_2_2_io_o_6_out[5] ,
    \cb_2_2_io_o_6_out[4] ,
    \cb_2_2_io_o_6_out[3] ,
    \cb_2_2_io_o_6_out[2] ,
    \cb_2_2_io_o_6_out[1] ,
    \cb_2_2_io_o_6_out[0] }),
    .io_i_7_in1({\cb_2_2_io_o_7_out[7] ,
    \cb_2_2_io_o_7_out[6] ,
    \cb_2_2_io_o_7_out[5] ,
    \cb_2_2_io_o_7_out[4] ,
    \cb_2_2_io_o_7_out[3] ,
    \cb_2_2_io_o_7_out[2] ,
    \cb_2_2_io_o_7_out[1] ,
    \cb_2_2_io_o_7_out[0] }),
    .io_o_0_out({\cb_2_3_io_o_0_out[7] ,
    \cb_2_3_io_o_0_out[6] ,
    \cb_2_3_io_o_0_out[5] ,
    \cb_2_3_io_o_0_out[4] ,
    \cb_2_3_io_o_0_out[3] ,
    \cb_2_3_io_o_0_out[2] ,
    \cb_2_3_io_o_0_out[1] ,
    \cb_2_3_io_o_0_out[0] }),
    .io_o_1_out({\cb_2_3_io_o_1_out[7] ,
    \cb_2_3_io_o_1_out[6] ,
    \cb_2_3_io_o_1_out[5] ,
    \cb_2_3_io_o_1_out[4] ,
    \cb_2_3_io_o_1_out[3] ,
    \cb_2_3_io_o_1_out[2] ,
    \cb_2_3_io_o_1_out[1] ,
    \cb_2_3_io_o_1_out[0] }),
    .io_o_2_out({\cb_2_3_io_o_2_out[7] ,
    \cb_2_3_io_o_2_out[6] ,
    \cb_2_3_io_o_2_out[5] ,
    \cb_2_3_io_o_2_out[4] ,
    \cb_2_3_io_o_2_out[3] ,
    \cb_2_3_io_o_2_out[2] ,
    \cb_2_3_io_o_2_out[1] ,
    \cb_2_3_io_o_2_out[0] }),
    .io_o_3_out({\cb_2_3_io_o_3_out[7] ,
    \cb_2_3_io_o_3_out[6] ,
    \cb_2_3_io_o_3_out[5] ,
    \cb_2_3_io_o_3_out[4] ,
    \cb_2_3_io_o_3_out[3] ,
    \cb_2_3_io_o_3_out[2] ,
    \cb_2_3_io_o_3_out[1] ,
    \cb_2_3_io_o_3_out[0] }),
    .io_o_4_out({\cb_2_3_io_o_4_out[7] ,
    \cb_2_3_io_o_4_out[6] ,
    \cb_2_3_io_o_4_out[5] ,
    \cb_2_3_io_o_4_out[4] ,
    \cb_2_3_io_o_4_out[3] ,
    \cb_2_3_io_o_4_out[2] ,
    \cb_2_3_io_o_4_out[1] ,
    \cb_2_3_io_o_4_out[0] }),
    .io_o_5_out({\cb_2_3_io_o_5_out[7] ,
    \cb_2_3_io_o_5_out[6] ,
    \cb_2_3_io_o_5_out[5] ,
    \cb_2_3_io_o_5_out[4] ,
    \cb_2_3_io_o_5_out[3] ,
    \cb_2_3_io_o_5_out[2] ,
    \cb_2_3_io_o_5_out[1] ,
    \cb_2_3_io_o_5_out[0] }),
    .io_o_6_out({\cb_2_3_io_o_6_out[7] ,
    \cb_2_3_io_o_6_out[6] ,
    \cb_2_3_io_o_6_out[5] ,
    \cb_2_3_io_o_6_out[4] ,
    \cb_2_3_io_o_6_out[3] ,
    \cb_2_3_io_o_6_out[2] ,
    \cb_2_3_io_o_6_out[1] ,
    \cb_2_3_io_o_6_out[0] }),
    .io_o_7_out({\cb_2_3_io_o_7_out[7] ,
    \cb_2_3_io_o_7_out[6] ,
    \cb_2_3_io_o_7_out[5] ,
    \cb_2_3_io_o_7_out[4] ,
    \cb_2_3_io_o_7_out[3] ,
    \cb_2_3_io_o_7_out[2] ,
    \cb_2_3_io_o_7_out[1] ,
    \cb_2_3_io_o_7_out[0] }),
    .io_wo({\cb_2_2_io_eo[63] ,
    \cb_2_2_io_eo[62] ,
    \cb_2_2_io_eo[61] ,
    \cb_2_2_io_eo[60] ,
    \cb_2_2_io_eo[59] ,
    \cb_2_2_io_eo[58] ,
    \cb_2_2_io_eo[57] ,
    \cb_2_2_io_eo[56] ,
    \cb_2_2_io_eo[55] ,
    \cb_2_2_io_eo[54] ,
    \cb_2_2_io_eo[53] ,
    \cb_2_2_io_eo[52] ,
    \cb_2_2_io_eo[51] ,
    \cb_2_2_io_eo[50] ,
    \cb_2_2_io_eo[49] ,
    \cb_2_2_io_eo[48] ,
    \cb_2_2_io_eo[47] ,
    \cb_2_2_io_eo[46] ,
    \cb_2_2_io_eo[45] ,
    \cb_2_2_io_eo[44] ,
    \cb_2_2_io_eo[43] ,
    \cb_2_2_io_eo[42] ,
    \cb_2_2_io_eo[41] ,
    \cb_2_2_io_eo[40] ,
    \cb_2_2_io_eo[39] ,
    \cb_2_2_io_eo[38] ,
    \cb_2_2_io_eo[37] ,
    \cb_2_2_io_eo[36] ,
    \cb_2_2_io_eo[35] ,
    \cb_2_2_io_eo[34] ,
    \cb_2_2_io_eo[33] ,
    \cb_2_2_io_eo[32] ,
    \cb_2_2_io_eo[31] ,
    \cb_2_2_io_eo[30] ,
    \cb_2_2_io_eo[29] ,
    \cb_2_2_io_eo[28] ,
    \cb_2_2_io_eo[27] ,
    \cb_2_2_io_eo[26] ,
    \cb_2_2_io_eo[25] ,
    \cb_2_2_io_eo[24] ,
    \cb_2_2_io_eo[23] ,
    \cb_2_2_io_eo[22] ,
    \cb_2_2_io_eo[21] ,
    \cb_2_2_io_eo[20] ,
    \cb_2_2_io_eo[19] ,
    \cb_2_2_io_eo[18] ,
    \cb_2_2_io_eo[17] ,
    \cb_2_2_io_eo[16] ,
    \cb_2_2_io_eo[15] ,
    \cb_2_2_io_eo[14] ,
    \cb_2_2_io_eo[13] ,
    \cb_2_2_io_eo[12] ,
    \cb_2_2_io_eo[11] ,
    \cb_2_2_io_eo[10] ,
    \cb_2_2_io_eo[9] ,
    \cb_2_2_io_eo[8] ,
    \cb_2_2_io_eo[7] ,
    \cb_2_2_io_eo[6] ,
    \cb_2_2_io_eo[5] ,
    \cb_2_2_io_eo[4] ,
    \cb_2_2_io_eo[3] ,
    \cb_2_2_io_eo[2] ,
    \cb_2_2_io_eo[1] ,
    \cb_2_2_io_eo[0] }));
 cic_block cb_2_4 (.io_cs_i(cb_2_4_io_cs_i),
    .io_i_0_ci(cb_2_3_io_o_0_co),
    .io_i_1_ci(cb_2_3_io_o_1_co),
    .io_i_2_ci(cb_2_3_io_o_2_co),
    .io_i_3_ci(cb_2_3_io_o_3_co),
    .io_i_4_ci(cb_2_3_io_o_4_co),
    .io_i_5_ci(cb_2_3_io_o_5_co),
    .io_i_6_ci(cb_2_3_io_o_6_co),
    .io_i_7_ci(cb_2_3_io_o_7_co),
    .io_o_0_co(cb_2_4_io_o_0_co),
    .io_o_1_co(cb_2_4_io_o_1_co),
    .io_o_2_co(cb_2_4_io_o_2_co),
    .io_o_3_co(cb_2_4_io_o_3_co),
    .io_o_4_co(cb_2_4_io_o_4_co),
    .io_o_5_co(cb_2_4_io_o_5_co),
    .io_o_6_co(cb_2_4_io_o_6_co),
    .io_o_7_co(cb_2_4_io_o_7_co),
    .io_vci(cb_2_3_io_vco),
    .io_vco(cb_2_4_io_vco),
    .io_vi(cb_2_4_io_vi),
    .io_we_i(cb_2_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_2_0_io_adr_i[1] ,
    \cb_2_0_io_adr_i[0] }),
    .io_dat_i({\cb_2_0_io_dat_i[15] ,
    \cb_2_0_io_dat_i[14] ,
    \cb_2_0_io_dat_i[13] ,
    \cb_2_0_io_dat_i[12] ,
    \cb_2_0_io_dat_i[11] ,
    \cb_2_0_io_dat_i[10] ,
    \cb_2_0_io_dat_i[9] ,
    \cb_2_0_io_dat_i[8] ,
    \cb_2_0_io_dat_i[7] ,
    \cb_2_0_io_dat_i[6] ,
    \cb_2_0_io_dat_i[5] ,
    \cb_2_0_io_dat_i[4] ,
    \cb_2_0_io_dat_i[3] ,
    \cb_2_0_io_dat_i[2] ,
    \cb_2_0_io_dat_i[1] ,
    \cb_2_0_io_dat_i[0] }),
    .io_dat_o({\cb_2_4_io_dat_o[15] ,
    \cb_2_4_io_dat_o[14] ,
    \cb_2_4_io_dat_o[13] ,
    \cb_2_4_io_dat_o[12] ,
    \cb_2_4_io_dat_o[11] ,
    \cb_2_4_io_dat_o[10] ,
    \cb_2_4_io_dat_o[9] ,
    \cb_2_4_io_dat_o[8] ,
    \cb_2_4_io_dat_o[7] ,
    \cb_2_4_io_dat_o[6] ,
    \cb_2_4_io_dat_o[5] ,
    \cb_2_4_io_dat_o[4] ,
    \cb_2_4_io_dat_o[3] ,
    \cb_2_4_io_dat_o[2] ,
    \cb_2_4_io_dat_o[1] ,
    \cb_2_4_io_dat_o[0] }),
    .io_eo({\cb_2_4_io_eo[63] ,
    \cb_2_4_io_eo[62] ,
    \cb_2_4_io_eo[61] ,
    \cb_2_4_io_eo[60] ,
    \cb_2_4_io_eo[59] ,
    \cb_2_4_io_eo[58] ,
    \cb_2_4_io_eo[57] ,
    \cb_2_4_io_eo[56] ,
    \cb_2_4_io_eo[55] ,
    \cb_2_4_io_eo[54] ,
    \cb_2_4_io_eo[53] ,
    \cb_2_4_io_eo[52] ,
    \cb_2_4_io_eo[51] ,
    \cb_2_4_io_eo[50] ,
    \cb_2_4_io_eo[49] ,
    \cb_2_4_io_eo[48] ,
    \cb_2_4_io_eo[47] ,
    \cb_2_4_io_eo[46] ,
    \cb_2_4_io_eo[45] ,
    \cb_2_4_io_eo[44] ,
    \cb_2_4_io_eo[43] ,
    \cb_2_4_io_eo[42] ,
    \cb_2_4_io_eo[41] ,
    \cb_2_4_io_eo[40] ,
    \cb_2_4_io_eo[39] ,
    \cb_2_4_io_eo[38] ,
    \cb_2_4_io_eo[37] ,
    \cb_2_4_io_eo[36] ,
    \cb_2_4_io_eo[35] ,
    \cb_2_4_io_eo[34] ,
    \cb_2_4_io_eo[33] ,
    \cb_2_4_io_eo[32] ,
    \cb_2_4_io_eo[31] ,
    \cb_2_4_io_eo[30] ,
    \cb_2_4_io_eo[29] ,
    \cb_2_4_io_eo[28] ,
    \cb_2_4_io_eo[27] ,
    \cb_2_4_io_eo[26] ,
    \cb_2_4_io_eo[25] ,
    \cb_2_4_io_eo[24] ,
    \cb_2_4_io_eo[23] ,
    \cb_2_4_io_eo[22] ,
    \cb_2_4_io_eo[21] ,
    \cb_2_4_io_eo[20] ,
    \cb_2_4_io_eo[19] ,
    \cb_2_4_io_eo[18] ,
    \cb_2_4_io_eo[17] ,
    \cb_2_4_io_eo[16] ,
    \cb_2_4_io_eo[15] ,
    \cb_2_4_io_eo[14] ,
    \cb_2_4_io_eo[13] ,
    \cb_2_4_io_eo[12] ,
    \cb_2_4_io_eo[11] ,
    \cb_2_4_io_eo[10] ,
    \cb_2_4_io_eo[9] ,
    \cb_2_4_io_eo[8] ,
    \cb_2_4_io_eo[7] ,
    \cb_2_4_io_eo[6] ,
    \cb_2_4_io_eo[5] ,
    \cb_2_4_io_eo[4] ,
    \cb_2_4_io_eo[3] ,
    \cb_2_4_io_eo[2] ,
    \cb_2_4_io_eo[1] ,
    \cb_2_4_io_eo[0] }),
    .io_i_0_in1({\cb_2_3_io_o_0_out[7] ,
    \cb_2_3_io_o_0_out[6] ,
    \cb_2_3_io_o_0_out[5] ,
    \cb_2_3_io_o_0_out[4] ,
    \cb_2_3_io_o_0_out[3] ,
    \cb_2_3_io_o_0_out[2] ,
    \cb_2_3_io_o_0_out[1] ,
    \cb_2_3_io_o_0_out[0] }),
    .io_i_1_in1({\cb_2_3_io_o_1_out[7] ,
    \cb_2_3_io_o_1_out[6] ,
    \cb_2_3_io_o_1_out[5] ,
    \cb_2_3_io_o_1_out[4] ,
    \cb_2_3_io_o_1_out[3] ,
    \cb_2_3_io_o_1_out[2] ,
    \cb_2_3_io_o_1_out[1] ,
    \cb_2_3_io_o_1_out[0] }),
    .io_i_2_in1({\cb_2_3_io_o_2_out[7] ,
    \cb_2_3_io_o_2_out[6] ,
    \cb_2_3_io_o_2_out[5] ,
    \cb_2_3_io_o_2_out[4] ,
    \cb_2_3_io_o_2_out[3] ,
    \cb_2_3_io_o_2_out[2] ,
    \cb_2_3_io_o_2_out[1] ,
    \cb_2_3_io_o_2_out[0] }),
    .io_i_3_in1({\cb_2_3_io_o_3_out[7] ,
    \cb_2_3_io_o_3_out[6] ,
    \cb_2_3_io_o_3_out[5] ,
    \cb_2_3_io_o_3_out[4] ,
    \cb_2_3_io_o_3_out[3] ,
    \cb_2_3_io_o_3_out[2] ,
    \cb_2_3_io_o_3_out[1] ,
    \cb_2_3_io_o_3_out[0] }),
    .io_i_4_in1({\cb_2_3_io_o_4_out[7] ,
    \cb_2_3_io_o_4_out[6] ,
    \cb_2_3_io_o_4_out[5] ,
    \cb_2_3_io_o_4_out[4] ,
    \cb_2_3_io_o_4_out[3] ,
    \cb_2_3_io_o_4_out[2] ,
    \cb_2_3_io_o_4_out[1] ,
    \cb_2_3_io_o_4_out[0] }),
    .io_i_5_in1({\cb_2_3_io_o_5_out[7] ,
    \cb_2_3_io_o_5_out[6] ,
    \cb_2_3_io_o_5_out[5] ,
    \cb_2_3_io_o_5_out[4] ,
    \cb_2_3_io_o_5_out[3] ,
    \cb_2_3_io_o_5_out[2] ,
    \cb_2_3_io_o_5_out[1] ,
    \cb_2_3_io_o_5_out[0] }),
    .io_i_6_in1({\cb_2_3_io_o_6_out[7] ,
    \cb_2_3_io_o_6_out[6] ,
    \cb_2_3_io_o_6_out[5] ,
    \cb_2_3_io_o_6_out[4] ,
    \cb_2_3_io_o_6_out[3] ,
    \cb_2_3_io_o_6_out[2] ,
    \cb_2_3_io_o_6_out[1] ,
    \cb_2_3_io_o_6_out[0] }),
    .io_i_7_in1({\cb_2_3_io_o_7_out[7] ,
    \cb_2_3_io_o_7_out[6] ,
    \cb_2_3_io_o_7_out[5] ,
    \cb_2_3_io_o_7_out[4] ,
    \cb_2_3_io_o_7_out[3] ,
    \cb_2_3_io_o_7_out[2] ,
    \cb_2_3_io_o_7_out[1] ,
    \cb_2_3_io_o_7_out[0] }),
    .io_o_0_out({\cb_2_4_io_o_0_out[7] ,
    \cb_2_4_io_o_0_out[6] ,
    \cb_2_4_io_o_0_out[5] ,
    \cb_2_4_io_o_0_out[4] ,
    \cb_2_4_io_o_0_out[3] ,
    \cb_2_4_io_o_0_out[2] ,
    \cb_2_4_io_o_0_out[1] ,
    \cb_2_4_io_o_0_out[0] }),
    .io_o_1_out({\cb_2_4_io_o_1_out[7] ,
    \cb_2_4_io_o_1_out[6] ,
    \cb_2_4_io_o_1_out[5] ,
    \cb_2_4_io_o_1_out[4] ,
    \cb_2_4_io_o_1_out[3] ,
    \cb_2_4_io_o_1_out[2] ,
    \cb_2_4_io_o_1_out[1] ,
    \cb_2_4_io_o_1_out[0] }),
    .io_o_2_out({\cb_2_4_io_o_2_out[7] ,
    \cb_2_4_io_o_2_out[6] ,
    \cb_2_4_io_o_2_out[5] ,
    \cb_2_4_io_o_2_out[4] ,
    \cb_2_4_io_o_2_out[3] ,
    \cb_2_4_io_o_2_out[2] ,
    \cb_2_4_io_o_2_out[1] ,
    \cb_2_4_io_o_2_out[0] }),
    .io_o_3_out({\cb_2_4_io_o_3_out[7] ,
    \cb_2_4_io_o_3_out[6] ,
    \cb_2_4_io_o_3_out[5] ,
    \cb_2_4_io_o_3_out[4] ,
    \cb_2_4_io_o_3_out[3] ,
    \cb_2_4_io_o_3_out[2] ,
    \cb_2_4_io_o_3_out[1] ,
    \cb_2_4_io_o_3_out[0] }),
    .io_o_4_out({\cb_2_4_io_o_4_out[7] ,
    \cb_2_4_io_o_4_out[6] ,
    \cb_2_4_io_o_4_out[5] ,
    \cb_2_4_io_o_4_out[4] ,
    \cb_2_4_io_o_4_out[3] ,
    \cb_2_4_io_o_4_out[2] ,
    \cb_2_4_io_o_4_out[1] ,
    \cb_2_4_io_o_4_out[0] }),
    .io_o_5_out({\cb_2_4_io_o_5_out[7] ,
    \cb_2_4_io_o_5_out[6] ,
    \cb_2_4_io_o_5_out[5] ,
    \cb_2_4_io_o_5_out[4] ,
    \cb_2_4_io_o_5_out[3] ,
    \cb_2_4_io_o_5_out[2] ,
    \cb_2_4_io_o_5_out[1] ,
    \cb_2_4_io_o_5_out[0] }),
    .io_o_6_out({\cb_2_4_io_o_6_out[7] ,
    \cb_2_4_io_o_6_out[6] ,
    \cb_2_4_io_o_6_out[5] ,
    \cb_2_4_io_o_6_out[4] ,
    \cb_2_4_io_o_6_out[3] ,
    \cb_2_4_io_o_6_out[2] ,
    \cb_2_4_io_o_6_out[1] ,
    \cb_2_4_io_o_6_out[0] }),
    .io_o_7_out({\cb_2_4_io_o_7_out[7] ,
    \cb_2_4_io_o_7_out[6] ,
    \cb_2_4_io_o_7_out[5] ,
    \cb_2_4_io_o_7_out[4] ,
    \cb_2_4_io_o_7_out[3] ,
    \cb_2_4_io_o_7_out[2] ,
    \cb_2_4_io_o_7_out[1] ,
    \cb_2_4_io_o_7_out[0] }),
    .io_wo({\cb_2_3_io_eo[63] ,
    \cb_2_3_io_eo[62] ,
    \cb_2_3_io_eo[61] ,
    \cb_2_3_io_eo[60] ,
    \cb_2_3_io_eo[59] ,
    \cb_2_3_io_eo[58] ,
    \cb_2_3_io_eo[57] ,
    \cb_2_3_io_eo[56] ,
    \cb_2_3_io_eo[55] ,
    \cb_2_3_io_eo[54] ,
    \cb_2_3_io_eo[53] ,
    \cb_2_3_io_eo[52] ,
    \cb_2_3_io_eo[51] ,
    \cb_2_3_io_eo[50] ,
    \cb_2_3_io_eo[49] ,
    \cb_2_3_io_eo[48] ,
    \cb_2_3_io_eo[47] ,
    \cb_2_3_io_eo[46] ,
    \cb_2_3_io_eo[45] ,
    \cb_2_3_io_eo[44] ,
    \cb_2_3_io_eo[43] ,
    \cb_2_3_io_eo[42] ,
    \cb_2_3_io_eo[41] ,
    \cb_2_3_io_eo[40] ,
    \cb_2_3_io_eo[39] ,
    \cb_2_3_io_eo[38] ,
    \cb_2_3_io_eo[37] ,
    \cb_2_3_io_eo[36] ,
    \cb_2_3_io_eo[35] ,
    \cb_2_3_io_eo[34] ,
    \cb_2_3_io_eo[33] ,
    \cb_2_3_io_eo[32] ,
    \cb_2_3_io_eo[31] ,
    \cb_2_3_io_eo[30] ,
    \cb_2_3_io_eo[29] ,
    \cb_2_3_io_eo[28] ,
    \cb_2_3_io_eo[27] ,
    \cb_2_3_io_eo[26] ,
    \cb_2_3_io_eo[25] ,
    \cb_2_3_io_eo[24] ,
    \cb_2_3_io_eo[23] ,
    \cb_2_3_io_eo[22] ,
    \cb_2_3_io_eo[21] ,
    \cb_2_3_io_eo[20] ,
    \cb_2_3_io_eo[19] ,
    \cb_2_3_io_eo[18] ,
    \cb_2_3_io_eo[17] ,
    \cb_2_3_io_eo[16] ,
    \cb_2_3_io_eo[15] ,
    \cb_2_3_io_eo[14] ,
    \cb_2_3_io_eo[13] ,
    \cb_2_3_io_eo[12] ,
    \cb_2_3_io_eo[11] ,
    \cb_2_3_io_eo[10] ,
    \cb_2_3_io_eo[9] ,
    \cb_2_3_io_eo[8] ,
    \cb_2_3_io_eo[7] ,
    \cb_2_3_io_eo[6] ,
    \cb_2_3_io_eo[5] ,
    \cb_2_3_io_eo[4] ,
    \cb_2_3_io_eo[3] ,
    \cb_2_3_io_eo[2] ,
    \cb_2_3_io_eo[1] ,
    \cb_2_3_io_eo[0] }));
 cic_block cb_2_5 (.io_cs_i(cb_2_5_io_cs_i),
    .io_i_0_ci(cb_2_4_io_o_0_co),
    .io_i_1_ci(cb_2_4_io_o_1_co),
    .io_i_2_ci(cb_2_4_io_o_2_co),
    .io_i_3_ci(cb_2_4_io_o_3_co),
    .io_i_4_ci(cb_2_4_io_o_4_co),
    .io_i_5_ci(cb_2_4_io_o_5_co),
    .io_i_6_ci(cb_2_4_io_o_6_co),
    .io_i_7_ci(cb_2_4_io_o_7_co),
    .io_o_0_co(cb_2_5_io_o_0_co),
    .io_o_1_co(cb_2_5_io_o_1_co),
    .io_o_2_co(cb_2_5_io_o_2_co),
    .io_o_3_co(cb_2_5_io_o_3_co),
    .io_o_4_co(cb_2_5_io_o_4_co),
    .io_o_5_co(cb_2_5_io_o_5_co),
    .io_o_6_co(cb_2_5_io_o_6_co),
    .io_o_7_co(cb_2_5_io_o_7_co),
    .io_vci(cb_2_4_io_vco),
    .io_vco(cb_2_5_io_vco),
    .io_vi(cb_2_5_io_vi),
    .io_we_i(cb_2_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_2_0_io_adr_i[1] ,
    \cb_2_0_io_adr_i[0] }),
    .io_dat_i({\cb_2_0_io_dat_i[15] ,
    \cb_2_0_io_dat_i[14] ,
    \cb_2_0_io_dat_i[13] ,
    \cb_2_0_io_dat_i[12] ,
    \cb_2_0_io_dat_i[11] ,
    \cb_2_0_io_dat_i[10] ,
    \cb_2_0_io_dat_i[9] ,
    \cb_2_0_io_dat_i[8] ,
    \cb_2_0_io_dat_i[7] ,
    \cb_2_0_io_dat_i[6] ,
    \cb_2_0_io_dat_i[5] ,
    \cb_2_0_io_dat_i[4] ,
    \cb_2_0_io_dat_i[3] ,
    \cb_2_0_io_dat_i[2] ,
    \cb_2_0_io_dat_i[1] ,
    \cb_2_0_io_dat_i[0] }),
    .io_dat_o({\cb_2_5_io_dat_o[15] ,
    \cb_2_5_io_dat_o[14] ,
    \cb_2_5_io_dat_o[13] ,
    \cb_2_5_io_dat_o[12] ,
    \cb_2_5_io_dat_o[11] ,
    \cb_2_5_io_dat_o[10] ,
    \cb_2_5_io_dat_o[9] ,
    \cb_2_5_io_dat_o[8] ,
    \cb_2_5_io_dat_o[7] ,
    \cb_2_5_io_dat_o[6] ,
    \cb_2_5_io_dat_o[5] ,
    \cb_2_5_io_dat_o[4] ,
    \cb_2_5_io_dat_o[3] ,
    \cb_2_5_io_dat_o[2] ,
    \cb_2_5_io_dat_o[1] ,
    \cb_2_5_io_dat_o[0] }),
    .io_eo({\cb_2_5_io_eo[63] ,
    \cb_2_5_io_eo[62] ,
    \cb_2_5_io_eo[61] ,
    \cb_2_5_io_eo[60] ,
    \cb_2_5_io_eo[59] ,
    \cb_2_5_io_eo[58] ,
    \cb_2_5_io_eo[57] ,
    \cb_2_5_io_eo[56] ,
    \cb_2_5_io_eo[55] ,
    \cb_2_5_io_eo[54] ,
    \cb_2_5_io_eo[53] ,
    \cb_2_5_io_eo[52] ,
    \cb_2_5_io_eo[51] ,
    \cb_2_5_io_eo[50] ,
    \cb_2_5_io_eo[49] ,
    \cb_2_5_io_eo[48] ,
    \cb_2_5_io_eo[47] ,
    \cb_2_5_io_eo[46] ,
    \cb_2_5_io_eo[45] ,
    \cb_2_5_io_eo[44] ,
    \cb_2_5_io_eo[43] ,
    \cb_2_5_io_eo[42] ,
    \cb_2_5_io_eo[41] ,
    \cb_2_5_io_eo[40] ,
    \cb_2_5_io_eo[39] ,
    \cb_2_5_io_eo[38] ,
    \cb_2_5_io_eo[37] ,
    \cb_2_5_io_eo[36] ,
    \cb_2_5_io_eo[35] ,
    \cb_2_5_io_eo[34] ,
    \cb_2_5_io_eo[33] ,
    \cb_2_5_io_eo[32] ,
    \cb_2_5_io_eo[31] ,
    \cb_2_5_io_eo[30] ,
    \cb_2_5_io_eo[29] ,
    \cb_2_5_io_eo[28] ,
    \cb_2_5_io_eo[27] ,
    \cb_2_5_io_eo[26] ,
    \cb_2_5_io_eo[25] ,
    \cb_2_5_io_eo[24] ,
    \cb_2_5_io_eo[23] ,
    \cb_2_5_io_eo[22] ,
    \cb_2_5_io_eo[21] ,
    \cb_2_5_io_eo[20] ,
    \cb_2_5_io_eo[19] ,
    \cb_2_5_io_eo[18] ,
    \cb_2_5_io_eo[17] ,
    \cb_2_5_io_eo[16] ,
    \cb_2_5_io_eo[15] ,
    \cb_2_5_io_eo[14] ,
    \cb_2_5_io_eo[13] ,
    \cb_2_5_io_eo[12] ,
    \cb_2_5_io_eo[11] ,
    \cb_2_5_io_eo[10] ,
    \cb_2_5_io_eo[9] ,
    \cb_2_5_io_eo[8] ,
    \cb_2_5_io_eo[7] ,
    \cb_2_5_io_eo[6] ,
    \cb_2_5_io_eo[5] ,
    \cb_2_5_io_eo[4] ,
    \cb_2_5_io_eo[3] ,
    \cb_2_5_io_eo[2] ,
    \cb_2_5_io_eo[1] ,
    \cb_2_5_io_eo[0] }),
    .io_i_0_in1({\cb_2_4_io_o_0_out[7] ,
    \cb_2_4_io_o_0_out[6] ,
    \cb_2_4_io_o_0_out[5] ,
    \cb_2_4_io_o_0_out[4] ,
    \cb_2_4_io_o_0_out[3] ,
    \cb_2_4_io_o_0_out[2] ,
    \cb_2_4_io_o_0_out[1] ,
    \cb_2_4_io_o_0_out[0] }),
    .io_i_1_in1({\cb_2_4_io_o_1_out[7] ,
    \cb_2_4_io_o_1_out[6] ,
    \cb_2_4_io_o_1_out[5] ,
    \cb_2_4_io_o_1_out[4] ,
    \cb_2_4_io_o_1_out[3] ,
    \cb_2_4_io_o_1_out[2] ,
    \cb_2_4_io_o_1_out[1] ,
    \cb_2_4_io_o_1_out[0] }),
    .io_i_2_in1({\cb_2_4_io_o_2_out[7] ,
    \cb_2_4_io_o_2_out[6] ,
    \cb_2_4_io_o_2_out[5] ,
    \cb_2_4_io_o_2_out[4] ,
    \cb_2_4_io_o_2_out[3] ,
    \cb_2_4_io_o_2_out[2] ,
    \cb_2_4_io_o_2_out[1] ,
    \cb_2_4_io_o_2_out[0] }),
    .io_i_3_in1({\cb_2_4_io_o_3_out[7] ,
    \cb_2_4_io_o_3_out[6] ,
    \cb_2_4_io_o_3_out[5] ,
    \cb_2_4_io_o_3_out[4] ,
    \cb_2_4_io_o_3_out[3] ,
    \cb_2_4_io_o_3_out[2] ,
    \cb_2_4_io_o_3_out[1] ,
    \cb_2_4_io_o_3_out[0] }),
    .io_i_4_in1({\cb_2_4_io_o_4_out[7] ,
    \cb_2_4_io_o_4_out[6] ,
    \cb_2_4_io_o_4_out[5] ,
    \cb_2_4_io_o_4_out[4] ,
    \cb_2_4_io_o_4_out[3] ,
    \cb_2_4_io_o_4_out[2] ,
    \cb_2_4_io_o_4_out[1] ,
    \cb_2_4_io_o_4_out[0] }),
    .io_i_5_in1({\cb_2_4_io_o_5_out[7] ,
    \cb_2_4_io_o_5_out[6] ,
    \cb_2_4_io_o_5_out[5] ,
    \cb_2_4_io_o_5_out[4] ,
    \cb_2_4_io_o_5_out[3] ,
    \cb_2_4_io_o_5_out[2] ,
    \cb_2_4_io_o_5_out[1] ,
    \cb_2_4_io_o_5_out[0] }),
    .io_i_6_in1({\cb_2_4_io_o_6_out[7] ,
    \cb_2_4_io_o_6_out[6] ,
    \cb_2_4_io_o_6_out[5] ,
    \cb_2_4_io_o_6_out[4] ,
    \cb_2_4_io_o_6_out[3] ,
    \cb_2_4_io_o_6_out[2] ,
    \cb_2_4_io_o_6_out[1] ,
    \cb_2_4_io_o_6_out[0] }),
    .io_i_7_in1({\cb_2_4_io_o_7_out[7] ,
    \cb_2_4_io_o_7_out[6] ,
    \cb_2_4_io_o_7_out[5] ,
    \cb_2_4_io_o_7_out[4] ,
    \cb_2_4_io_o_7_out[3] ,
    \cb_2_4_io_o_7_out[2] ,
    \cb_2_4_io_o_7_out[1] ,
    \cb_2_4_io_o_7_out[0] }),
    .io_o_0_out({\cb_2_5_io_o_0_out[7] ,
    \cb_2_5_io_o_0_out[6] ,
    \cb_2_5_io_o_0_out[5] ,
    \cb_2_5_io_o_0_out[4] ,
    \cb_2_5_io_o_0_out[3] ,
    \cb_2_5_io_o_0_out[2] ,
    \cb_2_5_io_o_0_out[1] ,
    \cb_2_5_io_o_0_out[0] }),
    .io_o_1_out({\cb_2_5_io_o_1_out[7] ,
    \cb_2_5_io_o_1_out[6] ,
    \cb_2_5_io_o_1_out[5] ,
    \cb_2_5_io_o_1_out[4] ,
    \cb_2_5_io_o_1_out[3] ,
    \cb_2_5_io_o_1_out[2] ,
    \cb_2_5_io_o_1_out[1] ,
    \cb_2_5_io_o_1_out[0] }),
    .io_o_2_out({\cb_2_5_io_o_2_out[7] ,
    \cb_2_5_io_o_2_out[6] ,
    \cb_2_5_io_o_2_out[5] ,
    \cb_2_5_io_o_2_out[4] ,
    \cb_2_5_io_o_2_out[3] ,
    \cb_2_5_io_o_2_out[2] ,
    \cb_2_5_io_o_2_out[1] ,
    \cb_2_5_io_o_2_out[0] }),
    .io_o_3_out({\cb_2_5_io_o_3_out[7] ,
    \cb_2_5_io_o_3_out[6] ,
    \cb_2_5_io_o_3_out[5] ,
    \cb_2_5_io_o_3_out[4] ,
    \cb_2_5_io_o_3_out[3] ,
    \cb_2_5_io_o_3_out[2] ,
    \cb_2_5_io_o_3_out[1] ,
    \cb_2_5_io_o_3_out[0] }),
    .io_o_4_out({\cb_2_5_io_o_4_out[7] ,
    \cb_2_5_io_o_4_out[6] ,
    \cb_2_5_io_o_4_out[5] ,
    \cb_2_5_io_o_4_out[4] ,
    \cb_2_5_io_o_4_out[3] ,
    \cb_2_5_io_o_4_out[2] ,
    \cb_2_5_io_o_4_out[1] ,
    \cb_2_5_io_o_4_out[0] }),
    .io_o_5_out({\cb_2_5_io_o_5_out[7] ,
    \cb_2_5_io_o_5_out[6] ,
    \cb_2_5_io_o_5_out[5] ,
    \cb_2_5_io_o_5_out[4] ,
    \cb_2_5_io_o_5_out[3] ,
    \cb_2_5_io_o_5_out[2] ,
    \cb_2_5_io_o_5_out[1] ,
    \cb_2_5_io_o_5_out[0] }),
    .io_o_6_out({\cb_2_5_io_o_6_out[7] ,
    \cb_2_5_io_o_6_out[6] ,
    \cb_2_5_io_o_6_out[5] ,
    \cb_2_5_io_o_6_out[4] ,
    \cb_2_5_io_o_6_out[3] ,
    \cb_2_5_io_o_6_out[2] ,
    \cb_2_5_io_o_6_out[1] ,
    \cb_2_5_io_o_6_out[0] }),
    .io_o_7_out({\cb_2_5_io_o_7_out[7] ,
    \cb_2_5_io_o_7_out[6] ,
    \cb_2_5_io_o_7_out[5] ,
    \cb_2_5_io_o_7_out[4] ,
    \cb_2_5_io_o_7_out[3] ,
    \cb_2_5_io_o_7_out[2] ,
    \cb_2_5_io_o_7_out[1] ,
    \cb_2_5_io_o_7_out[0] }),
    .io_wo({\cb_2_4_io_eo[63] ,
    \cb_2_4_io_eo[62] ,
    \cb_2_4_io_eo[61] ,
    \cb_2_4_io_eo[60] ,
    \cb_2_4_io_eo[59] ,
    \cb_2_4_io_eo[58] ,
    \cb_2_4_io_eo[57] ,
    \cb_2_4_io_eo[56] ,
    \cb_2_4_io_eo[55] ,
    \cb_2_4_io_eo[54] ,
    \cb_2_4_io_eo[53] ,
    \cb_2_4_io_eo[52] ,
    \cb_2_4_io_eo[51] ,
    \cb_2_4_io_eo[50] ,
    \cb_2_4_io_eo[49] ,
    \cb_2_4_io_eo[48] ,
    \cb_2_4_io_eo[47] ,
    \cb_2_4_io_eo[46] ,
    \cb_2_4_io_eo[45] ,
    \cb_2_4_io_eo[44] ,
    \cb_2_4_io_eo[43] ,
    \cb_2_4_io_eo[42] ,
    \cb_2_4_io_eo[41] ,
    \cb_2_4_io_eo[40] ,
    \cb_2_4_io_eo[39] ,
    \cb_2_4_io_eo[38] ,
    \cb_2_4_io_eo[37] ,
    \cb_2_4_io_eo[36] ,
    \cb_2_4_io_eo[35] ,
    \cb_2_4_io_eo[34] ,
    \cb_2_4_io_eo[33] ,
    \cb_2_4_io_eo[32] ,
    \cb_2_4_io_eo[31] ,
    \cb_2_4_io_eo[30] ,
    \cb_2_4_io_eo[29] ,
    \cb_2_4_io_eo[28] ,
    \cb_2_4_io_eo[27] ,
    \cb_2_4_io_eo[26] ,
    \cb_2_4_io_eo[25] ,
    \cb_2_4_io_eo[24] ,
    \cb_2_4_io_eo[23] ,
    \cb_2_4_io_eo[22] ,
    \cb_2_4_io_eo[21] ,
    \cb_2_4_io_eo[20] ,
    \cb_2_4_io_eo[19] ,
    \cb_2_4_io_eo[18] ,
    \cb_2_4_io_eo[17] ,
    \cb_2_4_io_eo[16] ,
    \cb_2_4_io_eo[15] ,
    \cb_2_4_io_eo[14] ,
    \cb_2_4_io_eo[13] ,
    \cb_2_4_io_eo[12] ,
    \cb_2_4_io_eo[11] ,
    \cb_2_4_io_eo[10] ,
    \cb_2_4_io_eo[9] ,
    \cb_2_4_io_eo[8] ,
    \cb_2_4_io_eo[7] ,
    \cb_2_4_io_eo[6] ,
    \cb_2_4_io_eo[5] ,
    \cb_2_4_io_eo[4] ,
    \cb_2_4_io_eo[3] ,
    \cb_2_4_io_eo[2] ,
    \cb_2_4_io_eo[1] ,
    \cb_2_4_io_eo[0] }));
 cic_block cb_2_6 (.io_cs_i(cb_2_6_io_cs_i),
    .io_i_0_ci(cb_2_5_io_o_0_co),
    .io_i_1_ci(cb_2_5_io_o_1_co),
    .io_i_2_ci(cb_2_5_io_o_2_co),
    .io_i_3_ci(cb_2_5_io_o_3_co),
    .io_i_4_ci(cb_2_5_io_o_4_co),
    .io_i_5_ci(cb_2_5_io_o_5_co),
    .io_i_6_ci(cb_2_5_io_o_6_co),
    .io_i_7_ci(cb_2_5_io_o_7_co),
    .io_o_0_co(cb_2_6_io_o_0_co),
    .io_o_1_co(cb_2_6_io_o_1_co),
    .io_o_2_co(cb_2_6_io_o_2_co),
    .io_o_3_co(cb_2_6_io_o_3_co),
    .io_o_4_co(cb_2_6_io_o_4_co),
    .io_o_5_co(cb_2_6_io_o_5_co),
    .io_o_6_co(cb_2_6_io_o_6_co),
    .io_o_7_co(cb_2_6_io_o_7_co),
    .io_vci(cb_2_5_io_vco),
    .io_vco(cb_2_6_io_vco),
    .io_vi(cb_2_6_io_vi),
    .io_we_i(cb_2_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_2_0_io_adr_i[1] ,
    \cb_2_0_io_adr_i[0] }),
    .io_dat_i({\cb_2_0_io_dat_i[15] ,
    \cb_2_0_io_dat_i[14] ,
    \cb_2_0_io_dat_i[13] ,
    \cb_2_0_io_dat_i[12] ,
    \cb_2_0_io_dat_i[11] ,
    \cb_2_0_io_dat_i[10] ,
    \cb_2_0_io_dat_i[9] ,
    \cb_2_0_io_dat_i[8] ,
    \cb_2_0_io_dat_i[7] ,
    \cb_2_0_io_dat_i[6] ,
    \cb_2_0_io_dat_i[5] ,
    \cb_2_0_io_dat_i[4] ,
    \cb_2_0_io_dat_i[3] ,
    \cb_2_0_io_dat_i[2] ,
    \cb_2_0_io_dat_i[1] ,
    \cb_2_0_io_dat_i[0] }),
    .io_dat_o({\cb_2_6_io_dat_o[15] ,
    \cb_2_6_io_dat_o[14] ,
    \cb_2_6_io_dat_o[13] ,
    \cb_2_6_io_dat_o[12] ,
    \cb_2_6_io_dat_o[11] ,
    \cb_2_6_io_dat_o[10] ,
    \cb_2_6_io_dat_o[9] ,
    \cb_2_6_io_dat_o[8] ,
    \cb_2_6_io_dat_o[7] ,
    \cb_2_6_io_dat_o[6] ,
    \cb_2_6_io_dat_o[5] ,
    \cb_2_6_io_dat_o[4] ,
    \cb_2_6_io_dat_o[3] ,
    \cb_2_6_io_dat_o[2] ,
    \cb_2_6_io_dat_o[1] ,
    \cb_2_6_io_dat_o[0] }),
    .io_eo({\cb_2_6_io_eo[63] ,
    \cb_2_6_io_eo[62] ,
    \cb_2_6_io_eo[61] ,
    \cb_2_6_io_eo[60] ,
    \cb_2_6_io_eo[59] ,
    \cb_2_6_io_eo[58] ,
    \cb_2_6_io_eo[57] ,
    \cb_2_6_io_eo[56] ,
    \cb_2_6_io_eo[55] ,
    \cb_2_6_io_eo[54] ,
    \cb_2_6_io_eo[53] ,
    \cb_2_6_io_eo[52] ,
    \cb_2_6_io_eo[51] ,
    \cb_2_6_io_eo[50] ,
    \cb_2_6_io_eo[49] ,
    \cb_2_6_io_eo[48] ,
    \cb_2_6_io_eo[47] ,
    \cb_2_6_io_eo[46] ,
    \cb_2_6_io_eo[45] ,
    \cb_2_6_io_eo[44] ,
    \cb_2_6_io_eo[43] ,
    \cb_2_6_io_eo[42] ,
    \cb_2_6_io_eo[41] ,
    \cb_2_6_io_eo[40] ,
    \cb_2_6_io_eo[39] ,
    \cb_2_6_io_eo[38] ,
    \cb_2_6_io_eo[37] ,
    \cb_2_6_io_eo[36] ,
    \cb_2_6_io_eo[35] ,
    \cb_2_6_io_eo[34] ,
    \cb_2_6_io_eo[33] ,
    \cb_2_6_io_eo[32] ,
    \cb_2_6_io_eo[31] ,
    \cb_2_6_io_eo[30] ,
    \cb_2_6_io_eo[29] ,
    \cb_2_6_io_eo[28] ,
    \cb_2_6_io_eo[27] ,
    \cb_2_6_io_eo[26] ,
    \cb_2_6_io_eo[25] ,
    \cb_2_6_io_eo[24] ,
    \cb_2_6_io_eo[23] ,
    \cb_2_6_io_eo[22] ,
    \cb_2_6_io_eo[21] ,
    \cb_2_6_io_eo[20] ,
    \cb_2_6_io_eo[19] ,
    \cb_2_6_io_eo[18] ,
    \cb_2_6_io_eo[17] ,
    \cb_2_6_io_eo[16] ,
    \cb_2_6_io_eo[15] ,
    \cb_2_6_io_eo[14] ,
    \cb_2_6_io_eo[13] ,
    \cb_2_6_io_eo[12] ,
    \cb_2_6_io_eo[11] ,
    \cb_2_6_io_eo[10] ,
    \cb_2_6_io_eo[9] ,
    \cb_2_6_io_eo[8] ,
    \cb_2_6_io_eo[7] ,
    \cb_2_6_io_eo[6] ,
    \cb_2_6_io_eo[5] ,
    \cb_2_6_io_eo[4] ,
    \cb_2_6_io_eo[3] ,
    \cb_2_6_io_eo[2] ,
    \cb_2_6_io_eo[1] ,
    \cb_2_6_io_eo[0] }),
    .io_i_0_in1({\cb_2_5_io_o_0_out[7] ,
    \cb_2_5_io_o_0_out[6] ,
    \cb_2_5_io_o_0_out[5] ,
    \cb_2_5_io_o_0_out[4] ,
    \cb_2_5_io_o_0_out[3] ,
    \cb_2_5_io_o_0_out[2] ,
    \cb_2_5_io_o_0_out[1] ,
    \cb_2_5_io_o_0_out[0] }),
    .io_i_1_in1({\cb_2_5_io_o_1_out[7] ,
    \cb_2_5_io_o_1_out[6] ,
    \cb_2_5_io_o_1_out[5] ,
    \cb_2_5_io_o_1_out[4] ,
    \cb_2_5_io_o_1_out[3] ,
    \cb_2_5_io_o_1_out[2] ,
    \cb_2_5_io_o_1_out[1] ,
    \cb_2_5_io_o_1_out[0] }),
    .io_i_2_in1({\cb_2_5_io_o_2_out[7] ,
    \cb_2_5_io_o_2_out[6] ,
    \cb_2_5_io_o_2_out[5] ,
    \cb_2_5_io_o_2_out[4] ,
    \cb_2_5_io_o_2_out[3] ,
    \cb_2_5_io_o_2_out[2] ,
    \cb_2_5_io_o_2_out[1] ,
    \cb_2_5_io_o_2_out[0] }),
    .io_i_3_in1({\cb_2_5_io_o_3_out[7] ,
    \cb_2_5_io_o_3_out[6] ,
    \cb_2_5_io_o_3_out[5] ,
    \cb_2_5_io_o_3_out[4] ,
    \cb_2_5_io_o_3_out[3] ,
    \cb_2_5_io_o_3_out[2] ,
    \cb_2_5_io_o_3_out[1] ,
    \cb_2_5_io_o_3_out[0] }),
    .io_i_4_in1({\cb_2_5_io_o_4_out[7] ,
    \cb_2_5_io_o_4_out[6] ,
    \cb_2_5_io_o_4_out[5] ,
    \cb_2_5_io_o_4_out[4] ,
    \cb_2_5_io_o_4_out[3] ,
    \cb_2_5_io_o_4_out[2] ,
    \cb_2_5_io_o_4_out[1] ,
    \cb_2_5_io_o_4_out[0] }),
    .io_i_5_in1({\cb_2_5_io_o_5_out[7] ,
    \cb_2_5_io_o_5_out[6] ,
    \cb_2_5_io_o_5_out[5] ,
    \cb_2_5_io_o_5_out[4] ,
    \cb_2_5_io_o_5_out[3] ,
    \cb_2_5_io_o_5_out[2] ,
    \cb_2_5_io_o_5_out[1] ,
    \cb_2_5_io_o_5_out[0] }),
    .io_i_6_in1({\cb_2_5_io_o_6_out[7] ,
    \cb_2_5_io_o_6_out[6] ,
    \cb_2_5_io_o_6_out[5] ,
    \cb_2_5_io_o_6_out[4] ,
    \cb_2_5_io_o_6_out[3] ,
    \cb_2_5_io_o_6_out[2] ,
    \cb_2_5_io_o_6_out[1] ,
    \cb_2_5_io_o_6_out[0] }),
    .io_i_7_in1({\cb_2_5_io_o_7_out[7] ,
    \cb_2_5_io_o_7_out[6] ,
    \cb_2_5_io_o_7_out[5] ,
    \cb_2_5_io_o_7_out[4] ,
    \cb_2_5_io_o_7_out[3] ,
    \cb_2_5_io_o_7_out[2] ,
    \cb_2_5_io_o_7_out[1] ,
    \cb_2_5_io_o_7_out[0] }),
    .io_o_0_out({\cb_2_6_io_o_0_out[7] ,
    \cb_2_6_io_o_0_out[6] ,
    \cb_2_6_io_o_0_out[5] ,
    \cb_2_6_io_o_0_out[4] ,
    \cb_2_6_io_o_0_out[3] ,
    \cb_2_6_io_o_0_out[2] ,
    \cb_2_6_io_o_0_out[1] ,
    \cb_2_6_io_o_0_out[0] }),
    .io_o_1_out({\cb_2_6_io_o_1_out[7] ,
    \cb_2_6_io_o_1_out[6] ,
    \cb_2_6_io_o_1_out[5] ,
    \cb_2_6_io_o_1_out[4] ,
    \cb_2_6_io_o_1_out[3] ,
    \cb_2_6_io_o_1_out[2] ,
    \cb_2_6_io_o_1_out[1] ,
    \cb_2_6_io_o_1_out[0] }),
    .io_o_2_out({\cb_2_6_io_o_2_out[7] ,
    \cb_2_6_io_o_2_out[6] ,
    \cb_2_6_io_o_2_out[5] ,
    \cb_2_6_io_o_2_out[4] ,
    \cb_2_6_io_o_2_out[3] ,
    \cb_2_6_io_o_2_out[2] ,
    \cb_2_6_io_o_2_out[1] ,
    \cb_2_6_io_o_2_out[0] }),
    .io_o_3_out({\cb_2_6_io_o_3_out[7] ,
    \cb_2_6_io_o_3_out[6] ,
    \cb_2_6_io_o_3_out[5] ,
    \cb_2_6_io_o_3_out[4] ,
    \cb_2_6_io_o_3_out[3] ,
    \cb_2_6_io_o_3_out[2] ,
    \cb_2_6_io_o_3_out[1] ,
    \cb_2_6_io_o_3_out[0] }),
    .io_o_4_out({\cb_2_6_io_o_4_out[7] ,
    \cb_2_6_io_o_4_out[6] ,
    \cb_2_6_io_o_4_out[5] ,
    \cb_2_6_io_o_4_out[4] ,
    \cb_2_6_io_o_4_out[3] ,
    \cb_2_6_io_o_4_out[2] ,
    \cb_2_6_io_o_4_out[1] ,
    \cb_2_6_io_o_4_out[0] }),
    .io_o_5_out({\cb_2_6_io_o_5_out[7] ,
    \cb_2_6_io_o_5_out[6] ,
    \cb_2_6_io_o_5_out[5] ,
    \cb_2_6_io_o_5_out[4] ,
    \cb_2_6_io_o_5_out[3] ,
    \cb_2_6_io_o_5_out[2] ,
    \cb_2_6_io_o_5_out[1] ,
    \cb_2_6_io_o_5_out[0] }),
    .io_o_6_out({\cb_2_6_io_o_6_out[7] ,
    \cb_2_6_io_o_6_out[6] ,
    \cb_2_6_io_o_6_out[5] ,
    \cb_2_6_io_o_6_out[4] ,
    \cb_2_6_io_o_6_out[3] ,
    \cb_2_6_io_o_6_out[2] ,
    \cb_2_6_io_o_6_out[1] ,
    \cb_2_6_io_o_6_out[0] }),
    .io_o_7_out({\cb_2_6_io_o_7_out[7] ,
    \cb_2_6_io_o_7_out[6] ,
    \cb_2_6_io_o_7_out[5] ,
    \cb_2_6_io_o_7_out[4] ,
    \cb_2_6_io_o_7_out[3] ,
    \cb_2_6_io_o_7_out[2] ,
    \cb_2_6_io_o_7_out[1] ,
    \cb_2_6_io_o_7_out[0] }),
    .io_wo({\cb_2_5_io_eo[63] ,
    \cb_2_5_io_eo[62] ,
    \cb_2_5_io_eo[61] ,
    \cb_2_5_io_eo[60] ,
    \cb_2_5_io_eo[59] ,
    \cb_2_5_io_eo[58] ,
    \cb_2_5_io_eo[57] ,
    \cb_2_5_io_eo[56] ,
    \cb_2_5_io_eo[55] ,
    \cb_2_5_io_eo[54] ,
    \cb_2_5_io_eo[53] ,
    \cb_2_5_io_eo[52] ,
    \cb_2_5_io_eo[51] ,
    \cb_2_5_io_eo[50] ,
    \cb_2_5_io_eo[49] ,
    \cb_2_5_io_eo[48] ,
    \cb_2_5_io_eo[47] ,
    \cb_2_5_io_eo[46] ,
    \cb_2_5_io_eo[45] ,
    \cb_2_5_io_eo[44] ,
    \cb_2_5_io_eo[43] ,
    \cb_2_5_io_eo[42] ,
    \cb_2_5_io_eo[41] ,
    \cb_2_5_io_eo[40] ,
    \cb_2_5_io_eo[39] ,
    \cb_2_5_io_eo[38] ,
    \cb_2_5_io_eo[37] ,
    \cb_2_5_io_eo[36] ,
    \cb_2_5_io_eo[35] ,
    \cb_2_5_io_eo[34] ,
    \cb_2_5_io_eo[33] ,
    \cb_2_5_io_eo[32] ,
    \cb_2_5_io_eo[31] ,
    \cb_2_5_io_eo[30] ,
    \cb_2_5_io_eo[29] ,
    \cb_2_5_io_eo[28] ,
    \cb_2_5_io_eo[27] ,
    \cb_2_5_io_eo[26] ,
    \cb_2_5_io_eo[25] ,
    \cb_2_5_io_eo[24] ,
    \cb_2_5_io_eo[23] ,
    \cb_2_5_io_eo[22] ,
    \cb_2_5_io_eo[21] ,
    \cb_2_5_io_eo[20] ,
    \cb_2_5_io_eo[19] ,
    \cb_2_5_io_eo[18] ,
    \cb_2_5_io_eo[17] ,
    \cb_2_5_io_eo[16] ,
    \cb_2_5_io_eo[15] ,
    \cb_2_5_io_eo[14] ,
    \cb_2_5_io_eo[13] ,
    \cb_2_5_io_eo[12] ,
    \cb_2_5_io_eo[11] ,
    \cb_2_5_io_eo[10] ,
    \cb_2_5_io_eo[9] ,
    \cb_2_5_io_eo[8] ,
    \cb_2_5_io_eo[7] ,
    \cb_2_5_io_eo[6] ,
    \cb_2_5_io_eo[5] ,
    \cb_2_5_io_eo[4] ,
    \cb_2_5_io_eo[3] ,
    \cb_2_5_io_eo[2] ,
    \cb_2_5_io_eo[1] ,
    \cb_2_5_io_eo[0] }));
 cic_block cb_2_7 (.io_cs_i(cb_2_7_io_cs_i),
    .io_i_0_ci(cb_2_6_io_o_0_co),
    .io_i_1_ci(cb_2_6_io_o_1_co),
    .io_i_2_ci(cb_2_6_io_o_2_co),
    .io_i_3_ci(cb_2_6_io_o_3_co),
    .io_i_4_ci(cb_2_6_io_o_4_co),
    .io_i_5_ci(cb_2_6_io_o_5_co),
    .io_i_6_ci(cb_2_6_io_o_6_co),
    .io_i_7_ci(cb_2_6_io_o_7_co),
    .io_o_0_co(cb_2_7_io_o_0_co),
    .io_o_1_co(cb_2_7_io_o_1_co),
    .io_o_2_co(cb_2_7_io_o_2_co),
    .io_o_3_co(cb_2_7_io_o_3_co),
    .io_o_4_co(cb_2_7_io_o_4_co),
    .io_o_5_co(cb_2_7_io_o_5_co),
    .io_o_6_co(cb_2_7_io_o_6_co),
    .io_o_7_co(cb_2_7_io_o_7_co),
    .io_vci(cb_2_6_io_vco),
    .io_vco(cb_2_7_io_vco),
    .io_vi(cb_2_7_io_vi),
    .io_we_i(cb_2_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_2_0_io_adr_i[1] ,
    \cb_2_0_io_adr_i[0] }),
    .io_dat_i({\cb_2_0_io_dat_i[15] ,
    \cb_2_0_io_dat_i[14] ,
    \cb_2_0_io_dat_i[13] ,
    \cb_2_0_io_dat_i[12] ,
    \cb_2_0_io_dat_i[11] ,
    \cb_2_0_io_dat_i[10] ,
    \cb_2_0_io_dat_i[9] ,
    \cb_2_0_io_dat_i[8] ,
    \cb_2_0_io_dat_i[7] ,
    \cb_2_0_io_dat_i[6] ,
    \cb_2_0_io_dat_i[5] ,
    \cb_2_0_io_dat_i[4] ,
    \cb_2_0_io_dat_i[3] ,
    \cb_2_0_io_dat_i[2] ,
    \cb_2_0_io_dat_i[1] ,
    \cb_2_0_io_dat_i[0] }),
    .io_dat_o({\cb_2_7_io_dat_o[15] ,
    \cb_2_7_io_dat_o[14] ,
    \cb_2_7_io_dat_o[13] ,
    \cb_2_7_io_dat_o[12] ,
    \cb_2_7_io_dat_o[11] ,
    \cb_2_7_io_dat_o[10] ,
    \cb_2_7_io_dat_o[9] ,
    \cb_2_7_io_dat_o[8] ,
    \cb_2_7_io_dat_o[7] ,
    \cb_2_7_io_dat_o[6] ,
    \cb_2_7_io_dat_o[5] ,
    \cb_2_7_io_dat_o[4] ,
    \cb_2_7_io_dat_o[3] ,
    \cb_2_7_io_dat_o[2] ,
    \cb_2_7_io_dat_o[1] ,
    \cb_2_7_io_dat_o[0] }),
    .io_eo({\cb_2_7_io_eo[63] ,
    \cb_2_7_io_eo[62] ,
    \cb_2_7_io_eo[61] ,
    \cb_2_7_io_eo[60] ,
    \cb_2_7_io_eo[59] ,
    \cb_2_7_io_eo[58] ,
    \cb_2_7_io_eo[57] ,
    \cb_2_7_io_eo[56] ,
    \cb_2_7_io_eo[55] ,
    \cb_2_7_io_eo[54] ,
    \cb_2_7_io_eo[53] ,
    \cb_2_7_io_eo[52] ,
    \cb_2_7_io_eo[51] ,
    \cb_2_7_io_eo[50] ,
    \cb_2_7_io_eo[49] ,
    \cb_2_7_io_eo[48] ,
    \cb_2_7_io_eo[47] ,
    \cb_2_7_io_eo[46] ,
    \cb_2_7_io_eo[45] ,
    \cb_2_7_io_eo[44] ,
    \cb_2_7_io_eo[43] ,
    \cb_2_7_io_eo[42] ,
    \cb_2_7_io_eo[41] ,
    \cb_2_7_io_eo[40] ,
    \cb_2_7_io_eo[39] ,
    \cb_2_7_io_eo[38] ,
    \cb_2_7_io_eo[37] ,
    \cb_2_7_io_eo[36] ,
    \cb_2_7_io_eo[35] ,
    \cb_2_7_io_eo[34] ,
    \cb_2_7_io_eo[33] ,
    \cb_2_7_io_eo[32] ,
    \cb_2_7_io_eo[31] ,
    \cb_2_7_io_eo[30] ,
    \cb_2_7_io_eo[29] ,
    \cb_2_7_io_eo[28] ,
    \cb_2_7_io_eo[27] ,
    \cb_2_7_io_eo[26] ,
    \cb_2_7_io_eo[25] ,
    \cb_2_7_io_eo[24] ,
    \cb_2_7_io_eo[23] ,
    \cb_2_7_io_eo[22] ,
    \cb_2_7_io_eo[21] ,
    \cb_2_7_io_eo[20] ,
    \cb_2_7_io_eo[19] ,
    \cb_2_7_io_eo[18] ,
    \cb_2_7_io_eo[17] ,
    \cb_2_7_io_eo[16] ,
    \cb_2_7_io_eo[15] ,
    \cb_2_7_io_eo[14] ,
    \cb_2_7_io_eo[13] ,
    \cb_2_7_io_eo[12] ,
    \cb_2_7_io_eo[11] ,
    \cb_2_7_io_eo[10] ,
    \cb_2_7_io_eo[9] ,
    \cb_2_7_io_eo[8] ,
    \cb_2_7_io_eo[7] ,
    \cb_2_7_io_eo[6] ,
    \cb_2_7_io_eo[5] ,
    \cb_2_7_io_eo[4] ,
    \cb_2_7_io_eo[3] ,
    \cb_2_7_io_eo[2] ,
    \cb_2_7_io_eo[1] ,
    \cb_2_7_io_eo[0] }),
    .io_i_0_in1({\cb_2_6_io_o_0_out[7] ,
    \cb_2_6_io_o_0_out[6] ,
    \cb_2_6_io_o_0_out[5] ,
    \cb_2_6_io_o_0_out[4] ,
    \cb_2_6_io_o_0_out[3] ,
    \cb_2_6_io_o_0_out[2] ,
    \cb_2_6_io_o_0_out[1] ,
    \cb_2_6_io_o_0_out[0] }),
    .io_i_1_in1({\cb_2_6_io_o_1_out[7] ,
    \cb_2_6_io_o_1_out[6] ,
    \cb_2_6_io_o_1_out[5] ,
    \cb_2_6_io_o_1_out[4] ,
    \cb_2_6_io_o_1_out[3] ,
    \cb_2_6_io_o_1_out[2] ,
    \cb_2_6_io_o_1_out[1] ,
    \cb_2_6_io_o_1_out[0] }),
    .io_i_2_in1({\cb_2_6_io_o_2_out[7] ,
    \cb_2_6_io_o_2_out[6] ,
    \cb_2_6_io_o_2_out[5] ,
    \cb_2_6_io_o_2_out[4] ,
    \cb_2_6_io_o_2_out[3] ,
    \cb_2_6_io_o_2_out[2] ,
    \cb_2_6_io_o_2_out[1] ,
    \cb_2_6_io_o_2_out[0] }),
    .io_i_3_in1({\cb_2_6_io_o_3_out[7] ,
    \cb_2_6_io_o_3_out[6] ,
    \cb_2_6_io_o_3_out[5] ,
    \cb_2_6_io_o_3_out[4] ,
    \cb_2_6_io_o_3_out[3] ,
    \cb_2_6_io_o_3_out[2] ,
    \cb_2_6_io_o_3_out[1] ,
    \cb_2_6_io_o_3_out[0] }),
    .io_i_4_in1({\cb_2_6_io_o_4_out[7] ,
    \cb_2_6_io_o_4_out[6] ,
    \cb_2_6_io_o_4_out[5] ,
    \cb_2_6_io_o_4_out[4] ,
    \cb_2_6_io_o_4_out[3] ,
    \cb_2_6_io_o_4_out[2] ,
    \cb_2_6_io_o_4_out[1] ,
    \cb_2_6_io_o_4_out[0] }),
    .io_i_5_in1({\cb_2_6_io_o_5_out[7] ,
    \cb_2_6_io_o_5_out[6] ,
    \cb_2_6_io_o_5_out[5] ,
    \cb_2_6_io_o_5_out[4] ,
    \cb_2_6_io_o_5_out[3] ,
    \cb_2_6_io_o_5_out[2] ,
    \cb_2_6_io_o_5_out[1] ,
    \cb_2_6_io_o_5_out[0] }),
    .io_i_6_in1({\cb_2_6_io_o_6_out[7] ,
    \cb_2_6_io_o_6_out[6] ,
    \cb_2_6_io_o_6_out[5] ,
    \cb_2_6_io_o_6_out[4] ,
    \cb_2_6_io_o_6_out[3] ,
    \cb_2_6_io_o_6_out[2] ,
    \cb_2_6_io_o_6_out[1] ,
    \cb_2_6_io_o_6_out[0] }),
    .io_i_7_in1({\cb_2_6_io_o_7_out[7] ,
    \cb_2_6_io_o_7_out[6] ,
    \cb_2_6_io_o_7_out[5] ,
    \cb_2_6_io_o_7_out[4] ,
    \cb_2_6_io_o_7_out[3] ,
    \cb_2_6_io_o_7_out[2] ,
    \cb_2_6_io_o_7_out[1] ,
    \cb_2_6_io_o_7_out[0] }),
    .io_o_0_out({\cb_2_7_io_o_0_out[7] ,
    \cb_2_7_io_o_0_out[6] ,
    \cb_2_7_io_o_0_out[5] ,
    \cb_2_7_io_o_0_out[4] ,
    \cb_2_7_io_o_0_out[3] ,
    \cb_2_7_io_o_0_out[2] ,
    \cb_2_7_io_o_0_out[1] ,
    \cb_2_7_io_o_0_out[0] }),
    .io_o_1_out({\cb_2_7_io_o_1_out[7] ,
    \cb_2_7_io_o_1_out[6] ,
    \cb_2_7_io_o_1_out[5] ,
    \cb_2_7_io_o_1_out[4] ,
    \cb_2_7_io_o_1_out[3] ,
    \cb_2_7_io_o_1_out[2] ,
    \cb_2_7_io_o_1_out[1] ,
    \cb_2_7_io_o_1_out[0] }),
    .io_o_2_out({\cb_2_7_io_o_2_out[7] ,
    \cb_2_7_io_o_2_out[6] ,
    \cb_2_7_io_o_2_out[5] ,
    \cb_2_7_io_o_2_out[4] ,
    \cb_2_7_io_o_2_out[3] ,
    \cb_2_7_io_o_2_out[2] ,
    \cb_2_7_io_o_2_out[1] ,
    \cb_2_7_io_o_2_out[0] }),
    .io_o_3_out({\cb_2_7_io_o_3_out[7] ,
    \cb_2_7_io_o_3_out[6] ,
    \cb_2_7_io_o_3_out[5] ,
    \cb_2_7_io_o_3_out[4] ,
    \cb_2_7_io_o_3_out[3] ,
    \cb_2_7_io_o_3_out[2] ,
    \cb_2_7_io_o_3_out[1] ,
    \cb_2_7_io_o_3_out[0] }),
    .io_o_4_out({\cb_2_7_io_o_4_out[7] ,
    \cb_2_7_io_o_4_out[6] ,
    \cb_2_7_io_o_4_out[5] ,
    \cb_2_7_io_o_4_out[4] ,
    \cb_2_7_io_o_4_out[3] ,
    \cb_2_7_io_o_4_out[2] ,
    \cb_2_7_io_o_4_out[1] ,
    \cb_2_7_io_o_4_out[0] }),
    .io_o_5_out({\cb_2_7_io_o_5_out[7] ,
    \cb_2_7_io_o_5_out[6] ,
    \cb_2_7_io_o_5_out[5] ,
    \cb_2_7_io_o_5_out[4] ,
    \cb_2_7_io_o_5_out[3] ,
    \cb_2_7_io_o_5_out[2] ,
    \cb_2_7_io_o_5_out[1] ,
    \cb_2_7_io_o_5_out[0] }),
    .io_o_6_out({\cb_2_7_io_o_6_out[7] ,
    \cb_2_7_io_o_6_out[6] ,
    \cb_2_7_io_o_6_out[5] ,
    \cb_2_7_io_o_6_out[4] ,
    \cb_2_7_io_o_6_out[3] ,
    \cb_2_7_io_o_6_out[2] ,
    \cb_2_7_io_o_6_out[1] ,
    \cb_2_7_io_o_6_out[0] }),
    .io_o_7_out({\cb_2_7_io_o_7_out[7] ,
    \cb_2_7_io_o_7_out[6] ,
    \cb_2_7_io_o_7_out[5] ,
    \cb_2_7_io_o_7_out[4] ,
    \cb_2_7_io_o_7_out[3] ,
    \cb_2_7_io_o_7_out[2] ,
    \cb_2_7_io_o_7_out[1] ,
    \cb_2_7_io_o_7_out[0] }),
    .io_wo({\cb_2_6_io_eo[63] ,
    \cb_2_6_io_eo[62] ,
    \cb_2_6_io_eo[61] ,
    \cb_2_6_io_eo[60] ,
    \cb_2_6_io_eo[59] ,
    \cb_2_6_io_eo[58] ,
    \cb_2_6_io_eo[57] ,
    \cb_2_6_io_eo[56] ,
    \cb_2_6_io_eo[55] ,
    \cb_2_6_io_eo[54] ,
    \cb_2_6_io_eo[53] ,
    \cb_2_6_io_eo[52] ,
    \cb_2_6_io_eo[51] ,
    \cb_2_6_io_eo[50] ,
    \cb_2_6_io_eo[49] ,
    \cb_2_6_io_eo[48] ,
    \cb_2_6_io_eo[47] ,
    \cb_2_6_io_eo[46] ,
    \cb_2_6_io_eo[45] ,
    \cb_2_6_io_eo[44] ,
    \cb_2_6_io_eo[43] ,
    \cb_2_6_io_eo[42] ,
    \cb_2_6_io_eo[41] ,
    \cb_2_6_io_eo[40] ,
    \cb_2_6_io_eo[39] ,
    \cb_2_6_io_eo[38] ,
    \cb_2_6_io_eo[37] ,
    \cb_2_6_io_eo[36] ,
    \cb_2_6_io_eo[35] ,
    \cb_2_6_io_eo[34] ,
    \cb_2_6_io_eo[33] ,
    \cb_2_6_io_eo[32] ,
    \cb_2_6_io_eo[31] ,
    \cb_2_6_io_eo[30] ,
    \cb_2_6_io_eo[29] ,
    \cb_2_6_io_eo[28] ,
    \cb_2_6_io_eo[27] ,
    \cb_2_6_io_eo[26] ,
    \cb_2_6_io_eo[25] ,
    \cb_2_6_io_eo[24] ,
    \cb_2_6_io_eo[23] ,
    \cb_2_6_io_eo[22] ,
    \cb_2_6_io_eo[21] ,
    \cb_2_6_io_eo[20] ,
    \cb_2_6_io_eo[19] ,
    \cb_2_6_io_eo[18] ,
    \cb_2_6_io_eo[17] ,
    \cb_2_6_io_eo[16] ,
    \cb_2_6_io_eo[15] ,
    \cb_2_6_io_eo[14] ,
    \cb_2_6_io_eo[13] ,
    \cb_2_6_io_eo[12] ,
    \cb_2_6_io_eo[11] ,
    \cb_2_6_io_eo[10] ,
    \cb_2_6_io_eo[9] ,
    \cb_2_6_io_eo[8] ,
    \cb_2_6_io_eo[7] ,
    \cb_2_6_io_eo[6] ,
    \cb_2_6_io_eo[5] ,
    \cb_2_6_io_eo[4] ,
    \cb_2_6_io_eo[3] ,
    \cb_2_6_io_eo[2] ,
    \cb_2_6_io_eo[1] ,
    \cb_2_6_io_eo[0] }));
 cic_block cb_2_8 (.io_cs_i(cb_2_8_io_cs_i),
    .io_i_0_ci(cb_2_7_io_o_0_co),
    .io_i_1_ci(cb_2_7_io_o_1_co),
    .io_i_2_ci(cb_2_7_io_o_2_co),
    .io_i_3_ci(cb_2_7_io_o_3_co),
    .io_i_4_ci(cb_2_7_io_o_4_co),
    .io_i_5_ci(cb_2_7_io_o_5_co),
    .io_i_6_ci(cb_2_7_io_o_6_co),
    .io_i_7_ci(cb_2_7_io_o_7_co),
    .io_o_0_co(cb_2_8_io_o_0_co),
    .io_o_1_co(cb_2_8_io_o_1_co),
    .io_o_2_co(cb_2_8_io_o_2_co),
    .io_o_3_co(cb_2_8_io_o_3_co),
    .io_o_4_co(cb_2_8_io_o_4_co),
    .io_o_5_co(cb_2_8_io_o_5_co),
    .io_o_6_co(cb_2_8_io_o_6_co),
    .io_o_7_co(cb_2_8_io_o_7_co),
    .io_vci(cb_2_7_io_vco),
    .io_vco(cb_2_8_io_vco),
    .io_vi(cb_2_8_io_vi),
    .io_we_i(cb_2_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_2_0_io_adr_i[1] ,
    \cb_2_0_io_adr_i[0] }),
    .io_dat_i({\cb_2_0_io_dat_i[15] ,
    \cb_2_0_io_dat_i[14] ,
    \cb_2_0_io_dat_i[13] ,
    \cb_2_0_io_dat_i[12] ,
    \cb_2_0_io_dat_i[11] ,
    \cb_2_0_io_dat_i[10] ,
    \cb_2_0_io_dat_i[9] ,
    \cb_2_0_io_dat_i[8] ,
    \cb_2_0_io_dat_i[7] ,
    \cb_2_0_io_dat_i[6] ,
    \cb_2_0_io_dat_i[5] ,
    \cb_2_0_io_dat_i[4] ,
    \cb_2_0_io_dat_i[3] ,
    \cb_2_0_io_dat_i[2] ,
    \cb_2_0_io_dat_i[1] ,
    \cb_2_0_io_dat_i[0] }),
    .io_dat_o({\cb_2_8_io_dat_o[15] ,
    \cb_2_8_io_dat_o[14] ,
    \cb_2_8_io_dat_o[13] ,
    \cb_2_8_io_dat_o[12] ,
    \cb_2_8_io_dat_o[11] ,
    \cb_2_8_io_dat_o[10] ,
    \cb_2_8_io_dat_o[9] ,
    \cb_2_8_io_dat_o[8] ,
    \cb_2_8_io_dat_o[7] ,
    \cb_2_8_io_dat_o[6] ,
    \cb_2_8_io_dat_o[5] ,
    \cb_2_8_io_dat_o[4] ,
    \cb_2_8_io_dat_o[3] ,
    \cb_2_8_io_dat_o[2] ,
    \cb_2_8_io_dat_o[1] ,
    \cb_2_8_io_dat_o[0] }),
    .io_eo({\cb_2_8_io_eo[63] ,
    \cb_2_8_io_eo[62] ,
    \cb_2_8_io_eo[61] ,
    \cb_2_8_io_eo[60] ,
    \cb_2_8_io_eo[59] ,
    \cb_2_8_io_eo[58] ,
    \cb_2_8_io_eo[57] ,
    \cb_2_8_io_eo[56] ,
    \cb_2_8_io_eo[55] ,
    \cb_2_8_io_eo[54] ,
    \cb_2_8_io_eo[53] ,
    \cb_2_8_io_eo[52] ,
    \cb_2_8_io_eo[51] ,
    \cb_2_8_io_eo[50] ,
    \cb_2_8_io_eo[49] ,
    \cb_2_8_io_eo[48] ,
    \cb_2_8_io_eo[47] ,
    \cb_2_8_io_eo[46] ,
    \cb_2_8_io_eo[45] ,
    \cb_2_8_io_eo[44] ,
    \cb_2_8_io_eo[43] ,
    \cb_2_8_io_eo[42] ,
    \cb_2_8_io_eo[41] ,
    \cb_2_8_io_eo[40] ,
    \cb_2_8_io_eo[39] ,
    \cb_2_8_io_eo[38] ,
    \cb_2_8_io_eo[37] ,
    \cb_2_8_io_eo[36] ,
    \cb_2_8_io_eo[35] ,
    \cb_2_8_io_eo[34] ,
    \cb_2_8_io_eo[33] ,
    \cb_2_8_io_eo[32] ,
    \cb_2_8_io_eo[31] ,
    \cb_2_8_io_eo[30] ,
    \cb_2_8_io_eo[29] ,
    \cb_2_8_io_eo[28] ,
    \cb_2_8_io_eo[27] ,
    \cb_2_8_io_eo[26] ,
    \cb_2_8_io_eo[25] ,
    \cb_2_8_io_eo[24] ,
    \cb_2_8_io_eo[23] ,
    \cb_2_8_io_eo[22] ,
    \cb_2_8_io_eo[21] ,
    \cb_2_8_io_eo[20] ,
    \cb_2_8_io_eo[19] ,
    \cb_2_8_io_eo[18] ,
    \cb_2_8_io_eo[17] ,
    \cb_2_8_io_eo[16] ,
    \cb_2_8_io_eo[15] ,
    \cb_2_8_io_eo[14] ,
    \cb_2_8_io_eo[13] ,
    \cb_2_8_io_eo[12] ,
    \cb_2_8_io_eo[11] ,
    \cb_2_8_io_eo[10] ,
    \cb_2_8_io_eo[9] ,
    \cb_2_8_io_eo[8] ,
    \cb_2_8_io_eo[7] ,
    \cb_2_8_io_eo[6] ,
    \cb_2_8_io_eo[5] ,
    \cb_2_8_io_eo[4] ,
    \cb_2_8_io_eo[3] ,
    \cb_2_8_io_eo[2] ,
    \cb_2_8_io_eo[1] ,
    \cb_2_8_io_eo[0] }),
    .io_i_0_in1({\cb_2_7_io_o_0_out[7] ,
    \cb_2_7_io_o_0_out[6] ,
    \cb_2_7_io_o_0_out[5] ,
    \cb_2_7_io_o_0_out[4] ,
    \cb_2_7_io_o_0_out[3] ,
    \cb_2_7_io_o_0_out[2] ,
    \cb_2_7_io_o_0_out[1] ,
    \cb_2_7_io_o_0_out[0] }),
    .io_i_1_in1({\cb_2_7_io_o_1_out[7] ,
    \cb_2_7_io_o_1_out[6] ,
    \cb_2_7_io_o_1_out[5] ,
    \cb_2_7_io_o_1_out[4] ,
    \cb_2_7_io_o_1_out[3] ,
    \cb_2_7_io_o_1_out[2] ,
    \cb_2_7_io_o_1_out[1] ,
    \cb_2_7_io_o_1_out[0] }),
    .io_i_2_in1({\cb_2_7_io_o_2_out[7] ,
    \cb_2_7_io_o_2_out[6] ,
    \cb_2_7_io_o_2_out[5] ,
    \cb_2_7_io_o_2_out[4] ,
    \cb_2_7_io_o_2_out[3] ,
    \cb_2_7_io_o_2_out[2] ,
    \cb_2_7_io_o_2_out[1] ,
    \cb_2_7_io_o_2_out[0] }),
    .io_i_3_in1({\cb_2_7_io_o_3_out[7] ,
    \cb_2_7_io_o_3_out[6] ,
    \cb_2_7_io_o_3_out[5] ,
    \cb_2_7_io_o_3_out[4] ,
    \cb_2_7_io_o_3_out[3] ,
    \cb_2_7_io_o_3_out[2] ,
    \cb_2_7_io_o_3_out[1] ,
    \cb_2_7_io_o_3_out[0] }),
    .io_i_4_in1({\cb_2_7_io_o_4_out[7] ,
    \cb_2_7_io_o_4_out[6] ,
    \cb_2_7_io_o_4_out[5] ,
    \cb_2_7_io_o_4_out[4] ,
    \cb_2_7_io_o_4_out[3] ,
    \cb_2_7_io_o_4_out[2] ,
    \cb_2_7_io_o_4_out[1] ,
    \cb_2_7_io_o_4_out[0] }),
    .io_i_5_in1({\cb_2_7_io_o_5_out[7] ,
    \cb_2_7_io_o_5_out[6] ,
    \cb_2_7_io_o_5_out[5] ,
    \cb_2_7_io_o_5_out[4] ,
    \cb_2_7_io_o_5_out[3] ,
    \cb_2_7_io_o_5_out[2] ,
    \cb_2_7_io_o_5_out[1] ,
    \cb_2_7_io_o_5_out[0] }),
    .io_i_6_in1({\cb_2_7_io_o_6_out[7] ,
    \cb_2_7_io_o_6_out[6] ,
    \cb_2_7_io_o_6_out[5] ,
    \cb_2_7_io_o_6_out[4] ,
    \cb_2_7_io_o_6_out[3] ,
    \cb_2_7_io_o_6_out[2] ,
    \cb_2_7_io_o_6_out[1] ,
    \cb_2_7_io_o_6_out[0] }),
    .io_i_7_in1({\cb_2_7_io_o_7_out[7] ,
    \cb_2_7_io_o_7_out[6] ,
    \cb_2_7_io_o_7_out[5] ,
    \cb_2_7_io_o_7_out[4] ,
    \cb_2_7_io_o_7_out[3] ,
    \cb_2_7_io_o_7_out[2] ,
    \cb_2_7_io_o_7_out[1] ,
    \cb_2_7_io_o_7_out[0] }),
    .io_o_0_out({\cb_2_8_io_o_0_out[7] ,
    \cb_2_8_io_o_0_out[6] ,
    \cb_2_8_io_o_0_out[5] ,
    \cb_2_8_io_o_0_out[4] ,
    \cb_2_8_io_o_0_out[3] ,
    \cb_2_8_io_o_0_out[2] ,
    \cb_2_8_io_o_0_out[1] ,
    \cb_2_8_io_o_0_out[0] }),
    .io_o_1_out({\cb_2_8_io_o_1_out[7] ,
    \cb_2_8_io_o_1_out[6] ,
    \cb_2_8_io_o_1_out[5] ,
    \cb_2_8_io_o_1_out[4] ,
    \cb_2_8_io_o_1_out[3] ,
    \cb_2_8_io_o_1_out[2] ,
    \cb_2_8_io_o_1_out[1] ,
    \cb_2_8_io_o_1_out[0] }),
    .io_o_2_out({\cb_2_8_io_o_2_out[7] ,
    \cb_2_8_io_o_2_out[6] ,
    \cb_2_8_io_o_2_out[5] ,
    \cb_2_8_io_o_2_out[4] ,
    \cb_2_8_io_o_2_out[3] ,
    \cb_2_8_io_o_2_out[2] ,
    \cb_2_8_io_o_2_out[1] ,
    \cb_2_8_io_o_2_out[0] }),
    .io_o_3_out({\cb_2_8_io_o_3_out[7] ,
    \cb_2_8_io_o_3_out[6] ,
    \cb_2_8_io_o_3_out[5] ,
    \cb_2_8_io_o_3_out[4] ,
    \cb_2_8_io_o_3_out[3] ,
    \cb_2_8_io_o_3_out[2] ,
    \cb_2_8_io_o_3_out[1] ,
    \cb_2_8_io_o_3_out[0] }),
    .io_o_4_out({\cb_2_8_io_o_4_out[7] ,
    \cb_2_8_io_o_4_out[6] ,
    \cb_2_8_io_o_4_out[5] ,
    \cb_2_8_io_o_4_out[4] ,
    \cb_2_8_io_o_4_out[3] ,
    \cb_2_8_io_o_4_out[2] ,
    \cb_2_8_io_o_4_out[1] ,
    \cb_2_8_io_o_4_out[0] }),
    .io_o_5_out({\cb_2_8_io_o_5_out[7] ,
    \cb_2_8_io_o_5_out[6] ,
    \cb_2_8_io_o_5_out[5] ,
    \cb_2_8_io_o_5_out[4] ,
    \cb_2_8_io_o_5_out[3] ,
    \cb_2_8_io_o_5_out[2] ,
    \cb_2_8_io_o_5_out[1] ,
    \cb_2_8_io_o_5_out[0] }),
    .io_o_6_out({\cb_2_8_io_o_6_out[7] ,
    \cb_2_8_io_o_6_out[6] ,
    \cb_2_8_io_o_6_out[5] ,
    \cb_2_8_io_o_6_out[4] ,
    \cb_2_8_io_o_6_out[3] ,
    \cb_2_8_io_o_6_out[2] ,
    \cb_2_8_io_o_6_out[1] ,
    \cb_2_8_io_o_6_out[0] }),
    .io_o_7_out({\cb_2_8_io_o_7_out[7] ,
    \cb_2_8_io_o_7_out[6] ,
    \cb_2_8_io_o_7_out[5] ,
    \cb_2_8_io_o_7_out[4] ,
    \cb_2_8_io_o_7_out[3] ,
    \cb_2_8_io_o_7_out[2] ,
    \cb_2_8_io_o_7_out[1] ,
    \cb_2_8_io_o_7_out[0] }),
    .io_wo({\cb_2_7_io_eo[63] ,
    \cb_2_7_io_eo[62] ,
    \cb_2_7_io_eo[61] ,
    \cb_2_7_io_eo[60] ,
    \cb_2_7_io_eo[59] ,
    \cb_2_7_io_eo[58] ,
    \cb_2_7_io_eo[57] ,
    \cb_2_7_io_eo[56] ,
    \cb_2_7_io_eo[55] ,
    \cb_2_7_io_eo[54] ,
    \cb_2_7_io_eo[53] ,
    \cb_2_7_io_eo[52] ,
    \cb_2_7_io_eo[51] ,
    \cb_2_7_io_eo[50] ,
    \cb_2_7_io_eo[49] ,
    \cb_2_7_io_eo[48] ,
    \cb_2_7_io_eo[47] ,
    \cb_2_7_io_eo[46] ,
    \cb_2_7_io_eo[45] ,
    \cb_2_7_io_eo[44] ,
    \cb_2_7_io_eo[43] ,
    \cb_2_7_io_eo[42] ,
    \cb_2_7_io_eo[41] ,
    \cb_2_7_io_eo[40] ,
    \cb_2_7_io_eo[39] ,
    \cb_2_7_io_eo[38] ,
    \cb_2_7_io_eo[37] ,
    \cb_2_7_io_eo[36] ,
    \cb_2_7_io_eo[35] ,
    \cb_2_7_io_eo[34] ,
    \cb_2_7_io_eo[33] ,
    \cb_2_7_io_eo[32] ,
    \cb_2_7_io_eo[31] ,
    \cb_2_7_io_eo[30] ,
    \cb_2_7_io_eo[29] ,
    \cb_2_7_io_eo[28] ,
    \cb_2_7_io_eo[27] ,
    \cb_2_7_io_eo[26] ,
    \cb_2_7_io_eo[25] ,
    \cb_2_7_io_eo[24] ,
    \cb_2_7_io_eo[23] ,
    \cb_2_7_io_eo[22] ,
    \cb_2_7_io_eo[21] ,
    \cb_2_7_io_eo[20] ,
    \cb_2_7_io_eo[19] ,
    \cb_2_7_io_eo[18] ,
    \cb_2_7_io_eo[17] ,
    \cb_2_7_io_eo[16] ,
    \cb_2_7_io_eo[15] ,
    \cb_2_7_io_eo[14] ,
    \cb_2_7_io_eo[13] ,
    \cb_2_7_io_eo[12] ,
    \cb_2_7_io_eo[11] ,
    \cb_2_7_io_eo[10] ,
    \cb_2_7_io_eo[9] ,
    \cb_2_7_io_eo[8] ,
    \cb_2_7_io_eo[7] ,
    \cb_2_7_io_eo[6] ,
    \cb_2_7_io_eo[5] ,
    \cb_2_7_io_eo[4] ,
    \cb_2_7_io_eo[3] ,
    \cb_2_7_io_eo[2] ,
    \cb_2_7_io_eo[1] ,
    \cb_2_7_io_eo[0] }));
 cic_block cb_2_9 (.io_cs_i(cb_2_9_io_cs_i),
    .io_i_0_ci(cb_2_8_io_o_0_co),
    .io_i_1_ci(cb_2_8_io_o_1_co),
    .io_i_2_ci(cb_2_8_io_o_2_co),
    .io_i_3_ci(cb_2_8_io_o_3_co),
    .io_i_4_ci(cb_2_8_io_o_4_co),
    .io_i_5_ci(cb_2_8_io_o_5_co),
    .io_i_6_ci(cb_2_8_io_o_6_co),
    .io_i_7_ci(cb_2_8_io_o_7_co),
    .io_o_0_co(cb_2_10_io_i_0_ci),
    .io_o_1_co(cb_2_10_io_i_1_ci),
    .io_o_2_co(cb_2_10_io_i_2_ci),
    .io_o_3_co(cb_2_10_io_i_3_ci),
    .io_o_4_co(cb_2_10_io_i_4_ci),
    .io_o_5_co(cb_2_10_io_i_5_ci),
    .io_o_6_co(cb_2_10_io_i_6_ci),
    .io_o_7_co(cb_2_10_io_i_7_ci),
    .io_vci(cb_2_8_io_vco),
    .io_vco(cb_2_10_io_vci),
    .io_vi(cb_2_9_io_vi),
    .io_we_i(cb_2_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_2_0_io_adr_i[1] ,
    \cb_2_0_io_adr_i[0] }),
    .io_dat_i({\cb_2_0_io_dat_i[15] ,
    \cb_2_0_io_dat_i[14] ,
    \cb_2_0_io_dat_i[13] ,
    \cb_2_0_io_dat_i[12] ,
    \cb_2_0_io_dat_i[11] ,
    \cb_2_0_io_dat_i[10] ,
    \cb_2_0_io_dat_i[9] ,
    \cb_2_0_io_dat_i[8] ,
    \cb_2_0_io_dat_i[7] ,
    \cb_2_0_io_dat_i[6] ,
    \cb_2_0_io_dat_i[5] ,
    \cb_2_0_io_dat_i[4] ,
    \cb_2_0_io_dat_i[3] ,
    \cb_2_0_io_dat_i[2] ,
    \cb_2_0_io_dat_i[1] ,
    \cb_2_0_io_dat_i[0] }),
    .io_dat_o({\cb_2_9_io_dat_o[15] ,
    \cb_2_9_io_dat_o[14] ,
    \cb_2_9_io_dat_o[13] ,
    \cb_2_9_io_dat_o[12] ,
    \cb_2_9_io_dat_o[11] ,
    \cb_2_9_io_dat_o[10] ,
    \cb_2_9_io_dat_o[9] ,
    \cb_2_9_io_dat_o[8] ,
    \cb_2_9_io_dat_o[7] ,
    \cb_2_9_io_dat_o[6] ,
    \cb_2_9_io_dat_o[5] ,
    \cb_2_9_io_dat_o[4] ,
    \cb_2_9_io_dat_o[3] ,
    \cb_2_9_io_dat_o[2] ,
    \cb_2_9_io_dat_o[1] ,
    \cb_2_9_io_dat_o[0] }),
    .io_eo({\cb_2_10_io_wo[63] ,
    \cb_2_10_io_wo[62] ,
    \cb_2_10_io_wo[61] ,
    \cb_2_10_io_wo[60] ,
    \cb_2_10_io_wo[59] ,
    \cb_2_10_io_wo[58] ,
    \cb_2_10_io_wo[57] ,
    \cb_2_10_io_wo[56] ,
    \cb_2_10_io_wo[55] ,
    \cb_2_10_io_wo[54] ,
    \cb_2_10_io_wo[53] ,
    \cb_2_10_io_wo[52] ,
    \cb_2_10_io_wo[51] ,
    \cb_2_10_io_wo[50] ,
    \cb_2_10_io_wo[49] ,
    \cb_2_10_io_wo[48] ,
    \cb_2_10_io_wo[47] ,
    \cb_2_10_io_wo[46] ,
    \cb_2_10_io_wo[45] ,
    \cb_2_10_io_wo[44] ,
    \cb_2_10_io_wo[43] ,
    \cb_2_10_io_wo[42] ,
    \cb_2_10_io_wo[41] ,
    \cb_2_10_io_wo[40] ,
    \cb_2_10_io_wo[39] ,
    \cb_2_10_io_wo[38] ,
    \cb_2_10_io_wo[37] ,
    \cb_2_10_io_wo[36] ,
    \cb_2_10_io_wo[35] ,
    \cb_2_10_io_wo[34] ,
    \cb_2_10_io_wo[33] ,
    \cb_2_10_io_wo[32] ,
    \cb_2_10_io_wo[31] ,
    \cb_2_10_io_wo[30] ,
    \cb_2_10_io_wo[29] ,
    \cb_2_10_io_wo[28] ,
    \cb_2_10_io_wo[27] ,
    \cb_2_10_io_wo[26] ,
    \cb_2_10_io_wo[25] ,
    \cb_2_10_io_wo[24] ,
    \cb_2_10_io_wo[23] ,
    \cb_2_10_io_wo[22] ,
    \cb_2_10_io_wo[21] ,
    \cb_2_10_io_wo[20] ,
    \cb_2_10_io_wo[19] ,
    \cb_2_10_io_wo[18] ,
    \cb_2_10_io_wo[17] ,
    \cb_2_10_io_wo[16] ,
    \cb_2_10_io_wo[15] ,
    \cb_2_10_io_wo[14] ,
    \cb_2_10_io_wo[13] ,
    \cb_2_10_io_wo[12] ,
    \cb_2_10_io_wo[11] ,
    \cb_2_10_io_wo[10] ,
    \cb_2_10_io_wo[9] ,
    \cb_2_10_io_wo[8] ,
    \cb_2_10_io_wo[7] ,
    \cb_2_10_io_wo[6] ,
    \cb_2_10_io_wo[5] ,
    \cb_2_10_io_wo[4] ,
    \cb_2_10_io_wo[3] ,
    \cb_2_10_io_wo[2] ,
    \cb_2_10_io_wo[1] ,
    \cb_2_10_io_wo[0] }),
    .io_i_0_in1({\cb_2_8_io_o_0_out[7] ,
    \cb_2_8_io_o_0_out[6] ,
    \cb_2_8_io_o_0_out[5] ,
    \cb_2_8_io_o_0_out[4] ,
    \cb_2_8_io_o_0_out[3] ,
    \cb_2_8_io_o_0_out[2] ,
    \cb_2_8_io_o_0_out[1] ,
    \cb_2_8_io_o_0_out[0] }),
    .io_i_1_in1({\cb_2_8_io_o_1_out[7] ,
    \cb_2_8_io_o_1_out[6] ,
    \cb_2_8_io_o_1_out[5] ,
    \cb_2_8_io_o_1_out[4] ,
    \cb_2_8_io_o_1_out[3] ,
    \cb_2_8_io_o_1_out[2] ,
    \cb_2_8_io_o_1_out[1] ,
    \cb_2_8_io_o_1_out[0] }),
    .io_i_2_in1({\cb_2_8_io_o_2_out[7] ,
    \cb_2_8_io_o_2_out[6] ,
    \cb_2_8_io_o_2_out[5] ,
    \cb_2_8_io_o_2_out[4] ,
    \cb_2_8_io_o_2_out[3] ,
    \cb_2_8_io_o_2_out[2] ,
    \cb_2_8_io_o_2_out[1] ,
    \cb_2_8_io_o_2_out[0] }),
    .io_i_3_in1({\cb_2_8_io_o_3_out[7] ,
    \cb_2_8_io_o_3_out[6] ,
    \cb_2_8_io_o_3_out[5] ,
    \cb_2_8_io_o_3_out[4] ,
    \cb_2_8_io_o_3_out[3] ,
    \cb_2_8_io_o_3_out[2] ,
    \cb_2_8_io_o_3_out[1] ,
    \cb_2_8_io_o_3_out[0] }),
    .io_i_4_in1({\cb_2_8_io_o_4_out[7] ,
    \cb_2_8_io_o_4_out[6] ,
    \cb_2_8_io_o_4_out[5] ,
    \cb_2_8_io_o_4_out[4] ,
    \cb_2_8_io_o_4_out[3] ,
    \cb_2_8_io_o_4_out[2] ,
    \cb_2_8_io_o_4_out[1] ,
    \cb_2_8_io_o_4_out[0] }),
    .io_i_5_in1({\cb_2_8_io_o_5_out[7] ,
    \cb_2_8_io_o_5_out[6] ,
    \cb_2_8_io_o_5_out[5] ,
    \cb_2_8_io_o_5_out[4] ,
    \cb_2_8_io_o_5_out[3] ,
    \cb_2_8_io_o_5_out[2] ,
    \cb_2_8_io_o_5_out[1] ,
    \cb_2_8_io_o_5_out[0] }),
    .io_i_6_in1({\cb_2_8_io_o_6_out[7] ,
    \cb_2_8_io_o_6_out[6] ,
    \cb_2_8_io_o_6_out[5] ,
    \cb_2_8_io_o_6_out[4] ,
    \cb_2_8_io_o_6_out[3] ,
    \cb_2_8_io_o_6_out[2] ,
    \cb_2_8_io_o_6_out[1] ,
    \cb_2_8_io_o_6_out[0] }),
    .io_i_7_in1({\cb_2_8_io_o_7_out[7] ,
    \cb_2_8_io_o_7_out[6] ,
    \cb_2_8_io_o_7_out[5] ,
    \cb_2_8_io_o_7_out[4] ,
    \cb_2_8_io_o_7_out[3] ,
    \cb_2_8_io_o_7_out[2] ,
    \cb_2_8_io_o_7_out[1] ,
    \cb_2_8_io_o_7_out[0] }),
    .io_o_0_out({\cb_2_10_io_i_0_in1[7] ,
    \cb_2_10_io_i_0_in1[6] ,
    \cb_2_10_io_i_0_in1[5] ,
    \cb_2_10_io_i_0_in1[4] ,
    \cb_2_10_io_i_0_in1[3] ,
    \cb_2_10_io_i_0_in1[2] ,
    \cb_2_10_io_i_0_in1[1] ,
    \cb_2_10_io_i_0_in1[0] }),
    .io_o_1_out({\cb_2_10_io_i_1_in1[7] ,
    \cb_2_10_io_i_1_in1[6] ,
    \cb_2_10_io_i_1_in1[5] ,
    \cb_2_10_io_i_1_in1[4] ,
    \cb_2_10_io_i_1_in1[3] ,
    \cb_2_10_io_i_1_in1[2] ,
    \cb_2_10_io_i_1_in1[1] ,
    \cb_2_10_io_i_1_in1[0] }),
    .io_o_2_out({\cb_2_10_io_i_2_in1[7] ,
    \cb_2_10_io_i_2_in1[6] ,
    \cb_2_10_io_i_2_in1[5] ,
    \cb_2_10_io_i_2_in1[4] ,
    \cb_2_10_io_i_2_in1[3] ,
    \cb_2_10_io_i_2_in1[2] ,
    \cb_2_10_io_i_2_in1[1] ,
    \cb_2_10_io_i_2_in1[0] }),
    .io_o_3_out({\cb_2_10_io_i_3_in1[7] ,
    \cb_2_10_io_i_3_in1[6] ,
    \cb_2_10_io_i_3_in1[5] ,
    \cb_2_10_io_i_3_in1[4] ,
    \cb_2_10_io_i_3_in1[3] ,
    \cb_2_10_io_i_3_in1[2] ,
    \cb_2_10_io_i_3_in1[1] ,
    \cb_2_10_io_i_3_in1[0] }),
    .io_o_4_out({\cb_2_10_io_i_4_in1[7] ,
    \cb_2_10_io_i_4_in1[6] ,
    \cb_2_10_io_i_4_in1[5] ,
    \cb_2_10_io_i_4_in1[4] ,
    \cb_2_10_io_i_4_in1[3] ,
    \cb_2_10_io_i_4_in1[2] ,
    \cb_2_10_io_i_4_in1[1] ,
    \cb_2_10_io_i_4_in1[0] }),
    .io_o_5_out({\cb_2_10_io_i_5_in1[7] ,
    \cb_2_10_io_i_5_in1[6] ,
    \cb_2_10_io_i_5_in1[5] ,
    \cb_2_10_io_i_5_in1[4] ,
    \cb_2_10_io_i_5_in1[3] ,
    \cb_2_10_io_i_5_in1[2] ,
    \cb_2_10_io_i_5_in1[1] ,
    \cb_2_10_io_i_5_in1[0] }),
    .io_o_6_out({\cb_2_10_io_i_6_in1[7] ,
    \cb_2_10_io_i_6_in1[6] ,
    \cb_2_10_io_i_6_in1[5] ,
    \cb_2_10_io_i_6_in1[4] ,
    \cb_2_10_io_i_6_in1[3] ,
    \cb_2_10_io_i_6_in1[2] ,
    \cb_2_10_io_i_6_in1[1] ,
    \cb_2_10_io_i_6_in1[0] }),
    .io_o_7_out({\cb_2_10_io_i_7_in1[7] ,
    \cb_2_10_io_i_7_in1[6] ,
    \cb_2_10_io_i_7_in1[5] ,
    \cb_2_10_io_i_7_in1[4] ,
    \cb_2_10_io_i_7_in1[3] ,
    \cb_2_10_io_i_7_in1[2] ,
    \cb_2_10_io_i_7_in1[1] ,
    \cb_2_10_io_i_7_in1[0] }),
    .io_wo({\cb_2_8_io_eo[63] ,
    \cb_2_8_io_eo[62] ,
    \cb_2_8_io_eo[61] ,
    \cb_2_8_io_eo[60] ,
    \cb_2_8_io_eo[59] ,
    \cb_2_8_io_eo[58] ,
    \cb_2_8_io_eo[57] ,
    \cb_2_8_io_eo[56] ,
    \cb_2_8_io_eo[55] ,
    \cb_2_8_io_eo[54] ,
    \cb_2_8_io_eo[53] ,
    \cb_2_8_io_eo[52] ,
    \cb_2_8_io_eo[51] ,
    \cb_2_8_io_eo[50] ,
    \cb_2_8_io_eo[49] ,
    \cb_2_8_io_eo[48] ,
    \cb_2_8_io_eo[47] ,
    \cb_2_8_io_eo[46] ,
    \cb_2_8_io_eo[45] ,
    \cb_2_8_io_eo[44] ,
    \cb_2_8_io_eo[43] ,
    \cb_2_8_io_eo[42] ,
    \cb_2_8_io_eo[41] ,
    \cb_2_8_io_eo[40] ,
    \cb_2_8_io_eo[39] ,
    \cb_2_8_io_eo[38] ,
    \cb_2_8_io_eo[37] ,
    \cb_2_8_io_eo[36] ,
    \cb_2_8_io_eo[35] ,
    \cb_2_8_io_eo[34] ,
    \cb_2_8_io_eo[33] ,
    \cb_2_8_io_eo[32] ,
    \cb_2_8_io_eo[31] ,
    \cb_2_8_io_eo[30] ,
    \cb_2_8_io_eo[29] ,
    \cb_2_8_io_eo[28] ,
    \cb_2_8_io_eo[27] ,
    \cb_2_8_io_eo[26] ,
    \cb_2_8_io_eo[25] ,
    \cb_2_8_io_eo[24] ,
    \cb_2_8_io_eo[23] ,
    \cb_2_8_io_eo[22] ,
    \cb_2_8_io_eo[21] ,
    \cb_2_8_io_eo[20] ,
    \cb_2_8_io_eo[19] ,
    \cb_2_8_io_eo[18] ,
    \cb_2_8_io_eo[17] ,
    \cb_2_8_io_eo[16] ,
    \cb_2_8_io_eo[15] ,
    \cb_2_8_io_eo[14] ,
    \cb_2_8_io_eo[13] ,
    \cb_2_8_io_eo[12] ,
    \cb_2_8_io_eo[11] ,
    \cb_2_8_io_eo[10] ,
    \cb_2_8_io_eo[9] ,
    \cb_2_8_io_eo[8] ,
    \cb_2_8_io_eo[7] ,
    \cb_2_8_io_eo[6] ,
    \cb_2_8_io_eo[5] ,
    \cb_2_8_io_eo[4] ,
    \cb_2_8_io_eo[3] ,
    \cb_2_8_io_eo[2] ,
    \cb_2_8_io_eo[1] ,
    \cb_2_8_io_eo[0] }));
 cic_block cb_3_0 (.io_cs_i(cb_3_0_io_cs_i),
    .io_i_0_ci(cb_3_0_io_i_0_ci),
    .io_o_0_co(cb_3_0_io_o_0_co),
    .io_o_1_co(cb_3_0_io_o_1_co),
    .io_o_2_co(cb_3_0_io_o_2_co),
    .io_o_3_co(cb_3_0_io_o_3_co),
    .io_o_4_co(cb_3_0_io_o_4_co),
    .io_o_5_co(cb_3_0_io_o_5_co),
    .io_o_6_co(cb_3_0_io_o_6_co),
    .io_o_7_co(cb_3_0_io_o_7_co),
    .io_vco(cb_3_0_io_vco),
    .io_vi(cb_3_0_io_vi),
    .io_we_i(cb_3_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_3_0_io_adr_i[1] ,
    \cb_3_0_io_adr_i[0] }),
    .io_dat_i({\cb_3_0_io_dat_i[15] ,
    \cb_3_0_io_dat_i[14] ,
    \cb_3_0_io_dat_i[13] ,
    \cb_3_0_io_dat_i[12] ,
    \cb_3_0_io_dat_i[11] ,
    \cb_3_0_io_dat_i[10] ,
    \cb_3_0_io_dat_i[9] ,
    \cb_3_0_io_dat_i[8] ,
    \cb_3_0_io_dat_i[7] ,
    \cb_3_0_io_dat_i[6] ,
    \cb_3_0_io_dat_i[5] ,
    \cb_3_0_io_dat_i[4] ,
    \cb_3_0_io_dat_i[3] ,
    \cb_3_0_io_dat_i[2] ,
    \cb_3_0_io_dat_i[1] ,
    \cb_3_0_io_dat_i[0] }),
    .io_dat_o({\cb_3_0_io_dat_o[15] ,
    \cb_3_0_io_dat_o[14] ,
    \cb_3_0_io_dat_o[13] ,
    \cb_3_0_io_dat_o[12] ,
    \cb_3_0_io_dat_o[11] ,
    \cb_3_0_io_dat_o[10] ,
    \cb_3_0_io_dat_o[9] ,
    \cb_3_0_io_dat_o[8] ,
    \cb_3_0_io_dat_o[7] ,
    \cb_3_0_io_dat_o[6] ,
    \cb_3_0_io_dat_o[5] ,
    \cb_3_0_io_dat_o[4] ,
    \cb_3_0_io_dat_o[3] ,
    \cb_3_0_io_dat_o[2] ,
    \cb_3_0_io_dat_o[1] ,
    \cb_3_0_io_dat_o[0] }),
    .io_eo({\cb_3_0_io_eo[63] ,
    \cb_3_0_io_eo[62] ,
    \cb_3_0_io_eo[61] ,
    \cb_3_0_io_eo[60] ,
    \cb_3_0_io_eo[59] ,
    \cb_3_0_io_eo[58] ,
    \cb_3_0_io_eo[57] ,
    \cb_3_0_io_eo[56] ,
    \cb_3_0_io_eo[55] ,
    \cb_3_0_io_eo[54] ,
    \cb_3_0_io_eo[53] ,
    \cb_3_0_io_eo[52] ,
    \cb_3_0_io_eo[51] ,
    \cb_3_0_io_eo[50] ,
    \cb_3_0_io_eo[49] ,
    \cb_3_0_io_eo[48] ,
    \cb_3_0_io_eo[47] ,
    \cb_3_0_io_eo[46] ,
    \cb_3_0_io_eo[45] ,
    \cb_3_0_io_eo[44] ,
    \cb_3_0_io_eo[43] ,
    \cb_3_0_io_eo[42] ,
    \cb_3_0_io_eo[41] ,
    \cb_3_0_io_eo[40] ,
    \cb_3_0_io_eo[39] ,
    \cb_3_0_io_eo[38] ,
    \cb_3_0_io_eo[37] ,
    \cb_3_0_io_eo[36] ,
    \cb_3_0_io_eo[35] ,
    \cb_3_0_io_eo[34] ,
    \cb_3_0_io_eo[33] ,
    \cb_3_0_io_eo[32] ,
    \cb_3_0_io_eo[31] ,
    \cb_3_0_io_eo[30] ,
    \cb_3_0_io_eo[29] ,
    \cb_3_0_io_eo[28] ,
    \cb_3_0_io_eo[27] ,
    \cb_3_0_io_eo[26] ,
    \cb_3_0_io_eo[25] ,
    \cb_3_0_io_eo[24] ,
    \cb_3_0_io_eo[23] ,
    \cb_3_0_io_eo[22] ,
    \cb_3_0_io_eo[21] ,
    \cb_3_0_io_eo[20] ,
    \cb_3_0_io_eo[19] ,
    \cb_3_0_io_eo[18] ,
    \cb_3_0_io_eo[17] ,
    \cb_3_0_io_eo[16] ,
    \cb_3_0_io_eo[15] ,
    \cb_3_0_io_eo[14] ,
    \cb_3_0_io_eo[13] ,
    \cb_3_0_io_eo[12] ,
    \cb_3_0_io_eo[11] ,
    \cb_3_0_io_eo[10] ,
    \cb_3_0_io_eo[9] ,
    \cb_3_0_io_eo[8] ,
    \cb_3_0_io_eo[7] ,
    \cb_3_0_io_eo[6] ,
    \cb_3_0_io_eo[5] ,
    \cb_3_0_io_eo[4] ,
    \cb_3_0_io_eo[3] ,
    \cb_3_0_io_eo[2] ,
    \cb_3_0_io_eo[1] ,
    \cb_3_0_io_eo[0] }),
    .io_i_0_in1({_NC193,
    _NC194,
    _NC195,
    _NC196,
    _NC197,
    _NC198,
    _NC199,
    _NC200}),
    .io_i_1_in1({_NC201,
    _NC202,
    _NC203,
    _NC204,
    _NC205,
    _NC206,
    _NC207,
    _NC208}),
    .io_i_2_in1({_NC209,
    _NC210,
    _NC211,
    _NC212,
    _NC213,
    _NC214,
    _NC215,
    _NC216}),
    .io_i_3_in1({_NC217,
    _NC218,
    _NC219,
    _NC220,
    _NC221,
    _NC222,
    _NC223,
    _NC224}),
    .io_i_4_in1({_NC225,
    _NC226,
    _NC227,
    _NC228,
    _NC229,
    _NC230,
    _NC231,
    _NC232}),
    .io_i_5_in1({_NC233,
    _NC234,
    _NC235,
    _NC236,
    _NC237,
    _NC238,
    _NC239,
    _NC240}),
    .io_i_6_in1({_NC241,
    _NC242,
    _NC243,
    _NC244,
    _NC245,
    _NC246,
    _NC247,
    _NC248}),
    .io_i_7_in1({_NC249,
    _NC250,
    _NC251,
    _NC252,
    _NC253,
    _NC254,
    _NC255,
    _NC256}),
    .io_o_0_out({\cb_3_0_io_o_0_out[7] ,
    \cb_3_0_io_o_0_out[6] ,
    \cb_3_0_io_o_0_out[5] ,
    \cb_3_0_io_o_0_out[4] ,
    \cb_3_0_io_o_0_out[3] ,
    \cb_3_0_io_o_0_out[2] ,
    \cb_3_0_io_o_0_out[1] ,
    \cb_3_0_io_o_0_out[0] }),
    .io_o_1_out({\cb_3_0_io_o_1_out[7] ,
    \cb_3_0_io_o_1_out[6] ,
    \cb_3_0_io_o_1_out[5] ,
    \cb_3_0_io_o_1_out[4] ,
    \cb_3_0_io_o_1_out[3] ,
    \cb_3_0_io_o_1_out[2] ,
    \cb_3_0_io_o_1_out[1] ,
    \cb_3_0_io_o_1_out[0] }),
    .io_o_2_out({\cb_3_0_io_o_2_out[7] ,
    \cb_3_0_io_o_2_out[6] ,
    \cb_3_0_io_o_2_out[5] ,
    \cb_3_0_io_o_2_out[4] ,
    \cb_3_0_io_o_2_out[3] ,
    \cb_3_0_io_o_2_out[2] ,
    \cb_3_0_io_o_2_out[1] ,
    \cb_3_0_io_o_2_out[0] }),
    .io_o_3_out({\cb_3_0_io_o_3_out[7] ,
    \cb_3_0_io_o_3_out[6] ,
    \cb_3_0_io_o_3_out[5] ,
    \cb_3_0_io_o_3_out[4] ,
    \cb_3_0_io_o_3_out[3] ,
    \cb_3_0_io_o_3_out[2] ,
    \cb_3_0_io_o_3_out[1] ,
    \cb_3_0_io_o_3_out[0] }),
    .io_o_4_out({\cb_3_0_io_o_4_out[7] ,
    \cb_3_0_io_o_4_out[6] ,
    \cb_3_0_io_o_4_out[5] ,
    \cb_3_0_io_o_4_out[4] ,
    \cb_3_0_io_o_4_out[3] ,
    \cb_3_0_io_o_4_out[2] ,
    \cb_3_0_io_o_4_out[1] ,
    \cb_3_0_io_o_4_out[0] }),
    .io_o_5_out({\cb_3_0_io_o_5_out[7] ,
    \cb_3_0_io_o_5_out[6] ,
    \cb_3_0_io_o_5_out[5] ,
    \cb_3_0_io_o_5_out[4] ,
    \cb_3_0_io_o_5_out[3] ,
    \cb_3_0_io_o_5_out[2] ,
    \cb_3_0_io_o_5_out[1] ,
    \cb_3_0_io_o_5_out[0] }),
    .io_o_6_out({\cb_3_0_io_o_6_out[7] ,
    \cb_3_0_io_o_6_out[6] ,
    \cb_3_0_io_o_6_out[5] ,
    \cb_3_0_io_o_6_out[4] ,
    \cb_3_0_io_o_6_out[3] ,
    \cb_3_0_io_o_6_out[2] ,
    \cb_3_0_io_o_6_out[1] ,
    \cb_3_0_io_o_6_out[0] }),
    .io_o_7_out({\cb_3_0_io_o_7_out[7] ,
    \cb_3_0_io_o_7_out[6] ,
    \cb_3_0_io_o_7_out[5] ,
    \cb_3_0_io_o_7_out[4] ,
    \cb_3_0_io_o_7_out[3] ,
    \cb_3_0_io_o_7_out[2] ,
    \cb_3_0_io_o_7_out[1] ,
    \cb_3_0_io_o_7_out[0] }),
    .io_wo({\cb_3_0_io_wo[63] ,
    \cb_3_0_io_wo[62] ,
    \cb_3_0_io_wo[61] ,
    \cb_3_0_io_wo[60] ,
    \cb_3_0_io_wo[59] ,
    \cb_3_0_io_wo[58] ,
    \cb_3_0_io_wo[57] ,
    \cb_3_0_io_wo[56] ,
    \cb_3_0_io_wo[55] ,
    \cb_3_0_io_wo[54] ,
    \cb_3_0_io_wo[53] ,
    \cb_3_0_io_wo[52] ,
    \cb_3_0_io_wo[51] ,
    \cb_3_0_io_wo[50] ,
    \cb_3_0_io_wo[49] ,
    \cb_3_0_io_wo[48] ,
    \cb_3_0_io_wo[47] ,
    \cb_3_0_io_wo[46] ,
    \cb_3_0_io_wo[45] ,
    \cb_3_0_io_wo[44] ,
    \cb_3_0_io_wo[43] ,
    \cb_3_0_io_wo[42] ,
    \cb_3_0_io_wo[41] ,
    \cb_3_0_io_wo[40] ,
    \cb_3_0_io_wo[39] ,
    \cb_3_0_io_wo[38] ,
    \cb_3_0_io_wo[37] ,
    \cb_3_0_io_wo[36] ,
    \cb_3_0_io_wo[35] ,
    \cb_3_0_io_wo[34] ,
    \cb_3_0_io_wo[33] ,
    \cb_3_0_io_wo[32] ,
    \cb_3_0_io_wo[31] ,
    \cb_3_0_io_wo[30] ,
    \cb_3_0_io_wo[29] ,
    \cb_3_0_io_wo[28] ,
    \cb_3_0_io_wo[27] ,
    \cb_3_0_io_wo[26] ,
    \cb_3_0_io_wo[25] ,
    \cb_3_0_io_wo[24] ,
    \cb_3_0_io_wo[23] ,
    \cb_3_0_io_wo[22] ,
    \cb_3_0_io_wo[21] ,
    \cb_3_0_io_wo[20] ,
    \cb_3_0_io_wo[19] ,
    \cb_3_0_io_wo[18] ,
    \cb_3_0_io_wo[17] ,
    \cb_3_0_io_wo[16] ,
    \cb_3_0_io_wo[15] ,
    \cb_3_0_io_wo[14] ,
    \cb_3_0_io_wo[13] ,
    \cb_3_0_io_wo[12] ,
    \cb_3_0_io_wo[11] ,
    \cb_3_0_io_wo[10] ,
    \cb_3_0_io_wo[9] ,
    \cb_3_0_io_wo[8] ,
    \cb_3_0_io_wo[7] ,
    \cb_3_0_io_wo[6] ,
    \cb_3_0_io_wo[5] ,
    \cb_3_0_io_wo[4] ,
    \cb_3_0_io_wo[3] ,
    \cb_3_0_io_wo[2] ,
    \cb_3_0_io_wo[1] ,
    \cb_3_0_io_wo[0] }));
 cic_block cb_3_1 (.io_cs_i(cb_3_1_io_cs_i),
    .io_i_0_ci(cb_3_0_io_o_0_co),
    .io_i_1_ci(cb_3_0_io_o_1_co),
    .io_i_2_ci(cb_3_0_io_o_2_co),
    .io_i_3_ci(cb_3_0_io_o_3_co),
    .io_i_4_ci(cb_3_0_io_o_4_co),
    .io_i_5_ci(cb_3_0_io_o_5_co),
    .io_i_6_ci(cb_3_0_io_o_6_co),
    .io_i_7_ci(cb_3_0_io_o_7_co),
    .io_o_0_co(cb_3_1_io_o_0_co),
    .io_o_1_co(cb_3_1_io_o_1_co),
    .io_o_2_co(cb_3_1_io_o_2_co),
    .io_o_3_co(cb_3_1_io_o_3_co),
    .io_o_4_co(cb_3_1_io_o_4_co),
    .io_o_5_co(cb_3_1_io_o_5_co),
    .io_o_6_co(cb_3_1_io_o_6_co),
    .io_o_7_co(cb_3_1_io_o_7_co),
    .io_vci(cb_3_0_io_vco),
    .io_vco(cb_3_1_io_vco),
    .io_vi(cb_3_1_io_vi),
    .io_we_i(cb_3_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_3_0_io_adr_i[1] ,
    \cb_3_0_io_adr_i[0] }),
    .io_dat_i({\cb_3_0_io_dat_i[15] ,
    \cb_3_0_io_dat_i[14] ,
    \cb_3_0_io_dat_i[13] ,
    \cb_3_0_io_dat_i[12] ,
    \cb_3_0_io_dat_i[11] ,
    \cb_3_0_io_dat_i[10] ,
    \cb_3_0_io_dat_i[9] ,
    \cb_3_0_io_dat_i[8] ,
    \cb_3_0_io_dat_i[7] ,
    \cb_3_0_io_dat_i[6] ,
    \cb_3_0_io_dat_i[5] ,
    \cb_3_0_io_dat_i[4] ,
    \cb_3_0_io_dat_i[3] ,
    \cb_3_0_io_dat_i[2] ,
    \cb_3_0_io_dat_i[1] ,
    \cb_3_0_io_dat_i[0] }),
    .io_dat_o({\cb_3_1_io_dat_o[15] ,
    \cb_3_1_io_dat_o[14] ,
    \cb_3_1_io_dat_o[13] ,
    \cb_3_1_io_dat_o[12] ,
    \cb_3_1_io_dat_o[11] ,
    \cb_3_1_io_dat_o[10] ,
    \cb_3_1_io_dat_o[9] ,
    \cb_3_1_io_dat_o[8] ,
    \cb_3_1_io_dat_o[7] ,
    \cb_3_1_io_dat_o[6] ,
    \cb_3_1_io_dat_o[5] ,
    \cb_3_1_io_dat_o[4] ,
    \cb_3_1_io_dat_o[3] ,
    \cb_3_1_io_dat_o[2] ,
    \cb_3_1_io_dat_o[1] ,
    \cb_3_1_io_dat_o[0] }),
    .io_eo({\cb_3_1_io_eo[63] ,
    \cb_3_1_io_eo[62] ,
    \cb_3_1_io_eo[61] ,
    \cb_3_1_io_eo[60] ,
    \cb_3_1_io_eo[59] ,
    \cb_3_1_io_eo[58] ,
    \cb_3_1_io_eo[57] ,
    \cb_3_1_io_eo[56] ,
    \cb_3_1_io_eo[55] ,
    \cb_3_1_io_eo[54] ,
    \cb_3_1_io_eo[53] ,
    \cb_3_1_io_eo[52] ,
    \cb_3_1_io_eo[51] ,
    \cb_3_1_io_eo[50] ,
    \cb_3_1_io_eo[49] ,
    \cb_3_1_io_eo[48] ,
    \cb_3_1_io_eo[47] ,
    \cb_3_1_io_eo[46] ,
    \cb_3_1_io_eo[45] ,
    \cb_3_1_io_eo[44] ,
    \cb_3_1_io_eo[43] ,
    \cb_3_1_io_eo[42] ,
    \cb_3_1_io_eo[41] ,
    \cb_3_1_io_eo[40] ,
    \cb_3_1_io_eo[39] ,
    \cb_3_1_io_eo[38] ,
    \cb_3_1_io_eo[37] ,
    \cb_3_1_io_eo[36] ,
    \cb_3_1_io_eo[35] ,
    \cb_3_1_io_eo[34] ,
    \cb_3_1_io_eo[33] ,
    \cb_3_1_io_eo[32] ,
    \cb_3_1_io_eo[31] ,
    \cb_3_1_io_eo[30] ,
    \cb_3_1_io_eo[29] ,
    \cb_3_1_io_eo[28] ,
    \cb_3_1_io_eo[27] ,
    \cb_3_1_io_eo[26] ,
    \cb_3_1_io_eo[25] ,
    \cb_3_1_io_eo[24] ,
    \cb_3_1_io_eo[23] ,
    \cb_3_1_io_eo[22] ,
    \cb_3_1_io_eo[21] ,
    \cb_3_1_io_eo[20] ,
    \cb_3_1_io_eo[19] ,
    \cb_3_1_io_eo[18] ,
    \cb_3_1_io_eo[17] ,
    \cb_3_1_io_eo[16] ,
    \cb_3_1_io_eo[15] ,
    \cb_3_1_io_eo[14] ,
    \cb_3_1_io_eo[13] ,
    \cb_3_1_io_eo[12] ,
    \cb_3_1_io_eo[11] ,
    \cb_3_1_io_eo[10] ,
    \cb_3_1_io_eo[9] ,
    \cb_3_1_io_eo[8] ,
    \cb_3_1_io_eo[7] ,
    \cb_3_1_io_eo[6] ,
    \cb_3_1_io_eo[5] ,
    \cb_3_1_io_eo[4] ,
    \cb_3_1_io_eo[3] ,
    \cb_3_1_io_eo[2] ,
    \cb_3_1_io_eo[1] ,
    \cb_3_1_io_eo[0] }),
    .io_i_0_in1({\cb_3_0_io_o_0_out[7] ,
    \cb_3_0_io_o_0_out[6] ,
    \cb_3_0_io_o_0_out[5] ,
    \cb_3_0_io_o_0_out[4] ,
    \cb_3_0_io_o_0_out[3] ,
    \cb_3_0_io_o_0_out[2] ,
    \cb_3_0_io_o_0_out[1] ,
    \cb_3_0_io_o_0_out[0] }),
    .io_i_1_in1({\cb_3_0_io_o_1_out[7] ,
    \cb_3_0_io_o_1_out[6] ,
    \cb_3_0_io_o_1_out[5] ,
    \cb_3_0_io_o_1_out[4] ,
    \cb_3_0_io_o_1_out[3] ,
    \cb_3_0_io_o_1_out[2] ,
    \cb_3_0_io_o_1_out[1] ,
    \cb_3_0_io_o_1_out[0] }),
    .io_i_2_in1({\cb_3_0_io_o_2_out[7] ,
    \cb_3_0_io_o_2_out[6] ,
    \cb_3_0_io_o_2_out[5] ,
    \cb_3_0_io_o_2_out[4] ,
    \cb_3_0_io_o_2_out[3] ,
    \cb_3_0_io_o_2_out[2] ,
    \cb_3_0_io_o_2_out[1] ,
    \cb_3_0_io_o_2_out[0] }),
    .io_i_3_in1({\cb_3_0_io_o_3_out[7] ,
    \cb_3_0_io_o_3_out[6] ,
    \cb_3_0_io_o_3_out[5] ,
    \cb_3_0_io_o_3_out[4] ,
    \cb_3_0_io_o_3_out[3] ,
    \cb_3_0_io_o_3_out[2] ,
    \cb_3_0_io_o_3_out[1] ,
    \cb_3_0_io_o_3_out[0] }),
    .io_i_4_in1({\cb_3_0_io_o_4_out[7] ,
    \cb_3_0_io_o_4_out[6] ,
    \cb_3_0_io_o_4_out[5] ,
    \cb_3_0_io_o_4_out[4] ,
    \cb_3_0_io_o_4_out[3] ,
    \cb_3_0_io_o_4_out[2] ,
    \cb_3_0_io_o_4_out[1] ,
    \cb_3_0_io_o_4_out[0] }),
    .io_i_5_in1({\cb_3_0_io_o_5_out[7] ,
    \cb_3_0_io_o_5_out[6] ,
    \cb_3_0_io_o_5_out[5] ,
    \cb_3_0_io_o_5_out[4] ,
    \cb_3_0_io_o_5_out[3] ,
    \cb_3_0_io_o_5_out[2] ,
    \cb_3_0_io_o_5_out[1] ,
    \cb_3_0_io_o_5_out[0] }),
    .io_i_6_in1({\cb_3_0_io_o_6_out[7] ,
    \cb_3_0_io_o_6_out[6] ,
    \cb_3_0_io_o_6_out[5] ,
    \cb_3_0_io_o_6_out[4] ,
    \cb_3_0_io_o_6_out[3] ,
    \cb_3_0_io_o_6_out[2] ,
    \cb_3_0_io_o_6_out[1] ,
    \cb_3_0_io_o_6_out[0] }),
    .io_i_7_in1({\cb_3_0_io_o_7_out[7] ,
    \cb_3_0_io_o_7_out[6] ,
    \cb_3_0_io_o_7_out[5] ,
    \cb_3_0_io_o_7_out[4] ,
    \cb_3_0_io_o_7_out[3] ,
    \cb_3_0_io_o_7_out[2] ,
    \cb_3_0_io_o_7_out[1] ,
    \cb_3_0_io_o_7_out[0] }),
    .io_o_0_out({\cb_3_1_io_o_0_out[7] ,
    \cb_3_1_io_o_0_out[6] ,
    \cb_3_1_io_o_0_out[5] ,
    \cb_3_1_io_o_0_out[4] ,
    \cb_3_1_io_o_0_out[3] ,
    \cb_3_1_io_o_0_out[2] ,
    \cb_3_1_io_o_0_out[1] ,
    \cb_3_1_io_o_0_out[0] }),
    .io_o_1_out({\cb_3_1_io_o_1_out[7] ,
    \cb_3_1_io_o_1_out[6] ,
    \cb_3_1_io_o_1_out[5] ,
    \cb_3_1_io_o_1_out[4] ,
    \cb_3_1_io_o_1_out[3] ,
    \cb_3_1_io_o_1_out[2] ,
    \cb_3_1_io_o_1_out[1] ,
    \cb_3_1_io_o_1_out[0] }),
    .io_o_2_out({\cb_3_1_io_o_2_out[7] ,
    \cb_3_1_io_o_2_out[6] ,
    \cb_3_1_io_o_2_out[5] ,
    \cb_3_1_io_o_2_out[4] ,
    \cb_3_1_io_o_2_out[3] ,
    \cb_3_1_io_o_2_out[2] ,
    \cb_3_1_io_o_2_out[1] ,
    \cb_3_1_io_o_2_out[0] }),
    .io_o_3_out({\cb_3_1_io_o_3_out[7] ,
    \cb_3_1_io_o_3_out[6] ,
    \cb_3_1_io_o_3_out[5] ,
    \cb_3_1_io_o_3_out[4] ,
    \cb_3_1_io_o_3_out[3] ,
    \cb_3_1_io_o_3_out[2] ,
    \cb_3_1_io_o_3_out[1] ,
    \cb_3_1_io_o_3_out[0] }),
    .io_o_4_out({\cb_3_1_io_o_4_out[7] ,
    \cb_3_1_io_o_4_out[6] ,
    \cb_3_1_io_o_4_out[5] ,
    \cb_3_1_io_o_4_out[4] ,
    \cb_3_1_io_o_4_out[3] ,
    \cb_3_1_io_o_4_out[2] ,
    \cb_3_1_io_o_4_out[1] ,
    \cb_3_1_io_o_4_out[0] }),
    .io_o_5_out({\cb_3_1_io_o_5_out[7] ,
    \cb_3_1_io_o_5_out[6] ,
    \cb_3_1_io_o_5_out[5] ,
    \cb_3_1_io_o_5_out[4] ,
    \cb_3_1_io_o_5_out[3] ,
    \cb_3_1_io_o_5_out[2] ,
    \cb_3_1_io_o_5_out[1] ,
    \cb_3_1_io_o_5_out[0] }),
    .io_o_6_out({\cb_3_1_io_o_6_out[7] ,
    \cb_3_1_io_o_6_out[6] ,
    \cb_3_1_io_o_6_out[5] ,
    \cb_3_1_io_o_6_out[4] ,
    \cb_3_1_io_o_6_out[3] ,
    \cb_3_1_io_o_6_out[2] ,
    \cb_3_1_io_o_6_out[1] ,
    \cb_3_1_io_o_6_out[0] }),
    .io_o_7_out({\cb_3_1_io_o_7_out[7] ,
    \cb_3_1_io_o_7_out[6] ,
    \cb_3_1_io_o_7_out[5] ,
    \cb_3_1_io_o_7_out[4] ,
    \cb_3_1_io_o_7_out[3] ,
    \cb_3_1_io_o_7_out[2] ,
    \cb_3_1_io_o_7_out[1] ,
    \cb_3_1_io_o_7_out[0] }),
    .io_wo({\cb_3_0_io_eo[63] ,
    \cb_3_0_io_eo[62] ,
    \cb_3_0_io_eo[61] ,
    \cb_3_0_io_eo[60] ,
    \cb_3_0_io_eo[59] ,
    \cb_3_0_io_eo[58] ,
    \cb_3_0_io_eo[57] ,
    \cb_3_0_io_eo[56] ,
    \cb_3_0_io_eo[55] ,
    \cb_3_0_io_eo[54] ,
    \cb_3_0_io_eo[53] ,
    \cb_3_0_io_eo[52] ,
    \cb_3_0_io_eo[51] ,
    \cb_3_0_io_eo[50] ,
    \cb_3_0_io_eo[49] ,
    \cb_3_0_io_eo[48] ,
    \cb_3_0_io_eo[47] ,
    \cb_3_0_io_eo[46] ,
    \cb_3_0_io_eo[45] ,
    \cb_3_0_io_eo[44] ,
    \cb_3_0_io_eo[43] ,
    \cb_3_0_io_eo[42] ,
    \cb_3_0_io_eo[41] ,
    \cb_3_0_io_eo[40] ,
    \cb_3_0_io_eo[39] ,
    \cb_3_0_io_eo[38] ,
    \cb_3_0_io_eo[37] ,
    \cb_3_0_io_eo[36] ,
    \cb_3_0_io_eo[35] ,
    \cb_3_0_io_eo[34] ,
    \cb_3_0_io_eo[33] ,
    \cb_3_0_io_eo[32] ,
    \cb_3_0_io_eo[31] ,
    \cb_3_0_io_eo[30] ,
    \cb_3_0_io_eo[29] ,
    \cb_3_0_io_eo[28] ,
    \cb_3_0_io_eo[27] ,
    \cb_3_0_io_eo[26] ,
    \cb_3_0_io_eo[25] ,
    \cb_3_0_io_eo[24] ,
    \cb_3_0_io_eo[23] ,
    \cb_3_0_io_eo[22] ,
    \cb_3_0_io_eo[21] ,
    \cb_3_0_io_eo[20] ,
    \cb_3_0_io_eo[19] ,
    \cb_3_0_io_eo[18] ,
    \cb_3_0_io_eo[17] ,
    \cb_3_0_io_eo[16] ,
    \cb_3_0_io_eo[15] ,
    \cb_3_0_io_eo[14] ,
    \cb_3_0_io_eo[13] ,
    \cb_3_0_io_eo[12] ,
    \cb_3_0_io_eo[11] ,
    \cb_3_0_io_eo[10] ,
    \cb_3_0_io_eo[9] ,
    \cb_3_0_io_eo[8] ,
    \cb_3_0_io_eo[7] ,
    \cb_3_0_io_eo[6] ,
    \cb_3_0_io_eo[5] ,
    \cb_3_0_io_eo[4] ,
    \cb_3_0_io_eo[3] ,
    \cb_3_0_io_eo[2] ,
    \cb_3_0_io_eo[1] ,
    \cb_3_0_io_eo[0] }));
 cic_block cb_3_10 (.io_cs_i(cb_3_10_io_cs_i),
    .io_i_0_ci(cb_3_10_io_i_0_ci),
    .io_i_1_ci(cb_3_10_io_i_1_ci),
    .io_i_2_ci(cb_3_10_io_i_2_ci),
    .io_i_3_ci(cb_3_10_io_i_3_ci),
    .io_i_4_ci(cb_3_10_io_i_4_ci),
    .io_i_5_ci(cb_3_10_io_i_5_ci),
    .io_i_6_ci(cb_3_10_io_i_6_ci),
    .io_i_7_ci(cb_3_10_io_i_7_ci),
    .io_o_0_co(cb_3_10_io_o_0_co),
    .io_o_1_co(cb_3_10_io_o_1_co),
    .io_o_2_co(cb_3_10_io_o_2_co),
    .io_o_3_co(cb_3_10_io_o_3_co),
    .io_o_4_co(cb_3_10_io_o_4_co),
    .io_o_5_co(cb_3_10_io_o_5_co),
    .io_o_6_co(cb_3_10_io_o_6_co),
    .io_o_7_co(cb_3_10_io_o_7_co),
    .io_vci(cb_3_10_io_vci),
    .io_vco(cb_3_10_io_vco),
    .io_vi(cb_3_10_io_vi),
    .io_we_i(cb_3_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_3_0_io_adr_i[1] ,
    \cb_3_0_io_adr_i[0] }),
    .io_dat_i({\cb_3_0_io_dat_i[15] ,
    \cb_3_0_io_dat_i[14] ,
    \cb_3_0_io_dat_i[13] ,
    \cb_3_0_io_dat_i[12] ,
    \cb_3_0_io_dat_i[11] ,
    \cb_3_0_io_dat_i[10] ,
    \cb_3_0_io_dat_i[9] ,
    \cb_3_0_io_dat_i[8] ,
    \cb_3_0_io_dat_i[7] ,
    \cb_3_0_io_dat_i[6] ,
    \cb_3_0_io_dat_i[5] ,
    \cb_3_0_io_dat_i[4] ,
    \cb_3_0_io_dat_i[3] ,
    \cb_3_0_io_dat_i[2] ,
    \cb_3_0_io_dat_i[1] ,
    \cb_3_0_io_dat_i[0] }),
    .io_dat_o({\cb_3_10_io_dat_o[15] ,
    \cb_3_10_io_dat_o[14] ,
    \cb_3_10_io_dat_o[13] ,
    \cb_3_10_io_dat_o[12] ,
    \cb_3_10_io_dat_o[11] ,
    \cb_3_10_io_dat_o[10] ,
    \cb_3_10_io_dat_o[9] ,
    \cb_3_10_io_dat_o[8] ,
    \cb_3_10_io_dat_o[7] ,
    \cb_3_10_io_dat_o[6] ,
    \cb_3_10_io_dat_o[5] ,
    \cb_3_10_io_dat_o[4] ,
    \cb_3_10_io_dat_o[3] ,
    \cb_3_10_io_dat_o[2] ,
    \cb_3_10_io_dat_o[1] ,
    \cb_3_10_io_dat_o[0] }),
    .io_eo({\_T_85[31] ,
    \_T_85[30] ,
    \_T_85[29] ,
    \_T_85[28] ,
    \_T_85[27] ,
    \_T_85[26] ,
    \_T_85[25] ,
    \_T_85[24] ,
    \_T_85[23] ,
    \_T_85[22] ,
    \_T_85[21] ,
    \_T_85[20] ,
    \_T_85[19] ,
    \_T_85[18] ,
    \_T_85[17] ,
    \_T_85[16] ,
    \_T_85[15] ,
    \_T_85[14] ,
    \_T_85[13] ,
    \_T_85[12] ,
    \_T_85[11] ,
    \_T_85[10] ,
    \_T_85[9] ,
    \_T_85[8] ,
    \_T_85[7] ,
    \_T_85[6] ,
    \_T_85[5] ,
    \_T_85[4] ,
    \_T_85[3] ,
    \_T_85[2] ,
    \_T_85[1] ,
    \_T_85[0] ,
    \_T_82[31] ,
    \_T_82[30] ,
    \_T_82[29] ,
    \_T_82[28] ,
    \_T_82[27] ,
    \_T_82[26] ,
    \_T_82[25] ,
    \_T_82[24] ,
    \_T_82[23] ,
    \_T_82[22] ,
    \_T_82[21] ,
    \_T_82[20] ,
    \_T_82[19] ,
    \_T_82[18] ,
    \_T_82[17] ,
    \_T_82[16] ,
    \_T_82[15] ,
    \_T_82[14] ,
    \_T_82[13] ,
    \_T_82[12] ,
    \_T_82[11] ,
    \_T_82[10] ,
    \_T_82[9] ,
    \_T_82[8] ,
    \_T_82[7] ,
    \_T_82[6] ,
    \_T_82[5] ,
    \_T_82[4] ,
    \_T_82[3] ,
    \_T_82[2] ,
    \_T_82[1] ,
    \_T_82[0] }),
    .io_i_0_in1({\cb_3_10_io_i_0_in1[7] ,
    \cb_3_10_io_i_0_in1[6] ,
    \cb_3_10_io_i_0_in1[5] ,
    \cb_3_10_io_i_0_in1[4] ,
    \cb_3_10_io_i_0_in1[3] ,
    \cb_3_10_io_i_0_in1[2] ,
    \cb_3_10_io_i_0_in1[1] ,
    \cb_3_10_io_i_0_in1[0] }),
    .io_i_1_in1({\cb_3_10_io_i_1_in1[7] ,
    \cb_3_10_io_i_1_in1[6] ,
    \cb_3_10_io_i_1_in1[5] ,
    \cb_3_10_io_i_1_in1[4] ,
    \cb_3_10_io_i_1_in1[3] ,
    \cb_3_10_io_i_1_in1[2] ,
    \cb_3_10_io_i_1_in1[1] ,
    \cb_3_10_io_i_1_in1[0] }),
    .io_i_2_in1({\cb_3_10_io_i_2_in1[7] ,
    \cb_3_10_io_i_2_in1[6] ,
    \cb_3_10_io_i_2_in1[5] ,
    \cb_3_10_io_i_2_in1[4] ,
    \cb_3_10_io_i_2_in1[3] ,
    \cb_3_10_io_i_2_in1[2] ,
    \cb_3_10_io_i_2_in1[1] ,
    \cb_3_10_io_i_2_in1[0] }),
    .io_i_3_in1({\cb_3_10_io_i_3_in1[7] ,
    \cb_3_10_io_i_3_in1[6] ,
    \cb_3_10_io_i_3_in1[5] ,
    \cb_3_10_io_i_3_in1[4] ,
    \cb_3_10_io_i_3_in1[3] ,
    \cb_3_10_io_i_3_in1[2] ,
    \cb_3_10_io_i_3_in1[1] ,
    \cb_3_10_io_i_3_in1[0] }),
    .io_i_4_in1({\cb_3_10_io_i_4_in1[7] ,
    \cb_3_10_io_i_4_in1[6] ,
    \cb_3_10_io_i_4_in1[5] ,
    \cb_3_10_io_i_4_in1[4] ,
    \cb_3_10_io_i_4_in1[3] ,
    \cb_3_10_io_i_4_in1[2] ,
    \cb_3_10_io_i_4_in1[1] ,
    \cb_3_10_io_i_4_in1[0] }),
    .io_i_5_in1({\cb_3_10_io_i_5_in1[7] ,
    \cb_3_10_io_i_5_in1[6] ,
    \cb_3_10_io_i_5_in1[5] ,
    \cb_3_10_io_i_5_in1[4] ,
    \cb_3_10_io_i_5_in1[3] ,
    \cb_3_10_io_i_5_in1[2] ,
    \cb_3_10_io_i_5_in1[1] ,
    \cb_3_10_io_i_5_in1[0] }),
    .io_i_6_in1({\cb_3_10_io_i_6_in1[7] ,
    \cb_3_10_io_i_6_in1[6] ,
    \cb_3_10_io_i_6_in1[5] ,
    \cb_3_10_io_i_6_in1[4] ,
    \cb_3_10_io_i_6_in1[3] ,
    \cb_3_10_io_i_6_in1[2] ,
    \cb_3_10_io_i_6_in1[1] ,
    \cb_3_10_io_i_6_in1[0] }),
    .io_i_7_in1({\cb_3_10_io_i_7_in1[7] ,
    \cb_3_10_io_i_7_in1[6] ,
    \cb_3_10_io_i_7_in1[5] ,
    \cb_3_10_io_i_7_in1[4] ,
    \cb_3_10_io_i_7_in1[3] ,
    \cb_3_10_io_i_7_in1[2] ,
    \cb_3_10_io_i_7_in1[1] ,
    \cb_3_10_io_i_7_in1[0] }),
    .io_o_0_out({\_T_82[7] ,
    \_T_82[6] ,
    \_T_82[5] ,
    \_T_82[4] ,
    \_T_82[3] ,
    \_T_82[2] ,
    \_T_82[1] ,
    \_T_82[0] }),
    .io_o_1_out({\_T_82[15] ,
    \_T_82[14] ,
    \_T_82[13] ,
    \_T_82[12] ,
    \_T_82[11] ,
    \_T_82[10] ,
    \_T_82[9] ,
    \_T_82[8] }),
    .io_o_2_out({\_T_82[23] ,
    \_T_82[22] ,
    \_T_82[21] ,
    \_T_82[20] ,
    \_T_82[19] ,
    \_T_82[18] ,
    \_T_82[17] ,
    \_T_82[16] }),
    .io_o_3_out({\_T_82[31] ,
    \_T_82[30] ,
    \_T_82[29] ,
    \_T_82[28] ,
    \_T_82[27] ,
    \_T_82[26] ,
    \_T_82[25] ,
    \_T_82[24] }),
    .io_o_4_out({\_T_85[7] ,
    \_T_85[6] ,
    \_T_85[5] ,
    \_T_85[4] ,
    \_T_85[3] ,
    \_T_85[2] ,
    \_T_85[1] ,
    \_T_85[0] }),
    .io_o_5_out({\_T_85[15] ,
    \_T_85[14] ,
    \_T_85[13] ,
    \_T_85[12] ,
    \_T_85[11] ,
    \_T_85[10] ,
    \_T_85[9] ,
    \_T_85[8] }),
    .io_o_6_out({\_T_85[23] ,
    \_T_85[22] ,
    \_T_85[21] ,
    \_T_85[20] ,
    \_T_85[19] ,
    \_T_85[18] ,
    \_T_85[17] ,
    \_T_85[16] }),
    .io_o_7_out({\_T_85[31] ,
    \_T_85[30] ,
    \_T_85[29] ,
    \_T_85[28] ,
    \_T_85[27] ,
    \_T_85[26] ,
    \_T_85[25] ,
    \_T_85[24] }),
    .io_wo({\cb_3_10_io_wo[63] ,
    \cb_3_10_io_wo[62] ,
    \cb_3_10_io_wo[61] ,
    \cb_3_10_io_wo[60] ,
    \cb_3_10_io_wo[59] ,
    \cb_3_10_io_wo[58] ,
    \cb_3_10_io_wo[57] ,
    \cb_3_10_io_wo[56] ,
    \cb_3_10_io_wo[55] ,
    \cb_3_10_io_wo[54] ,
    \cb_3_10_io_wo[53] ,
    \cb_3_10_io_wo[52] ,
    \cb_3_10_io_wo[51] ,
    \cb_3_10_io_wo[50] ,
    \cb_3_10_io_wo[49] ,
    \cb_3_10_io_wo[48] ,
    \cb_3_10_io_wo[47] ,
    \cb_3_10_io_wo[46] ,
    \cb_3_10_io_wo[45] ,
    \cb_3_10_io_wo[44] ,
    \cb_3_10_io_wo[43] ,
    \cb_3_10_io_wo[42] ,
    \cb_3_10_io_wo[41] ,
    \cb_3_10_io_wo[40] ,
    \cb_3_10_io_wo[39] ,
    \cb_3_10_io_wo[38] ,
    \cb_3_10_io_wo[37] ,
    \cb_3_10_io_wo[36] ,
    \cb_3_10_io_wo[35] ,
    \cb_3_10_io_wo[34] ,
    \cb_3_10_io_wo[33] ,
    \cb_3_10_io_wo[32] ,
    \cb_3_10_io_wo[31] ,
    \cb_3_10_io_wo[30] ,
    \cb_3_10_io_wo[29] ,
    \cb_3_10_io_wo[28] ,
    \cb_3_10_io_wo[27] ,
    \cb_3_10_io_wo[26] ,
    \cb_3_10_io_wo[25] ,
    \cb_3_10_io_wo[24] ,
    \cb_3_10_io_wo[23] ,
    \cb_3_10_io_wo[22] ,
    \cb_3_10_io_wo[21] ,
    \cb_3_10_io_wo[20] ,
    \cb_3_10_io_wo[19] ,
    \cb_3_10_io_wo[18] ,
    \cb_3_10_io_wo[17] ,
    \cb_3_10_io_wo[16] ,
    \cb_3_10_io_wo[15] ,
    \cb_3_10_io_wo[14] ,
    \cb_3_10_io_wo[13] ,
    \cb_3_10_io_wo[12] ,
    \cb_3_10_io_wo[11] ,
    \cb_3_10_io_wo[10] ,
    \cb_3_10_io_wo[9] ,
    \cb_3_10_io_wo[8] ,
    \cb_3_10_io_wo[7] ,
    \cb_3_10_io_wo[6] ,
    \cb_3_10_io_wo[5] ,
    \cb_3_10_io_wo[4] ,
    \cb_3_10_io_wo[3] ,
    \cb_3_10_io_wo[2] ,
    \cb_3_10_io_wo[1] ,
    \cb_3_10_io_wo[0] }));
 cic_block cb_3_2 (.io_cs_i(cb_3_2_io_cs_i),
    .io_i_0_ci(cb_3_1_io_o_0_co),
    .io_i_1_ci(cb_3_1_io_o_1_co),
    .io_i_2_ci(cb_3_1_io_o_2_co),
    .io_i_3_ci(cb_3_1_io_o_3_co),
    .io_i_4_ci(cb_3_1_io_o_4_co),
    .io_i_5_ci(cb_3_1_io_o_5_co),
    .io_i_6_ci(cb_3_1_io_o_6_co),
    .io_i_7_ci(cb_3_1_io_o_7_co),
    .io_o_0_co(cb_3_2_io_o_0_co),
    .io_o_1_co(cb_3_2_io_o_1_co),
    .io_o_2_co(cb_3_2_io_o_2_co),
    .io_o_3_co(cb_3_2_io_o_3_co),
    .io_o_4_co(cb_3_2_io_o_4_co),
    .io_o_5_co(cb_3_2_io_o_5_co),
    .io_o_6_co(cb_3_2_io_o_6_co),
    .io_o_7_co(cb_3_2_io_o_7_co),
    .io_vci(cb_3_1_io_vco),
    .io_vco(cb_3_2_io_vco),
    .io_vi(cb_3_2_io_vi),
    .io_we_i(cb_3_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_3_0_io_adr_i[1] ,
    \cb_3_0_io_adr_i[0] }),
    .io_dat_i({\cb_3_0_io_dat_i[15] ,
    \cb_3_0_io_dat_i[14] ,
    \cb_3_0_io_dat_i[13] ,
    \cb_3_0_io_dat_i[12] ,
    \cb_3_0_io_dat_i[11] ,
    \cb_3_0_io_dat_i[10] ,
    \cb_3_0_io_dat_i[9] ,
    \cb_3_0_io_dat_i[8] ,
    \cb_3_0_io_dat_i[7] ,
    \cb_3_0_io_dat_i[6] ,
    \cb_3_0_io_dat_i[5] ,
    \cb_3_0_io_dat_i[4] ,
    \cb_3_0_io_dat_i[3] ,
    \cb_3_0_io_dat_i[2] ,
    \cb_3_0_io_dat_i[1] ,
    \cb_3_0_io_dat_i[0] }),
    .io_dat_o({\cb_3_2_io_dat_o[15] ,
    \cb_3_2_io_dat_o[14] ,
    \cb_3_2_io_dat_o[13] ,
    \cb_3_2_io_dat_o[12] ,
    \cb_3_2_io_dat_o[11] ,
    \cb_3_2_io_dat_o[10] ,
    \cb_3_2_io_dat_o[9] ,
    \cb_3_2_io_dat_o[8] ,
    \cb_3_2_io_dat_o[7] ,
    \cb_3_2_io_dat_o[6] ,
    \cb_3_2_io_dat_o[5] ,
    \cb_3_2_io_dat_o[4] ,
    \cb_3_2_io_dat_o[3] ,
    \cb_3_2_io_dat_o[2] ,
    \cb_3_2_io_dat_o[1] ,
    \cb_3_2_io_dat_o[0] }),
    .io_eo({\cb_3_2_io_eo[63] ,
    \cb_3_2_io_eo[62] ,
    \cb_3_2_io_eo[61] ,
    \cb_3_2_io_eo[60] ,
    \cb_3_2_io_eo[59] ,
    \cb_3_2_io_eo[58] ,
    \cb_3_2_io_eo[57] ,
    \cb_3_2_io_eo[56] ,
    \cb_3_2_io_eo[55] ,
    \cb_3_2_io_eo[54] ,
    \cb_3_2_io_eo[53] ,
    \cb_3_2_io_eo[52] ,
    \cb_3_2_io_eo[51] ,
    \cb_3_2_io_eo[50] ,
    \cb_3_2_io_eo[49] ,
    \cb_3_2_io_eo[48] ,
    \cb_3_2_io_eo[47] ,
    \cb_3_2_io_eo[46] ,
    \cb_3_2_io_eo[45] ,
    \cb_3_2_io_eo[44] ,
    \cb_3_2_io_eo[43] ,
    \cb_3_2_io_eo[42] ,
    \cb_3_2_io_eo[41] ,
    \cb_3_2_io_eo[40] ,
    \cb_3_2_io_eo[39] ,
    \cb_3_2_io_eo[38] ,
    \cb_3_2_io_eo[37] ,
    \cb_3_2_io_eo[36] ,
    \cb_3_2_io_eo[35] ,
    \cb_3_2_io_eo[34] ,
    \cb_3_2_io_eo[33] ,
    \cb_3_2_io_eo[32] ,
    \cb_3_2_io_eo[31] ,
    \cb_3_2_io_eo[30] ,
    \cb_3_2_io_eo[29] ,
    \cb_3_2_io_eo[28] ,
    \cb_3_2_io_eo[27] ,
    \cb_3_2_io_eo[26] ,
    \cb_3_2_io_eo[25] ,
    \cb_3_2_io_eo[24] ,
    \cb_3_2_io_eo[23] ,
    \cb_3_2_io_eo[22] ,
    \cb_3_2_io_eo[21] ,
    \cb_3_2_io_eo[20] ,
    \cb_3_2_io_eo[19] ,
    \cb_3_2_io_eo[18] ,
    \cb_3_2_io_eo[17] ,
    \cb_3_2_io_eo[16] ,
    \cb_3_2_io_eo[15] ,
    \cb_3_2_io_eo[14] ,
    \cb_3_2_io_eo[13] ,
    \cb_3_2_io_eo[12] ,
    \cb_3_2_io_eo[11] ,
    \cb_3_2_io_eo[10] ,
    \cb_3_2_io_eo[9] ,
    \cb_3_2_io_eo[8] ,
    \cb_3_2_io_eo[7] ,
    \cb_3_2_io_eo[6] ,
    \cb_3_2_io_eo[5] ,
    \cb_3_2_io_eo[4] ,
    \cb_3_2_io_eo[3] ,
    \cb_3_2_io_eo[2] ,
    \cb_3_2_io_eo[1] ,
    \cb_3_2_io_eo[0] }),
    .io_i_0_in1({\cb_3_1_io_o_0_out[7] ,
    \cb_3_1_io_o_0_out[6] ,
    \cb_3_1_io_o_0_out[5] ,
    \cb_3_1_io_o_0_out[4] ,
    \cb_3_1_io_o_0_out[3] ,
    \cb_3_1_io_o_0_out[2] ,
    \cb_3_1_io_o_0_out[1] ,
    \cb_3_1_io_o_0_out[0] }),
    .io_i_1_in1({\cb_3_1_io_o_1_out[7] ,
    \cb_3_1_io_o_1_out[6] ,
    \cb_3_1_io_o_1_out[5] ,
    \cb_3_1_io_o_1_out[4] ,
    \cb_3_1_io_o_1_out[3] ,
    \cb_3_1_io_o_1_out[2] ,
    \cb_3_1_io_o_1_out[1] ,
    \cb_3_1_io_o_1_out[0] }),
    .io_i_2_in1({\cb_3_1_io_o_2_out[7] ,
    \cb_3_1_io_o_2_out[6] ,
    \cb_3_1_io_o_2_out[5] ,
    \cb_3_1_io_o_2_out[4] ,
    \cb_3_1_io_o_2_out[3] ,
    \cb_3_1_io_o_2_out[2] ,
    \cb_3_1_io_o_2_out[1] ,
    \cb_3_1_io_o_2_out[0] }),
    .io_i_3_in1({\cb_3_1_io_o_3_out[7] ,
    \cb_3_1_io_o_3_out[6] ,
    \cb_3_1_io_o_3_out[5] ,
    \cb_3_1_io_o_3_out[4] ,
    \cb_3_1_io_o_3_out[3] ,
    \cb_3_1_io_o_3_out[2] ,
    \cb_3_1_io_o_3_out[1] ,
    \cb_3_1_io_o_3_out[0] }),
    .io_i_4_in1({\cb_3_1_io_o_4_out[7] ,
    \cb_3_1_io_o_4_out[6] ,
    \cb_3_1_io_o_4_out[5] ,
    \cb_3_1_io_o_4_out[4] ,
    \cb_3_1_io_o_4_out[3] ,
    \cb_3_1_io_o_4_out[2] ,
    \cb_3_1_io_o_4_out[1] ,
    \cb_3_1_io_o_4_out[0] }),
    .io_i_5_in1({\cb_3_1_io_o_5_out[7] ,
    \cb_3_1_io_o_5_out[6] ,
    \cb_3_1_io_o_5_out[5] ,
    \cb_3_1_io_o_5_out[4] ,
    \cb_3_1_io_o_5_out[3] ,
    \cb_3_1_io_o_5_out[2] ,
    \cb_3_1_io_o_5_out[1] ,
    \cb_3_1_io_o_5_out[0] }),
    .io_i_6_in1({\cb_3_1_io_o_6_out[7] ,
    \cb_3_1_io_o_6_out[6] ,
    \cb_3_1_io_o_6_out[5] ,
    \cb_3_1_io_o_6_out[4] ,
    \cb_3_1_io_o_6_out[3] ,
    \cb_3_1_io_o_6_out[2] ,
    \cb_3_1_io_o_6_out[1] ,
    \cb_3_1_io_o_6_out[0] }),
    .io_i_7_in1({\cb_3_1_io_o_7_out[7] ,
    \cb_3_1_io_o_7_out[6] ,
    \cb_3_1_io_o_7_out[5] ,
    \cb_3_1_io_o_7_out[4] ,
    \cb_3_1_io_o_7_out[3] ,
    \cb_3_1_io_o_7_out[2] ,
    \cb_3_1_io_o_7_out[1] ,
    \cb_3_1_io_o_7_out[0] }),
    .io_o_0_out({\cb_3_2_io_o_0_out[7] ,
    \cb_3_2_io_o_0_out[6] ,
    \cb_3_2_io_o_0_out[5] ,
    \cb_3_2_io_o_0_out[4] ,
    \cb_3_2_io_o_0_out[3] ,
    \cb_3_2_io_o_0_out[2] ,
    \cb_3_2_io_o_0_out[1] ,
    \cb_3_2_io_o_0_out[0] }),
    .io_o_1_out({\cb_3_2_io_o_1_out[7] ,
    \cb_3_2_io_o_1_out[6] ,
    \cb_3_2_io_o_1_out[5] ,
    \cb_3_2_io_o_1_out[4] ,
    \cb_3_2_io_o_1_out[3] ,
    \cb_3_2_io_o_1_out[2] ,
    \cb_3_2_io_o_1_out[1] ,
    \cb_3_2_io_o_1_out[0] }),
    .io_o_2_out({\cb_3_2_io_o_2_out[7] ,
    \cb_3_2_io_o_2_out[6] ,
    \cb_3_2_io_o_2_out[5] ,
    \cb_3_2_io_o_2_out[4] ,
    \cb_3_2_io_o_2_out[3] ,
    \cb_3_2_io_o_2_out[2] ,
    \cb_3_2_io_o_2_out[1] ,
    \cb_3_2_io_o_2_out[0] }),
    .io_o_3_out({\cb_3_2_io_o_3_out[7] ,
    \cb_3_2_io_o_3_out[6] ,
    \cb_3_2_io_o_3_out[5] ,
    \cb_3_2_io_o_3_out[4] ,
    \cb_3_2_io_o_3_out[3] ,
    \cb_3_2_io_o_3_out[2] ,
    \cb_3_2_io_o_3_out[1] ,
    \cb_3_2_io_o_3_out[0] }),
    .io_o_4_out({\cb_3_2_io_o_4_out[7] ,
    \cb_3_2_io_o_4_out[6] ,
    \cb_3_2_io_o_4_out[5] ,
    \cb_3_2_io_o_4_out[4] ,
    \cb_3_2_io_o_4_out[3] ,
    \cb_3_2_io_o_4_out[2] ,
    \cb_3_2_io_o_4_out[1] ,
    \cb_3_2_io_o_4_out[0] }),
    .io_o_5_out({\cb_3_2_io_o_5_out[7] ,
    \cb_3_2_io_o_5_out[6] ,
    \cb_3_2_io_o_5_out[5] ,
    \cb_3_2_io_o_5_out[4] ,
    \cb_3_2_io_o_5_out[3] ,
    \cb_3_2_io_o_5_out[2] ,
    \cb_3_2_io_o_5_out[1] ,
    \cb_3_2_io_o_5_out[0] }),
    .io_o_6_out({\cb_3_2_io_o_6_out[7] ,
    \cb_3_2_io_o_6_out[6] ,
    \cb_3_2_io_o_6_out[5] ,
    \cb_3_2_io_o_6_out[4] ,
    \cb_3_2_io_o_6_out[3] ,
    \cb_3_2_io_o_6_out[2] ,
    \cb_3_2_io_o_6_out[1] ,
    \cb_3_2_io_o_6_out[0] }),
    .io_o_7_out({\cb_3_2_io_o_7_out[7] ,
    \cb_3_2_io_o_7_out[6] ,
    \cb_3_2_io_o_7_out[5] ,
    \cb_3_2_io_o_7_out[4] ,
    \cb_3_2_io_o_7_out[3] ,
    \cb_3_2_io_o_7_out[2] ,
    \cb_3_2_io_o_7_out[1] ,
    \cb_3_2_io_o_7_out[0] }),
    .io_wo({\cb_3_1_io_eo[63] ,
    \cb_3_1_io_eo[62] ,
    \cb_3_1_io_eo[61] ,
    \cb_3_1_io_eo[60] ,
    \cb_3_1_io_eo[59] ,
    \cb_3_1_io_eo[58] ,
    \cb_3_1_io_eo[57] ,
    \cb_3_1_io_eo[56] ,
    \cb_3_1_io_eo[55] ,
    \cb_3_1_io_eo[54] ,
    \cb_3_1_io_eo[53] ,
    \cb_3_1_io_eo[52] ,
    \cb_3_1_io_eo[51] ,
    \cb_3_1_io_eo[50] ,
    \cb_3_1_io_eo[49] ,
    \cb_3_1_io_eo[48] ,
    \cb_3_1_io_eo[47] ,
    \cb_3_1_io_eo[46] ,
    \cb_3_1_io_eo[45] ,
    \cb_3_1_io_eo[44] ,
    \cb_3_1_io_eo[43] ,
    \cb_3_1_io_eo[42] ,
    \cb_3_1_io_eo[41] ,
    \cb_3_1_io_eo[40] ,
    \cb_3_1_io_eo[39] ,
    \cb_3_1_io_eo[38] ,
    \cb_3_1_io_eo[37] ,
    \cb_3_1_io_eo[36] ,
    \cb_3_1_io_eo[35] ,
    \cb_3_1_io_eo[34] ,
    \cb_3_1_io_eo[33] ,
    \cb_3_1_io_eo[32] ,
    \cb_3_1_io_eo[31] ,
    \cb_3_1_io_eo[30] ,
    \cb_3_1_io_eo[29] ,
    \cb_3_1_io_eo[28] ,
    \cb_3_1_io_eo[27] ,
    \cb_3_1_io_eo[26] ,
    \cb_3_1_io_eo[25] ,
    \cb_3_1_io_eo[24] ,
    \cb_3_1_io_eo[23] ,
    \cb_3_1_io_eo[22] ,
    \cb_3_1_io_eo[21] ,
    \cb_3_1_io_eo[20] ,
    \cb_3_1_io_eo[19] ,
    \cb_3_1_io_eo[18] ,
    \cb_3_1_io_eo[17] ,
    \cb_3_1_io_eo[16] ,
    \cb_3_1_io_eo[15] ,
    \cb_3_1_io_eo[14] ,
    \cb_3_1_io_eo[13] ,
    \cb_3_1_io_eo[12] ,
    \cb_3_1_io_eo[11] ,
    \cb_3_1_io_eo[10] ,
    \cb_3_1_io_eo[9] ,
    \cb_3_1_io_eo[8] ,
    \cb_3_1_io_eo[7] ,
    \cb_3_1_io_eo[6] ,
    \cb_3_1_io_eo[5] ,
    \cb_3_1_io_eo[4] ,
    \cb_3_1_io_eo[3] ,
    \cb_3_1_io_eo[2] ,
    \cb_3_1_io_eo[1] ,
    \cb_3_1_io_eo[0] }));
 cic_block cb_3_3 (.io_cs_i(cb_3_3_io_cs_i),
    .io_i_0_ci(cb_3_2_io_o_0_co),
    .io_i_1_ci(cb_3_2_io_o_1_co),
    .io_i_2_ci(cb_3_2_io_o_2_co),
    .io_i_3_ci(cb_3_2_io_o_3_co),
    .io_i_4_ci(cb_3_2_io_o_4_co),
    .io_i_5_ci(cb_3_2_io_o_5_co),
    .io_i_6_ci(cb_3_2_io_o_6_co),
    .io_i_7_ci(cb_3_2_io_o_7_co),
    .io_o_0_co(cb_3_3_io_o_0_co),
    .io_o_1_co(cb_3_3_io_o_1_co),
    .io_o_2_co(cb_3_3_io_o_2_co),
    .io_o_3_co(cb_3_3_io_o_3_co),
    .io_o_4_co(cb_3_3_io_o_4_co),
    .io_o_5_co(cb_3_3_io_o_5_co),
    .io_o_6_co(cb_3_3_io_o_6_co),
    .io_o_7_co(cb_3_3_io_o_7_co),
    .io_vci(cb_3_2_io_vco),
    .io_vco(cb_3_3_io_vco),
    .io_vi(cb_3_3_io_vi),
    .io_we_i(cb_3_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_3_0_io_adr_i[1] ,
    \cb_3_0_io_adr_i[0] }),
    .io_dat_i({\cb_3_0_io_dat_i[15] ,
    \cb_3_0_io_dat_i[14] ,
    \cb_3_0_io_dat_i[13] ,
    \cb_3_0_io_dat_i[12] ,
    \cb_3_0_io_dat_i[11] ,
    \cb_3_0_io_dat_i[10] ,
    \cb_3_0_io_dat_i[9] ,
    \cb_3_0_io_dat_i[8] ,
    \cb_3_0_io_dat_i[7] ,
    \cb_3_0_io_dat_i[6] ,
    \cb_3_0_io_dat_i[5] ,
    \cb_3_0_io_dat_i[4] ,
    \cb_3_0_io_dat_i[3] ,
    \cb_3_0_io_dat_i[2] ,
    \cb_3_0_io_dat_i[1] ,
    \cb_3_0_io_dat_i[0] }),
    .io_dat_o({\cb_3_3_io_dat_o[15] ,
    \cb_3_3_io_dat_o[14] ,
    \cb_3_3_io_dat_o[13] ,
    \cb_3_3_io_dat_o[12] ,
    \cb_3_3_io_dat_o[11] ,
    \cb_3_3_io_dat_o[10] ,
    \cb_3_3_io_dat_o[9] ,
    \cb_3_3_io_dat_o[8] ,
    \cb_3_3_io_dat_o[7] ,
    \cb_3_3_io_dat_o[6] ,
    \cb_3_3_io_dat_o[5] ,
    \cb_3_3_io_dat_o[4] ,
    \cb_3_3_io_dat_o[3] ,
    \cb_3_3_io_dat_o[2] ,
    \cb_3_3_io_dat_o[1] ,
    \cb_3_3_io_dat_o[0] }),
    .io_eo({\cb_3_3_io_eo[63] ,
    \cb_3_3_io_eo[62] ,
    \cb_3_3_io_eo[61] ,
    \cb_3_3_io_eo[60] ,
    \cb_3_3_io_eo[59] ,
    \cb_3_3_io_eo[58] ,
    \cb_3_3_io_eo[57] ,
    \cb_3_3_io_eo[56] ,
    \cb_3_3_io_eo[55] ,
    \cb_3_3_io_eo[54] ,
    \cb_3_3_io_eo[53] ,
    \cb_3_3_io_eo[52] ,
    \cb_3_3_io_eo[51] ,
    \cb_3_3_io_eo[50] ,
    \cb_3_3_io_eo[49] ,
    \cb_3_3_io_eo[48] ,
    \cb_3_3_io_eo[47] ,
    \cb_3_3_io_eo[46] ,
    \cb_3_3_io_eo[45] ,
    \cb_3_3_io_eo[44] ,
    \cb_3_3_io_eo[43] ,
    \cb_3_3_io_eo[42] ,
    \cb_3_3_io_eo[41] ,
    \cb_3_3_io_eo[40] ,
    \cb_3_3_io_eo[39] ,
    \cb_3_3_io_eo[38] ,
    \cb_3_3_io_eo[37] ,
    \cb_3_3_io_eo[36] ,
    \cb_3_3_io_eo[35] ,
    \cb_3_3_io_eo[34] ,
    \cb_3_3_io_eo[33] ,
    \cb_3_3_io_eo[32] ,
    \cb_3_3_io_eo[31] ,
    \cb_3_3_io_eo[30] ,
    \cb_3_3_io_eo[29] ,
    \cb_3_3_io_eo[28] ,
    \cb_3_3_io_eo[27] ,
    \cb_3_3_io_eo[26] ,
    \cb_3_3_io_eo[25] ,
    \cb_3_3_io_eo[24] ,
    \cb_3_3_io_eo[23] ,
    \cb_3_3_io_eo[22] ,
    \cb_3_3_io_eo[21] ,
    \cb_3_3_io_eo[20] ,
    \cb_3_3_io_eo[19] ,
    \cb_3_3_io_eo[18] ,
    \cb_3_3_io_eo[17] ,
    \cb_3_3_io_eo[16] ,
    \cb_3_3_io_eo[15] ,
    \cb_3_3_io_eo[14] ,
    \cb_3_3_io_eo[13] ,
    \cb_3_3_io_eo[12] ,
    \cb_3_3_io_eo[11] ,
    \cb_3_3_io_eo[10] ,
    \cb_3_3_io_eo[9] ,
    \cb_3_3_io_eo[8] ,
    \cb_3_3_io_eo[7] ,
    \cb_3_3_io_eo[6] ,
    \cb_3_3_io_eo[5] ,
    \cb_3_3_io_eo[4] ,
    \cb_3_3_io_eo[3] ,
    \cb_3_3_io_eo[2] ,
    \cb_3_3_io_eo[1] ,
    \cb_3_3_io_eo[0] }),
    .io_i_0_in1({\cb_3_2_io_o_0_out[7] ,
    \cb_3_2_io_o_0_out[6] ,
    \cb_3_2_io_o_0_out[5] ,
    \cb_3_2_io_o_0_out[4] ,
    \cb_3_2_io_o_0_out[3] ,
    \cb_3_2_io_o_0_out[2] ,
    \cb_3_2_io_o_0_out[1] ,
    \cb_3_2_io_o_0_out[0] }),
    .io_i_1_in1({\cb_3_2_io_o_1_out[7] ,
    \cb_3_2_io_o_1_out[6] ,
    \cb_3_2_io_o_1_out[5] ,
    \cb_3_2_io_o_1_out[4] ,
    \cb_3_2_io_o_1_out[3] ,
    \cb_3_2_io_o_1_out[2] ,
    \cb_3_2_io_o_1_out[1] ,
    \cb_3_2_io_o_1_out[0] }),
    .io_i_2_in1({\cb_3_2_io_o_2_out[7] ,
    \cb_3_2_io_o_2_out[6] ,
    \cb_3_2_io_o_2_out[5] ,
    \cb_3_2_io_o_2_out[4] ,
    \cb_3_2_io_o_2_out[3] ,
    \cb_3_2_io_o_2_out[2] ,
    \cb_3_2_io_o_2_out[1] ,
    \cb_3_2_io_o_2_out[0] }),
    .io_i_3_in1({\cb_3_2_io_o_3_out[7] ,
    \cb_3_2_io_o_3_out[6] ,
    \cb_3_2_io_o_3_out[5] ,
    \cb_3_2_io_o_3_out[4] ,
    \cb_3_2_io_o_3_out[3] ,
    \cb_3_2_io_o_3_out[2] ,
    \cb_3_2_io_o_3_out[1] ,
    \cb_3_2_io_o_3_out[0] }),
    .io_i_4_in1({\cb_3_2_io_o_4_out[7] ,
    \cb_3_2_io_o_4_out[6] ,
    \cb_3_2_io_o_4_out[5] ,
    \cb_3_2_io_o_4_out[4] ,
    \cb_3_2_io_o_4_out[3] ,
    \cb_3_2_io_o_4_out[2] ,
    \cb_3_2_io_o_4_out[1] ,
    \cb_3_2_io_o_4_out[0] }),
    .io_i_5_in1({\cb_3_2_io_o_5_out[7] ,
    \cb_3_2_io_o_5_out[6] ,
    \cb_3_2_io_o_5_out[5] ,
    \cb_3_2_io_o_5_out[4] ,
    \cb_3_2_io_o_5_out[3] ,
    \cb_3_2_io_o_5_out[2] ,
    \cb_3_2_io_o_5_out[1] ,
    \cb_3_2_io_o_5_out[0] }),
    .io_i_6_in1({\cb_3_2_io_o_6_out[7] ,
    \cb_3_2_io_o_6_out[6] ,
    \cb_3_2_io_o_6_out[5] ,
    \cb_3_2_io_o_6_out[4] ,
    \cb_3_2_io_o_6_out[3] ,
    \cb_3_2_io_o_6_out[2] ,
    \cb_3_2_io_o_6_out[1] ,
    \cb_3_2_io_o_6_out[0] }),
    .io_i_7_in1({\cb_3_2_io_o_7_out[7] ,
    \cb_3_2_io_o_7_out[6] ,
    \cb_3_2_io_o_7_out[5] ,
    \cb_3_2_io_o_7_out[4] ,
    \cb_3_2_io_o_7_out[3] ,
    \cb_3_2_io_o_7_out[2] ,
    \cb_3_2_io_o_7_out[1] ,
    \cb_3_2_io_o_7_out[0] }),
    .io_o_0_out({\cb_3_3_io_o_0_out[7] ,
    \cb_3_3_io_o_0_out[6] ,
    \cb_3_3_io_o_0_out[5] ,
    \cb_3_3_io_o_0_out[4] ,
    \cb_3_3_io_o_0_out[3] ,
    \cb_3_3_io_o_0_out[2] ,
    \cb_3_3_io_o_0_out[1] ,
    \cb_3_3_io_o_0_out[0] }),
    .io_o_1_out({\cb_3_3_io_o_1_out[7] ,
    \cb_3_3_io_o_1_out[6] ,
    \cb_3_3_io_o_1_out[5] ,
    \cb_3_3_io_o_1_out[4] ,
    \cb_3_3_io_o_1_out[3] ,
    \cb_3_3_io_o_1_out[2] ,
    \cb_3_3_io_o_1_out[1] ,
    \cb_3_3_io_o_1_out[0] }),
    .io_o_2_out({\cb_3_3_io_o_2_out[7] ,
    \cb_3_3_io_o_2_out[6] ,
    \cb_3_3_io_o_2_out[5] ,
    \cb_3_3_io_o_2_out[4] ,
    \cb_3_3_io_o_2_out[3] ,
    \cb_3_3_io_o_2_out[2] ,
    \cb_3_3_io_o_2_out[1] ,
    \cb_3_3_io_o_2_out[0] }),
    .io_o_3_out({\cb_3_3_io_o_3_out[7] ,
    \cb_3_3_io_o_3_out[6] ,
    \cb_3_3_io_o_3_out[5] ,
    \cb_3_3_io_o_3_out[4] ,
    \cb_3_3_io_o_3_out[3] ,
    \cb_3_3_io_o_3_out[2] ,
    \cb_3_3_io_o_3_out[1] ,
    \cb_3_3_io_o_3_out[0] }),
    .io_o_4_out({\cb_3_3_io_o_4_out[7] ,
    \cb_3_3_io_o_4_out[6] ,
    \cb_3_3_io_o_4_out[5] ,
    \cb_3_3_io_o_4_out[4] ,
    \cb_3_3_io_o_4_out[3] ,
    \cb_3_3_io_o_4_out[2] ,
    \cb_3_3_io_o_4_out[1] ,
    \cb_3_3_io_o_4_out[0] }),
    .io_o_5_out({\cb_3_3_io_o_5_out[7] ,
    \cb_3_3_io_o_5_out[6] ,
    \cb_3_3_io_o_5_out[5] ,
    \cb_3_3_io_o_5_out[4] ,
    \cb_3_3_io_o_5_out[3] ,
    \cb_3_3_io_o_5_out[2] ,
    \cb_3_3_io_o_5_out[1] ,
    \cb_3_3_io_o_5_out[0] }),
    .io_o_6_out({\cb_3_3_io_o_6_out[7] ,
    \cb_3_3_io_o_6_out[6] ,
    \cb_3_3_io_o_6_out[5] ,
    \cb_3_3_io_o_6_out[4] ,
    \cb_3_3_io_o_6_out[3] ,
    \cb_3_3_io_o_6_out[2] ,
    \cb_3_3_io_o_6_out[1] ,
    \cb_3_3_io_o_6_out[0] }),
    .io_o_7_out({\cb_3_3_io_o_7_out[7] ,
    \cb_3_3_io_o_7_out[6] ,
    \cb_3_3_io_o_7_out[5] ,
    \cb_3_3_io_o_7_out[4] ,
    \cb_3_3_io_o_7_out[3] ,
    \cb_3_3_io_o_7_out[2] ,
    \cb_3_3_io_o_7_out[1] ,
    \cb_3_3_io_o_7_out[0] }),
    .io_wo({\cb_3_2_io_eo[63] ,
    \cb_3_2_io_eo[62] ,
    \cb_3_2_io_eo[61] ,
    \cb_3_2_io_eo[60] ,
    \cb_3_2_io_eo[59] ,
    \cb_3_2_io_eo[58] ,
    \cb_3_2_io_eo[57] ,
    \cb_3_2_io_eo[56] ,
    \cb_3_2_io_eo[55] ,
    \cb_3_2_io_eo[54] ,
    \cb_3_2_io_eo[53] ,
    \cb_3_2_io_eo[52] ,
    \cb_3_2_io_eo[51] ,
    \cb_3_2_io_eo[50] ,
    \cb_3_2_io_eo[49] ,
    \cb_3_2_io_eo[48] ,
    \cb_3_2_io_eo[47] ,
    \cb_3_2_io_eo[46] ,
    \cb_3_2_io_eo[45] ,
    \cb_3_2_io_eo[44] ,
    \cb_3_2_io_eo[43] ,
    \cb_3_2_io_eo[42] ,
    \cb_3_2_io_eo[41] ,
    \cb_3_2_io_eo[40] ,
    \cb_3_2_io_eo[39] ,
    \cb_3_2_io_eo[38] ,
    \cb_3_2_io_eo[37] ,
    \cb_3_2_io_eo[36] ,
    \cb_3_2_io_eo[35] ,
    \cb_3_2_io_eo[34] ,
    \cb_3_2_io_eo[33] ,
    \cb_3_2_io_eo[32] ,
    \cb_3_2_io_eo[31] ,
    \cb_3_2_io_eo[30] ,
    \cb_3_2_io_eo[29] ,
    \cb_3_2_io_eo[28] ,
    \cb_3_2_io_eo[27] ,
    \cb_3_2_io_eo[26] ,
    \cb_3_2_io_eo[25] ,
    \cb_3_2_io_eo[24] ,
    \cb_3_2_io_eo[23] ,
    \cb_3_2_io_eo[22] ,
    \cb_3_2_io_eo[21] ,
    \cb_3_2_io_eo[20] ,
    \cb_3_2_io_eo[19] ,
    \cb_3_2_io_eo[18] ,
    \cb_3_2_io_eo[17] ,
    \cb_3_2_io_eo[16] ,
    \cb_3_2_io_eo[15] ,
    \cb_3_2_io_eo[14] ,
    \cb_3_2_io_eo[13] ,
    \cb_3_2_io_eo[12] ,
    \cb_3_2_io_eo[11] ,
    \cb_3_2_io_eo[10] ,
    \cb_3_2_io_eo[9] ,
    \cb_3_2_io_eo[8] ,
    \cb_3_2_io_eo[7] ,
    \cb_3_2_io_eo[6] ,
    \cb_3_2_io_eo[5] ,
    \cb_3_2_io_eo[4] ,
    \cb_3_2_io_eo[3] ,
    \cb_3_2_io_eo[2] ,
    \cb_3_2_io_eo[1] ,
    \cb_3_2_io_eo[0] }));
 cic_block cb_3_4 (.io_cs_i(cb_3_4_io_cs_i),
    .io_i_0_ci(cb_3_3_io_o_0_co),
    .io_i_1_ci(cb_3_3_io_o_1_co),
    .io_i_2_ci(cb_3_3_io_o_2_co),
    .io_i_3_ci(cb_3_3_io_o_3_co),
    .io_i_4_ci(cb_3_3_io_o_4_co),
    .io_i_5_ci(cb_3_3_io_o_5_co),
    .io_i_6_ci(cb_3_3_io_o_6_co),
    .io_i_7_ci(cb_3_3_io_o_7_co),
    .io_o_0_co(cb_3_4_io_o_0_co),
    .io_o_1_co(cb_3_4_io_o_1_co),
    .io_o_2_co(cb_3_4_io_o_2_co),
    .io_o_3_co(cb_3_4_io_o_3_co),
    .io_o_4_co(cb_3_4_io_o_4_co),
    .io_o_5_co(cb_3_4_io_o_5_co),
    .io_o_6_co(cb_3_4_io_o_6_co),
    .io_o_7_co(cb_3_4_io_o_7_co),
    .io_vci(cb_3_3_io_vco),
    .io_vco(cb_3_4_io_vco),
    .io_vi(cb_3_4_io_vi),
    .io_we_i(cb_3_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_3_0_io_adr_i[1] ,
    \cb_3_0_io_adr_i[0] }),
    .io_dat_i({\cb_3_0_io_dat_i[15] ,
    \cb_3_0_io_dat_i[14] ,
    \cb_3_0_io_dat_i[13] ,
    \cb_3_0_io_dat_i[12] ,
    \cb_3_0_io_dat_i[11] ,
    \cb_3_0_io_dat_i[10] ,
    \cb_3_0_io_dat_i[9] ,
    \cb_3_0_io_dat_i[8] ,
    \cb_3_0_io_dat_i[7] ,
    \cb_3_0_io_dat_i[6] ,
    \cb_3_0_io_dat_i[5] ,
    \cb_3_0_io_dat_i[4] ,
    \cb_3_0_io_dat_i[3] ,
    \cb_3_0_io_dat_i[2] ,
    \cb_3_0_io_dat_i[1] ,
    \cb_3_0_io_dat_i[0] }),
    .io_dat_o({\cb_3_4_io_dat_o[15] ,
    \cb_3_4_io_dat_o[14] ,
    \cb_3_4_io_dat_o[13] ,
    \cb_3_4_io_dat_o[12] ,
    \cb_3_4_io_dat_o[11] ,
    \cb_3_4_io_dat_o[10] ,
    \cb_3_4_io_dat_o[9] ,
    \cb_3_4_io_dat_o[8] ,
    \cb_3_4_io_dat_o[7] ,
    \cb_3_4_io_dat_o[6] ,
    \cb_3_4_io_dat_o[5] ,
    \cb_3_4_io_dat_o[4] ,
    \cb_3_4_io_dat_o[3] ,
    \cb_3_4_io_dat_o[2] ,
    \cb_3_4_io_dat_o[1] ,
    \cb_3_4_io_dat_o[0] }),
    .io_eo({\cb_3_4_io_eo[63] ,
    \cb_3_4_io_eo[62] ,
    \cb_3_4_io_eo[61] ,
    \cb_3_4_io_eo[60] ,
    \cb_3_4_io_eo[59] ,
    \cb_3_4_io_eo[58] ,
    \cb_3_4_io_eo[57] ,
    \cb_3_4_io_eo[56] ,
    \cb_3_4_io_eo[55] ,
    \cb_3_4_io_eo[54] ,
    \cb_3_4_io_eo[53] ,
    \cb_3_4_io_eo[52] ,
    \cb_3_4_io_eo[51] ,
    \cb_3_4_io_eo[50] ,
    \cb_3_4_io_eo[49] ,
    \cb_3_4_io_eo[48] ,
    \cb_3_4_io_eo[47] ,
    \cb_3_4_io_eo[46] ,
    \cb_3_4_io_eo[45] ,
    \cb_3_4_io_eo[44] ,
    \cb_3_4_io_eo[43] ,
    \cb_3_4_io_eo[42] ,
    \cb_3_4_io_eo[41] ,
    \cb_3_4_io_eo[40] ,
    \cb_3_4_io_eo[39] ,
    \cb_3_4_io_eo[38] ,
    \cb_3_4_io_eo[37] ,
    \cb_3_4_io_eo[36] ,
    \cb_3_4_io_eo[35] ,
    \cb_3_4_io_eo[34] ,
    \cb_3_4_io_eo[33] ,
    \cb_3_4_io_eo[32] ,
    \cb_3_4_io_eo[31] ,
    \cb_3_4_io_eo[30] ,
    \cb_3_4_io_eo[29] ,
    \cb_3_4_io_eo[28] ,
    \cb_3_4_io_eo[27] ,
    \cb_3_4_io_eo[26] ,
    \cb_3_4_io_eo[25] ,
    \cb_3_4_io_eo[24] ,
    \cb_3_4_io_eo[23] ,
    \cb_3_4_io_eo[22] ,
    \cb_3_4_io_eo[21] ,
    \cb_3_4_io_eo[20] ,
    \cb_3_4_io_eo[19] ,
    \cb_3_4_io_eo[18] ,
    \cb_3_4_io_eo[17] ,
    \cb_3_4_io_eo[16] ,
    \cb_3_4_io_eo[15] ,
    \cb_3_4_io_eo[14] ,
    \cb_3_4_io_eo[13] ,
    \cb_3_4_io_eo[12] ,
    \cb_3_4_io_eo[11] ,
    \cb_3_4_io_eo[10] ,
    \cb_3_4_io_eo[9] ,
    \cb_3_4_io_eo[8] ,
    \cb_3_4_io_eo[7] ,
    \cb_3_4_io_eo[6] ,
    \cb_3_4_io_eo[5] ,
    \cb_3_4_io_eo[4] ,
    \cb_3_4_io_eo[3] ,
    \cb_3_4_io_eo[2] ,
    \cb_3_4_io_eo[1] ,
    \cb_3_4_io_eo[0] }),
    .io_i_0_in1({\cb_3_3_io_o_0_out[7] ,
    \cb_3_3_io_o_0_out[6] ,
    \cb_3_3_io_o_0_out[5] ,
    \cb_3_3_io_o_0_out[4] ,
    \cb_3_3_io_o_0_out[3] ,
    \cb_3_3_io_o_0_out[2] ,
    \cb_3_3_io_o_0_out[1] ,
    \cb_3_3_io_o_0_out[0] }),
    .io_i_1_in1({\cb_3_3_io_o_1_out[7] ,
    \cb_3_3_io_o_1_out[6] ,
    \cb_3_3_io_o_1_out[5] ,
    \cb_3_3_io_o_1_out[4] ,
    \cb_3_3_io_o_1_out[3] ,
    \cb_3_3_io_o_1_out[2] ,
    \cb_3_3_io_o_1_out[1] ,
    \cb_3_3_io_o_1_out[0] }),
    .io_i_2_in1({\cb_3_3_io_o_2_out[7] ,
    \cb_3_3_io_o_2_out[6] ,
    \cb_3_3_io_o_2_out[5] ,
    \cb_3_3_io_o_2_out[4] ,
    \cb_3_3_io_o_2_out[3] ,
    \cb_3_3_io_o_2_out[2] ,
    \cb_3_3_io_o_2_out[1] ,
    \cb_3_3_io_o_2_out[0] }),
    .io_i_3_in1({\cb_3_3_io_o_3_out[7] ,
    \cb_3_3_io_o_3_out[6] ,
    \cb_3_3_io_o_3_out[5] ,
    \cb_3_3_io_o_3_out[4] ,
    \cb_3_3_io_o_3_out[3] ,
    \cb_3_3_io_o_3_out[2] ,
    \cb_3_3_io_o_3_out[1] ,
    \cb_3_3_io_o_3_out[0] }),
    .io_i_4_in1({\cb_3_3_io_o_4_out[7] ,
    \cb_3_3_io_o_4_out[6] ,
    \cb_3_3_io_o_4_out[5] ,
    \cb_3_3_io_o_4_out[4] ,
    \cb_3_3_io_o_4_out[3] ,
    \cb_3_3_io_o_4_out[2] ,
    \cb_3_3_io_o_4_out[1] ,
    \cb_3_3_io_o_4_out[0] }),
    .io_i_5_in1({\cb_3_3_io_o_5_out[7] ,
    \cb_3_3_io_o_5_out[6] ,
    \cb_3_3_io_o_5_out[5] ,
    \cb_3_3_io_o_5_out[4] ,
    \cb_3_3_io_o_5_out[3] ,
    \cb_3_3_io_o_5_out[2] ,
    \cb_3_3_io_o_5_out[1] ,
    \cb_3_3_io_o_5_out[0] }),
    .io_i_6_in1({\cb_3_3_io_o_6_out[7] ,
    \cb_3_3_io_o_6_out[6] ,
    \cb_3_3_io_o_6_out[5] ,
    \cb_3_3_io_o_6_out[4] ,
    \cb_3_3_io_o_6_out[3] ,
    \cb_3_3_io_o_6_out[2] ,
    \cb_3_3_io_o_6_out[1] ,
    \cb_3_3_io_o_6_out[0] }),
    .io_i_7_in1({\cb_3_3_io_o_7_out[7] ,
    \cb_3_3_io_o_7_out[6] ,
    \cb_3_3_io_o_7_out[5] ,
    \cb_3_3_io_o_7_out[4] ,
    \cb_3_3_io_o_7_out[3] ,
    \cb_3_3_io_o_7_out[2] ,
    \cb_3_3_io_o_7_out[1] ,
    \cb_3_3_io_o_7_out[0] }),
    .io_o_0_out({\cb_3_4_io_o_0_out[7] ,
    \cb_3_4_io_o_0_out[6] ,
    \cb_3_4_io_o_0_out[5] ,
    \cb_3_4_io_o_0_out[4] ,
    \cb_3_4_io_o_0_out[3] ,
    \cb_3_4_io_o_0_out[2] ,
    \cb_3_4_io_o_0_out[1] ,
    \cb_3_4_io_o_0_out[0] }),
    .io_o_1_out({\cb_3_4_io_o_1_out[7] ,
    \cb_3_4_io_o_1_out[6] ,
    \cb_3_4_io_o_1_out[5] ,
    \cb_3_4_io_o_1_out[4] ,
    \cb_3_4_io_o_1_out[3] ,
    \cb_3_4_io_o_1_out[2] ,
    \cb_3_4_io_o_1_out[1] ,
    \cb_3_4_io_o_1_out[0] }),
    .io_o_2_out({\cb_3_4_io_o_2_out[7] ,
    \cb_3_4_io_o_2_out[6] ,
    \cb_3_4_io_o_2_out[5] ,
    \cb_3_4_io_o_2_out[4] ,
    \cb_3_4_io_o_2_out[3] ,
    \cb_3_4_io_o_2_out[2] ,
    \cb_3_4_io_o_2_out[1] ,
    \cb_3_4_io_o_2_out[0] }),
    .io_o_3_out({\cb_3_4_io_o_3_out[7] ,
    \cb_3_4_io_o_3_out[6] ,
    \cb_3_4_io_o_3_out[5] ,
    \cb_3_4_io_o_3_out[4] ,
    \cb_3_4_io_o_3_out[3] ,
    \cb_3_4_io_o_3_out[2] ,
    \cb_3_4_io_o_3_out[1] ,
    \cb_3_4_io_o_3_out[0] }),
    .io_o_4_out({\cb_3_4_io_o_4_out[7] ,
    \cb_3_4_io_o_4_out[6] ,
    \cb_3_4_io_o_4_out[5] ,
    \cb_3_4_io_o_4_out[4] ,
    \cb_3_4_io_o_4_out[3] ,
    \cb_3_4_io_o_4_out[2] ,
    \cb_3_4_io_o_4_out[1] ,
    \cb_3_4_io_o_4_out[0] }),
    .io_o_5_out({\cb_3_4_io_o_5_out[7] ,
    \cb_3_4_io_o_5_out[6] ,
    \cb_3_4_io_o_5_out[5] ,
    \cb_3_4_io_o_5_out[4] ,
    \cb_3_4_io_o_5_out[3] ,
    \cb_3_4_io_o_5_out[2] ,
    \cb_3_4_io_o_5_out[1] ,
    \cb_3_4_io_o_5_out[0] }),
    .io_o_6_out({\cb_3_4_io_o_6_out[7] ,
    \cb_3_4_io_o_6_out[6] ,
    \cb_3_4_io_o_6_out[5] ,
    \cb_3_4_io_o_6_out[4] ,
    \cb_3_4_io_o_6_out[3] ,
    \cb_3_4_io_o_6_out[2] ,
    \cb_3_4_io_o_6_out[1] ,
    \cb_3_4_io_o_6_out[0] }),
    .io_o_7_out({\cb_3_4_io_o_7_out[7] ,
    \cb_3_4_io_o_7_out[6] ,
    \cb_3_4_io_o_7_out[5] ,
    \cb_3_4_io_o_7_out[4] ,
    \cb_3_4_io_o_7_out[3] ,
    \cb_3_4_io_o_7_out[2] ,
    \cb_3_4_io_o_7_out[1] ,
    \cb_3_4_io_o_7_out[0] }),
    .io_wo({\cb_3_3_io_eo[63] ,
    \cb_3_3_io_eo[62] ,
    \cb_3_3_io_eo[61] ,
    \cb_3_3_io_eo[60] ,
    \cb_3_3_io_eo[59] ,
    \cb_3_3_io_eo[58] ,
    \cb_3_3_io_eo[57] ,
    \cb_3_3_io_eo[56] ,
    \cb_3_3_io_eo[55] ,
    \cb_3_3_io_eo[54] ,
    \cb_3_3_io_eo[53] ,
    \cb_3_3_io_eo[52] ,
    \cb_3_3_io_eo[51] ,
    \cb_3_3_io_eo[50] ,
    \cb_3_3_io_eo[49] ,
    \cb_3_3_io_eo[48] ,
    \cb_3_3_io_eo[47] ,
    \cb_3_3_io_eo[46] ,
    \cb_3_3_io_eo[45] ,
    \cb_3_3_io_eo[44] ,
    \cb_3_3_io_eo[43] ,
    \cb_3_3_io_eo[42] ,
    \cb_3_3_io_eo[41] ,
    \cb_3_3_io_eo[40] ,
    \cb_3_3_io_eo[39] ,
    \cb_3_3_io_eo[38] ,
    \cb_3_3_io_eo[37] ,
    \cb_3_3_io_eo[36] ,
    \cb_3_3_io_eo[35] ,
    \cb_3_3_io_eo[34] ,
    \cb_3_3_io_eo[33] ,
    \cb_3_3_io_eo[32] ,
    \cb_3_3_io_eo[31] ,
    \cb_3_3_io_eo[30] ,
    \cb_3_3_io_eo[29] ,
    \cb_3_3_io_eo[28] ,
    \cb_3_3_io_eo[27] ,
    \cb_3_3_io_eo[26] ,
    \cb_3_3_io_eo[25] ,
    \cb_3_3_io_eo[24] ,
    \cb_3_3_io_eo[23] ,
    \cb_3_3_io_eo[22] ,
    \cb_3_3_io_eo[21] ,
    \cb_3_3_io_eo[20] ,
    \cb_3_3_io_eo[19] ,
    \cb_3_3_io_eo[18] ,
    \cb_3_3_io_eo[17] ,
    \cb_3_3_io_eo[16] ,
    \cb_3_3_io_eo[15] ,
    \cb_3_3_io_eo[14] ,
    \cb_3_3_io_eo[13] ,
    \cb_3_3_io_eo[12] ,
    \cb_3_3_io_eo[11] ,
    \cb_3_3_io_eo[10] ,
    \cb_3_3_io_eo[9] ,
    \cb_3_3_io_eo[8] ,
    \cb_3_3_io_eo[7] ,
    \cb_3_3_io_eo[6] ,
    \cb_3_3_io_eo[5] ,
    \cb_3_3_io_eo[4] ,
    \cb_3_3_io_eo[3] ,
    \cb_3_3_io_eo[2] ,
    \cb_3_3_io_eo[1] ,
    \cb_3_3_io_eo[0] }));
 cic_block cb_3_5 (.io_cs_i(cb_3_5_io_cs_i),
    .io_i_0_ci(cb_3_4_io_o_0_co),
    .io_i_1_ci(cb_3_4_io_o_1_co),
    .io_i_2_ci(cb_3_4_io_o_2_co),
    .io_i_3_ci(cb_3_4_io_o_3_co),
    .io_i_4_ci(cb_3_4_io_o_4_co),
    .io_i_5_ci(cb_3_4_io_o_5_co),
    .io_i_6_ci(cb_3_4_io_o_6_co),
    .io_i_7_ci(cb_3_4_io_o_7_co),
    .io_o_0_co(cb_3_5_io_o_0_co),
    .io_o_1_co(cb_3_5_io_o_1_co),
    .io_o_2_co(cb_3_5_io_o_2_co),
    .io_o_3_co(cb_3_5_io_o_3_co),
    .io_o_4_co(cb_3_5_io_o_4_co),
    .io_o_5_co(cb_3_5_io_o_5_co),
    .io_o_6_co(cb_3_5_io_o_6_co),
    .io_o_7_co(cb_3_5_io_o_7_co),
    .io_vci(cb_3_4_io_vco),
    .io_vco(cb_3_5_io_vco),
    .io_vi(cb_3_5_io_vi),
    .io_we_i(cb_3_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_3_0_io_adr_i[1] ,
    \cb_3_0_io_adr_i[0] }),
    .io_dat_i({\cb_3_0_io_dat_i[15] ,
    \cb_3_0_io_dat_i[14] ,
    \cb_3_0_io_dat_i[13] ,
    \cb_3_0_io_dat_i[12] ,
    \cb_3_0_io_dat_i[11] ,
    \cb_3_0_io_dat_i[10] ,
    \cb_3_0_io_dat_i[9] ,
    \cb_3_0_io_dat_i[8] ,
    \cb_3_0_io_dat_i[7] ,
    \cb_3_0_io_dat_i[6] ,
    \cb_3_0_io_dat_i[5] ,
    \cb_3_0_io_dat_i[4] ,
    \cb_3_0_io_dat_i[3] ,
    \cb_3_0_io_dat_i[2] ,
    \cb_3_0_io_dat_i[1] ,
    \cb_3_0_io_dat_i[0] }),
    .io_dat_o({\cb_3_5_io_dat_o[15] ,
    \cb_3_5_io_dat_o[14] ,
    \cb_3_5_io_dat_o[13] ,
    \cb_3_5_io_dat_o[12] ,
    \cb_3_5_io_dat_o[11] ,
    \cb_3_5_io_dat_o[10] ,
    \cb_3_5_io_dat_o[9] ,
    \cb_3_5_io_dat_o[8] ,
    \cb_3_5_io_dat_o[7] ,
    \cb_3_5_io_dat_o[6] ,
    \cb_3_5_io_dat_o[5] ,
    \cb_3_5_io_dat_o[4] ,
    \cb_3_5_io_dat_o[3] ,
    \cb_3_5_io_dat_o[2] ,
    \cb_3_5_io_dat_o[1] ,
    \cb_3_5_io_dat_o[0] }),
    .io_eo({\cb_3_5_io_eo[63] ,
    \cb_3_5_io_eo[62] ,
    \cb_3_5_io_eo[61] ,
    \cb_3_5_io_eo[60] ,
    \cb_3_5_io_eo[59] ,
    \cb_3_5_io_eo[58] ,
    \cb_3_5_io_eo[57] ,
    \cb_3_5_io_eo[56] ,
    \cb_3_5_io_eo[55] ,
    \cb_3_5_io_eo[54] ,
    \cb_3_5_io_eo[53] ,
    \cb_3_5_io_eo[52] ,
    \cb_3_5_io_eo[51] ,
    \cb_3_5_io_eo[50] ,
    \cb_3_5_io_eo[49] ,
    \cb_3_5_io_eo[48] ,
    \cb_3_5_io_eo[47] ,
    \cb_3_5_io_eo[46] ,
    \cb_3_5_io_eo[45] ,
    \cb_3_5_io_eo[44] ,
    \cb_3_5_io_eo[43] ,
    \cb_3_5_io_eo[42] ,
    \cb_3_5_io_eo[41] ,
    \cb_3_5_io_eo[40] ,
    \cb_3_5_io_eo[39] ,
    \cb_3_5_io_eo[38] ,
    \cb_3_5_io_eo[37] ,
    \cb_3_5_io_eo[36] ,
    \cb_3_5_io_eo[35] ,
    \cb_3_5_io_eo[34] ,
    \cb_3_5_io_eo[33] ,
    \cb_3_5_io_eo[32] ,
    \cb_3_5_io_eo[31] ,
    \cb_3_5_io_eo[30] ,
    \cb_3_5_io_eo[29] ,
    \cb_3_5_io_eo[28] ,
    \cb_3_5_io_eo[27] ,
    \cb_3_5_io_eo[26] ,
    \cb_3_5_io_eo[25] ,
    \cb_3_5_io_eo[24] ,
    \cb_3_5_io_eo[23] ,
    \cb_3_5_io_eo[22] ,
    \cb_3_5_io_eo[21] ,
    \cb_3_5_io_eo[20] ,
    \cb_3_5_io_eo[19] ,
    \cb_3_5_io_eo[18] ,
    \cb_3_5_io_eo[17] ,
    \cb_3_5_io_eo[16] ,
    \cb_3_5_io_eo[15] ,
    \cb_3_5_io_eo[14] ,
    \cb_3_5_io_eo[13] ,
    \cb_3_5_io_eo[12] ,
    \cb_3_5_io_eo[11] ,
    \cb_3_5_io_eo[10] ,
    \cb_3_5_io_eo[9] ,
    \cb_3_5_io_eo[8] ,
    \cb_3_5_io_eo[7] ,
    \cb_3_5_io_eo[6] ,
    \cb_3_5_io_eo[5] ,
    \cb_3_5_io_eo[4] ,
    \cb_3_5_io_eo[3] ,
    \cb_3_5_io_eo[2] ,
    \cb_3_5_io_eo[1] ,
    \cb_3_5_io_eo[0] }),
    .io_i_0_in1({\cb_3_4_io_o_0_out[7] ,
    \cb_3_4_io_o_0_out[6] ,
    \cb_3_4_io_o_0_out[5] ,
    \cb_3_4_io_o_0_out[4] ,
    \cb_3_4_io_o_0_out[3] ,
    \cb_3_4_io_o_0_out[2] ,
    \cb_3_4_io_o_0_out[1] ,
    \cb_3_4_io_o_0_out[0] }),
    .io_i_1_in1({\cb_3_4_io_o_1_out[7] ,
    \cb_3_4_io_o_1_out[6] ,
    \cb_3_4_io_o_1_out[5] ,
    \cb_3_4_io_o_1_out[4] ,
    \cb_3_4_io_o_1_out[3] ,
    \cb_3_4_io_o_1_out[2] ,
    \cb_3_4_io_o_1_out[1] ,
    \cb_3_4_io_o_1_out[0] }),
    .io_i_2_in1({\cb_3_4_io_o_2_out[7] ,
    \cb_3_4_io_o_2_out[6] ,
    \cb_3_4_io_o_2_out[5] ,
    \cb_3_4_io_o_2_out[4] ,
    \cb_3_4_io_o_2_out[3] ,
    \cb_3_4_io_o_2_out[2] ,
    \cb_3_4_io_o_2_out[1] ,
    \cb_3_4_io_o_2_out[0] }),
    .io_i_3_in1({\cb_3_4_io_o_3_out[7] ,
    \cb_3_4_io_o_3_out[6] ,
    \cb_3_4_io_o_3_out[5] ,
    \cb_3_4_io_o_3_out[4] ,
    \cb_3_4_io_o_3_out[3] ,
    \cb_3_4_io_o_3_out[2] ,
    \cb_3_4_io_o_3_out[1] ,
    \cb_3_4_io_o_3_out[0] }),
    .io_i_4_in1({\cb_3_4_io_o_4_out[7] ,
    \cb_3_4_io_o_4_out[6] ,
    \cb_3_4_io_o_4_out[5] ,
    \cb_3_4_io_o_4_out[4] ,
    \cb_3_4_io_o_4_out[3] ,
    \cb_3_4_io_o_4_out[2] ,
    \cb_3_4_io_o_4_out[1] ,
    \cb_3_4_io_o_4_out[0] }),
    .io_i_5_in1({\cb_3_4_io_o_5_out[7] ,
    \cb_3_4_io_o_5_out[6] ,
    \cb_3_4_io_o_5_out[5] ,
    \cb_3_4_io_o_5_out[4] ,
    \cb_3_4_io_o_5_out[3] ,
    \cb_3_4_io_o_5_out[2] ,
    \cb_3_4_io_o_5_out[1] ,
    \cb_3_4_io_o_5_out[0] }),
    .io_i_6_in1({\cb_3_4_io_o_6_out[7] ,
    \cb_3_4_io_o_6_out[6] ,
    \cb_3_4_io_o_6_out[5] ,
    \cb_3_4_io_o_6_out[4] ,
    \cb_3_4_io_o_6_out[3] ,
    \cb_3_4_io_o_6_out[2] ,
    \cb_3_4_io_o_6_out[1] ,
    \cb_3_4_io_o_6_out[0] }),
    .io_i_7_in1({\cb_3_4_io_o_7_out[7] ,
    \cb_3_4_io_o_7_out[6] ,
    \cb_3_4_io_o_7_out[5] ,
    \cb_3_4_io_o_7_out[4] ,
    \cb_3_4_io_o_7_out[3] ,
    \cb_3_4_io_o_7_out[2] ,
    \cb_3_4_io_o_7_out[1] ,
    \cb_3_4_io_o_7_out[0] }),
    .io_o_0_out({\cb_3_5_io_o_0_out[7] ,
    \cb_3_5_io_o_0_out[6] ,
    \cb_3_5_io_o_0_out[5] ,
    \cb_3_5_io_o_0_out[4] ,
    \cb_3_5_io_o_0_out[3] ,
    \cb_3_5_io_o_0_out[2] ,
    \cb_3_5_io_o_0_out[1] ,
    \cb_3_5_io_o_0_out[0] }),
    .io_o_1_out({\cb_3_5_io_o_1_out[7] ,
    \cb_3_5_io_o_1_out[6] ,
    \cb_3_5_io_o_1_out[5] ,
    \cb_3_5_io_o_1_out[4] ,
    \cb_3_5_io_o_1_out[3] ,
    \cb_3_5_io_o_1_out[2] ,
    \cb_3_5_io_o_1_out[1] ,
    \cb_3_5_io_o_1_out[0] }),
    .io_o_2_out({\cb_3_5_io_o_2_out[7] ,
    \cb_3_5_io_o_2_out[6] ,
    \cb_3_5_io_o_2_out[5] ,
    \cb_3_5_io_o_2_out[4] ,
    \cb_3_5_io_o_2_out[3] ,
    \cb_3_5_io_o_2_out[2] ,
    \cb_3_5_io_o_2_out[1] ,
    \cb_3_5_io_o_2_out[0] }),
    .io_o_3_out({\cb_3_5_io_o_3_out[7] ,
    \cb_3_5_io_o_3_out[6] ,
    \cb_3_5_io_o_3_out[5] ,
    \cb_3_5_io_o_3_out[4] ,
    \cb_3_5_io_o_3_out[3] ,
    \cb_3_5_io_o_3_out[2] ,
    \cb_3_5_io_o_3_out[1] ,
    \cb_3_5_io_o_3_out[0] }),
    .io_o_4_out({\cb_3_5_io_o_4_out[7] ,
    \cb_3_5_io_o_4_out[6] ,
    \cb_3_5_io_o_4_out[5] ,
    \cb_3_5_io_o_4_out[4] ,
    \cb_3_5_io_o_4_out[3] ,
    \cb_3_5_io_o_4_out[2] ,
    \cb_3_5_io_o_4_out[1] ,
    \cb_3_5_io_o_4_out[0] }),
    .io_o_5_out({\cb_3_5_io_o_5_out[7] ,
    \cb_3_5_io_o_5_out[6] ,
    \cb_3_5_io_o_5_out[5] ,
    \cb_3_5_io_o_5_out[4] ,
    \cb_3_5_io_o_5_out[3] ,
    \cb_3_5_io_o_5_out[2] ,
    \cb_3_5_io_o_5_out[1] ,
    \cb_3_5_io_o_5_out[0] }),
    .io_o_6_out({\cb_3_5_io_o_6_out[7] ,
    \cb_3_5_io_o_6_out[6] ,
    \cb_3_5_io_o_6_out[5] ,
    \cb_3_5_io_o_6_out[4] ,
    \cb_3_5_io_o_6_out[3] ,
    \cb_3_5_io_o_6_out[2] ,
    \cb_3_5_io_o_6_out[1] ,
    \cb_3_5_io_o_6_out[0] }),
    .io_o_7_out({\cb_3_5_io_o_7_out[7] ,
    \cb_3_5_io_o_7_out[6] ,
    \cb_3_5_io_o_7_out[5] ,
    \cb_3_5_io_o_7_out[4] ,
    \cb_3_5_io_o_7_out[3] ,
    \cb_3_5_io_o_7_out[2] ,
    \cb_3_5_io_o_7_out[1] ,
    \cb_3_5_io_o_7_out[0] }),
    .io_wo({\cb_3_4_io_eo[63] ,
    \cb_3_4_io_eo[62] ,
    \cb_3_4_io_eo[61] ,
    \cb_3_4_io_eo[60] ,
    \cb_3_4_io_eo[59] ,
    \cb_3_4_io_eo[58] ,
    \cb_3_4_io_eo[57] ,
    \cb_3_4_io_eo[56] ,
    \cb_3_4_io_eo[55] ,
    \cb_3_4_io_eo[54] ,
    \cb_3_4_io_eo[53] ,
    \cb_3_4_io_eo[52] ,
    \cb_3_4_io_eo[51] ,
    \cb_3_4_io_eo[50] ,
    \cb_3_4_io_eo[49] ,
    \cb_3_4_io_eo[48] ,
    \cb_3_4_io_eo[47] ,
    \cb_3_4_io_eo[46] ,
    \cb_3_4_io_eo[45] ,
    \cb_3_4_io_eo[44] ,
    \cb_3_4_io_eo[43] ,
    \cb_3_4_io_eo[42] ,
    \cb_3_4_io_eo[41] ,
    \cb_3_4_io_eo[40] ,
    \cb_3_4_io_eo[39] ,
    \cb_3_4_io_eo[38] ,
    \cb_3_4_io_eo[37] ,
    \cb_3_4_io_eo[36] ,
    \cb_3_4_io_eo[35] ,
    \cb_3_4_io_eo[34] ,
    \cb_3_4_io_eo[33] ,
    \cb_3_4_io_eo[32] ,
    \cb_3_4_io_eo[31] ,
    \cb_3_4_io_eo[30] ,
    \cb_3_4_io_eo[29] ,
    \cb_3_4_io_eo[28] ,
    \cb_3_4_io_eo[27] ,
    \cb_3_4_io_eo[26] ,
    \cb_3_4_io_eo[25] ,
    \cb_3_4_io_eo[24] ,
    \cb_3_4_io_eo[23] ,
    \cb_3_4_io_eo[22] ,
    \cb_3_4_io_eo[21] ,
    \cb_3_4_io_eo[20] ,
    \cb_3_4_io_eo[19] ,
    \cb_3_4_io_eo[18] ,
    \cb_3_4_io_eo[17] ,
    \cb_3_4_io_eo[16] ,
    \cb_3_4_io_eo[15] ,
    \cb_3_4_io_eo[14] ,
    \cb_3_4_io_eo[13] ,
    \cb_3_4_io_eo[12] ,
    \cb_3_4_io_eo[11] ,
    \cb_3_4_io_eo[10] ,
    \cb_3_4_io_eo[9] ,
    \cb_3_4_io_eo[8] ,
    \cb_3_4_io_eo[7] ,
    \cb_3_4_io_eo[6] ,
    \cb_3_4_io_eo[5] ,
    \cb_3_4_io_eo[4] ,
    \cb_3_4_io_eo[3] ,
    \cb_3_4_io_eo[2] ,
    \cb_3_4_io_eo[1] ,
    \cb_3_4_io_eo[0] }));
 cic_block cb_3_6 (.io_cs_i(cb_3_6_io_cs_i),
    .io_i_0_ci(cb_3_5_io_o_0_co),
    .io_i_1_ci(cb_3_5_io_o_1_co),
    .io_i_2_ci(cb_3_5_io_o_2_co),
    .io_i_3_ci(cb_3_5_io_o_3_co),
    .io_i_4_ci(cb_3_5_io_o_4_co),
    .io_i_5_ci(cb_3_5_io_o_5_co),
    .io_i_6_ci(cb_3_5_io_o_6_co),
    .io_i_7_ci(cb_3_5_io_o_7_co),
    .io_o_0_co(cb_3_6_io_o_0_co),
    .io_o_1_co(cb_3_6_io_o_1_co),
    .io_o_2_co(cb_3_6_io_o_2_co),
    .io_o_3_co(cb_3_6_io_o_3_co),
    .io_o_4_co(cb_3_6_io_o_4_co),
    .io_o_5_co(cb_3_6_io_o_5_co),
    .io_o_6_co(cb_3_6_io_o_6_co),
    .io_o_7_co(cb_3_6_io_o_7_co),
    .io_vci(cb_3_5_io_vco),
    .io_vco(cb_3_6_io_vco),
    .io_vi(cb_3_6_io_vi),
    .io_we_i(cb_3_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_3_0_io_adr_i[1] ,
    \cb_3_0_io_adr_i[0] }),
    .io_dat_i({\cb_3_0_io_dat_i[15] ,
    \cb_3_0_io_dat_i[14] ,
    \cb_3_0_io_dat_i[13] ,
    \cb_3_0_io_dat_i[12] ,
    \cb_3_0_io_dat_i[11] ,
    \cb_3_0_io_dat_i[10] ,
    \cb_3_0_io_dat_i[9] ,
    \cb_3_0_io_dat_i[8] ,
    \cb_3_0_io_dat_i[7] ,
    \cb_3_0_io_dat_i[6] ,
    \cb_3_0_io_dat_i[5] ,
    \cb_3_0_io_dat_i[4] ,
    \cb_3_0_io_dat_i[3] ,
    \cb_3_0_io_dat_i[2] ,
    \cb_3_0_io_dat_i[1] ,
    \cb_3_0_io_dat_i[0] }),
    .io_dat_o({\cb_3_6_io_dat_o[15] ,
    \cb_3_6_io_dat_o[14] ,
    \cb_3_6_io_dat_o[13] ,
    \cb_3_6_io_dat_o[12] ,
    \cb_3_6_io_dat_o[11] ,
    \cb_3_6_io_dat_o[10] ,
    \cb_3_6_io_dat_o[9] ,
    \cb_3_6_io_dat_o[8] ,
    \cb_3_6_io_dat_o[7] ,
    \cb_3_6_io_dat_o[6] ,
    \cb_3_6_io_dat_o[5] ,
    \cb_3_6_io_dat_o[4] ,
    \cb_3_6_io_dat_o[3] ,
    \cb_3_6_io_dat_o[2] ,
    \cb_3_6_io_dat_o[1] ,
    \cb_3_6_io_dat_o[0] }),
    .io_eo({\cb_3_6_io_eo[63] ,
    \cb_3_6_io_eo[62] ,
    \cb_3_6_io_eo[61] ,
    \cb_3_6_io_eo[60] ,
    \cb_3_6_io_eo[59] ,
    \cb_3_6_io_eo[58] ,
    \cb_3_6_io_eo[57] ,
    \cb_3_6_io_eo[56] ,
    \cb_3_6_io_eo[55] ,
    \cb_3_6_io_eo[54] ,
    \cb_3_6_io_eo[53] ,
    \cb_3_6_io_eo[52] ,
    \cb_3_6_io_eo[51] ,
    \cb_3_6_io_eo[50] ,
    \cb_3_6_io_eo[49] ,
    \cb_3_6_io_eo[48] ,
    \cb_3_6_io_eo[47] ,
    \cb_3_6_io_eo[46] ,
    \cb_3_6_io_eo[45] ,
    \cb_3_6_io_eo[44] ,
    \cb_3_6_io_eo[43] ,
    \cb_3_6_io_eo[42] ,
    \cb_3_6_io_eo[41] ,
    \cb_3_6_io_eo[40] ,
    \cb_3_6_io_eo[39] ,
    \cb_3_6_io_eo[38] ,
    \cb_3_6_io_eo[37] ,
    \cb_3_6_io_eo[36] ,
    \cb_3_6_io_eo[35] ,
    \cb_3_6_io_eo[34] ,
    \cb_3_6_io_eo[33] ,
    \cb_3_6_io_eo[32] ,
    \cb_3_6_io_eo[31] ,
    \cb_3_6_io_eo[30] ,
    \cb_3_6_io_eo[29] ,
    \cb_3_6_io_eo[28] ,
    \cb_3_6_io_eo[27] ,
    \cb_3_6_io_eo[26] ,
    \cb_3_6_io_eo[25] ,
    \cb_3_6_io_eo[24] ,
    \cb_3_6_io_eo[23] ,
    \cb_3_6_io_eo[22] ,
    \cb_3_6_io_eo[21] ,
    \cb_3_6_io_eo[20] ,
    \cb_3_6_io_eo[19] ,
    \cb_3_6_io_eo[18] ,
    \cb_3_6_io_eo[17] ,
    \cb_3_6_io_eo[16] ,
    \cb_3_6_io_eo[15] ,
    \cb_3_6_io_eo[14] ,
    \cb_3_6_io_eo[13] ,
    \cb_3_6_io_eo[12] ,
    \cb_3_6_io_eo[11] ,
    \cb_3_6_io_eo[10] ,
    \cb_3_6_io_eo[9] ,
    \cb_3_6_io_eo[8] ,
    \cb_3_6_io_eo[7] ,
    \cb_3_6_io_eo[6] ,
    \cb_3_6_io_eo[5] ,
    \cb_3_6_io_eo[4] ,
    \cb_3_6_io_eo[3] ,
    \cb_3_6_io_eo[2] ,
    \cb_3_6_io_eo[1] ,
    \cb_3_6_io_eo[0] }),
    .io_i_0_in1({\cb_3_5_io_o_0_out[7] ,
    \cb_3_5_io_o_0_out[6] ,
    \cb_3_5_io_o_0_out[5] ,
    \cb_3_5_io_o_0_out[4] ,
    \cb_3_5_io_o_0_out[3] ,
    \cb_3_5_io_o_0_out[2] ,
    \cb_3_5_io_o_0_out[1] ,
    \cb_3_5_io_o_0_out[0] }),
    .io_i_1_in1({\cb_3_5_io_o_1_out[7] ,
    \cb_3_5_io_o_1_out[6] ,
    \cb_3_5_io_o_1_out[5] ,
    \cb_3_5_io_o_1_out[4] ,
    \cb_3_5_io_o_1_out[3] ,
    \cb_3_5_io_o_1_out[2] ,
    \cb_3_5_io_o_1_out[1] ,
    \cb_3_5_io_o_1_out[0] }),
    .io_i_2_in1({\cb_3_5_io_o_2_out[7] ,
    \cb_3_5_io_o_2_out[6] ,
    \cb_3_5_io_o_2_out[5] ,
    \cb_3_5_io_o_2_out[4] ,
    \cb_3_5_io_o_2_out[3] ,
    \cb_3_5_io_o_2_out[2] ,
    \cb_3_5_io_o_2_out[1] ,
    \cb_3_5_io_o_2_out[0] }),
    .io_i_3_in1({\cb_3_5_io_o_3_out[7] ,
    \cb_3_5_io_o_3_out[6] ,
    \cb_3_5_io_o_3_out[5] ,
    \cb_3_5_io_o_3_out[4] ,
    \cb_3_5_io_o_3_out[3] ,
    \cb_3_5_io_o_3_out[2] ,
    \cb_3_5_io_o_3_out[1] ,
    \cb_3_5_io_o_3_out[0] }),
    .io_i_4_in1({\cb_3_5_io_o_4_out[7] ,
    \cb_3_5_io_o_4_out[6] ,
    \cb_3_5_io_o_4_out[5] ,
    \cb_3_5_io_o_4_out[4] ,
    \cb_3_5_io_o_4_out[3] ,
    \cb_3_5_io_o_4_out[2] ,
    \cb_3_5_io_o_4_out[1] ,
    \cb_3_5_io_o_4_out[0] }),
    .io_i_5_in1({\cb_3_5_io_o_5_out[7] ,
    \cb_3_5_io_o_5_out[6] ,
    \cb_3_5_io_o_5_out[5] ,
    \cb_3_5_io_o_5_out[4] ,
    \cb_3_5_io_o_5_out[3] ,
    \cb_3_5_io_o_5_out[2] ,
    \cb_3_5_io_o_5_out[1] ,
    \cb_3_5_io_o_5_out[0] }),
    .io_i_6_in1({\cb_3_5_io_o_6_out[7] ,
    \cb_3_5_io_o_6_out[6] ,
    \cb_3_5_io_o_6_out[5] ,
    \cb_3_5_io_o_6_out[4] ,
    \cb_3_5_io_o_6_out[3] ,
    \cb_3_5_io_o_6_out[2] ,
    \cb_3_5_io_o_6_out[1] ,
    \cb_3_5_io_o_6_out[0] }),
    .io_i_7_in1({\cb_3_5_io_o_7_out[7] ,
    \cb_3_5_io_o_7_out[6] ,
    \cb_3_5_io_o_7_out[5] ,
    \cb_3_5_io_o_7_out[4] ,
    \cb_3_5_io_o_7_out[3] ,
    \cb_3_5_io_o_7_out[2] ,
    \cb_3_5_io_o_7_out[1] ,
    \cb_3_5_io_o_7_out[0] }),
    .io_o_0_out({\cb_3_6_io_o_0_out[7] ,
    \cb_3_6_io_o_0_out[6] ,
    \cb_3_6_io_o_0_out[5] ,
    \cb_3_6_io_o_0_out[4] ,
    \cb_3_6_io_o_0_out[3] ,
    \cb_3_6_io_o_0_out[2] ,
    \cb_3_6_io_o_0_out[1] ,
    \cb_3_6_io_o_0_out[0] }),
    .io_o_1_out({\cb_3_6_io_o_1_out[7] ,
    \cb_3_6_io_o_1_out[6] ,
    \cb_3_6_io_o_1_out[5] ,
    \cb_3_6_io_o_1_out[4] ,
    \cb_3_6_io_o_1_out[3] ,
    \cb_3_6_io_o_1_out[2] ,
    \cb_3_6_io_o_1_out[1] ,
    \cb_3_6_io_o_1_out[0] }),
    .io_o_2_out({\cb_3_6_io_o_2_out[7] ,
    \cb_3_6_io_o_2_out[6] ,
    \cb_3_6_io_o_2_out[5] ,
    \cb_3_6_io_o_2_out[4] ,
    \cb_3_6_io_o_2_out[3] ,
    \cb_3_6_io_o_2_out[2] ,
    \cb_3_6_io_o_2_out[1] ,
    \cb_3_6_io_o_2_out[0] }),
    .io_o_3_out({\cb_3_6_io_o_3_out[7] ,
    \cb_3_6_io_o_3_out[6] ,
    \cb_3_6_io_o_3_out[5] ,
    \cb_3_6_io_o_3_out[4] ,
    \cb_3_6_io_o_3_out[3] ,
    \cb_3_6_io_o_3_out[2] ,
    \cb_3_6_io_o_3_out[1] ,
    \cb_3_6_io_o_3_out[0] }),
    .io_o_4_out({\cb_3_6_io_o_4_out[7] ,
    \cb_3_6_io_o_4_out[6] ,
    \cb_3_6_io_o_4_out[5] ,
    \cb_3_6_io_o_4_out[4] ,
    \cb_3_6_io_o_4_out[3] ,
    \cb_3_6_io_o_4_out[2] ,
    \cb_3_6_io_o_4_out[1] ,
    \cb_3_6_io_o_4_out[0] }),
    .io_o_5_out({\cb_3_6_io_o_5_out[7] ,
    \cb_3_6_io_o_5_out[6] ,
    \cb_3_6_io_o_5_out[5] ,
    \cb_3_6_io_o_5_out[4] ,
    \cb_3_6_io_o_5_out[3] ,
    \cb_3_6_io_o_5_out[2] ,
    \cb_3_6_io_o_5_out[1] ,
    \cb_3_6_io_o_5_out[0] }),
    .io_o_6_out({\cb_3_6_io_o_6_out[7] ,
    \cb_3_6_io_o_6_out[6] ,
    \cb_3_6_io_o_6_out[5] ,
    \cb_3_6_io_o_6_out[4] ,
    \cb_3_6_io_o_6_out[3] ,
    \cb_3_6_io_o_6_out[2] ,
    \cb_3_6_io_o_6_out[1] ,
    \cb_3_6_io_o_6_out[0] }),
    .io_o_7_out({\cb_3_6_io_o_7_out[7] ,
    \cb_3_6_io_o_7_out[6] ,
    \cb_3_6_io_o_7_out[5] ,
    \cb_3_6_io_o_7_out[4] ,
    \cb_3_6_io_o_7_out[3] ,
    \cb_3_6_io_o_7_out[2] ,
    \cb_3_6_io_o_7_out[1] ,
    \cb_3_6_io_o_7_out[0] }),
    .io_wo({\cb_3_5_io_eo[63] ,
    \cb_3_5_io_eo[62] ,
    \cb_3_5_io_eo[61] ,
    \cb_3_5_io_eo[60] ,
    \cb_3_5_io_eo[59] ,
    \cb_3_5_io_eo[58] ,
    \cb_3_5_io_eo[57] ,
    \cb_3_5_io_eo[56] ,
    \cb_3_5_io_eo[55] ,
    \cb_3_5_io_eo[54] ,
    \cb_3_5_io_eo[53] ,
    \cb_3_5_io_eo[52] ,
    \cb_3_5_io_eo[51] ,
    \cb_3_5_io_eo[50] ,
    \cb_3_5_io_eo[49] ,
    \cb_3_5_io_eo[48] ,
    \cb_3_5_io_eo[47] ,
    \cb_3_5_io_eo[46] ,
    \cb_3_5_io_eo[45] ,
    \cb_3_5_io_eo[44] ,
    \cb_3_5_io_eo[43] ,
    \cb_3_5_io_eo[42] ,
    \cb_3_5_io_eo[41] ,
    \cb_3_5_io_eo[40] ,
    \cb_3_5_io_eo[39] ,
    \cb_3_5_io_eo[38] ,
    \cb_3_5_io_eo[37] ,
    \cb_3_5_io_eo[36] ,
    \cb_3_5_io_eo[35] ,
    \cb_3_5_io_eo[34] ,
    \cb_3_5_io_eo[33] ,
    \cb_3_5_io_eo[32] ,
    \cb_3_5_io_eo[31] ,
    \cb_3_5_io_eo[30] ,
    \cb_3_5_io_eo[29] ,
    \cb_3_5_io_eo[28] ,
    \cb_3_5_io_eo[27] ,
    \cb_3_5_io_eo[26] ,
    \cb_3_5_io_eo[25] ,
    \cb_3_5_io_eo[24] ,
    \cb_3_5_io_eo[23] ,
    \cb_3_5_io_eo[22] ,
    \cb_3_5_io_eo[21] ,
    \cb_3_5_io_eo[20] ,
    \cb_3_5_io_eo[19] ,
    \cb_3_5_io_eo[18] ,
    \cb_3_5_io_eo[17] ,
    \cb_3_5_io_eo[16] ,
    \cb_3_5_io_eo[15] ,
    \cb_3_5_io_eo[14] ,
    \cb_3_5_io_eo[13] ,
    \cb_3_5_io_eo[12] ,
    \cb_3_5_io_eo[11] ,
    \cb_3_5_io_eo[10] ,
    \cb_3_5_io_eo[9] ,
    \cb_3_5_io_eo[8] ,
    \cb_3_5_io_eo[7] ,
    \cb_3_5_io_eo[6] ,
    \cb_3_5_io_eo[5] ,
    \cb_3_5_io_eo[4] ,
    \cb_3_5_io_eo[3] ,
    \cb_3_5_io_eo[2] ,
    \cb_3_5_io_eo[1] ,
    \cb_3_5_io_eo[0] }));
 cic_block cb_3_7 (.io_cs_i(cb_3_7_io_cs_i),
    .io_i_0_ci(cb_3_6_io_o_0_co),
    .io_i_1_ci(cb_3_6_io_o_1_co),
    .io_i_2_ci(cb_3_6_io_o_2_co),
    .io_i_3_ci(cb_3_6_io_o_3_co),
    .io_i_4_ci(cb_3_6_io_o_4_co),
    .io_i_5_ci(cb_3_6_io_o_5_co),
    .io_i_6_ci(cb_3_6_io_o_6_co),
    .io_i_7_ci(cb_3_6_io_o_7_co),
    .io_o_0_co(cb_3_7_io_o_0_co),
    .io_o_1_co(cb_3_7_io_o_1_co),
    .io_o_2_co(cb_3_7_io_o_2_co),
    .io_o_3_co(cb_3_7_io_o_3_co),
    .io_o_4_co(cb_3_7_io_o_4_co),
    .io_o_5_co(cb_3_7_io_o_5_co),
    .io_o_6_co(cb_3_7_io_o_6_co),
    .io_o_7_co(cb_3_7_io_o_7_co),
    .io_vci(cb_3_6_io_vco),
    .io_vco(cb_3_7_io_vco),
    .io_vi(cb_3_7_io_vi),
    .io_we_i(cb_3_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_3_0_io_adr_i[1] ,
    \cb_3_0_io_adr_i[0] }),
    .io_dat_i({\cb_3_0_io_dat_i[15] ,
    \cb_3_0_io_dat_i[14] ,
    \cb_3_0_io_dat_i[13] ,
    \cb_3_0_io_dat_i[12] ,
    \cb_3_0_io_dat_i[11] ,
    \cb_3_0_io_dat_i[10] ,
    \cb_3_0_io_dat_i[9] ,
    \cb_3_0_io_dat_i[8] ,
    \cb_3_0_io_dat_i[7] ,
    \cb_3_0_io_dat_i[6] ,
    \cb_3_0_io_dat_i[5] ,
    \cb_3_0_io_dat_i[4] ,
    \cb_3_0_io_dat_i[3] ,
    \cb_3_0_io_dat_i[2] ,
    \cb_3_0_io_dat_i[1] ,
    \cb_3_0_io_dat_i[0] }),
    .io_dat_o({\cb_3_7_io_dat_o[15] ,
    \cb_3_7_io_dat_o[14] ,
    \cb_3_7_io_dat_o[13] ,
    \cb_3_7_io_dat_o[12] ,
    \cb_3_7_io_dat_o[11] ,
    \cb_3_7_io_dat_o[10] ,
    \cb_3_7_io_dat_o[9] ,
    \cb_3_7_io_dat_o[8] ,
    \cb_3_7_io_dat_o[7] ,
    \cb_3_7_io_dat_o[6] ,
    \cb_3_7_io_dat_o[5] ,
    \cb_3_7_io_dat_o[4] ,
    \cb_3_7_io_dat_o[3] ,
    \cb_3_7_io_dat_o[2] ,
    \cb_3_7_io_dat_o[1] ,
    \cb_3_7_io_dat_o[0] }),
    .io_eo({\cb_3_7_io_eo[63] ,
    \cb_3_7_io_eo[62] ,
    \cb_3_7_io_eo[61] ,
    \cb_3_7_io_eo[60] ,
    \cb_3_7_io_eo[59] ,
    \cb_3_7_io_eo[58] ,
    \cb_3_7_io_eo[57] ,
    \cb_3_7_io_eo[56] ,
    \cb_3_7_io_eo[55] ,
    \cb_3_7_io_eo[54] ,
    \cb_3_7_io_eo[53] ,
    \cb_3_7_io_eo[52] ,
    \cb_3_7_io_eo[51] ,
    \cb_3_7_io_eo[50] ,
    \cb_3_7_io_eo[49] ,
    \cb_3_7_io_eo[48] ,
    \cb_3_7_io_eo[47] ,
    \cb_3_7_io_eo[46] ,
    \cb_3_7_io_eo[45] ,
    \cb_3_7_io_eo[44] ,
    \cb_3_7_io_eo[43] ,
    \cb_3_7_io_eo[42] ,
    \cb_3_7_io_eo[41] ,
    \cb_3_7_io_eo[40] ,
    \cb_3_7_io_eo[39] ,
    \cb_3_7_io_eo[38] ,
    \cb_3_7_io_eo[37] ,
    \cb_3_7_io_eo[36] ,
    \cb_3_7_io_eo[35] ,
    \cb_3_7_io_eo[34] ,
    \cb_3_7_io_eo[33] ,
    \cb_3_7_io_eo[32] ,
    \cb_3_7_io_eo[31] ,
    \cb_3_7_io_eo[30] ,
    \cb_3_7_io_eo[29] ,
    \cb_3_7_io_eo[28] ,
    \cb_3_7_io_eo[27] ,
    \cb_3_7_io_eo[26] ,
    \cb_3_7_io_eo[25] ,
    \cb_3_7_io_eo[24] ,
    \cb_3_7_io_eo[23] ,
    \cb_3_7_io_eo[22] ,
    \cb_3_7_io_eo[21] ,
    \cb_3_7_io_eo[20] ,
    \cb_3_7_io_eo[19] ,
    \cb_3_7_io_eo[18] ,
    \cb_3_7_io_eo[17] ,
    \cb_3_7_io_eo[16] ,
    \cb_3_7_io_eo[15] ,
    \cb_3_7_io_eo[14] ,
    \cb_3_7_io_eo[13] ,
    \cb_3_7_io_eo[12] ,
    \cb_3_7_io_eo[11] ,
    \cb_3_7_io_eo[10] ,
    \cb_3_7_io_eo[9] ,
    \cb_3_7_io_eo[8] ,
    \cb_3_7_io_eo[7] ,
    \cb_3_7_io_eo[6] ,
    \cb_3_7_io_eo[5] ,
    \cb_3_7_io_eo[4] ,
    \cb_3_7_io_eo[3] ,
    \cb_3_7_io_eo[2] ,
    \cb_3_7_io_eo[1] ,
    \cb_3_7_io_eo[0] }),
    .io_i_0_in1({\cb_3_6_io_o_0_out[7] ,
    \cb_3_6_io_o_0_out[6] ,
    \cb_3_6_io_o_0_out[5] ,
    \cb_3_6_io_o_0_out[4] ,
    \cb_3_6_io_o_0_out[3] ,
    \cb_3_6_io_o_0_out[2] ,
    \cb_3_6_io_o_0_out[1] ,
    \cb_3_6_io_o_0_out[0] }),
    .io_i_1_in1({\cb_3_6_io_o_1_out[7] ,
    \cb_3_6_io_o_1_out[6] ,
    \cb_3_6_io_o_1_out[5] ,
    \cb_3_6_io_o_1_out[4] ,
    \cb_3_6_io_o_1_out[3] ,
    \cb_3_6_io_o_1_out[2] ,
    \cb_3_6_io_o_1_out[1] ,
    \cb_3_6_io_o_1_out[0] }),
    .io_i_2_in1({\cb_3_6_io_o_2_out[7] ,
    \cb_3_6_io_o_2_out[6] ,
    \cb_3_6_io_o_2_out[5] ,
    \cb_3_6_io_o_2_out[4] ,
    \cb_3_6_io_o_2_out[3] ,
    \cb_3_6_io_o_2_out[2] ,
    \cb_3_6_io_o_2_out[1] ,
    \cb_3_6_io_o_2_out[0] }),
    .io_i_3_in1({\cb_3_6_io_o_3_out[7] ,
    \cb_3_6_io_o_3_out[6] ,
    \cb_3_6_io_o_3_out[5] ,
    \cb_3_6_io_o_3_out[4] ,
    \cb_3_6_io_o_3_out[3] ,
    \cb_3_6_io_o_3_out[2] ,
    \cb_3_6_io_o_3_out[1] ,
    \cb_3_6_io_o_3_out[0] }),
    .io_i_4_in1({\cb_3_6_io_o_4_out[7] ,
    \cb_3_6_io_o_4_out[6] ,
    \cb_3_6_io_o_4_out[5] ,
    \cb_3_6_io_o_4_out[4] ,
    \cb_3_6_io_o_4_out[3] ,
    \cb_3_6_io_o_4_out[2] ,
    \cb_3_6_io_o_4_out[1] ,
    \cb_3_6_io_o_4_out[0] }),
    .io_i_5_in1({\cb_3_6_io_o_5_out[7] ,
    \cb_3_6_io_o_5_out[6] ,
    \cb_3_6_io_o_5_out[5] ,
    \cb_3_6_io_o_5_out[4] ,
    \cb_3_6_io_o_5_out[3] ,
    \cb_3_6_io_o_5_out[2] ,
    \cb_3_6_io_o_5_out[1] ,
    \cb_3_6_io_o_5_out[0] }),
    .io_i_6_in1({\cb_3_6_io_o_6_out[7] ,
    \cb_3_6_io_o_6_out[6] ,
    \cb_3_6_io_o_6_out[5] ,
    \cb_3_6_io_o_6_out[4] ,
    \cb_3_6_io_o_6_out[3] ,
    \cb_3_6_io_o_6_out[2] ,
    \cb_3_6_io_o_6_out[1] ,
    \cb_3_6_io_o_6_out[0] }),
    .io_i_7_in1({\cb_3_6_io_o_7_out[7] ,
    \cb_3_6_io_o_7_out[6] ,
    \cb_3_6_io_o_7_out[5] ,
    \cb_3_6_io_o_7_out[4] ,
    \cb_3_6_io_o_7_out[3] ,
    \cb_3_6_io_o_7_out[2] ,
    \cb_3_6_io_o_7_out[1] ,
    \cb_3_6_io_o_7_out[0] }),
    .io_o_0_out({\cb_3_7_io_o_0_out[7] ,
    \cb_3_7_io_o_0_out[6] ,
    \cb_3_7_io_o_0_out[5] ,
    \cb_3_7_io_o_0_out[4] ,
    \cb_3_7_io_o_0_out[3] ,
    \cb_3_7_io_o_0_out[2] ,
    \cb_3_7_io_o_0_out[1] ,
    \cb_3_7_io_o_0_out[0] }),
    .io_o_1_out({\cb_3_7_io_o_1_out[7] ,
    \cb_3_7_io_o_1_out[6] ,
    \cb_3_7_io_o_1_out[5] ,
    \cb_3_7_io_o_1_out[4] ,
    \cb_3_7_io_o_1_out[3] ,
    \cb_3_7_io_o_1_out[2] ,
    \cb_3_7_io_o_1_out[1] ,
    \cb_3_7_io_o_1_out[0] }),
    .io_o_2_out({\cb_3_7_io_o_2_out[7] ,
    \cb_3_7_io_o_2_out[6] ,
    \cb_3_7_io_o_2_out[5] ,
    \cb_3_7_io_o_2_out[4] ,
    \cb_3_7_io_o_2_out[3] ,
    \cb_3_7_io_o_2_out[2] ,
    \cb_3_7_io_o_2_out[1] ,
    \cb_3_7_io_o_2_out[0] }),
    .io_o_3_out({\cb_3_7_io_o_3_out[7] ,
    \cb_3_7_io_o_3_out[6] ,
    \cb_3_7_io_o_3_out[5] ,
    \cb_3_7_io_o_3_out[4] ,
    \cb_3_7_io_o_3_out[3] ,
    \cb_3_7_io_o_3_out[2] ,
    \cb_3_7_io_o_3_out[1] ,
    \cb_3_7_io_o_3_out[0] }),
    .io_o_4_out({\cb_3_7_io_o_4_out[7] ,
    \cb_3_7_io_o_4_out[6] ,
    \cb_3_7_io_o_4_out[5] ,
    \cb_3_7_io_o_4_out[4] ,
    \cb_3_7_io_o_4_out[3] ,
    \cb_3_7_io_o_4_out[2] ,
    \cb_3_7_io_o_4_out[1] ,
    \cb_3_7_io_o_4_out[0] }),
    .io_o_5_out({\cb_3_7_io_o_5_out[7] ,
    \cb_3_7_io_o_5_out[6] ,
    \cb_3_7_io_o_5_out[5] ,
    \cb_3_7_io_o_5_out[4] ,
    \cb_3_7_io_o_5_out[3] ,
    \cb_3_7_io_o_5_out[2] ,
    \cb_3_7_io_o_5_out[1] ,
    \cb_3_7_io_o_5_out[0] }),
    .io_o_6_out({\cb_3_7_io_o_6_out[7] ,
    \cb_3_7_io_o_6_out[6] ,
    \cb_3_7_io_o_6_out[5] ,
    \cb_3_7_io_o_6_out[4] ,
    \cb_3_7_io_o_6_out[3] ,
    \cb_3_7_io_o_6_out[2] ,
    \cb_3_7_io_o_6_out[1] ,
    \cb_3_7_io_o_6_out[0] }),
    .io_o_7_out({\cb_3_7_io_o_7_out[7] ,
    \cb_3_7_io_o_7_out[6] ,
    \cb_3_7_io_o_7_out[5] ,
    \cb_3_7_io_o_7_out[4] ,
    \cb_3_7_io_o_7_out[3] ,
    \cb_3_7_io_o_7_out[2] ,
    \cb_3_7_io_o_7_out[1] ,
    \cb_3_7_io_o_7_out[0] }),
    .io_wo({\cb_3_6_io_eo[63] ,
    \cb_3_6_io_eo[62] ,
    \cb_3_6_io_eo[61] ,
    \cb_3_6_io_eo[60] ,
    \cb_3_6_io_eo[59] ,
    \cb_3_6_io_eo[58] ,
    \cb_3_6_io_eo[57] ,
    \cb_3_6_io_eo[56] ,
    \cb_3_6_io_eo[55] ,
    \cb_3_6_io_eo[54] ,
    \cb_3_6_io_eo[53] ,
    \cb_3_6_io_eo[52] ,
    \cb_3_6_io_eo[51] ,
    \cb_3_6_io_eo[50] ,
    \cb_3_6_io_eo[49] ,
    \cb_3_6_io_eo[48] ,
    \cb_3_6_io_eo[47] ,
    \cb_3_6_io_eo[46] ,
    \cb_3_6_io_eo[45] ,
    \cb_3_6_io_eo[44] ,
    \cb_3_6_io_eo[43] ,
    \cb_3_6_io_eo[42] ,
    \cb_3_6_io_eo[41] ,
    \cb_3_6_io_eo[40] ,
    \cb_3_6_io_eo[39] ,
    \cb_3_6_io_eo[38] ,
    \cb_3_6_io_eo[37] ,
    \cb_3_6_io_eo[36] ,
    \cb_3_6_io_eo[35] ,
    \cb_3_6_io_eo[34] ,
    \cb_3_6_io_eo[33] ,
    \cb_3_6_io_eo[32] ,
    \cb_3_6_io_eo[31] ,
    \cb_3_6_io_eo[30] ,
    \cb_3_6_io_eo[29] ,
    \cb_3_6_io_eo[28] ,
    \cb_3_6_io_eo[27] ,
    \cb_3_6_io_eo[26] ,
    \cb_3_6_io_eo[25] ,
    \cb_3_6_io_eo[24] ,
    \cb_3_6_io_eo[23] ,
    \cb_3_6_io_eo[22] ,
    \cb_3_6_io_eo[21] ,
    \cb_3_6_io_eo[20] ,
    \cb_3_6_io_eo[19] ,
    \cb_3_6_io_eo[18] ,
    \cb_3_6_io_eo[17] ,
    \cb_3_6_io_eo[16] ,
    \cb_3_6_io_eo[15] ,
    \cb_3_6_io_eo[14] ,
    \cb_3_6_io_eo[13] ,
    \cb_3_6_io_eo[12] ,
    \cb_3_6_io_eo[11] ,
    \cb_3_6_io_eo[10] ,
    \cb_3_6_io_eo[9] ,
    \cb_3_6_io_eo[8] ,
    \cb_3_6_io_eo[7] ,
    \cb_3_6_io_eo[6] ,
    \cb_3_6_io_eo[5] ,
    \cb_3_6_io_eo[4] ,
    \cb_3_6_io_eo[3] ,
    \cb_3_6_io_eo[2] ,
    \cb_3_6_io_eo[1] ,
    \cb_3_6_io_eo[0] }));
 cic_block cb_3_8 (.io_cs_i(cb_3_8_io_cs_i),
    .io_i_0_ci(cb_3_7_io_o_0_co),
    .io_i_1_ci(cb_3_7_io_o_1_co),
    .io_i_2_ci(cb_3_7_io_o_2_co),
    .io_i_3_ci(cb_3_7_io_o_3_co),
    .io_i_4_ci(cb_3_7_io_o_4_co),
    .io_i_5_ci(cb_3_7_io_o_5_co),
    .io_i_6_ci(cb_3_7_io_o_6_co),
    .io_i_7_ci(cb_3_7_io_o_7_co),
    .io_o_0_co(cb_3_8_io_o_0_co),
    .io_o_1_co(cb_3_8_io_o_1_co),
    .io_o_2_co(cb_3_8_io_o_2_co),
    .io_o_3_co(cb_3_8_io_o_3_co),
    .io_o_4_co(cb_3_8_io_o_4_co),
    .io_o_5_co(cb_3_8_io_o_5_co),
    .io_o_6_co(cb_3_8_io_o_6_co),
    .io_o_7_co(cb_3_8_io_o_7_co),
    .io_vci(cb_3_7_io_vco),
    .io_vco(cb_3_8_io_vco),
    .io_vi(cb_3_8_io_vi),
    .io_we_i(cb_3_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_3_0_io_adr_i[1] ,
    \cb_3_0_io_adr_i[0] }),
    .io_dat_i({\cb_3_0_io_dat_i[15] ,
    \cb_3_0_io_dat_i[14] ,
    \cb_3_0_io_dat_i[13] ,
    \cb_3_0_io_dat_i[12] ,
    \cb_3_0_io_dat_i[11] ,
    \cb_3_0_io_dat_i[10] ,
    \cb_3_0_io_dat_i[9] ,
    \cb_3_0_io_dat_i[8] ,
    \cb_3_0_io_dat_i[7] ,
    \cb_3_0_io_dat_i[6] ,
    \cb_3_0_io_dat_i[5] ,
    \cb_3_0_io_dat_i[4] ,
    \cb_3_0_io_dat_i[3] ,
    \cb_3_0_io_dat_i[2] ,
    \cb_3_0_io_dat_i[1] ,
    \cb_3_0_io_dat_i[0] }),
    .io_dat_o({\cb_3_8_io_dat_o[15] ,
    \cb_3_8_io_dat_o[14] ,
    \cb_3_8_io_dat_o[13] ,
    \cb_3_8_io_dat_o[12] ,
    \cb_3_8_io_dat_o[11] ,
    \cb_3_8_io_dat_o[10] ,
    \cb_3_8_io_dat_o[9] ,
    \cb_3_8_io_dat_o[8] ,
    \cb_3_8_io_dat_o[7] ,
    \cb_3_8_io_dat_o[6] ,
    \cb_3_8_io_dat_o[5] ,
    \cb_3_8_io_dat_o[4] ,
    \cb_3_8_io_dat_o[3] ,
    \cb_3_8_io_dat_o[2] ,
    \cb_3_8_io_dat_o[1] ,
    \cb_3_8_io_dat_o[0] }),
    .io_eo({\cb_3_8_io_eo[63] ,
    \cb_3_8_io_eo[62] ,
    \cb_3_8_io_eo[61] ,
    \cb_3_8_io_eo[60] ,
    \cb_3_8_io_eo[59] ,
    \cb_3_8_io_eo[58] ,
    \cb_3_8_io_eo[57] ,
    \cb_3_8_io_eo[56] ,
    \cb_3_8_io_eo[55] ,
    \cb_3_8_io_eo[54] ,
    \cb_3_8_io_eo[53] ,
    \cb_3_8_io_eo[52] ,
    \cb_3_8_io_eo[51] ,
    \cb_3_8_io_eo[50] ,
    \cb_3_8_io_eo[49] ,
    \cb_3_8_io_eo[48] ,
    \cb_3_8_io_eo[47] ,
    \cb_3_8_io_eo[46] ,
    \cb_3_8_io_eo[45] ,
    \cb_3_8_io_eo[44] ,
    \cb_3_8_io_eo[43] ,
    \cb_3_8_io_eo[42] ,
    \cb_3_8_io_eo[41] ,
    \cb_3_8_io_eo[40] ,
    \cb_3_8_io_eo[39] ,
    \cb_3_8_io_eo[38] ,
    \cb_3_8_io_eo[37] ,
    \cb_3_8_io_eo[36] ,
    \cb_3_8_io_eo[35] ,
    \cb_3_8_io_eo[34] ,
    \cb_3_8_io_eo[33] ,
    \cb_3_8_io_eo[32] ,
    \cb_3_8_io_eo[31] ,
    \cb_3_8_io_eo[30] ,
    \cb_3_8_io_eo[29] ,
    \cb_3_8_io_eo[28] ,
    \cb_3_8_io_eo[27] ,
    \cb_3_8_io_eo[26] ,
    \cb_3_8_io_eo[25] ,
    \cb_3_8_io_eo[24] ,
    \cb_3_8_io_eo[23] ,
    \cb_3_8_io_eo[22] ,
    \cb_3_8_io_eo[21] ,
    \cb_3_8_io_eo[20] ,
    \cb_3_8_io_eo[19] ,
    \cb_3_8_io_eo[18] ,
    \cb_3_8_io_eo[17] ,
    \cb_3_8_io_eo[16] ,
    \cb_3_8_io_eo[15] ,
    \cb_3_8_io_eo[14] ,
    \cb_3_8_io_eo[13] ,
    \cb_3_8_io_eo[12] ,
    \cb_3_8_io_eo[11] ,
    \cb_3_8_io_eo[10] ,
    \cb_3_8_io_eo[9] ,
    \cb_3_8_io_eo[8] ,
    \cb_3_8_io_eo[7] ,
    \cb_3_8_io_eo[6] ,
    \cb_3_8_io_eo[5] ,
    \cb_3_8_io_eo[4] ,
    \cb_3_8_io_eo[3] ,
    \cb_3_8_io_eo[2] ,
    \cb_3_8_io_eo[1] ,
    \cb_3_8_io_eo[0] }),
    .io_i_0_in1({\cb_3_7_io_o_0_out[7] ,
    \cb_3_7_io_o_0_out[6] ,
    \cb_3_7_io_o_0_out[5] ,
    \cb_3_7_io_o_0_out[4] ,
    \cb_3_7_io_o_0_out[3] ,
    \cb_3_7_io_o_0_out[2] ,
    \cb_3_7_io_o_0_out[1] ,
    \cb_3_7_io_o_0_out[0] }),
    .io_i_1_in1({\cb_3_7_io_o_1_out[7] ,
    \cb_3_7_io_o_1_out[6] ,
    \cb_3_7_io_o_1_out[5] ,
    \cb_3_7_io_o_1_out[4] ,
    \cb_3_7_io_o_1_out[3] ,
    \cb_3_7_io_o_1_out[2] ,
    \cb_3_7_io_o_1_out[1] ,
    \cb_3_7_io_o_1_out[0] }),
    .io_i_2_in1({\cb_3_7_io_o_2_out[7] ,
    \cb_3_7_io_o_2_out[6] ,
    \cb_3_7_io_o_2_out[5] ,
    \cb_3_7_io_o_2_out[4] ,
    \cb_3_7_io_o_2_out[3] ,
    \cb_3_7_io_o_2_out[2] ,
    \cb_3_7_io_o_2_out[1] ,
    \cb_3_7_io_o_2_out[0] }),
    .io_i_3_in1({\cb_3_7_io_o_3_out[7] ,
    \cb_3_7_io_o_3_out[6] ,
    \cb_3_7_io_o_3_out[5] ,
    \cb_3_7_io_o_3_out[4] ,
    \cb_3_7_io_o_3_out[3] ,
    \cb_3_7_io_o_3_out[2] ,
    \cb_3_7_io_o_3_out[1] ,
    \cb_3_7_io_o_3_out[0] }),
    .io_i_4_in1({\cb_3_7_io_o_4_out[7] ,
    \cb_3_7_io_o_4_out[6] ,
    \cb_3_7_io_o_4_out[5] ,
    \cb_3_7_io_o_4_out[4] ,
    \cb_3_7_io_o_4_out[3] ,
    \cb_3_7_io_o_4_out[2] ,
    \cb_3_7_io_o_4_out[1] ,
    \cb_3_7_io_o_4_out[0] }),
    .io_i_5_in1({\cb_3_7_io_o_5_out[7] ,
    \cb_3_7_io_o_5_out[6] ,
    \cb_3_7_io_o_5_out[5] ,
    \cb_3_7_io_o_5_out[4] ,
    \cb_3_7_io_o_5_out[3] ,
    \cb_3_7_io_o_5_out[2] ,
    \cb_3_7_io_o_5_out[1] ,
    \cb_3_7_io_o_5_out[0] }),
    .io_i_6_in1({\cb_3_7_io_o_6_out[7] ,
    \cb_3_7_io_o_6_out[6] ,
    \cb_3_7_io_o_6_out[5] ,
    \cb_3_7_io_o_6_out[4] ,
    \cb_3_7_io_o_6_out[3] ,
    \cb_3_7_io_o_6_out[2] ,
    \cb_3_7_io_o_6_out[1] ,
    \cb_3_7_io_o_6_out[0] }),
    .io_i_7_in1({\cb_3_7_io_o_7_out[7] ,
    \cb_3_7_io_o_7_out[6] ,
    \cb_3_7_io_o_7_out[5] ,
    \cb_3_7_io_o_7_out[4] ,
    \cb_3_7_io_o_7_out[3] ,
    \cb_3_7_io_o_7_out[2] ,
    \cb_3_7_io_o_7_out[1] ,
    \cb_3_7_io_o_7_out[0] }),
    .io_o_0_out({\cb_3_8_io_o_0_out[7] ,
    \cb_3_8_io_o_0_out[6] ,
    \cb_3_8_io_o_0_out[5] ,
    \cb_3_8_io_o_0_out[4] ,
    \cb_3_8_io_o_0_out[3] ,
    \cb_3_8_io_o_0_out[2] ,
    \cb_3_8_io_o_0_out[1] ,
    \cb_3_8_io_o_0_out[0] }),
    .io_o_1_out({\cb_3_8_io_o_1_out[7] ,
    \cb_3_8_io_o_1_out[6] ,
    \cb_3_8_io_o_1_out[5] ,
    \cb_3_8_io_o_1_out[4] ,
    \cb_3_8_io_o_1_out[3] ,
    \cb_3_8_io_o_1_out[2] ,
    \cb_3_8_io_o_1_out[1] ,
    \cb_3_8_io_o_1_out[0] }),
    .io_o_2_out({\cb_3_8_io_o_2_out[7] ,
    \cb_3_8_io_o_2_out[6] ,
    \cb_3_8_io_o_2_out[5] ,
    \cb_3_8_io_o_2_out[4] ,
    \cb_3_8_io_o_2_out[3] ,
    \cb_3_8_io_o_2_out[2] ,
    \cb_3_8_io_o_2_out[1] ,
    \cb_3_8_io_o_2_out[0] }),
    .io_o_3_out({\cb_3_8_io_o_3_out[7] ,
    \cb_3_8_io_o_3_out[6] ,
    \cb_3_8_io_o_3_out[5] ,
    \cb_3_8_io_o_3_out[4] ,
    \cb_3_8_io_o_3_out[3] ,
    \cb_3_8_io_o_3_out[2] ,
    \cb_3_8_io_o_3_out[1] ,
    \cb_3_8_io_o_3_out[0] }),
    .io_o_4_out({\cb_3_8_io_o_4_out[7] ,
    \cb_3_8_io_o_4_out[6] ,
    \cb_3_8_io_o_4_out[5] ,
    \cb_3_8_io_o_4_out[4] ,
    \cb_3_8_io_o_4_out[3] ,
    \cb_3_8_io_o_4_out[2] ,
    \cb_3_8_io_o_4_out[1] ,
    \cb_3_8_io_o_4_out[0] }),
    .io_o_5_out({\cb_3_8_io_o_5_out[7] ,
    \cb_3_8_io_o_5_out[6] ,
    \cb_3_8_io_o_5_out[5] ,
    \cb_3_8_io_o_5_out[4] ,
    \cb_3_8_io_o_5_out[3] ,
    \cb_3_8_io_o_5_out[2] ,
    \cb_3_8_io_o_5_out[1] ,
    \cb_3_8_io_o_5_out[0] }),
    .io_o_6_out({\cb_3_8_io_o_6_out[7] ,
    \cb_3_8_io_o_6_out[6] ,
    \cb_3_8_io_o_6_out[5] ,
    \cb_3_8_io_o_6_out[4] ,
    \cb_3_8_io_o_6_out[3] ,
    \cb_3_8_io_o_6_out[2] ,
    \cb_3_8_io_o_6_out[1] ,
    \cb_3_8_io_o_6_out[0] }),
    .io_o_7_out({\cb_3_8_io_o_7_out[7] ,
    \cb_3_8_io_o_7_out[6] ,
    \cb_3_8_io_o_7_out[5] ,
    \cb_3_8_io_o_7_out[4] ,
    \cb_3_8_io_o_7_out[3] ,
    \cb_3_8_io_o_7_out[2] ,
    \cb_3_8_io_o_7_out[1] ,
    \cb_3_8_io_o_7_out[0] }),
    .io_wo({\cb_3_7_io_eo[63] ,
    \cb_3_7_io_eo[62] ,
    \cb_3_7_io_eo[61] ,
    \cb_3_7_io_eo[60] ,
    \cb_3_7_io_eo[59] ,
    \cb_3_7_io_eo[58] ,
    \cb_3_7_io_eo[57] ,
    \cb_3_7_io_eo[56] ,
    \cb_3_7_io_eo[55] ,
    \cb_3_7_io_eo[54] ,
    \cb_3_7_io_eo[53] ,
    \cb_3_7_io_eo[52] ,
    \cb_3_7_io_eo[51] ,
    \cb_3_7_io_eo[50] ,
    \cb_3_7_io_eo[49] ,
    \cb_3_7_io_eo[48] ,
    \cb_3_7_io_eo[47] ,
    \cb_3_7_io_eo[46] ,
    \cb_3_7_io_eo[45] ,
    \cb_3_7_io_eo[44] ,
    \cb_3_7_io_eo[43] ,
    \cb_3_7_io_eo[42] ,
    \cb_3_7_io_eo[41] ,
    \cb_3_7_io_eo[40] ,
    \cb_3_7_io_eo[39] ,
    \cb_3_7_io_eo[38] ,
    \cb_3_7_io_eo[37] ,
    \cb_3_7_io_eo[36] ,
    \cb_3_7_io_eo[35] ,
    \cb_3_7_io_eo[34] ,
    \cb_3_7_io_eo[33] ,
    \cb_3_7_io_eo[32] ,
    \cb_3_7_io_eo[31] ,
    \cb_3_7_io_eo[30] ,
    \cb_3_7_io_eo[29] ,
    \cb_3_7_io_eo[28] ,
    \cb_3_7_io_eo[27] ,
    \cb_3_7_io_eo[26] ,
    \cb_3_7_io_eo[25] ,
    \cb_3_7_io_eo[24] ,
    \cb_3_7_io_eo[23] ,
    \cb_3_7_io_eo[22] ,
    \cb_3_7_io_eo[21] ,
    \cb_3_7_io_eo[20] ,
    \cb_3_7_io_eo[19] ,
    \cb_3_7_io_eo[18] ,
    \cb_3_7_io_eo[17] ,
    \cb_3_7_io_eo[16] ,
    \cb_3_7_io_eo[15] ,
    \cb_3_7_io_eo[14] ,
    \cb_3_7_io_eo[13] ,
    \cb_3_7_io_eo[12] ,
    \cb_3_7_io_eo[11] ,
    \cb_3_7_io_eo[10] ,
    \cb_3_7_io_eo[9] ,
    \cb_3_7_io_eo[8] ,
    \cb_3_7_io_eo[7] ,
    \cb_3_7_io_eo[6] ,
    \cb_3_7_io_eo[5] ,
    \cb_3_7_io_eo[4] ,
    \cb_3_7_io_eo[3] ,
    \cb_3_7_io_eo[2] ,
    \cb_3_7_io_eo[1] ,
    \cb_3_7_io_eo[0] }));
 cic_block cb_3_9 (.io_cs_i(cb_3_9_io_cs_i),
    .io_i_0_ci(cb_3_8_io_o_0_co),
    .io_i_1_ci(cb_3_8_io_o_1_co),
    .io_i_2_ci(cb_3_8_io_o_2_co),
    .io_i_3_ci(cb_3_8_io_o_3_co),
    .io_i_4_ci(cb_3_8_io_o_4_co),
    .io_i_5_ci(cb_3_8_io_o_5_co),
    .io_i_6_ci(cb_3_8_io_o_6_co),
    .io_i_7_ci(cb_3_8_io_o_7_co),
    .io_o_0_co(cb_3_10_io_i_0_ci),
    .io_o_1_co(cb_3_10_io_i_1_ci),
    .io_o_2_co(cb_3_10_io_i_2_ci),
    .io_o_3_co(cb_3_10_io_i_3_ci),
    .io_o_4_co(cb_3_10_io_i_4_ci),
    .io_o_5_co(cb_3_10_io_i_5_ci),
    .io_o_6_co(cb_3_10_io_i_6_ci),
    .io_o_7_co(cb_3_10_io_i_7_ci),
    .io_vci(cb_3_8_io_vco),
    .io_vco(cb_3_10_io_vci),
    .io_vi(cb_3_9_io_vi),
    .io_we_i(cb_3_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_3_0_io_adr_i[1] ,
    \cb_3_0_io_adr_i[0] }),
    .io_dat_i({\cb_3_0_io_dat_i[15] ,
    \cb_3_0_io_dat_i[14] ,
    \cb_3_0_io_dat_i[13] ,
    \cb_3_0_io_dat_i[12] ,
    \cb_3_0_io_dat_i[11] ,
    \cb_3_0_io_dat_i[10] ,
    \cb_3_0_io_dat_i[9] ,
    \cb_3_0_io_dat_i[8] ,
    \cb_3_0_io_dat_i[7] ,
    \cb_3_0_io_dat_i[6] ,
    \cb_3_0_io_dat_i[5] ,
    \cb_3_0_io_dat_i[4] ,
    \cb_3_0_io_dat_i[3] ,
    \cb_3_0_io_dat_i[2] ,
    \cb_3_0_io_dat_i[1] ,
    \cb_3_0_io_dat_i[0] }),
    .io_dat_o({\cb_3_9_io_dat_o[15] ,
    \cb_3_9_io_dat_o[14] ,
    \cb_3_9_io_dat_o[13] ,
    \cb_3_9_io_dat_o[12] ,
    \cb_3_9_io_dat_o[11] ,
    \cb_3_9_io_dat_o[10] ,
    \cb_3_9_io_dat_o[9] ,
    \cb_3_9_io_dat_o[8] ,
    \cb_3_9_io_dat_o[7] ,
    \cb_3_9_io_dat_o[6] ,
    \cb_3_9_io_dat_o[5] ,
    \cb_3_9_io_dat_o[4] ,
    \cb_3_9_io_dat_o[3] ,
    \cb_3_9_io_dat_o[2] ,
    \cb_3_9_io_dat_o[1] ,
    \cb_3_9_io_dat_o[0] }),
    .io_eo({\cb_3_10_io_wo[63] ,
    \cb_3_10_io_wo[62] ,
    \cb_3_10_io_wo[61] ,
    \cb_3_10_io_wo[60] ,
    \cb_3_10_io_wo[59] ,
    \cb_3_10_io_wo[58] ,
    \cb_3_10_io_wo[57] ,
    \cb_3_10_io_wo[56] ,
    \cb_3_10_io_wo[55] ,
    \cb_3_10_io_wo[54] ,
    \cb_3_10_io_wo[53] ,
    \cb_3_10_io_wo[52] ,
    \cb_3_10_io_wo[51] ,
    \cb_3_10_io_wo[50] ,
    \cb_3_10_io_wo[49] ,
    \cb_3_10_io_wo[48] ,
    \cb_3_10_io_wo[47] ,
    \cb_3_10_io_wo[46] ,
    \cb_3_10_io_wo[45] ,
    \cb_3_10_io_wo[44] ,
    \cb_3_10_io_wo[43] ,
    \cb_3_10_io_wo[42] ,
    \cb_3_10_io_wo[41] ,
    \cb_3_10_io_wo[40] ,
    \cb_3_10_io_wo[39] ,
    \cb_3_10_io_wo[38] ,
    \cb_3_10_io_wo[37] ,
    \cb_3_10_io_wo[36] ,
    \cb_3_10_io_wo[35] ,
    \cb_3_10_io_wo[34] ,
    \cb_3_10_io_wo[33] ,
    \cb_3_10_io_wo[32] ,
    \cb_3_10_io_wo[31] ,
    \cb_3_10_io_wo[30] ,
    \cb_3_10_io_wo[29] ,
    \cb_3_10_io_wo[28] ,
    \cb_3_10_io_wo[27] ,
    \cb_3_10_io_wo[26] ,
    \cb_3_10_io_wo[25] ,
    \cb_3_10_io_wo[24] ,
    \cb_3_10_io_wo[23] ,
    \cb_3_10_io_wo[22] ,
    \cb_3_10_io_wo[21] ,
    \cb_3_10_io_wo[20] ,
    \cb_3_10_io_wo[19] ,
    \cb_3_10_io_wo[18] ,
    \cb_3_10_io_wo[17] ,
    \cb_3_10_io_wo[16] ,
    \cb_3_10_io_wo[15] ,
    \cb_3_10_io_wo[14] ,
    \cb_3_10_io_wo[13] ,
    \cb_3_10_io_wo[12] ,
    \cb_3_10_io_wo[11] ,
    \cb_3_10_io_wo[10] ,
    \cb_3_10_io_wo[9] ,
    \cb_3_10_io_wo[8] ,
    \cb_3_10_io_wo[7] ,
    \cb_3_10_io_wo[6] ,
    \cb_3_10_io_wo[5] ,
    \cb_3_10_io_wo[4] ,
    \cb_3_10_io_wo[3] ,
    \cb_3_10_io_wo[2] ,
    \cb_3_10_io_wo[1] ,
    \cb_3_10_io_wo[0] }),
    .io_i_0_in1({\cb_3_8_io_o_0_out[7] ,
    \cb_3_8_io_o_0_out[6] ,
    \cb_3_8_io_o_0_out[5] ,
    \cb_3_8_io_o_0_out[4] ,
    \cb_3_8_io_o_0_out[3] ,
    \cb_3_8_io_o_0_out[2] ,
    \cb_3_8_io_o_0_out[1] ,
    \cb_3_8_io_o_0_out[0] }),
    .io_i_1_in1({\cb_3_8_io_o_1_out[7] ,
    \cb_3_8_io_o_1_out[6] ,
    \cb_3_8_io_o_1_out[5] ,
    \cb_3_8_io_o_1_out[4] ,
    \cb_3_8_io_o_1_out[3] ,
    \cb_3_8_io_o_1_out[2] ,
    \cb_3_8_io_o_1_out[1] ,
    \cb_3_8_io_o_1_out[0] }),
    .io_i_2_in1({\cb_3_8_io_o_2_out[7] ,
    \cb_3_8_io_o_2_out[6] ,
    \cb_3_8_io_o_2_out[5] ,
    \cb_3_8_io_o_2_out[4] ,
    \cb_3_8_io_o_2_out[3] ,
    \cb_3_8_io_o_2_out[2] ,
    \cb_3_8_io_o_2_out[1] ,
    \cb_3_8_io_o_2_out[0] }),
    .io_i_3_in1({\cb_3_8_io_o_3_out[7] ,
    \cb_3_8_io_o_3_out[6] ,
    \cb_3_8_io_o_3_out[5] ,
    \cb_3_8_io_o_3_out[4] ,
    \cb_3_8_io_o_3_out[3] ,
    \cb_3_8_io_o_3_out[2] ,
    \cb_3_8_io_o_3_out[1] ,
    \cb_3_8_io_o_3_out[0] }),
    .io_i_4_in1({\cb_3_8_io_o_4_out[7] ,
    \cb_3_8_io_o_4_out[6] ,
    \cb_3_8_io_o_4_out[5] ,
    \cb_3_8_io_o_4_out[4] ,
    \cb_3_8_io_o_4_out[3] ,
    \cb_3_8_io_o_4_out[2] ,
    \cb_3_8_io_o_4_out[1] ,
    \cb_3_8_io_o_4_out[0] }),
    .io_i_5_in1({\cb_3_8_io_o_5_out[7] ,
    \cb_3_8_io_o_5_out[6] ,
    \cb_3_8_io_o_5_out[5] ,
    \cb_3_8_io_o_5_out[4] ,
    \cb_3_8_io_o_5_out[3] ,
    \cb_3_8_io_o_5_out[2] ,
    \cb_3_8_io_o_5_out[1] ,
    \cb_3_8_io_o_5_out[0] }),
    .io_i_6_in1({\cb_3_8_io_o_6_out[7] ,
    \cb_3_8_io_o_6_out[6] ,
    \cb_3_8_io_o_6_out[5] ,
    \cb_3_8_io_o_6_out[4] ,
    \cb_3_8_io_o_6_out[3] ,
    \cb_3_8_io_o_6_out[2] ,
    \cb_3_8_io_o_6_out[1] ,
    \cb_3_8_io_o_6_out[0] }),
    .io_i_7_in1({\cb_3_8_io_o_7_out[7] ,
    \cb_3_8_io_o_7_out[6] ,
    \cb_3_8_io_o_7_out[5] ,
    \cb_3_8_io_o_7_out[4] ,
    \cb_3_8_io_o_7_out[3] ,
    \cb_3_8_io_o_7_out[2] ,
    \cb_3_8_io_o_7_out[1] ,
    \cb_3_8_io_o_7_out[0] }),
    .io_o_0_out({\cb_3_10_io_i_0_in1[7] ,
    \cb_3_10_io_i_0_in1[6] ,
    \cb_3_10_io_i_0_in1[5] ,
    \cb_3_10_io_i_0_in1[4] ,
    \cb_3_10_io_i_0_in1[3] ,
    \cb_3_10_io_i_0_in1[2] ,
    \cb_3_10_io_i_0_in1[1] ,
    \cb_3_10_io_i_0_in1[0] }),
    .io_o_1_out({\cb_3_10_io_i_1_in1[7] ,
    \cb_3_10_io_i_1_in1[6] ,
    \cb_3_10_io_i_1_in1[5] ,
    \cb_3_10_io_i_1_in1[4] ,
    \cb_3_10_io_i_1_in1[3] ,
    \cb_3_10_io_i_1_in1[2] ,
    \cb_3_10_io_i_1_in1[1] ,
    \cb_3_10_io_i_1_in1[0] }),
    .io_o_2_out({\cb_3_10_io_i_2_in1[7] ,
    \cb_3_10_io_i_2_in1[6] ,
    \cb_3_10_io_i_2_in1[5] ,
    \cb_3_10_io_i_2_in1[4] ,
    \cb_3_10_io_i_2_in1[3] ,
    \cb_3_10_io_i_2_in1[2] ,
    \cb_3_10_io_i_2_in1[1] ,
    \cb_3_10_io_i_2_in1[0] }),
    .io_o_3_out({\cb_3_10_io_i_3_in1[7] ,
    \cb_3_10_io_i_3_in1[6] ,
    \cb_3_10_io_i_3_in1[5] ,
    \cb_3_10_io_i_3_in1[4] ,
    \cb_3_10_io_i_3_in1[3] ,
    \cb_3_10_io_i_3_in1[2] ,
    \cb_3_10_io_i_3_in1[1] ,
    \cb_3_10_io_i_3_in1[0] }),
    .io_o_4_out({\cb_3_10_io_i_4_in1[7] ,
    \cb_3_10_io_i_4_in1[6] ,
    \cb_3_10_io_i_4_in1[5] ,
    \cb_3_10_io_i_4_in1[4] ,
    \cb_3_10_io_i_4_in1[3] ,
    \cb_3_10_io_i_4_in1[2] ,
    \cb_3_10_io_i_4_in1[1] ,
    \cb_3_10_io_i_4_in1[0] }),
    .io_o_5_out({\cb_3_10_io_i_5_in1[7] ,
    \cb_3_10_io_i_5_in1[6] ,
    \cb_3_10_io_i_5_in1[5] ,
    \cb_3_10_io_i_5_in1[4] ,
    \cb_3_10_io_i_5_in1[3] ,
    \cb_3_10_io_i_5_in1[2] ,
    \cb_3_10_io_i_5_in1[1] ,
    \cb_3_10_io_i_5_in1[0] }),
    .io_o_6_out({\cb_3_10_io_i_6_in1[7] ,
    \cb_3_10_io_i_6_in1[6] ,
    \cb_3_10_io_i_6_in1[5] ,
    \cb_3_10_io_i_6_in1[4] ,
    \cb_3_10_io_i_6_in1[3] ,
    \cb_3_10_io_i_6_in1[2] ,
    \cb_3_10_io_i_6_in1[1] ,
    \cb_3_10_io_i_6_in1[0] }),
    .io_o_7_out({\cb_3_10_io_i_7_in1[7] ,
    \cb_3_10_io_i_7_in1[6] ,
    \cb_3_10_io_i_7_in1[5] ,
    \cb_3_10_io_i_7_in1[4] ,
    \cb_3_10_io_i_7_in1[3] ,
    \cb_3_10_io_i_7_in1[2] ,
    \cb_3_10_io_i_7_in1[1] ,
    \cb_3_10_io_i_7_in1[0] }),
    .io_wo({\cb_3_8_io_eo[63] ,
    \cb_3_8_io_eo[62] ,
    \cb_3_8_io_eo[61] ,
    \cb_3_8_io_eo[60] ,
    \cb_3_8_io_eo[59] ,
    \cb_3_8_io_eo[58] ,
    \cb_3_8_io_eo[57] ,
    \cb_3_8_io_eo[56] ,
    \cb_3_8_io_eo[55] ,
    \cb_3_8_io_eo[54] ,
    \cb_3_8_io_eo[53] ,
    \cb_3_8_io_eo[52] ,
    \cb_3_8_io_eo[51] ,
    \cb_3_8_io_eo[50] ,
    \cb_3_8_io_eo[49] ,
    \cb_3_8_io_eo[48] ,
    \cb_3_8_io_eo[47] ,
    \cb_3_8_io_eo[46] ,
    \cb_3_8_io_eo[45] ,
    \cb_3_8_io_eo[44] ,
    \cb_3_8_io_eo[43] ,
    \cb_3_8_io_eo[42] ,
    \cb_3_8_io_eo[41] ,
    \cb_3_8_io_eo[40] ,
    \cb_3_8_io_eo[39] ,
    \cb_3_8_io_eo[38] ,
    \cb_3_8_io_eo[37] ,
    \cb_3_8_io_eo[36] ,
    \cb_3_8_io_eo[35] ,
    \cb_3_8_io_eo[34] ,
    \cb_3_8_io_eo[33] ,
    \cb_3_8_io_eo[32] ,
    \cb_3_8_io_eo[31] ,
    \cb_3_8_io_eo[30] ,
    \cb_3_8_io_eo[29] ,
    \cb_3_8_io_eo[28] ,
    \cb_3_8_io_eo[27] ,
    \cb_3_8_io_eo[26] ,
    \cb_3_8_io_eo[25] ,
    \cb_3_8_io_eo[24] ,
    \cb_3_8_io_eo[23] ,
    \cb_3_8_io_eo[22] ,
    \cb_3_8_io_eo[21] ,
    \cb_3_8_io_eo[20] ,
    \cb_3_8_io_eo[19] ,
    \cb_3_8_io_eo[18] ,
    \cb_3_8_io_eo[17] ,
    \cb_3_8_io_eo[16] ,
    \cb_3_8_io_eo[15] ,
    \cb_3_8_io_eo[14] ,
    \cb_3_8_io_eo[13] ,
    \cb_3_8_io_eo[12] ,
    \cb_3_8_io_eo[11] ,
    \cb_3_8_io_eo[10] ,
    \cb_3_8_io_eo[9] ,
    \cb_3_8_io_eo[8] ,
    \cb_3_8_io_eo[7] ,
    \cb_3_8_io_eo[6] ,
    \cb_3_8_io_eo[5] ,
    \cb_3_8_io_eo[4] ,
    \cb_3_8_io_eo[3] ,
    \cb_3_8_io_eo[2] ,
    \cb_3_8_io_eo[1] ,
    \cb_3_8_io_eo[0] }));
 cic_block cb_4_0 (.io_cs_i(cb_4_0_io_cs_i),
    .io_i_0_ci(cb_4_0_io_i_0_ci),
    .io_o_0_co(cb_4_0_io_o_0_co),
    .io_o_1_co(cb_4_0_io_o_1_co),
    .io_o_2_co(cb_4_0_io_o_2_co),
    .io_o_3_co(cb_4_0_io_o_3_co),
    .io_o_4_co(cb_4_0_io_o_4_co),
    .io_o_5_co(cb_4_0_io_o_5_co),
    .io_o_6_co(cb_4_0_io_o_6_co),
    .io_o_7_co(cb_4_0_io_o_7_co),
    .io_vco(cb_4_0_io_vco),
    .io_vi(cb_4_0_io_vi),
    .io_we_i(cb_4_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_4_0_io_adr_i[1] ,
    \cb_4_0_io_adr_i[0] }),
    .io_dat_i({\cb_4_0_io_dat_i[15] ,
    \cb_4_0_io_dat_i[14] ,
    \cb_4_0_io_dat_i[13] ,
    \cb_4_0_io_dat_i[12] ,
    \cb_4_0_io_dat_i[11] ,
    \cb_4_0_io_dat_i[10] ,
    \cb_4_0_io_dat_i[9] ,
    \cb_4_0_io_dat_i[8] ,
    \cb_4_0_io_dat_i[7] ,
    \cb_4_0_io_dat_i[6] ,
    \cb_4_0_io_dat_i[5] ,
    \cb_4_0_io_dat_i[4] ,
    \cb_4_0_io_dat_i[3] ,
    \cb_4_0_io_dat_i[2] ,
    \cb_4_0_io_dat_i[1] ,
    \cb_4_0_io_dat_i[0] }),
    .io_dat_o({\cb_4_0_io_dat_o[15] ,
    \cb_4_0_io_dat_o[14] ,
    \cb_4_0_io_dat_o[13] ,
    \cb_4_0_io_dat_o[12] ,
    \cb_4_0_io_dat_o[11] ,
    \cb_4_0_io_dat_o[10] ,
    \cb_4_0_io_dat_o[9] ,
    \cb_4_0_io_dat_o[8] ,
    \cb_4_0_io_dat_o[7] ,
    \cb_4_0_io_dat_o[6] ,
    \cb_4_0_io_dat_o[5] ,
    \cb_4_0_io_dat_o[4] ,
    \cb_4_0_io_dat_o[3] ,
    \cb_4_0_io_dat_o[2] ,
    \cb_4_0_io_dat_o[1] ,
    \cb_4_0_io_dat_o[0] }),
    .io_eo({\cb_4_0_io_eo[63] ,
    \cb_4_0_io_eo[62] ,
    \cb_4_0_io_eo[61] ,
    \cb_4_0_io_eo[60] ,
    \cb_4_0_io_eo[59] ,
    \cb_4_0_io_eo[58] ,
    \cb_4_0_io_eo[57] ,
    \cb_4_0_io_eo[56] ,
    \cb_4_0_io_eo[55] ,
    \cb_4_0_io_eo[54] ,
    \cb_4_0_io_eo[53] ,
    \cb_4_0_io_eo[52] ,
    \cb_4_0_io_eo[51] ,
    \cb_4_0_io_eo[50] ,
    \cb_4_0_io_eo[49] ,
    \cb_4_0_io_eo[48] ,
    \cb_4_0_io_eo[47] ,
    \cb_4_0_io_eo[46] ,
    \cb_4_0_io_eo[45] ,
    \cb_4_0_io_eo[44] ,
    \cb_4_0_io_eo[43] ,
    \cb_4_0_io_eo[42] ,
    \cb_4_0_io_eo[41] ,
    \cb_4_0_io_eo[40] ,
    \cb_4_0_io_eo[39] ,
    \cb_4_0_io_eo[38] ,
    \cb_4_0_io_eo[37] ,
    \cb_4_0_io_eo[36] ,
    \cb_4_0_io_eo[35] ,
    \cb_4_0_io_eo[34] ,
    \cb_4_0_io_eo[33] ,
    \cb_4_0_io_eo[32] ,
    \cb_4_0_io_eo[31] ,
    \cb_4_0_io_eo[30] ,
    \cb_4_0_io_eo[29] ,
    \cb_4_0_io_eo[28] ,
    \cb_4_0_io_eo[27] ,
    \cb_4_0_io_eo[26] ,
    \cb_4_0_io_eo[25] ,
    \cb_4_0_io_eo[24] ,
    \cb_4_0_io_eo[23] ,
    \cb_4_0_io_eo[22] ,
    \cb_4_0_io_eo[21] ,
    \cb_4_0_io_eo[20] ,
    \cb_4_0_io_eo[19] ,
    \cb_4_0_io_eo[18] ,
    \cb_4_0_io_eo[17] ,
    \cb_4_0_io_eo[16] ,
    \cb_4_0_io_eo[15] ,
    \cb_4_0_io_eo[14] ,
    \cb_4_0_io_eo[13] ,
    \cb_4_0_io_eo[12] ,
    \cb_4_0_io_eo[11] ,
    \cb_4_0_io_eo[10] ,
    \cb_4_0_io_eo[9] ,
    \cb_4_0_io_eo[8] ,
    \cb_4_0_io_eo[7] ,
    \cb_4_0_io_eo[6] ,
    \cb_4_0_io_eo[5] ,
    \cb_4_0_io_eo[4] ,
    \cb_4_0_io_eo[3] ,
    \cb_4_0_io_eo[2] ,
    \cb_4_0_io_eo[1] ,
    \cb_4_0_io_eo[0] }),
    .io_i_0_in1({_NC257,
    _NC258,
    _NC259,
    _NC260,
    _NC261,
    _NC262,
    _NC263,
    _NC264}),
    .io_i_1_in1({_NC265,
    _NC266,
    _NC267,
    _NC268,
    _NC269,
    _NC270,
    _NC271,
    _NC272}),
    .io_i_2_in1({_NC273,
    _NC274,
    _NC275,
    _NC276,
    _NC277,
    _NC278,
    _NC279,
    _NC280}),
    .io_i_3_in1({_NC281,
    _NC282,
    _NC283,
    _NC284,
    _NC285,
    _NC286,
    _NC287,
    _NC288}),
    .io_i_4_in1({_NC289,
    _NC290,
    _NC291,
    _NC292,
    _NC293,
    _NC294,
    _NC295,
    _NC296}),
    .io_i_5_in1({_NC297,
    _NC298,
    _NC299,
    _NC300,
    _NC301,
    _NC302,
    _NC303,
    _NC304}),
    .io_i_6_in1({_NC305,
    _NC306,
    _NC307,
    _NC308,
    _NC309,
    _NC310,
    _NC311,
    _NC312}),
    .io_i_7_in1({_NC313,
    _NC314,
    _NC315,
    _NC316,
    _NC317,
    _NC318,
    _NC319,
    _NC320}),
    .io_o_0_out({\cb_4_0_io_o_0_out[7] ,
    \cb_4_0_io_o_0_out[6] ,
    \cb_4_0_io_o_0_out[5] ,
    \cb_4_0_io_o_0_out[4] ,
    \cb_4_0_io_o_0_out[3] ,
    \cb_4_0_io_o_0_out[2] ,
    \cb_4_0_io_o_0_out[1] ,
    \cb_4_0_io_o_0_out[0] }),
    .io_o_1_out({\cb_4_0_io_o_1_out[7] ,
    \cb_4_0_io_o_1_out[6] ,
    \cb_4_0_io_o_1_out[5] ,
    \cb_4_0_io_o_1_out[4] ,
    \cb_4_0_io_o_1_out[3] ,
    \cb_4_0_io_o_1_out[2] ,
    \cb_4_0_io_o_1_out[1] ,
    \cb_4_0_io_o_1_out[0] }),
    .io_o_2_out({\cb_4_0_io_o_2_out[7] ,
    \cb_4_0_io_o_2_out[6] ,
    \cb_4_0_io_o_2_out[5] ,
    \cb_4_0_io_o_2_out[4] ,
    \cb_4_0_io_o_2_out[3] ,
    \cb_4_0_io_o_2_out[2] ,
    \cb_4_0_io_o_2_out[1] ,
    \cb_4_0_io_o_2_out[0] }),
    .io_o_3_out({\cb_4_0_io_o_3_out[7] ,
    \cb_4_0_io_o_3_out[6] ,
    \cb_4_0_io_o_3_out[5] ,
    \cb_4_0_io_o_3_out[4] ,
    \cb_4_0_io_o_3_out[3] ,
    \cb_4_0_io_o_3_out[2] ,
    \cb_4_0_io_o_3_out[1] ,
    \cb_4_0_io_o_3_out[0] }),
    .io_o_4_out({\cb_4_0_io_o_4_out[7] ,
    \cb_4_0_io_o_4_out[6] ,
    \cb_4_0_io_o_4_out[5] ,
    \cb_4_0_io_o_4_out[4] ,
    \cb_4_0_io_o_4_out[3] ,
    \cb_4_0_io_o_4_out[2] ,
    \cb_4_0_io_o_4_out[1] ,
    \cb_4_0_io_o_4_out[0] }),
    .io_o_5_out({\cb_4_0_io_o_5_out[7] ,
    \cb_4_0_io_o_5_out[6] ,
    \cb_4_0_io_o_5_out[5] ,
    \cb_4_0_io_o_5_out[4] ,
    \cb_4_0_io_o_5_out[3] ,
    \cb_4_0_io_o_5_out[2] ,
    \cb_4_0_io_o_5_out[1] ,
    \cb_4_0_io_o_5_out[0] }),
    .io_o_6_out({\cb_4_0_io_o_6_out[7] ,
    \cb_4_0_io_o_6_out[6] ,
    \cb_4_0_io_o_6_out[5] ,
    \cb_4_0_io_o_6_out[4] ,
    \cb_4_0_io_o_6_out[3] ,
    \cb_4_0_io_o_6_out[2] ,
    \cb_4_0_io_o_6_out[1] ,
    \cb_4_0_io_o_6_out[0] }),
    .io_o_7_out({\cb_4_0_io_o_7_out[7] ,
    \cb_4_0_io_o_7_out[6] ,
    \cb_4_0_io_o_7_out[5] ,
    \cb_4_0_io_o_7_out[4] ,
    \cb_4_0_io_o_7_out[3] ,
    \cb_4_0_io_o_7_out[2] ,
    \cb_4_0_io_o_7_out[1] ,
    \cb_4_0_io_o_7_out[0] }),
    .io_wo({\cb_4_0_io_wo[63] ,
    \cb_4_0_io_wo[62] ,
    \cb_4_0_io_wo[61] ,
    \cb_4_0_io_wo[60] ,
    \cb_4_0_io_wo[59] ,
    \cb_4_0_io_wo[58] ,
    \cb_4_0_io_wo[57] ,
    \cb_4_0_io_wo[56] ,
    \cb_4_0_io_wo[55] ,
    \cb_4_0_io_wo[54] ,
    \cb_4_0_io_wo[53] ,
    \cb_4_0_io_wo[52] ,
    \cb_4_0_io_wo[51] ,
    \cb_4_0_io_wo[50] ,
    \cb_4_0_io_wo[49] ,
    \cb_4_0_io_wo[48] ,
    \cb_4_0_io_wo[47] ,
    \cb_4_0_io_wo[46] ,
    \cb_4_0_io_wo[45] ,
    \cb_4_0_io_wo[44] ,
    \cb_4_0_io_wo[43] ,
    \cb_4_0_io_wo[42] ,
    \cb_4_0_io_wo[41] ,
    \cb_4_0_io_wo[40] ,
    \cb_4_0_io_wo[39] ,
    \cb_4_0_io_wo[38] ,
    \cb_4_0_io_wo[37] ,
    \cb_4_0_io_wo[36] ,
    \cb_4_0_io_wo[35] ,
    \cb_4_0_io_wo[34] ,
    \cb_4_0_io_wo[33] ,
    \cb_4_0_io_wo[32] ,
    \cb_4_0_io_wo[31] ,
    \cb_4_0_io_wo[30] ,
    \cb_4_0_io_wo[29] ,
    \cb_4_0_io_wo[28] ,
    \cb_4_0_io_wo[27] ,
    \cb_4_0_io_wo[26] ,
    \cb_4_0_io_wo[25] ,
    \cb_4_0_io_wo[24] ,
    \cb_4_0_io_wo[23] ,
    \cb_4_0_io_wo[22] ,
    \cb_4_0_io_wo[21] ,
    \cb_4_0_io_wo[20] ,
    \cb_4_0_io_wo[19] ,
    \cb_4_0_io_wo[18] ,
    \cb_4_0_io_wo[17] ,
    \cb_4_0_io_wo[16] ,
    \cb_4_0_io_wo[15] ,
    \cb_4_0_io_wo[14] ,
    \cb_4_0_io_wo[13] ,
    \cb_4_0_io_wo[12] ,
    \cb_4_0_io_wo[11] ,
    \cb_4_0_io_wo[10] ,
    \cb_4_0_io_wo[9] ,
    \cb_4_0_io_wo[8] ,
    \cb_4_0_io_wo[7] ,
    \cb_4_0_io_wo[6] ,
    \cb_4_0_io_wo[5] ,
    \cb_4_0_io_wo[4] ,
    \cb_4_0_io_wo[3] ,
    \cb_4_0_io_wo[2] ,
    \cb_4_0_io_wo[1] ,
    \cb_4_0_io_wo[0] }));
 cic_block cb_4_1 (.io_cs_i(cb_4_1_io_cs_i),
    .io_i_0_ci(cb_4_0_io_o_0_co),
    .io_i_1_ci(cb_4_0_io_o_1_co),
    .io_i_2_ci(cb_4_0_io_o_2_co),
    .io_i_3_ci(cb_4_0_io_o_3_co),
    .io_i_4_ci(cb_4_0_io_o_4_co),
    .io_i_5_ci(cb_4_0_io_o_5_co),
    .io_i_6_ci(cb_4_0_io_o_6_co),
    .io_i_7_ci(cb_4_0_io_o_7_co),
    .io_o_0_co(cb_4_1_io_o_0_co),
    .io_o_1_co(cb_4_1_io_o_1_co),
    .io_o_2_co(cb_4_1_io_o_2_co),
    .io_o_3_co(cb_4_1_io_o_3_co),
    .io_o_4_co(cb_4_1_io_o_4_co),
    .io_o_5_co(cb_4_1_io_o_5_co),
    .io_o_6_co(cb_4_1_io_o_6_co),
    .io_o_7_co(cb_4_1_io_o_7_co),
    .io_vci(cb_4_0_io_vco),
    .io_vco(cb_4_1_io_vco),
    .io_vi(cb_4_1_io_vi),
    .io_we_i(cb_4_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_4_0_io_adr_i[1] ,
    \cb_4_0_io_adr_i[0] }),
    .io_dat_i({\cb_4_0_io_dat_i[15] ,
    \cb_4_0_io_dat_i[14] ,
    \cb_4_0_io_dat_i[13] ,
    \cb_4_0_io_dat_i[12] ,
    \cb_4_0_io_dat_i[11] ,
    \cb_4_0_io_dat_i[10] ,
    \cb_4_0_io_dat_i[9] ,
    \cb_4_0_io_dat_i[8] ,
    \cb_4_0_io_dat_i[7] ,
    \cb_4_0_io_dat_i[6] ,
    \cb_4_0_io_dat_i[5] ,
    \cb_4_0_io_dat_i[4] ,
    \cb_4_0_io_dat_i[3] ,
    \cb_4_0_io_dat_i[2] ,
    \cb_4_0_io_dat_i[1] ,
    \cb_4_0_io_dat_i[0] }),
    .io_dat_o({\cb_4_1_io_dat_o[15] ,
    \cb_4_1_io_dat_o[14] ,
    \cb_4_1_io_dat_o[13] ,
    \cb_4_1_io_dat_o[12] ,
    \cb_4_1_io_dat_o[11] ,
    \cb_4_1_io_dat_o[10] ,
    \cb_4_1_io_dat_o[9] ,
    \cb_4_1_io_dat_o[8] ,
    \cb_4_1_io_dat_o[7] ,
    \cb_4_1_io_dat_o[6] ,
    \cb_4_1_io_dat_o[5] ,
    \cb_4_1_io_dat_o[4] ,
    \cb_4_1_io_dat_o[3] ,
    \cb_4_1_io_dat_o[2] ,
    \cb_4_1_io_dat_o[1] ,
    \cb_4_1_io_dat_o[0] }),
    .io_eo({\cb_4_1_io_eo[63] ,
    \cb_4_1_io_eo[62] ,
    \cb_4_1_io_eo[61] ,
    \cb_4_1_io_eo[60] ,
    \cb_4_1_io_eo[59] ,
    \cb_4_1_io_eo[58] ,
    \cb_4_1_io_eo[57] ,
    \cb_4_1_io_eo[56] ,
    \cb_4_1_io_eo[55] ,
    \cb_4_1_io_eo[54] ,
    \cb_4_1_io_eo[53] ,
    \cb_4_1_io_eo[52] ,
    \cb_4_1_io_eo[51] ,
    \cb_4_1_io_eo[50] ,
    \cb_4_1_io_eo[49] ,
    \cb_4_1_io_eo[48] ,
    \cb_4_1_io_eo[47] ,
    \cb_4_1_io_eo[46] ,
    \cb_4_1_io_eo[45] ,
    \cb_4_1_io_eo[44] ,
    \cb_4_1_io_eo[43] ,
    \cb_4_1_io_eo[42] ,
    \cb_4_1_io_eo[41] ,
    \cb_4_1_io_eo[40] ,
    \cb_4_1_io_eo[39] ,
    \cb_4_1_io_eo[38] ,
    \cb_4_1_io_eo[37] ,
    \cb_4_1_io_eo[36] ,
    \cb_4_1_io_eo[35] ,
    \cb_4_1_io_eo[34] ,
    \cb_4_1_io_eo[33] ,
    \cb_4_1_io_eo[32] ,
    \cb_4_1_io_eo[31] ,
    \cb_4_1_io_eo[30] ,
    \cb_4_1_io_eo[29] ,
    \cb_4_1_io_eo[28] ,
    \cb_4_1_io_eo[27] ,
    \cb_4_1_io_eo[26] ,
    \cb_4_1_io_eo[25] ,
    \cb_4_1_io_eo[24] ,
    \cb_4_1_io_eo[23] ,
    \cb_4_1_io_eo[22] ,
    \cb_4_1_io_eo[21] ,
    \cb_4_1_io_eo[20] ,
    \cb_4_1_io_eo[19] ,
    \cb_4_1_io_eo[18] ,
    \cb_4_1_io_eo[17] ,
    \cb_4_1_io_eo[16] ,
    \cb_4_1_io_eo[15] ,
    \cb_4_1_io_eo[14] ,
    \cb_4_1_io_eo[13] ,
    \cb_4_1_io_eo[12] ,
    \cb_4_1_io_eo[11] ,
    \cb_4_1_io_eo[10] ,
    \cb_4_1_io_eo[9] ,
    \cb_4_1_io_eo[8] ,
    \cb_4_1_io_eo[7] ,
    \cb_4_1_io_eo[6] ,
    \cb_4_1_io_eo[5] ,
    \cb_4_1_io_eo[4] ,
    \cb_4_1_io_eo[3] ,
    \cb_4_1_io_eo[2] ,
    \cb_4_1_io_eo[1] ,
    \cb_4_1_io_eo[0] }),
    .io_i_0_in1({\cb_4_0_io_o_0_out[7] ,
    \cb_4_0_io_o_0_out[6] ,
    \cb_4_0_io_o_0_out[5] ,
    \cb_4_0_io_o_0_out[4] ,
    \cb_4_0_io_o_0_out[3] ,
    \cb_4_0_io_o_0_out[2] ,
    \cb_4_0_io_o_0_out[1] ,
    \cb_4_0_io_o_0_out[0] }),
    .io_i_1_in1({\cb_4_0_io_o_1_out[7] ,
    \cb_4_0_io_o_1_out[6] ,
    \cb_4_0_io_o_1_out[5] ,
    \cb_4_0_io_o_1_out[4] ,
    \cb_4_0_io_o_1_out[3] ,
    \cb_4_0_io_o_1_out[2] ,
    \cb_4_0_io_o_1_out[1] ,
    \cb_4_0_io_o_1_out[0] }),
    .io_i_2_in1({\cb_4_0_io_o_2_out[7] ,
    \cb_4_0_io_o_2_out[6] ,
    \cb_4_0_io_o_2_out[5] ,
    \cb_4_0_io_o_2_out[4] ,
    \cb_4_0_io_o_2_out[3] ,
    \cb_4_0_io_o_2_out[2] ,
    \cb_4_0_io_o_2_out[1] ,
    \cb_4_0_io_o_2_out[0] }),
    .io_i_3_in1({\cb_4_0_io_o_3_out[7] ,
    \cb_4_0_io_o_3_out[6] ,
    \cb_4_0_io_o_3_out[5] ,
    \cb_4_0_io_o_3_out[4] ,
    \cb_4_0_io_o_3_out[3] ,
    \cb_4_0_io_o_3_out[2] ,
    \cb_4_0_io_o_3_out[1] ,
    \cb_4_0_io_o_3_out[0] }),
    .io_i_4_in1({\cb_4_0_io_o_4_out[7] ,
    \cb_4_0_io_o_4_out[6] ,
    \cb_4_0_io_o_4_out[5] ,
    \cb_4_0_io_o_4_out[4] ,
    \cb_4_0_io_o_4_out[3] ,
    \cb_4_0_io_o_4_out[2] ,
    \cb_4_0_io_o_4_out[1] ,
    \cb_4_0_io_o_4_out[0] }),
    .io_i_5_in1({\cb_4_0_io_o_5_out[7] ,
    \cb_4_0_io_o_5_out[6] ,
    \cb_4_0_io_o_5_out[5] ,
    \cb_4_0_io_o_5_out[4] ,
    \cb_4_0_io_o_5_out[3] ,
    \cb_4_0_io_o_5_out[2] ,
    \cb_4_0_io_o_5_out[1] ,
    \cb_4_0_io_o_5_out[0] }),
    .io_i_6_in1({\cb_4_0_io_o_6_out[7] ,
    \cb_4_0_io_o_6_out[6] ,
    \cb_4_0_io_o_6_out[5] ,
    \cb_4_0_io_o_6_out[4] ,
    \cb_4_0_io_o_6_out[3] ,
    \cb_4_0_io_o_6_out[2] ,
    \cb_4_0_io_o_6_out[1] ,
    \cb_4_0_io_o_6_out[0] }),
    .io_i_7_in1({\cb_4_0_io_o_7_out[7] ,
    \cb_4_0_io_o_7_out[6] ,
    \cb_4_0_io_o_7_out[5] ,
    \cb_4_0_io_o_7_out[4] ,
    \cb_4_0_io_o_7_out[3] ,
    \cb_4_0_io_o_7_out[2] ,
    \cb_4_0_io_o_7_out[1] ,
    \cb_4_0_io_o_7_out[0] }),
    .io_o_0_out({\cb_4_1_io_o_0_out[7] ,
    \cb_4_1_io_o_0_out[6] ,
    \cb_4_1_io_o_0_out[5] ,
    \cb_4_1_io_o_0_out[4] ,
    \cb_4_1_io_o_0_out[3] ,
    \cb_4_1_io_o_0_out[2] ,
    \cb_4_1_io_o_0_out[1] ,
    \cb_4_1_io_o_0_out[0] }),
    .io_o_1_out({\cb_4_1_io_o_1_out[7] ,
    \cb_4_1_io_o_1_out[6] ,
    \cb_4_1_io_o_1_out[5] ,
    \cb_4_1_io_o_1_out[4] ,
    \cb_4_1_io_o_1_out[3] ,
    \cb_4_1_io_o_1_out[2] ,
    \cb_4_1_io_o_1_out[1] ,
    \cb_4_1_io_o_1_out[0] }),
    .io_o_2_out({\cb_4_1_io_o_2_out[7] ,
    \cb_4_1_io_o_2_out[6] ,
    \cb_4_1_io_o_2_out[5] ,
    \cb_4_1_io_o_2_out[4] ,
    \cb_4_1_io_o_2_out[3] ,
    \cb_4_1_io_o_2_out[2] ,
    \cb_4_1_io_o_2_out[1] ,
    \cb_4_1_io_o_2_out[0] }),
    .io_o_3_out({\cb_4_1_io_o_3_out[7] ,
    \cb_4_1_io_o_3_out[6] ,
    \cb_4_1_io_o_3_out[5] ,
    \cb_4_1_io_o_3_out[4] ,
    \cb_4_1_io_o_3_out[3] ,
    \cb_4_1_io_o_3_out[2] ,
    \cb_4_1_io_o_3_out[1] ,
    \cb_4_1_io_o_3_out[0] }),
    .io_o_4_out({\cb_4_1_io_o_4_out[7] ,
    \cb_4_1_io_o_4_out[6] ,
    \cb_4_1_io_o_4_out[5] ,
    \cb_4_1_io_o_4_out[4] ,
    \cb_4_1_io_o_4_out[3] ,
    \cb_4_1_io_o_4_out[2] ,
    \cb_4_1_io_o_4_out[1] ,
    \cb_4_1_io_o_4_out[0] }),
    .io_o_5_out({\cb_4_1_io_o_5_out[7] ,
    \cb_4_1_io_o_5_out[6] ,
    \cb_4_1_io_o_5_out[5] ,
    \cb_4_1_io_o_5_out[4] ,
    \cb_4_1_io_o_5_out[3] ,
    \cb_4_1_io_o_5_out[2] ,
    \cb_4_1_io_o_5_out[1] ,
    \cb_4_1_io_o_5_out[0] }),
    .io_o_6_out({\cb_4_1_io_o_6_out[7] ,
    \cb_4_1_io_o_6_out[6] ,
    \cb_4_1_io_o_6_out[5] ,
    \cb_4_1_io_o_6_out[4] ,
    \cb_4_1_io_o_6_out[3] ,
    \cb_4_1_io_o_6_out[2] ,
    \cb_4_1_io_o_6_out[1] ,
    \cb_4_1_io_o_6_out[0] }),
    .io_o_7_out({\cb_4_1_io_o_7_out[7] ,
    \cb_4_1_io_o_7_out[6] ,
    \cb_4_1_io_o_7_out[5] ,
    \cb_4_1_io_o_7_out[4] ,
    \cb_4_1_io_o_7_out[3] ,
    \cb_4_1_io_o_7_out[2] ,
    \cb_4_1_io_o_7_out[1] ,
    \cb_4_1_io_o_7_out[0] }),
    .io_wo({\cb_4_0_io_eo[63] ,
    \cb_4_0_io_eo[62] ,
    \cb_4_0_io_eo[61] ,
    \cb_4_0_io_eo[60] ,
    \cb_4_0_io_eo[59] ,
    \cb_4_0_io_eo[58] ,
    \cb_4_0_io_eo[57] ,
    \cb_4_0_io_eo[56] ,
    \cb_4_0_io_eo[55] ,
    \cb_4_0_io_eo[54] ,
    \cb_4_0_io_eo[53] ,
    \cb_4_0_io_eo[52] ,
    \cb_4_0_io_eo[51] ,
    \cb_4_0_io_eo[50] ,
    \cb_4_0_io_eo[49] ,
    \cb_4_0_io_eo[48] ,
    \cb_4_0_io_eo[47] ,
    \cb_4_0_io_eo[46] ,
    \cb_4_0_io_eo[45] ,
    \cb_4_0_io_eo[44] ,
    \cb_4_0_io_eo[43] ,
    \cb_4_0_io_eo[42] ,
    \cb_4_0_io_eo[41] ,
    \cb_4_0_io_eo[40] ,
    \cb_4_0_io_eo[39] ,
    \cb_4_0_io_eo[38] ,
    \cb_4_0_io_eo[37] ,
    \cb_4_0_io_eo[36] ,
    \cb_4_0_io_eo[35] ,
    \cb_4_0_io_eo[34] ,
    \cb_4_0_io_eo[33] ,
    \cb_4_0_io_eo[32] ,
    \cb_4_0_io_eo[31] ,
    \cb_4_0_io_eo[30] ,
    \cb_4_0_io_eo[29] ,
    \cb_4_0_io_eo[28] ,
    \cb_4_0_io_eo[27] ,
    \cb_4_0_io_eo[26] ,
    \cb_4_0_io_eo[25] ,
    \cb_4_0_io_eo[24] ,
    \cb_4_0_io_eo[23] ,
    \cb_4_0_io_eo[22] ,
    \cb_4_0_io_eo[21] ,
    \cb_4_0_io_eo[20] ,
    \cb_4_0_io_eo[19] ,
    \cb_4_0_io_eo[18] ,
    \cb_4_0_io_eo[17] ,
    \cb_4_0_io_eo[16] ,
    \cb_4_0_io_eo[15] ,
    \cb_4_0_io_eo[14] ,
    \cb_4_0_io_eo[13] ,
    \cb_4_0_io_eo[12] ,
    \cb_4_0_io_eo[11] ,
    \cb_4_0_io_eo[10] ,
    \cb_4_0_io_eo[9] ,
    \cb_4_0_io_eo[8] ,
    \cb_4_0_io_eo[7] ,
    \cb_4_0_io_eo[6] ,
    \cb_4_0_io_eo[5] ,
    \cb_4_0_io_eo[4] ,
    \cb_4_0_io_eo[3] ,
    \cb_4_0_io_eo[2] ,
    \cb_4_0_io_eo[1] ,
    \cb_4_0_io_eo[0] }));
 cic_block cb_4_10 (.io_cs_i(cb_4_10_io_cs_i),
    .io_i_0_ci(cb_4_10_io_i_0_ci),
    .io_i_1_ci(cb_4_10_io_i_1_ci),
    .io_i_2_ci(cb_4_10_io_i_2_ci),
    .io_i_3_ci(cb_4_10_io_i_3_ci),
    .io_i_4_ci(cb_4_10_io_i_4_ci),
    .io_i_5_ci(cb_4_10_io_i_5_ci),
    .io_i_6_ci(cb_4_10_io_i_6_ci),
    .io_i_7_ci(cb_4_10_io_i_7_ci),
    .io_o_0_co(cb_4_10_io_o_0_co),
    .io_o_1_co(cb_4_10_io_o_1_co),
    .io_o_2_co(cb_4_10_io_o_2_co),
    .io_o_3_co(cb_4_10_io_o_3_co),
    .io_o_4_co(cb_4_10_io_o_4_co),
    .io_o_5_co(cb_4_10_io_o_5_co),
    .io_o_6_co(cb_4_10_io_o_6_co),
    .io_o_7_co(cb_4_10_io_o_7_co),
    .io_vci(cb_4_10_io_vci),
    .io_vco(cb_4_10_io_vco),
    .io_vi(cb_4_10_io_vi),
    .io_we_i(cb_4_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_4_0_io_adr_i[1] ,
    \cb_4_0_io_adr_i[0] }),
    .io_dat_i({\cb_4_0_io_dat_i[15] ,
    \cb_4_0_io_dat_i[14] ,
    \cb_4_0_io_dat_i[13] ,
    \cb_4_0_io_dat_i[12] ,
    \cb_4_0_io_dat_i[11] ,
    \cb_4_0_io_dat_i[10] ,
    \cb_4_0_io_dat_i[9] ,
    \cb_4_0_io_dat_i[8] ,
    \cb_4_0_io_dat_i[7] ,
    \cb_4_0_io_dat_i[6] ,
    \cb_4_0_io_dat_i[5] ,
    \cb_4_0_io_dat_i[4] ,
    \cb_4_0_io_dat_i[3] ,
    \cb_4_0_io_dat_i[2] ,
    \cb_4_0_io_dat_i[1] ,
    \cb_4_0_io_dat_i[0] }),
    .io_dat_o({\cb_4_10_io_dat_o[15] ,
    \cb_4_10_io_dat_o[14] ,
    \cb_4_10_io_dat_o[13] ,
    \cb_4_10_io_dat_o[12] ,
    \cb_4_10_io_dat_o[11] ,
    \cb_4_10_io_dat_o[10] ,
    \cb_4_10_io_dat_o[9] ,
    \cb_4_10_io_dat_o[8] ,
    \cb_4_10_io_dat_o[7] ,
    \cb_4_10_io_dat_o[6] ,
    \cb_4_10_io_dat_o[5] ,
    \cb_4_10_io_dat_o[4] ,
    \cb_4_10_io_dat_o[3] ,
    \cb_4_10_io_dat_o[2] ,
    \cb_4_10_io_dat_o[1] ,
    \cb_4_10_io_dat_o[0] }),
    .io_eo({\_T_104[31] ,
    \_T_104[30] ,
    \_T_104[29] ,
    \_T_104[28] ,
    \_T_104[27] ,
    \_T_104[26] ,
    \_T_104[25] ,
    \_T_104[24] ,
    \_T_104[23] ,
    \_T_104[22] ,
    \_T_104[21] ,
    \_T_104[20] ,
    \_T_104[19] ,
    \_T_104[18] ,
    \_T_104[17] ,
    \_T_104[16] ,
    \_T_104[15] ,
    \_T_104[14] ,
    \_T_104[13] ,
    \_T_104[12] ,
    \_T_104[11] ,
    \_T_104[10] ,
    \_T_104[9] ,
    \_T_104[8] ,
    \_T_104[7] ,
    \_T_104[6] ,
    \_T_104[5] ,
    \_T_104[4] ,
    \_T_104[3] ,
    \_T_104[2] ,
    \_T_104[1] ,
    \_T_104[0] ,
    \_T_101[31] ,
    \_T_101[30] ,
    \_T_101[29] ,
    \_T_101[28] ,
    \_T_101[27] ,
    \_T_101[26] ,
    \_T_101[25] ,
    \_T_101[24] ,
    \_T_101[23] ,
    \_T_101[22] ,
    \_T_101[21] ,
    \_T_101[20] ,
    \_T_101[19] ,
    \_T_101[18] ,
    \_T_101[17] ,
    \_T_101[16] ,
    \_T_101[15] ,
    \_T_101[14] ,
    \_T_101[13] ,
    \_T_101[12] ,
    \_T_101[11] ,
    \_T_101[10] ,
    \_T_101[9] ,
    \_T_101[8] ,
    \_T_101[7] ,
    \_T_101[6] ,
    \_T_101[5] ,
    \_T_101[4] ,
    \_T_101[3] ,
    \_T_101[2] ,
    \_T_101[1] ,
    \_T_101[0] }),
    .io_i_0_in1({\cb_4_10_io_i_0_in1[7] ,
    \cb_4_10_io_i_0_in1[6] ,
    \cb_4_10_io_i_0_in1[5] ,
    \cb_4_10_io_i_0_in1[4] ,
    \cb_4_10_io_i_0_in1[3] ,
    \cb_4_10_io_i_0_in1[2] ,
    \cb_4_10_io_i_0_in1[1] ,
    \cb_4_10_io_i_0_in1[0] }),
    .io_i_1_in1({\cb_4_10_io_i_1_in1[7] ,
    \cb_4_10_io_i_1_in1[6] ,
    \cb_4_10_io_i_1_in1[5] ,
    \cb_4_10_io_i_1_in1[4] ,
    \cb_4_10_io_i_1_in1[3] ,
    \cb_4_10_io_i_1_in1[2] ,
    \cb_4_10_io_i_1_in1[1] ,
    \cb_4_10_io_i_1_in1[0] }),
    .io_i_2_in1({\cb_4_10_io_i_2_in1[7] ,
    \cb_4_10_io_i_2_in1[6] ,
    \cb_4_10_io_i_2_in1[5] ,
    \cb_4_10_io_i_2_in1[4] ,
    \cb_4_10_io_i_2_in1[3] ,
    \cb_4_10_io_i_2_in1[2] ,
    \cb_4_10_io_i_2_in1[1] ,
    \cb_4_10_io_i_2_in1[0] }),
    .io_i_3_in1({\cb_4_10_io_i_3_in1[7] ,
    \cb_4_10_io_i_3_in1[6] ,
    \cb_4_10_io_i_3_in1[5] ,
    \cb_4_10_io_i_3_in1[4] ,
    \cb_4_10_io_i_3_in1[3] ,
    \cb_4_10_io_i_3_in1[2] ,
    \cb_4_10_io_i_3_in1[1] ,
    \cb_4_10_io_i_3_in1[0] }),
    .io_i_4_in1({\cb_4_10_io_i_4_in1[7] ,
    \cb_4_10_io_i_4_in1[6] ,
    \cb_4_10_io_i_4_in1[5] ,
    \cb_4_10_io_i_4_in1[4] ,
    \cb_4_10_io_i_4_in1[3] ,
    \cb_4_10_io_i_4_in1[2] ,
    \cb_4_10_io_i_4_in1[1] ,
    \cb_4_10_io_i_4_in1[0] }),
    .io_i_5_in1({\cb_4_10_io_i_5_in1[7] ,
    \cb_4_10_io_i_5_in1[6] ,
    \cb_4_10_io_i_5_in1[5] ,
    \cb_4_10_io_i_5_in1[4] ,
    \cb_4_10_io_i_5_in1[3] ,
    \cb_4_10_io_i_5_in1[2] ,
    \cb_4_10_io_i_5_in1[1] ,
    \cb_4_10_io_i_5_in1[0] }),
    .io_i_6_in1({\cb_4_10_io_i_6_in1[7] ,
    \cb_4_10_io_i_6_in1[6] ,
    \cb_4_10_io_i_6_in1[5] ,
    \cb_4_10_io_i_6_in1[4] ,
    \cb_4_10_io_i_6_in1[3] ,
    \cb_4_10_io_i_6_in1[2] ,
    \cb_4_10_io_i_6_in1[1] ,
    \cb_4_10_io_i_6_in1[0] }),
    .io_i_7_in1({\cb_4_10_io_i_7_in1[7] ,
    \cb_4_10_io_i_7_in1[6] ,
    \cb_4_10_io_i_7_in1[5] ,
    \cb_4_10_io_i_7_in1[4] ,
    \cb_4_10_io_i_7_in1[3] ,
    \cb_4_10_io_i_7_in1[2] ,
    \cb_4_10_io_i_7_in1[1] ,
    \cb_4_10_io_i_7_in1[0] }),
    .io_o_0_out({\_T_101[7] ,
    \_T_101[6] ,
    \_T_101[5] ,
    \_T_101[4] ,
    \_T_101[3] ,
    \_T_101[2] ,
    \_T_101[1] ,
    \_T_101[0] }),
    .io_o_1_out({\_T_101[15] ,
    \_T_101[14] ,
    \_T_101[13] ,
    \_T_101[12] ,
    \_T_101[11] ,
    \_T_101[10] ,
    \_T_101[9] ,
    \_T_101[8] }),
    .io_o_2_out({\_T_101[23] ,
    \_T_101[22] ,
    \_T_101[21] ,
    \_T_101[20] ,
    \_T_101[19] ,
    \_T_101[18] ,
    \_T_101[17] ,
    \_T_101[16] }),
    .io_o_3_out({\_T_101[31] ,
    \_T_101[30] ,
    \_T_101[29] ,
    \_T_101[28] ,
    \_T_101[27] ,
    \_T_101[26] ,
    \_T_101[25] ,
    \_T_101[24] }),
    .io_o_4_out({\_T_104[7] ,
    \_T_104[6] ,
    \_T_104[5] ,
    \_T_104[4] ,
    \_T_104[3] ,
    \_T_104[2] ,
    \_T_104[1] ,
    \_T_104[0] }),
    .io_o_5_out({\_T_104[15] ,
    \_T_104[14] ,
    \_T_104[13] ,
    \_T_104[12] ,
    \_T_104[11] ,
    \_T_104[10] ,
    \_T_104[9] ,
    \_T_104[8] }),
    .io_o_6_out({\_T_104[23] ,
    \_T_104[22] ,
    \_T_104[21] ,
    \_T_104[20] ,
    \_T_104[19] ,
    \_T_104[18] ,
    \_T_104[17] ,
    \_T_104[16] }),
    .io_o_7_out({\_T_104[31] ,
    \_T_104[30] ,
    \_T_104[29] ,
    \_T_104[28] ,
    \_T_104[27] ,
    \_T_104[26] ,
    \_T_104[25] ,
    \_T_104[24] }),
    .io_wo({\cb_4_10_io_wo[63] ,
    \cb_4_10_io_wo[62] ,
    \cb_4_10_io_wo[61] ,
    \cb_4_10_io_wo[60] ,
    \cb_4_10_io_wo[59] ,
    \cb_4_10_io_wo[58] ,
    \cb_4_10_io_wo[57] ,
    \cb_4_10_io_wo[56] ,
    \cb_4_10_io_wo[55] ,
    \cb_4_10_io_wo[54] ,
    \cb_4_10_io_wo[53] ,
    \cb_4_10_io_wo[52] ,
    \cb_4_10_io_wo[51] ,
    \cb_4_10_io_wo[50] ,
    \cb_4_10_io_wo[49] ,
    \cb_4_10_io_wo[48] ,
    \cb_4_10_io_wo[47] ,
    \cb_4_10_io_wo[46] ,
    \cb_4_10_io_wo[45] ,
    \cb_4_10_io_wo[44] ,
    \cb_4_10_io_wo[43] ,
    \cb_4_10_io_wo[42] ,
    \cb_4_10_io_wo[41] ,
    \cb_4_10_io_wo[40] ,
    \cb_4_10_io_wo[39] ,
    \cb_4_10_io_wo[38] ,
    \cb_4_10_io_wo[37] ,
    \cb_4_10_io_wo[36] ,
    \cb_4_10_io_wo[35] ,
    \cb_4_10_io_wo[34] ,
    \cb_4_10_io_wo[33] ,
    \cb_4_10_io_wo[32] ,
    \cb_4_10_io_wo[31] ,
    \cb_4_10_io_wo[30] ,
    \cb_4_10_io_wo[29] ,
    \cb_4_10_io_wo[28] ,
    \cb_4_10_io_wo[27] ,
    \cb_4_10_io_wo[26] ,
    \cb_4_10_io_wo[25] ,
    \cb_4_10_io_wo[24] ,
    \cb_4_10_io_wo[23] ,
    \cb_4_10_io_wo[22] ,
    \cb_4_10_io_wo[21] ,
    \cb_4_10_io_wo[20] ,
    \cb_4_10_io_wo[19] ,
    \cb_4_10_io_wo[18] ,
    \cb_4_10_io_wo[17] ,
    \cb_4_10_io_wo[16] ,
    \cb_4_10_io_wo[15] ,
    \cb_4_10_io_wo[14] ,
    \cb_4_10_io_wo[13] ,
    \cb_4_10_io_wo[12] ,
    \cb_4_10_io_wo[11] ,
    \cb_4_10_io_wo[10] ,
    \cb_4_10_io_wo[9] ,
    \cb_4_10_io_wo[8] ,
    \cb_4_10_io_wo[7] ,
    \cb_4_10_io_wo[6] ,
    \cb_4_10_io_wo[5] ,
    \cb_4_10_io_wo[4] ,
    \cb_4_10_io_wo[3] ,
    \cb_4_10_io_wo[2] ,
    \cb_4_10_io_wo[1] ,
    \cb_4_10_io_wo[0] }));
 cic_block cb_4_2 (.io_cs_i(cb_4_2_io_cs_i),
    .io_i_0_ci(cb_4_1_io_o_0_co),
    .io_i_1_ci(cb_4_1_io_o_1_co),
    .io_i_2_ci(cb_4_1_io_o_2_co),
    .io_i_3_ci(cb_4_1_io_o_3_co),
    .io_i_4_ci(cb_4_1_io_o_4_co),
    .io_i_5_ci(cb_4_1_io_o_5_co),
    .io_i_6_ci(cb_4_1_io_o_6_co),
    .io_i_7_ci(cb_4_1_io_o_7_co),
    .io_o_0_co(cb_4_2_io_o_0_co),
    .io_o_1_co(cb_4_2_io_o_1_co),
    .io_o_2_co(cb_4_2_io_o_2_co),
    .io_o_3_co(cb_4_2_io_o_3_co),
    .io_o_4_co(cb_4_2_io_o_4_co),
    .io_o_5_co(cb_4_2_io_o_5_co),
    .io_o_6_co(cb_4_2_io_o_6_co),
    .io_o_7_co(cb_4_2_io_o_7_co),
    .io_vci(cb_4_1_io_vco),
    .io_vco(cb_4_2_io_vco),
    .io_vi(cb_4_2_io_vi),
    .io_we_i(cb_4_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_4_0_io_adr_i[1] ,
    \cb_4_0_io_adr_i[0] }),
    .io_dat_i({\cb_4_0_io_dat_i[15] ,
    \cb_4_0_io_dat_i[14] ,
    \cb_4_0_io_dat_i[13] ,
    \cb_4_0_io_dat_i[12] ,
    \cb_4_0_io_dat_i[11] ,
    \cb_4_0_io_dat_i[10] ,
    \cb_4_0_io_dat_i[9] ,
    \cb_4_0_io_dat_i[8] ,
    \cb_4_0_io_dat_i[7] ,
    \cb_4_0_io_dat_i[6] ,
    \cb_4_0_io_dat_i[5] ,
    \cb_4_0_io_dat_i[4] ,
    \cb_4_0_io_dat_i[3] ,
    \cb_4_0_io_dat_i[2] ,
    \cb_4_0_io_dat_i[1] ,
    \cb_4_0_io_dat_i[0] }),
    .io_dat_o({\cb_4_2_io_dat_o[15] ,
    \cb_4_2_io_dat_o[14] ,
    \cb_4_2_io_dat_o[13] ,
    \cb_4_2_io_dat_o[12] ,
    \cb_4_2_io_dat_o[11] ,
    \cb_4_2_io_dat_o[10] ,
    \cb_4_2_io_dat_o[9] ,
    \cb_4_2_io_dat_o[8] ,
    \cb_4_2_io_dat_o[7] ,
    \cb_4_2_io_dat_o[6] ,
    \cb_4_2_io_dat_o[5] ,
    \cb_4_2_io_dat_o[4] ,
    \cb_4_2_io_dat_o[3] ,
    \cb_4_2_io_dat_o[2] ,
    \cb_4_2_io_dat_o[1] ,
    \cb_4_2_io_dat_o[0] }),
    .io_eo({\cb_4_2_io_eo[63] ,
    \cb_4_2_io_eo[62] ,
    \cb_4_2_io_eo[61] ,
    \cb_4_2_io_eo[60] ,
    \cb_4_2_io_eo[59] ,
    \cb_4_2_io_eo[58] ,
    \cb_4_2_io_eo[57] ,
    \cb_4_2_io_eo[56] ,
    \cb_4_2_io_eo[55] ,
    \cb_4_2_io_eo[54] ,
    \cb_4_2_io_eo[53] ,
    \cb_4_2_io_eo[52] ,
    \cb_4_2_io_eo[51] ,
    \cb_4_2_io_eo[50] ,
    \cb_4_2_io_eo[49] ,
    \cb_4_2_io_eo[48] ,
    \cb_4_2_io_eo[47] ,
    \cb_4_2_io_eo[46] ,
    \cb_4_2_io_eo[45] ,
    \cb_4_2_io_eo[44] ,
    \cb_4_2_io_eo[43] ,
    \cb_4_2_io_eo[42] ,
    \cb_4_2_io_eo[41] ,
    \cb_4_2_io_eo[40] ,
    \cb_4_2_io_eo[39] ,
    \cb_4_2_io_eo[38] ,
    \cb_4_2_io_eo[37] ,
    \cb_4_2_io_eo[36] ,
    \cb_4_2_io_eo[35] ,
    \cb_4_2_io_eo[34] ,
    \cb_4_2_io_eo[33] ,
    \cb_4_2_io_eo[32] ,
    \cb_4_2_io_eo[31] ,
    \cb_4_2_io_eo[30] ,
    \cb_4_2_io_eo[29] ,
    \cb_4_2_io_eo[28] ,
    \cb_4_2_io_eo[27] ,
    \cb_4_2_io_eo[26] ,
    \cb_4_2_io_eo[25] ,
    \cb_4_2_io_eo[24] ,
    \cb_4_2_io_eo[23] ,
    \cb_4_2_io_eo[22] ,
    \cb_4_2_io_eo[21] ,
    \cb_4_2_io_eo[20] ,
    \cb_4_2_io_eo[19] ,
    \cb_4_2_io_eo[18] ,
    \cb_4_2_io_eo[17] ,
    \cb_4_2_io_eo[16] ,
    \cb_4_2_io_eo[15] ,
    \cb_4_2_io_eo[14] ,
    \cb_4_2_io_eo[13] ,
    \cb_4_2_io_eo[12] ,
    \cb_4_2_io_eo[11] ,
    \cb_4_2_io_eo[10] ,
    \cb_4_2_io_eo[9] ,
    \cb_4_2_io_eo[8] ,
    \cb_4_2_io_eo[7] ,
    \cb_4_2_io_eo[6] ,
    \cb_4_2_io_eo[5] ,
    \cb_4_2_io_eo[4] ,
    \cb_4_2_io_eo[3] ,
    \cb_4_2_io_eo[2] ,
    \cb_4_2_io_eo[1] ,
    \cb_4_2_io_eo[0] }),
    .io_i_0_in1({\cb_4_1_io_o_0_out[7] ,
    \cb_4_1_io_o_0_out[6] ,
    \cb_4_1_io_o_0_out[5] ,
    \cb_4_1_io_o_0_out[4] ,
    \cb_4_1_io_o_0_out[3] ,
    \cb_4_1_io_o_0_out[2] ,
    \cb_4_1_io_o_0_out[1] ,
    \cb_4_1_io_o_0_out[0] }),
    .io_i_1_in1({\cb_4_1_io_o_1_out[7] ,
    \cb_4_1_io_o_1_out[6] ,
    \cb_4_1_io_o_1_out[5] ,
    \cb_4_1_io_o_1_out[4] ,
    \cb_4_1_io_o_1_out[3] ,
    \cb_4_1_io_o_1_out[2] ,
    \cb_4_1_io_o_1_out[1] ,
    \cb_4_1_io_o_1_out[0] }),
    .io_i_2_in1({\cb_4_1_io_o_2_out[7] ,
    \cb_4_1_io_o_2_out[6] ,
    \cb_4_1_io_o_2_out[5] ,
    \cb_4_1_io_o_2_out[4] ,
    \cb_4_1_io_o_2_out[3] ,
    \cb_4_1_io_o_2_out[2] ,
    \cb_4_1_io_o_2_out[1] ,
    \cb_4_1_io_o_2_out[0] }),
    .io_i_3_in1({\cb_4_1_io_o_3_out[7] ,
    \cb_4_1_io_o_3_out[6] ,
    \cb_4_1_io_o_3_out[5] ,
    \cb_4_1_io_o_3_out[4] ,
    \cb_4_1_io_o_3_out[3] ,
    \cb_4_1_io_o_3_out[2] ,
    \cb_4_1_io_o_3_out[1] ,
    \cb_4_1_io_o_3_out[0] }),
    .io_i_4_in1({\cb_4_1_io_o_4_out[7] ,
    \cb_4_1_io_o_4_out[6] ,
    \cb_4_1_io_o_4_out[5] ,
    \cb_4_1_io_o_4_out[4] ,
    \cb_4_1_io_o_4_out[3] ,
    \cb_4_1_io_o_4_out[2] ,
    \cb_4_1_io_o_4_out[1] ,
    \cb_4_1_io_o_4_out[0] }),
    .io_i_5_in1({\cb_4_1_io_o_5_out[7] ,
    \cb_4_1_io_o_5_out[6] ,
    \cb_4_1_io_o_5_out[5] ,
    \cb_4_1_io_o_5_out[4] ,
    \cb_4_1_io_o_5_out[3] ,
    \cb_4_1_io_o_5_out[2] ,
    \cb_4_1_io_o_5_out[1] ,
    \cb_4_1_io_o_5_out[0] }),
    .io_i_6_in1({\cb_4_1_io_o_6_out[7] ,
    \cb_4_1_io_o_6_out[6] ,
    \cb_4_1_io_o_6_out[5] ,
    \cb_4_1_io_o_6_out[4] ,
    \cb_4_1_io_o_6_out[3] ,
    \cb_4_1_io_o_6_out[2] ,
    \cb_4_1_io_o_6_out[1] ,
    \cb_4_1_io_o_6_out[0] }),
    .io_i_7_in1({\cb_4_1_io_o_7_out[7] ,
    \cb_4_1_io_o_7_out[6] ,
    \cb_4_1_io_o_7_out[5] ,
    \cb_4_1_io_o_7_out[4] ,
    \cb_4_1_io_o_7_out[3] ,
    \cb_4_1_io_o_7_out[2] ,
    \cb_4_1_io_o_7_out[1] ,
    \cb_4_1_io_o_7_out[0] }),
    .io_o_0_out({\cb_4_2_io_o_0_out[7] ,
    \cb_4_2_io_o_0_out[6] ,
    \cb_4_2_io_o_0_out[5] ,
    \cb_4_2_io_o_0_out[4] ,
    \cb_4_2_io_o_0_out[3] ,
    \cb_4_2_io_o_0_out[2] ,
    \cb_4_2_io_o_0_out[1] ,
    \cb_4_2_io_o_0_out[0] }),
    .io_o_1_out({\cb_4_2_io_o_1_out[7] ,
    \cb_4_2_io_o_1_out[6] ,
    \cb_4_2_io_o_1_out[5] ,
    \cb_4_2_io_o_1_out[4] ,
    \cb_4_2_io_o_1_out[3] ,
    \cb_4_2_io_o_1_out[2] ,
    \cb_4_2_io_o_1_out[1] ,
    \cb_4_2_io_o_1_out[0] }),
    .io_o_2_out({\cb_4_2_io_o_2_out[7] ,
    \cb_4_2_io_o_2_out[6] ,
    \cb_4_2_io_o_2_out[5] ,
    \cb_4_2_io_o_2_out[4] ,
    \cb_4_2_io_o_2_out[3] ,
    \cb_4_2_io_o_2_out[2] ,
    \cb_4_2_io_o_2_out[1] ,
    \cb_4_2_io_o_2_out[0] }),
    .io_o_3_out({\cb_4_2_io_o_3_out[7] ,
    \cb_4_2_io_o_3_out[6] ,
    \cb_4_2_io_o_3_out[5] ,
    \cb_4_2_io_o_3_out[4] ,
    \cb_4_2_io_o_3_out[3] ,
    \cb_4_2_io_o_3_out[2] ,
    \cb_4_2_io_o_3_out[1] ,
    \cb_4_2_io_o_3_out[0] }),
    .io_o_4_out({\cb_4_2_io_o_4_out[7] ,
    \cb_4_2_io_o_4_out[6] ,
    \cb_4_2_io_o_4_out[5] ,
    \cb_4_2_io_o_4_out[4] ,
    \cb_4_2_io_o_4_out[3] ,
    \cb_4_2_io_o_4_out[2] ,
    \cb_4_2_io_o_4_out[1] ,
    \cb_4_2_io_o_4_out[0] }),
    .io_o_5_out({\cb_4_2_io_o_5_out[7] ,
    \cb_4_2_io_o_5_out[6] ,
    \cb_4_2_io_o_5_out[5] ,
    \cb_4_2_io_o_5_out[4] ,
    \cb_4_2_io_o_5_out[3] ,
    \cb_4_2_io_o_5_out[2] ,
    \cb_4_2_io_o_5_out[1] ,
    \cb_4_2_io_o_5_out[0] }),
    .io_o_6_out({\cb_4_2_io_o_6_out[7] ,
    \cb_4_2_io_o_6_out[6] ,
    \cb_4_2_io_o_6_out[5] ,
    \cb_4_2_io_o_6_out[4] ,
    \cb_4_2_io_o_6_out[3] ,
    \cb_4_2_io_o_6_out[2] ,
    \cb_4_2_io_o_6_out[1] ,
    \cb_4_2_io_o_6_out[0] }),
    .io_o_7_out({\cb_4_2_io_o_7_out[7] ,
    \cb_4_2_io_o_7_out[6] ,
    \cb_4_2_io_o_7_out[5] ,
    \cb_4_2_io_o_7_out[4] ,
    \cb_4_2_io_o_7_out[3] ,
    \cb_4_2_io_o_7_out[2] ,
    \cb_4_2_io_o_7_out[1] ,
    \cb_4_2_io_o_7_out[0] }),
    .io_wo({\cb_4_1_io_eo[63] ,
    \cb_4_1_io_eo[62] ,
    \cb_4_1_io_eo[61] ,
    \cb_4_1_io_eo[60] ,
    \cb_4_1_io_eo[59] ,
    \cb_4_1_io_eo[58] ,
    \cb_4_1_io_eo[57] ,
    \cb_4_1_io_eo[56] ,
    \cb_4_1_io_eo[55] ,
    \cb_4_1_io_eo[54] ,
    \cb_4_1_io_eo[53] ,
    \cb_4_1_io_eo[52] ,
    \cb_4_1_io_eo[51] ,
    \cb_4_1_io_eo[50] ,
    \cb_4_1_io_eo[49] ,
    \cb_4_1_io_eo[48] ,
    \cb_4_1_io_eo[47] ,
    \cb_4_1_io_eo[46] ,
    \cb_4_1_io_eo[45] ,
    \cb_4_1_io_eo[44] ,
    \cb_4_1_io_eo[43] ,
    \cb_4_1_io_eo[42] ,
    \cb_4_1_io_eo[41] ,
    \cb_4_1_io_eo[40] ,
    \cb_4_1_io_eo[39] ,
    \cb_4_1_io_eo[38] ,
    \cb_4_1_io_eo[37] ,
    \cb_4_1_io_eo[36] ,
    \cb_4_1_io_eo[35] ,
    \cb_4_1_io_eo[34] ,
    \cb_4_1_io_eo[33] ,
    \cb_4_1_io_eo[32] ,
    \cb_4_1_io_eo[31] ,
    \cb_4_1_io_eo[30] ,
    \cb_4_1_io_eo[29] ,
    \cb_4_1_io_eo[28] ,
    \cb_4_1_io_eo[27] ,
    \cb_4_1_io_eo[26] ,
    \cb_4_1_io_eo[25] ,
    \cb_4_1_io_eo[24] ,
    \cb_4_1_io_eo[23] ,
    \cb_4_1_io_eo[22] ,
    \cb_4_1_io_eo[21] ,
    \cb_4_1_io_eo[20] ,
    \cb_4_1_io_eo[19] ,
    \cb_4_1_io_eo[18] ,
    \cb_4_1_io_eo[17] ,
    \cb_4_1_io_eo[16] ,
    \cb_4_1_io_eo[15] ,
    \cb_4_1_io_eo[14] ,
    \cb_4_1_io_eo[13] ,
    \cb_4_1_io_eo[12] ,
    \cb_4_1_io_eo[11] ,
    \cb_4_1_io_eo[10] ,
    \cb_4_1_io_eo[9] ,
    \cb_4_1_io_eo[8] ,
    \cb_4_1_io_eo[7] ,
    \cb_4_1_io_eo[6] ,
    \cb_4_1_io_eo[5] ,
    \cb_4_1_io_eo[4] ,
    \cb_4_1_io_eo[3] ,
    \cb_4_1_io_eo[2] ,
    \cb_4_1_io_eo[1] ,
    \cb_4_1_io_eo[0] }));
 cic_block cb_4_3 (.io_cs_i(cb_4_3_io_cs_i),
    .io_i_0_ci(cb_4_2_io_o_0_co),
    .io_i_1_ci(cb_4_2_io_o_1_co),
    .io_i_2_ci(cb_4_2_io_o_2_co),
    .io_i_3_ci(cb_4_2_io_o_3_co),
    .io_i_4_ci(cb_4_2_io_o_4_co),
    .io_i_5_ci(cb_4_2_io_o_5_co),
    .io_i_6_ci(cb_4_2_io_o_6_co),
    .io_i_7_ci(cb_4_2_io_o_7_co),
    .io_o_0_co(cb_4_3_io_o_0_co),
    .io_o_1_co(cb_4_3_io_o_1_co),
    .io_o_2_co(cb_4_3_io_o_2_co),
    .io_o_3_co(cb_4_3_io_o_3_co),
    .io_o_4_co(cb_4_3_io_o_4_co),
    .io_o_5_co(cb_4_3_io_o_5_co),
    .io_o_6_co(cb_4_3_io_o_6_co),
    .io_o_7_co(cb_4_3_io_o_7_co),
    .io_vci(cb_4_2_io_vco),
    .io_vco(cb_4_3_io_vco),
    .io_vi(cb_4_3_io_vi),
    .io_we_i(cb_4_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_4_0_io_adr_i[1] ,
    \cb_4_0_io_adr_i[0] }),
    .io_dat_i({\cb_4_0_io_dat_i[15] ,
    \cb_4_0_io_dat_i[14] ,
    \cb_4_0_io_dat_i[13] ,
    \cb_4_0_io_dat_i[12] ,
    \cb_4_0_io_dat_i[11] ,
    \cb_4_0_io_dat_i[10] ,
    \cb_4_0_io_dat_i[9] ,
    \cb_4_0_io_dat_i[8] ,
    \cb_4_0_io_dat_i[7] ,
    \cb_4_0_io_dat_i[6] ,
    \cb_4_0_io_dat_i[5] ,
    \cb_4_0_io_dat_i[4] ,
    \cb_4_0_io_dat_i[3] ,
    \cb_4_0_io_dat_i[2] ,
    \cb_4_0_io_dat_i[1] ,
    \cb_4_0_io_dat_i[0] }),
    .io_dat_o({\cb_4_3_io_dat_o[15] ,
    \cb_4_3_io_dat_o[14] ,
    \cb_4_3_io_dat_o[13] ,
    \cb_4_3_io_dat_o[12] ,
    \cb_4_3_io_dat_o[11] ,
    \cb_4_3_io_dat_o[10] ,
    \cb_4_3_io_dat_o[9] ,
    \cb_4_3_io_dat_o[8] ,
    \cb_4_3_io_dat_o[7] ,
    \cb_4_3_io_dat_o[6] ,
    \cb_4_3_io_dat_o[5] ,
    \cb_4_3_io_dat_o[4] ,
    \cb_4_3_io_dat_o[3] ,
    \cb_4_3_io_dat_o[2] ,
    \cb_4_3_io_dat_o[1] ,
    \cb_4_3_io_dat_o[0] }),
    .io_eo({\cb_4_3_io_eo[63] ,
    \cb_4_3_io_eo[62] ,
    \cb_4_3_io_eo[61] ,
    \cb_4_3_io_eo[60] ,
    \cb_4_3_io_eo[59] ,
    \cb_4_3_io_eo[58] ,
    \cb_4_3_io_eo[57] ,
    \cb_4_3_io_eo[56] ,
    \cb_4_3_io_eo[55] ,
    \cb_4_3_io_eo[54] ,
    \cb_4_3_io_eo[53] ,
    \cb_4_3_io_eo[52] ,
    \cb_4_3_io_eo[51] ,
    \cb_4_3_io_eo[50] ,
    \cb_4_3_io_eo[49] ,
    \cb_4_3_io_eo[48] ,
    \cb_4_3_io_eo[47] ,
    \cb_4_3_io_eo[46] ,
    \cb_4_3_io_eo[45] ,
    \cb_4_3_io_eo[44] ,
    \cb_4_3_io_eo[43] ,
    \cb_4_3_io_eo[42] ,
    \cb_4_3_io_eo[41] ,
    \cb_4_3_io_eo[40] ,
    \cb_4_3_io_eo[39] ,
    \cb_4_3_io_eo[38] ,
    \cb_4_3_io_eo[37] ,
    \cb_4_3_io_eo[36] ,
    \cb_4_3_io_eo[35] ,
    \cb_4_3_io_eo[34] ,
    \cb_4_3_io_eo[33] ,
    \cb_4_3_io_eo[32] ,
    \cb_4_3_io_eo[31] ,
    \cb_4_3_io_eo[30] ,
    \cb_4_3_io_eo[29] ,
    \cb_4_3_io_eo[28] ,
    \cb_4_3_io_eo[27] ,
    \cb_4_3_io_eo[26] ,
    \cb_4_3_io_eo[25] ,
    \cb_4_3_io_eo[24] ,
    \cb_4_3_io_eo[23] ,
    \cb_4_3_io_eo[22] ,
    \cb_4_3_io_eo[21] ,
    \cb_4_3_io_eo[20] ,
    \cb_4_3_io_eo[19] ,
    \cb_4_3_io_eo[18] ,
    \cb_4_3_io_eo[17] ,
    \cb_4_3_io_eo[16] ,
    \cb_4_3_io_eo[15] ,
    \cb_4_3_io_eo[14] ,
    \cb_4_3_io_eo[13] ,
    \cb_4_3_io_eo[12] ,
    \cb_4_3_io_eo[11] ,
    \cb_4_3_io_eo[10] ,
    \cb_4_3_io_eo[9] ,
    \cb_4_3_io_eo[8] ,
    \cb_4_3_io_eo[7] ,
    \cb_4_3_io_eo[6] ,
    \cb_4_3_io_eo[5] ,
    \cb_4_3_io_eo[4] ,
    \cb_4_3_io_eo[3] ,
    \cb_4_3_io_eo[2] ,
    \cb_4_3_io_eo[1] ,
    \cb_4_3_io_eo[0] }),
    .io_i_0_in1({\cb_4_2_io_o_0_out[7] ,
    \cb_4_2_io_o_0_out[6] ,
    \cb_4_2_io_o_0_out[5] ,
    \cb_4_2_io_o_0_out[4] ,
    \cb_4_2_io_o_0_out[3] ,
    \cb_4_2_io_o_0_out[2] ,
    \cb_4_2_io_o_0_out[1] ,
    \cb_4_2_io_o_0_out[0] }),
    .io_i_1_in1({\cb_4_2_io_o_1_out[7] ,
    \cb_4_2_io_o_1_out[6] ,
    \cb_4_2_io_o_1_out[5] ,
    \cb_4_2_io_o_1_out[4] ,
    \cb_4_2_io_o_1_out[3] ,
    \cb_4_2_io_o_1_out[2] ,
    \cb_4_2_io_o_1_out[1] ,
    \cb_4_2_io_o_1_out[0] }),
    .io_i_2_in1({\cb_4_2_io_o_2_out[7] ,
    \cb_4_2_io_o_2_out[6] ,
    \cb_4_2_io_o_2_out[5] ,
    \cb_4_2_io_o_2_out[4] ,
    \cb_4_2_io_o_2_out[3] ,
    \cb_4_2_io_o_2_out[2] ,
    \cb_4_2_io_o_2_out[1] ,
    \cb_4_2_io_o_2_out[0] }),
    .io_i_3_in1({\cb_4_2_io_o_3_out[7] ,
    \cb_4_2_io_o_3_out[6] ,
    \cb_4_2_io_o_3_out[5] ,
    \cb_4_2_io_o_3_out[4] ,
    \cb_4_2_io_o_3_out[3] ,
    \cb_4_2_io_o_3_out[2] ,
    \cb_4_2_io_o_3_out[1] ,
    \cb_4_2_io_o_3_out[0] }),
    .io_i_4_in1({\cb_4_2_io_o_4_out[7] ,
    \cb_4_2_io_o_4_out[6] ,
    \cb_4_2_io_o_4_out[5] ,
    \cb_4_2_io_o_4_out[4] ,
    \cb_4_2_io_o_4_out[3] ,
    \cb_4_2_io_o_4_out[2] ,
    \cb_4_2_io_o_4_out[1] ,
    \cb_4_2_io_o_4_out[0] }),
    .io_i_5_in1({\cb_4_2_io_o_5_out[7] ,
    \cb_4_2_io_o_5_out[6] ,
    \cb_4_2_io_o_5_out[5] ,
    \cb_4_2_io_o_5_out[4] ,
    \cb_4_2_io_o_5_out[3] ,
    \cb_4_2_io_o_5_out[2] ,
    \cb_4_2_io_o_5_out[1] ,
    \cb_4_2_io_o_5_out[0] }),
    .io_i_6_in1({\cb_4_2_io_o_6_out[7] ,
    \cb_4_2_io_o_6_out[6] ,
    \cb_4_2_io_o_6_out[5] ,
    \cb_4_2_io_o_6_out[4] ,
    \cb_4_2_io_o_6_out[3] ,
    \cb_4_2_io_o_6_out[2] ,
    \cb_4_2_io_o_6_out[1] ,
    \cb_4_2_io_o_6_out[0] }),
    .io_i_7_in1({\cb_4_2_io_o_7_out[7] ,
    \cb_4_2_io_o_7_out[6] ,
    \cb_4_2_io_o_7_out[5] ,
    \cb_4_2_io_o_7_out[4] ,
    \cb_4_2_io_o_7_out[3] ,
    \cb_4_2_io_o_7_out[2] ,
    \cb_4_2_io_o_7_out[1] ,
    \cb_4_2_io_o_7_out[0] }),
    .io_o_0_out({\cb_4_3_io_o_0_out[7] ,
    \cb_4_3_io_o_0_out[6] ,
    \cb_4_3_io_o_0_out[5] ,
    \cb_4_3_io_o_0_out[4] ,
    \cb_4_3_io_o_0_out[3] ,
    \cb_4_3_io_o_0_out[2] ,
    \cb_4_3_io_o_0_out[1] ,
    \cb_4_3_io_o_0_out[0] }),
    .io_o_1_out({\cb_4_3_io_o_1_out[7] ,
    \cb_4_3_io_o_1_out[6] ,
    \cb_4_3_io_o_1_out[5] ,
    \cb_4_3_io_o_1_out[4] ,
    \cb_4_3_io_o_1_out[3] ,
    \cb_4_3_io_o_1_out[2] ,
    \cb_4_3_io_o_1_out[1] ,
    \cb_4_3_io_o_1_out[0] }),
    .io_o_2_out({\cb_4_3_io_o_2_out[7] ,
    \cb_4_3_io_o_2_out[6] ,
    \cb_4_3_io_o_2_out[5] ,
    \cb_4_3_io_o_2_out[4] ,
    \cb_4_3_io_o_2_out[3] ,
    \cb_4_3_io_o_2_out[2] ,
    \cb_4_3_io_o_2_out[1] ,
    \cb_4_3_io_o_2_out[0] }),
    .io_o_3_out({\cb_4_3_io_o_3_out[7] ,
    \cb_4_3_io_o_3_out[6] ,
    \cb_4_3_io_o_3_out[5] ,
    \cb_4_3_io_o_3_out[4] ,
    \cb_4_3_io_o_3_out[3] ,
    \cb_4_3_io_o_3_out[2] ,
    \cb_4_3_io_o_3_out[1] ,
    \cb_4_3_io_o_3_out[0] }),
    .io_o_4_out({\cb_4_3_io_o_4_out[7] ,
    \cb_4_3_io_o_4_out[6] ,
    \cb_4_3_io_o_4_out[5] ,
    \cb_4_3_io_o_4_out[4] ,
    \cb_4_3_io_o_4_out[3] ,
    \cb_4_3_io_o_4_out[2] ,
    \cb_4_3_io_o_4_out[1] ,
    \cb_4_3_io_o_4_out[0] }),
    .io_o_5_out({\cb_4_3_io_o_5_out[7] ,
    \cb_4_3_io_o_5_out[6] ,
    \cb_4_3_io_o_5_out[5] ,
    \cb_4_3_io_o_5_out[4] ,
    \cb_4_3_io_o_5_out[3] ,
    \cb_4_3_io_o_5_out[2] ,
    \cb_4_3_io_o_5_out[1] ,
    \cb_4_3_io_o_5_out[0] }),
    .io_o_6_out({\cb_4_3_io_o_6_out[7] ,
    \cb_4_3_io_o_6_out[6] ,
    \cb_4_3_io_o_6_out[5] ,
    \cb_4_3_io_o_6_out[4] ,
    \cb_4_3_io_o_6_out[3] ,
    \cb_4_3_io_o_6_out[2] ,
    \cb_4_3_io_o_6_out[1] ,
    \cb_4_3_io_o_6_out[0] }),
    .io_o_7_out({\cb_4_3_io_o_7_out[7] ,
    \cb_4_3_io_o_7_out[6] ,
    \cb_4_3_io_o_7_out[5] ,
    \cb_4_3_io_o_7_out[4] ,
    \cb_4_3_io_o_7_out[3] ,
    \cb_4_3_io_o_7_out[2] ,
    \cb_4_3_io_o_7_out[1] ,
    \cb_4_3_io_o_7_out[0] }),
    .io_wo({\cb_4_2_io_eo[63] ,
    \cb_4_2_io_eo[62] ,
    \cb_4_2_io_eo[61] ,
    \cb_4_2_io_eo[60] ,
    \cb_4_2_io_eo[59] ,
    \cb_4_2_io_eo[58] ,
    \cb_4_2_io_eo[57] ,
    \cb_4_2_io_eo[56] ,
    \cb_4_2_io_eo[55] ,
    \cb_4_2_io_eo[54] ,
    \cb_4_2_io_eo[53] ,
    \cb_4_2_io_eo[52] ,
    \cb_4_2_io_eo[51] ,
    \cb_4_2_io_eo[50] ,
    \cb_4_2_io_eo[49] ,
    \cb_4_2_io_eo[48] ,
    \cb_4_2_io_eo[47] ,
    \cb_4_2_io_eo[46] ,
    \cb_4_2_io_eo[45] ,
    \cb_4_2_io_eo[44] ,
    \cb_4_2_io_eo[43] ,
    \cb_4_2_io_eo[42] ,
    \cb_4_2_io_eo[41] ,
    \cb_4_2_io_eo[40] ,
    \cb_4_2_io_eo[39] ,
    \cb_4_2_io_eo[38] ,
    \cb_4_2_io_eo[37] ,
    \cb_4_2_io_eo[36] ,
    \cb_4_2_io_eo[35] ,
    \cb_4_2_io_eo[34] ,
    \cb_4_2_io_eo[33] ,
    \cb_4_2_io_eo[32] ,
    \cb_4_2_io_eo[31] ,
    \cb_4_2_io_eo[30] ,
    \cb_4_2_io_eo[29] ,
    \cb_4_2_io_eo[28] ,
    \cb_4_2_io_eo[27] ,
    \cb_4_2_io_eo[26] ,
    \cb_4_2_io_eo[25] ,
    \cb_4_2_io_eo[24] ,
    \cb_4_2_io_eo[23] ,
    \cb_4_2_io_eo[22] ,
    \cb_4_2_io_eo[21] ,
    \cb_4_2_io_eo[20] ,
    \cb_4_2_io_eo[19] ,
    \cb_4_2_io_eo[18] ,
    \cb_4_2_io_eo[17] ,
    \cb_4_2_io_eo[16] ,
    \cb_4_2_io_eo[15] ,
    \cb_4_2_io_eo[14] ,
    \cb_4_2_io_eo[13] ,
    \cb_4_2_io_eo[12] ,
    \cb_4_2_io_eo[11] ,
    \cb_4_2_io_eo[10] ,
    \cb_4_2_io_eo[9] ,
    \cb_4_2_io_eo[8] ,
    \cb_4_2_io_eo[7] ,
    \cb_4_2_io_eo[6] ,
    \cb_4_2_io_eo[5] ,
    \cb_4_2_io_eo[4] ,
    \cb_4_2_io_eo[3] ,
    \cb_4_2_io_eo[2] ,
    \cb_4_2_io_eo[1] ,
    \cb_4_2_io_eo[0] }));
 cic_block cb_4_4 (.io_cs_i(cb_4_4_io_cs_i),
    .io_i_0_ci(cb_4_3_io_o_0_co),
    .io_i_1_ci(cb_4_3_io_o_1_co),
    .io_i_2_ci(cb_4_3_io_o_2_co),
    .io_i_3_ci(cb_4_3_io_o_3_co),
    .io_i_4_ci(cb_4_3_io_o_4_co),
    .io_i_5_ci(cb_4_3_io_o_5_co),
    .io_i_6_ci(cb_4_3_io_o_6_co),
    .io_i_7_ci(cb_4_3_io_o_7_co),
    .io_o_0_co(cb_4_4_io_o_0_co),
    .io_o_1_co(cb_4_4_io_o_1_co),
    .io_o_2_co(cb_4_4_io_o_2_co),
    .io_o_3_co(cb_4_4_io_o_3_co),
    .io_o_4_co(cb_4_4_io_o_4_co),
    .io_o_5_co(cb_4_4_io_o_5_co),
    .io_o_6_co(cb_4_4_io_o_6_co),
    .io_o_7_co(cb_4_4_io_o_7_co),
    .io_vci(cb_4_3_io_vco),
    .io_vco(cb_4_4_io_vco),
    .io_vi(cb_4_4_io_vi),
    .io_we_i(cb_4_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_4_0_io_adr_i[1] ,
    \cb_4_0_io_adr_i[0] }),
    .io_dat_i({\cb_4_0_io_dat_i[15] ,
    \cb_4_0_io_dat_i[14] ,
    \cb_4_0_io_dat_i[13] ,
    \cb_4_0_io_dat_i[12] ,
    \cb_4_0_io_dat_i[11] ,
    \cb_4_0_io_dat_i[10] ,
    \cb_4_0_io_dat_i[9] ,
    \cb_4_0_io_dat_i[8] ,
    \cb_4_0_io_dat_i[7] ,
    \cb_4_0_io_dat_i[6] ,
    \cb_4_0_io_dat_i[5] ,
    \cb_4_0_io_dat_i[4] ,
    \cb_4_0_io_dat_i[3] ,
    \cb_4_0_io_dat_i[2] ,
    \cb_4_0_io_dat_i[1] ,
    \cb_4_0_io_dat_i[0] }),
    .io_dat_o({\cb_4_4_io_dat_o[15] ,
    \cb_4_4_io_dat_o[14] ,
    \cb_4_4_io_dat_o[13] ,
    \cb_4_4_io_dat_o[12] ,
    \cb_4_4_io_dat_o[11] ,
    \cb_4_4_io_dat_o[10] ,
    \cb_4_4_io_dat_o[9] ,
    \cb_4_4_io_dat_o[8] ,
    \cb_4_4_io_dat_o[7] ,
    \cb_4_4_io_dat_o[6] ,
    \cb_4_4_io_dat_o[5] ,
    \cb_4_4_io_dat_o[4] ,
    \cb_4_4_io_dat_o[3] ,
    \cb_4_4_io_dat_o[2] ,
    \cb_4_4_io_dat_o[1] ,
    \cb_4_4_io_dat_o[0] }),
    .io_eo({\cb_4_4_io_eo[63] ,
    \cb_4_4_io_eo[62] ,
    \cb_4_4_io_eo[61] ,
    \cb_4_4_io_eo[60] ,
    \cb_4_4_io_eo[59] ,
    \cb_4_4_io_eo[58] ,
    \cb_4_4_io_eo[57] ,
    \cb_4_4_io_eo[56] ,
    \cb_4_4_io_eo[55] ,
    \cb_4_4_io_eo[54] ,
    \cb_4_4_io_eo[53] ,
    \cb_4_4_io_eo[52] ,
    \cb_4_4_io_eo[51] ,
    \cb_4_4_io_eo[50] ,
    \cb_4_4_io_eo[49] ,
    \cb_4_4_io_eo[48] ,
    \cb_4_4_io_eo[47] ,
    \cb_4_4_io_eo[46] ,
    \cb_4_4_io_eo[45] ,
    \cb_4_4_io_eo[44] ,
    \cb_4_4_io_eo[43] ,
    \cb_4_4_io_eo[42] ,
    \cb_4_4_io_eo[41] ,
    \cb_4_4_io_eo[40] ,
    \cb_4_4_io_eo[39] ,
    \cb_4_4_io_eo[38] ,
    \cb_4_4_io_eo[37] ,
    \cb_4_4_io_eo[36] ,
    \cb_4_4_io_eo[35] ,
    \cb_4_4_io_eo[34] ,
    \cb_4_4_io_eo[33] ,
    \cb_4_4_io_eo[32] ,
    \cb_4_4_io_eo[31] ,
    \cb_4_4_io_eo[30] ,
    \cb_4_4_io_eo[29] ,
    \cb_4_4_io_eo[28] ,
    \cb_4_4_io_eo[27] ,
    \cb_4_4_io_eo[26] ,
    \cb_4_4_io_eo[25] ,
    \cb_4_4_io_eo[24] ,
    \cb_4_4_io_eo[23] ,
    \cb_4_4_io_eo[22] ,
    \cb_4_4_io_eo[21] ,
    \cb_4_4_io_eo[20] ,
    \cb_4_4_io_eo[19] ,
    \cb_4_4_io_eo[18] ,
    \cb_4_4_io_eo[17] ,
    \cb_4_4_io_eo[16] ,
    \cb_4_4_io_eo[15] ,
    \cb_4_4_io_eo[14] ,
    \cb_4_4_io_eo[13] ,
    \cb_4_4_io_eo[12] ,
    \cb_4_4_io_eo[11] ,
    \cb_4_4_io_eo[10] ,
    \cb_4_4_io_eo[9] ,
    \cb_4_4_io_eo[8] ,
    \cb_4_4_io_eo[7] ,
    \cb_4_4_io_eo[6] ,
    \cb_4_4_io_eo[5] ,
    \cb_4_4_io_eo[4] ,
    \cb_4_4_io_eo[3] ,
    \cb_4_4_io_eo[2] ,
    \cb_4_4_io_eo[1] ,
    \cb_4_4_io_eo[0] }),
    .io_i_0_in1({\cb_4_3_io_o_0_out[7] ,
    \cb_4_3_io_o_0_out[6] ,
    \cb_4_3_io_o_0_out[5] ,
    \cb_4_3_io_o_0_out[4] ,
    \cb_4_3_io_o_0_out[3] ,
    \cb_4_3_io_o_0_out[2] ,
    \cb_4_3_io_o_0_out[1] ,
    \cb_4_3_io_o_0_out[0] }),
    .io_i_1_in1({\cb_4_3_io_o_1_out[7] ,
    \cb_4_3_io_o_1_out[6] ,
    \cb_4_3_io_o_1_out[5] ,
    \cb_4_3_io_o_1_out[4] ,
    \cb_4_3_io_o_1_out[3] ,
    \cb_4_3_io_o_1_out[2] ,
    \cb_4_3_io_o_1_out[1] ,
    \cb_4_3_io_o_1_out[0] }),
    .io_i_2_in1({\cb_4_3_io_o_2_out[7] ,
    \cb_4_3_io_o_2_out[6] ,
    \cb_4_3_io_o_2_out[5] ,
    \cb_4_3_io_o_2_out[4] ,
    \cb_4_3_io_o_2_out[3] ,
    \cb_4_3_io_o_2_out[2] ,
    \cb_4_3_io_o_2_out[1] ,
    \cb_4_3_io_o_2_out[0] }),
    .io_i_3_in1({\cb_4_3_io_o_3_out[7] ,
    \cb_4_3_io_o_3_out[6] ,
    \cb_4_3_io_o_3_out[5] ,
    \cb_4_3_io_o_3_out[4] ,
    \cb_4_3_io_o_3_out[3] ,
    \cb_4_3_io_o_3_out[2] ,
    \cb_4_3_io_o_3_out[1] ,
    \cb_4_3_io_o_3_out[0] }),
    .io_i_4_in1({\cb_4_3_io_o_4_out[7] ,
    \cb_4_3_io_o_4_out[6] ,
    \cb_4_3_io_o_4_out[5] ,
    \cb_4_3_io_o_4_out[4] ,
    \cb_4_3_io_o_4_out[3] ,
    \cb_4_3_io_o_4_out[2] ,
    \cb_4_3_io_o_4_out[1] ,
    \cb_4_3_io_o_4_out[0] }),
    .io_i_5_in1({\cb_4_3_io_o_5_out[7] ,
    \cb_4_3_io_o_5_out[6] ,
    \cb_4_3_io_o_5_out[5] ,
    \cb_4_3_io_o_5_out[4] ,
    \cb_4_3_io_o_5_out[3] ,
    \cb_4_3_io_o_5_out[2] ,
    \cb_4_3_io_o_5_out[1] ,
    \cb_4_3_io_o_5_out[0] }),
    .io_i_6_in1({\cb_4_3_io_o_6_out[7] ,
    \cb_4_3_io_o_6_out[6] ,
    \cb_4_3_io_o_6_out[5] ,
    \cb_4_3_io_o_6_out[4] ,
    \cb_4_3_io_o_6_out[3] ,
    \cb_4_3_io_o_6_out[2] ,
    \cb_4_3_io_o_6_out[1] ,
    \cb_4_3_io_o_6_out[0] }),
    .io_i_7_in1({\cb_4_3_io_o_7_out[7] ,
    \cb_4_3_io_o_7_out[6] ,
    \cb_4_3_io_o_7_out[5] ,
    \cb_4_3_io_o_7_out[4] ,
    \cb_4_3_io_o_7_out[3] ,
    \cb_4_3_io_o_7_out[2] ,
    \cb_4_3_io_o_7_out[1] ,
    \cb_4_3_io_o_7_out[0] }),
    .io_o_0_out({\cb_4_4_io_o_0_out[7] ,
    \cb_4_4_io_o_0_out[6] ,
    \cb_4_4_io_o_0_out[5] ,
    \cb_4_4_io_o_0_out[4] ,
    \cb_4_4_io_o_0_out[3] ,
    \cb_4_4_io_o_0_out[2] ,
    \cb_4_4_io_o_0_out[1] ,
    \cb_4_4_io_o_0_out[0] }),
    .io_o_1_out({\cb_4_4_io_o_1_out[7] ,
    \cb_4_4_io_o_1_out[6] ,
    \cb_4_4_io_o_1_out[5] ,
    \cb_4_4_io_o_1_out[4] ,
    \cb_4_4_io_o_1_out[3] ,
    \cb_4_4_io_o_1_out[2] ,
    \cb_4_4_io_o_1_out[1] ,
    \cb_4_4_io_o_1_out[0] }),
    .io_o_2_out({\cb_4_4_io_o_2_out[7] ,
    \cb_4_4_io_o_2_out[6] ,
    \cb_4_4_io_o_2_out[5] ,
    \cb_4_4_io_o_2_out[4] ,
    \cb_4_4_io_o_2_out[3] ,
    \cb_4_4_io_o_2_out[2] ,
    \cb_4_4_io_o_2_out[1] ,
    \cb_4_4_io_o_2_out[0] }),
    .io_o_3_out({\cb_4_4_io_o_3_out[7] ,
    \cb_4_4_io_o_3_out[6] ,
    \cb_4_4_io_o_3_out[5] ,
    \cb_4_4_io_o_3_out[4] ,
    \cb_4_4_io_o_3_out[3] ,
    \cb_4_4_io_o_3_out[2] ,
    \cb_4_4_io_o_3_out[1] ,
    \cb_4_4_io_o_3_out[0] }),
    .io_o_4_out({\cb_4_4_io_o_4_out[7] ,
    \cb_4_4_io_o_4_out[6] ,
    \cb_4_4_io_o_4_out[5] ,
    \cb_4_4_io_o_4_out[4] ,
    \cb_4_4_io_o_4_out[3] ,
    \cb_4_4_io_o_4_out[2] ,
    \cb_4_4_io_o_4_out[1] ,
    \cb_4_4_io_o_4_out[0] }),
    .io_o_5_out({\cb_4_4_io_o_5_out[7] ,
    \cb_4_4_io_o_5_out[6] ,
    \cb_4_4_io_o_5_out[5] ,
    \cb_4_4_io_o_5_out[4] ,
    \cb_4_4_io_o_5_out[3] ,
    \cb_4_4_io_o_5_out[2] ,
    \cb_4_4_io_o_5_out[1] ,
    \cb_4_4_io_o_5_out[0] }),
    .io_o_6_out({\cb_4_4_io_o_6_out[7] ,
    \cb_4_4_io_o_6_out[6] ,
    \cb_4_4_io_o_6_out[5] ,
    \cb_4_4_io_o_6_out[4] ,
    \cb_4_4_io_o_6_out[3] ,
    \cb_4_4_io_o_6_out[2] ,
    \cb_4_4_io_o_6_out[1] ,
    \cb_4_4_io_o_6_out[0] }),
    .io_o_7_out({\cb_4_4_io_o_7_out[7] ,
    \cb_4_4_io_o_7_out[6] ,
    \cb_4_4_io_o_7_out[5] ,
    \cb_4_4_io_o_7_out[4] ,
    \cb_4_4_io_o_7_out[3] ,
    \cb_4_4_io_o_7_out[2] ,
    \cb_4_4_io_o_7_out[1] ,
    \cb_4_4_io_o_7_out[0] }),
    .io_wo({\cb_4_3_io_eo[63] ,
    \cb_4_3_io_eo[62] ,
    \cb_4_3_io_eo[61] ,
    \cb_4_3_io_eo[60] ,
    \cb_4_3_io_eo[59] ,
    \cb_4_3_io_eo[58] ,
    \cb_4_3_io_eo[57] ,
    \cb_4_3_io_eo[56] ,
    \cb_4_3_io_eo[55] ,
    \cb_4_3_io_eo[54] ,
    \cb_4_3_io_eo[53] ,
    \cb_4_3_io_eo[52] ,
    \cb_4_3_io_eo[51] ,
    \cb_4_3_io_eo[50] ,
    \cb_4_3_io_eo[49] ,
    \cb_4_3_io_eo[48] ,
    \cb_4_3_io_eo[47] ,
    \cb_4_3_io_eo[46] ,
    \cb_4_3_io_eo[45] ,
    \cb_4_3_io_eo[44] ,
    \cb_4_3_io_eo[43] ,
    \cb_4_3_io_eo[42] ,
    \cb_4_3_io_eo[41] ,
    \cb_4_3_io_eo[40] ,
    \cb_4_3_io_eo[39] ,
    \cb_4_3_io_eo[38] ,
    \cb_4_3_io_eo[37] ,
    \cb_4_3_io_eo[36] ,
    \cb_4_3_io_eo[35] ,
    \cb_4_3_io_eo[34] ,
    \cb_4_3_io_eo[33] ,
    \cb_4_3_io_eo[32] ,
    \cb_4_3_io_eo[31] ,
    \cb_4_3_io_eo[30] ,
    \cb_4_3_io_eo[29] ,
    \cb_4_3_io_eo[28] ,
    \cb_4_3_io_eo[27] ,
    \cb_4_3_io_eo[26] ,
    \cb_4_3_io_eo[25] ,
    \cb_4_3_io_eo[24] ,
    \cb_4_3_io_eo[23] ,
    \cb_4_3_io_eo[22] ,
    \cb_4_3_io_eo[21] ,
    \cb_4_3_io_eo[20] ,
    \cb_4_3_io_eo[19] ,
    \cb_4_3_io_eo[18] ,
    \cb_4_3_io_eo[17] ,
    \cb_4_3_io_eo[16] ,
    \cb_4_3_io_eo[15] ,
    \cb_4_3_io_eo[14] ,
    \cb_4_3_io_eo[13] ,
    \cb_4_3_io_eo[12] ,
    \cb_4_3_io_eo[11] ,
    \cb_4_3_io_eo[10] ,
    \cb_4_3_io_eo[9] ,
    \cb_4_3_io_eo[8] ,
    \cb_4_3_io_eo[7] ,
    \cb_4_3_io_eo[6] ,
    \cb_4_3_io_eo[5] ,
    \cb_4_3_io_eo[4] ,
    \cb_4_3_io_eo[3] ,
    \cb_4_3_io_eo[2] ,
    \cb_4_3_io_eo[1] ,
    \cb_4_3_io_eo[0] }));
 cic_block cb_4_5 (.io_cs_i(cb_4_5_io_cs_i),
    .io_i_0_ci(cb_4_4_io_o_0_co),
    .io_i_1_ci(cb_4_4_io_o_1_co),
    .io_i_2_ci(cb_4_4_io_o_2_co),
    .io_i_3_ci(cb_4_4_io_o_3_co),
    .io_i_4_ci(cb_4_4_io_o_4_co),
    .io_i_5_ci(cb_4_4_io_o_5_co),
    .io_i_6_ci(cb_4_4_io_o_6_co),
    .io_i_7_ci(cb_4_4_io_o_7_co),
    .io_o_0_co(cb_4_5_io_o_0_co),
    .io_o_1_co(cb_4_5_io_o_1_co),
    .io_o_2_co(cb_4_5_io_o_2_co),
    .io_o_3_co(cb_4_5_io_o_3_co),
    .io_o_4_co(cb_4_5_io_o_4_co),
    .io_o_5_co(cb_4_5_io_o_5_co),
    .io_o_6_co(cb_4_5_io_o_6_co),
    .io_o_7_co(cb_4_5_io_o_7_co),
    .io_vci(cb_4_4_io_vco),
    .io_vco(cb_4_5_io_vco),
    .io_vi(cb_4_5_io_vi),
    .io_we_i(cb_4_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_4_0_io_adr_i[1] ,
    \cb_4_0_io_adr_i[0] }),
    .io_dat_i({\cb_4_0_io_dat_i[15] ,
    \cb_4_0_io_dat_i[14] ,
    \cb_4_0_io_dat_i[13] ,
    \cb_4_0_io_dat_i[12] ,
    \cb_4_0_io_dat_i[11] ,
    \cb_4_0_io_dat_i[10] ,
    \cb_4_0_io_dat_i[9] ,
    \cb_4_0_io_dat_i[8] ,
    \cb_4_0_io_dat_i[7] ,
    \cb_4_0_io_dat_i[6] ,
    \cb_4_0_io_dat_i[5] ,
    \cb_4_0_io_dat_i[4] ,
    \cb_4_0_io_dat_i[3] ,
    \cb_4_0_io_dat_i[2] ,
    \cb_4_0_io_dat_i[1] ,
    \cb_4_0_io_dat_i[0] }),
    .io_dat_o({\cb_4_5_io_dat_o[15] ,
    \cb_4_5_io_dat_o[14] ,
    \cb_4_5_io_dat_o[13] ,
    \cb_4_5_io_dat_o[12] ,
    \cb_4_5_io_dat_o[11] ,
    \cb_4_5_io_dat_o[10] ,
    \cb_4_5_io_dat_o[9] ,
    \cb_4_5_io_dat_o[8] ,
    \cb_4_5_io_dat_o[7] ,
    \cb_4_5_io_dat_o[6] ,
    \cb_4_5_io_dat_o[5] ,
    \cb_4_5_io_dat_o[4] ,
    \cb_4_5_io_dat_o[3] ,
    \cb_4_5_io_dat_o[2] ,
    \cb_4_5_io_dat_o[1] ,
    \cb_4_5_io_dat_o[0] }),
    .io_eo({\cb_4_5_io_eo[63] ,
    \cb_4_5_io_eo[62] ,
    \cb_4_5_io_eo[61] ,
    \cb_4_5_io_eo[60] ,
    \cb_4_5_io_eo[59] ,
    \cb_4_5_io_eo[58] ,
    \cb_4_5_io_eo[57] ,
    \cb_4_5_io_eo[56] ,
    \cb_4_5_io_eo[55] ,
    \cb_4_5_io_eo[54] ,
    \cb_4_5_io_eo[53] ,
    \cb_4_5_io_eo[52] ,
    \cb_4_5_io_eo[51] ,
    \cb_4_5_io_eo[50] ,
    \cb_4_5_io_eo[49] ,
    \cb_4_5_io_eo[48] ,
    \cb_4_5_io_eo[47] ,
    \cb_4_5_io_eo[46] ,
    \cb_4_5_io_eo[45] ,
    \cb_4_5_io_eo[44] ,
    \cb_4_5_io_eo[43] ,
    \cb_4_5_io_eo[42] ,
    \cb_4_5_io_eo[41] ,
    \cb_4_5_io_eo[40] ,
    \cb_4_5_io_eo[39] ,
    \cb_4_5_io_eo[38] ,
    \cb_4_5_io_eo[37] ,
    \cb_4_5_io_eo[36] ,
    \cb_4_5_io_eo[35] ,
    \cb_4_5_io_eo[34] ,
    \cb_4_5_io_eo[33] ,
    \cb_4_5_io_eo[32] ,
    \cb_4_5_io_eo[31] ,
    \cb_4_5_io_eo[30] ,
    \cb_4_5_io_eo[29] ,
    \cb_4_5_io_eo[28] ,
    \cb_4_5_io_eo[27] ,
    \cb_4_5_io_eo[26] ,
    \cb_4_5_io_eo[25] ,
    \cb_4_5_io_eo[24] ,
    \cb_4_5_io_eo[23] ,
    \cb_4_5_io_eo[22] ,
    \cb_4_5_io_eo[21] ,
    \cb_4_5_io_eo[20] ,
    \cb_4_5_io_eo[19] ,
    \cb_4_5_io_eo[18] ,
    \cb_4_5_io_eo[17] ,
    \cb_4_5_io_eo[16] ,
    \cb_4_5_io_eo[15] ,
    \cb_4_5_io_eo[14] ,
    \cb_4_5_io_eo[13] ,
    \cb_4_5_io_eo[12] ,
    \cb_4_5_io_eo[11] ,
    \cb_4_5_io_eo[10] ,
    \cb_4_5_io_eo[9] ,
    \cb_4_5_io_eo[8] ,
    \cb_4_5_io_eo[7] ,
    \cb_4_5_io_eo[6] ,
    \cb_4_5_io_eo[5] ,
    \cb_4_5_io_eo[4] ,
    \cb_4_5_io_eo[3] ,
    \cb_4_5_io_eo[2] ,
    \cb_4_5_io_eo[1] ,
    \cb_4_5_io_eo[0] }),
    .io_i_0_in1({\cb_4_4_io_o_0_out[7] ,
    \cb_4_4_io_o_0_out[6] ,
    \cb_4_4_io_o_0_out[5] ,
    \cb_4_4_io_o_0_out[4] ,
    \cb_4_4_io_o_0_out[3] ,
    \cb_4_4_io_o_0_out[2] ,
    \cb_4_4_io_o_0_out[1] ,
    \cb_4_4_io_o_0_out[0] }),
    .io_i_1_in1({\cb_4_4_io_o_1_out[7] ,
    \cb_4_4_io_o_1_out[6] ,
    \cb_4_4_io_o_1_out[5] ,
    \cb_4_4_io_o_1_out[4] ,
    \cb_4_4_io_o_1_out[3] ,
    \cb_4_4_io_o_1_out[2] ,
    \cb_4_4_io_o_1_out[1] ,
    \cb_4_4_io_o_1_out[0] }),
    .io_i_2_in1({\cb_4_4_io_o_2_out[7] ,
    \cb_4_4_io_o_2_out[6] ,
    \cb_4_4_io_o_2_out[5] ,
    \cb_4_4_io_o_2_out[4] ,
    \cb_4_4_io_o_2_out[3] ,
    \cb_4_4_io_o_2_out[2] ,
    \cb_4_4_io_o_2_out[1] ,
    \cb_4_4_io_o_2_out[0] }),
    .io_i_3_in1({\cb_4_4_io_o_3_out[7] ,
    \cb_4_4_io_o_3_out[6] ,
    \cb_4_4_io_o_3_out[5] ,
    \cb_4_4_io_o_3_out[4] ,
    \cb_4_4_io_o_3_out[3] ,
    \cb_4_4_io_o_3_out[2] ,
    \cb_4_4_io_o_3_out[1] ,
    \cb_4_4_io_o_3_out[0] }),
    .io_i_4_in1({\cb_4_4_io_o_4_out[7] ,
    \cb_4_4_io_o_4_out[6] ,
    \cb_4_4_io_o_4_out[5] ,
    \cb_4_4_io_o_4_out[4] ,
    \cb_4_4_io_o_4_out[3] ,
    \cb_4_4_io_o_4_out[2] ,
    \cb_4_4_io_o_4_out[1] ,
    \cb_4_4_io_o_4_out[0] }),
    .io_i_5_in1({\cb_4_4_io_o_5_out[7] ,
    \cb_4_4_io_o_5_out[6] ,
    \cb_4_4_io_o_5_out[5] ,
    \cb_4_4_io_o_5_out[4] ,
    \cb_4_4_io_o_5_out[3] ,
    \cb_4_4_io_o_5_out[2] ,
    \cb_4_4_io_o_5_out[1] ,
    \cb_4_4_io_o_5_out[0] }),
    .io_i_6_in1({\cb_4_4_io_o_6_out[7] ,
    \cb_4_4_io_o_6_out[6] ,
    \cb_4_4_io_o_6_out[5] ,
    \cb_4_4_io_o_6_out[4] ,
    \cb_4_4_io_o_6_out[3] ,
    \cb_4_4_io_o_6_out[2] ,
    \cb_4_4_io_o_6_out[1] ,
    \cb_4_4_io_o_6_out[0] }),
    .io_i_7_in1({\cb_4_4_io_o_7_out[7] ,
    \cb_4_4_io_o_7_out[6] ,
    \cb_4_4_io_o_7_out[5] ,
    \cb_4_4_io_o_7_out[4] ,
    \cb_4_4_io_o_7_out[3] ,
    \cb_4_4_io_o_7_out[2] ,
    \cb_4_4_io_o_7_out[1] ,
    \cb_4_4_io_o_7_out[0] }),
    .io_o_0_out({\cb_4_5_io_o_0_out[7] ,
    \cb_4_5_io_o_0_out[6] ,
    \cb_4_5_io_o_0_out[5] ,
    \cb_4_5_io_o_0_out[4] ,
    \cb_4_5_io_o_0_out[3] ,
    \cb_4_5_io_o_0_out[2] ,
    \cb_4_5_io_o_0_out[1] ,
    \cb_4_5_io_o_0_out[0] }),
    .io_o_1_out({\cb_4_5_io_o_1_out[7] ,
    \cb_4_5_io_o_1_out[6] ,
    \cb_4_5_io_o_1_out[5] ,
    \cb_4_5_io_o_1_out[4] ,
    \cb_4_5_io_o_1_out[3] ,
    \cb_4_5_io_o_1_out[2] ,
    \cb_4_5_io_o_1_out[1] ,
    \cb_4_5_io_o_1_out[0] }),
    .io_o_2_out({\cb_4_5_io_o_2_out[7] ,
    \cb_4_5_io_o_2_out[6] ,
    \cb_4_5_io_o_2_out[5] ,
    \cb_4_5_io_o_2_out[4] ,
    \cb_4_5_io_o_2_out[3] ,
    \cb_4_5_io_o_2_out[2] ,
    \cb_4_5_io_o_2_out[1] ,
    \cb_4_5_io_o_2_out[0] }),
    .io_o_3_out({\cb_4_5_io_o_3_out[7] ,
    \cb_4_5_io_o_3_out[6] ,
    \cb_4_5_io_o_3_out[5] ,
    \cb_4_5_io_o_3_out[4] ,
    \cb_4_5_io_o_3_out[3] ,
    \cb_4_5_io_o_3_out[2] ,
    \cb_4_5_io_o_3_out[1] ,
    \cb_4_5_io_o_3_out[0] }),
    .io_o_4_out({\cb_4_5_io_o_4_out[7] ,
    \cb_4_5_io_o_4_out[6] ,
    \cb_4_5_io_o_4_out[5] ,
    \cb_4_5_io_o_4_out[4] ,
    \cb_4_5_io_o_4_out[3] ,
    \cb_4_5_io_o_4_out[2] ,
    \cb_4_5_io_o_4_out[1] ,
    \cb_4_5_io_o_4_out[0] }),
    .io_o_5_out({\cb_4_5_io_o_5_out[7] ,
    \cb_4_5_io_o_5_out[6] ,
    \cb_4_5_io_o_5_out[5] ,
    \cb_4_5_io_o_5_out[4] ,
    \cb_4_5_io_o_5_out[3] ,
    \cb_4_5_io_o_5_out[2] ,
    \cb_4_5_io_o_5_out[1] ,
    \cb_4_5_io_o_5_out[0] }),
    .io_o_6_out({\cb_4_5_io_o_6_out[7] ,
    \cb_4_5_io_o_6_out[6] ,
    \cb_4_5_io_o_6_out[5] ,
    \cb_4_5_io_o_6_out[4] ,
    \cb_4_5_io_o_6_out[3] ,
    \cb_4_5_io_o_6_out[2] ,
    \cb_4_5_io_o_6_out[1] ,
    \cb_4_5_io_o_6_out[0] }),
    .io_o_7_out({\cb_4_5_io_o_7_out[7] ,
    \cb_4_5_io_o_7_out[6] ,
    \cb_4_5_io_o_7_out[5] ,
    \cb_4_5_io_o_7_out[4] ,
    \cb_4_5_io_o_7_out[3] ,
    \cb_4_5_io_o_7_out[2] ,
    \cb_4_5_io_o_7_out[1] ,
    \cb_4_5_io_o_7_out[0] }),
    .io_wo({\cb_4_4_io_eo[63] ,
    \cb_4_4_io_eo[62] ,
    \cb_4_4_io_eo[61] ,
    \cb_4_4_io_eo[60] ,
    \cb_4_4_io_eo[59] ,
    \cb_4_4_io_eo[58] ,
    \cb_4_4_io_eo[57] ,
    \cb_4_4_io_eo[56] ,
    \cb_4_4_io_eo[55] ,
    \cb_4_4_io_eo[54] ,
    \cb_4_4_io_eo[53] ,
    \cb_4_4_io_eo[52] ,
    \cb_4_4_io_eo[51] ,
    \cb_4_4_io_eo[50] ,
    \cb_4_4_io_eo[49] ,
    \cb_4_4_io_eo[48] ,
    \cb_4_4_io_eo[47] ,
    \cb_4_4_io_eo[46] ,
    \cb_4_4_io_eo[45] ,
    \cb_4_4_io_eo[44] ,
    \cb_4_4_io_eo[43] ,
    \cb_4_4_io_eo[42] ,
    \cb_4_4_io_eo[41] ,
    \cb_4_4_io_eo[40] ,
    \cb_4_4_io_eo[39] ,
    \cb_4_4_io_eo[38] ,
    \cb_4_4_io_eo[37] ,
    \cb_4_4_io_eo[36] ,
    \cb_4_4_io_eo[35] ,
    \cb_4_4_io_eo[34] ,
    \cb_4_4_io_eo[33] ,
    \cb_4_4_io_eo[32] ,
    \cb_4_4_io_eo[31] ,
    \cb_4_4_io_eo[30] ,
    \cb_4_4_io_eo[29] ,
    \cb_4_4_io_eo[28] ,
    \cb_4_4_io_eo[27] ,
    \cb_4_4_io_eo[26] ,
    \cb_4_4_io_eo[25] ,
    \cb_4_4_io_eo[24] ,
    \cb_4_4_io_eo[23] ,
    \cb_4_4_io_eo[22] ,
    \cb_4_4_io_eo[21] ,
    \cb_4_4_io_eo[20] ,
    \cb_4_4_io_eo[19] ,
    \cb_4_4_io_eo[18] ,
    \cb_4_4_io_eo[17] ,
    \cb_4_4_io_eo[16] ,
    \cb_4_4_io_eo[15] ,
    \cb_4_4_io_eo[14] ,
    \cb_4_4_io_eo[13] ,
    \cb_4_4_io_eo[12] ,
    \cb_4_4_io_eo[11] ,
    \cb_4_4_io_eo[10] ,
    \cb_4_4_io_eo[9] ,
    \cb_4_4_io_eo[8] ,
    \cb_4_4_io_eo[7] ,
    \cb_4_4_io_eo[6] ,
    \cb_4_4_io_eo[5] ,
    \cb_4_4_io_eo[4] ,
    \cb_4_4_io_eo[3] ,
    \cb_4_4_io_eo[2] ,
    \cb_4_4_io_eo[1] ,
    \cb_4_4_io_eo[0] }));
 cic_block cb_4_6 (.io_cs_i(cb_4_6_io_cs_i),
    .io_i_0_ci(cb_4_5_io_o_0_co),
    .io_i_1_ci(cb_4_5_io_o_1_co),
    .io_i_2_ci(cb_4_5_io_o_2_co),
    .io_i_3_ci(cb_4_5_io_o_3_co),
    .io_i_4_ci(cb_4_5_io_o_4_co),
    .io_i_5_ci(cb_4_5_io_o_5_co),
    .io_i_6_ci(cb_4_5_io_o_6_co),
    .io_i_7_ci(cb_4_5_io_o_7_co),
    .io_o_0_co(cb_4_6_io_o_0_co),
    .io_o_1_co(cb_4_6_io_o_1_co),
    .io_o_2_co(cb_4_6_io_o_2_co),
    .io_o_3_co(cb_4_6_io_o_3_co),
    .io_o_4_co(cb_4_6_io_o_4_co),
    .io_o_5_co(cb_4_6_io_o_5_co),
    .io_o_6_co(cb_4_6_io_o_6_co),
    .io_o_7_co(cb_4_6_io_o_7_co),
    .io_vci(cb_4_5_io_vco),
    .io_vco(cb_4_6_io_vco),
    .io_vi(cb_4_6_io_vi),
    .io_we_i(cb_4_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_4_0_io_adr_i[1] ,
    \cb_4_0_io_adr_i[0] }),
    .io_dat_i({\cb_4_0_io_dat_i[15] ,
    \cb_4_0_io_dat_i[14] ,
    \cb_4_0_io_dat_i[13] ,
    \cb_4_0_io_dat_i[12] ,
    \cb_4_0_io_dat_i[11] ,
    \cb_4_0_io_dat_i[10] ,
    \cb_4_0_io_dat_i[9] ,
    \cb_4_0_io_dat_i[8] ,
    \cb_4_0_io_dat_i[7] ,
    \cb_4_0_io_dat_i[6] ,
    \cb_4_0_io_dat_i[5] ,
    \cb_4_0_io_dat_i[4] ,
    \cb_4_0_io_dat_i[3] ,
    \cb_4_0_io_dat_i[2] ,
    \cb_4_0_io_dat_i[1] ,
    \cb_4_0_io_dat_i[0] }),
    .io_dat_o({\cb_4_6_io_dat_o[15] ,
    \cb_4_6_io_dat_o[14] ,
    \cb_4_6_io_dat_o[13] ,
    \cb_4_6_io_dat_o[12] ,
    \cb_4_6_io_dat_o[11] ,
    \cb_4_6_io_dat_o[10] ,
    \cb_4_6_io_dat_o[9] ,
    \cb_4_6_io_dat_o[8] ,
    \cb_4_6_io_dat_o[7] ,
    \cb_4_6_io_dat_o[6] ,
    \cb_4_6_io_dat_o[5] ,
    \cb_4_6_io_dat_o[4] ,
    \cb_4_6_io_dat_o[3] ,
    \cb_4_6_io_dat_o[2] ,
    \cb_4_6_io_dat_o[1] ,
    \cb_4_6_io_dat_o[0] }),
    .io_eo({\cb_4_6_io_eo[63] ,
    \cb_4_6_io_eo[62] ,
    \cb_4_6_io_eo[61] ,
    \cb_4_6_io_eo[60] ,
    \cb_4_6_io_eo[59] ,
    \cb_4_6_io_eo[58] ,
    \cb_4_6_io_eo[57] ,
    \cb_4_6_io_eo[56] ,
    \cb_4_6_io_eo[55] ,
    \cb_4_6_io_eo[54] ,
    \cb_4_6_io_eo[53] ,
    \cb_4_6_io_eo[52] ,
    \cb_4_6_io_eo[51] ,
    \cb_4_6_io_eo[50] ,
    \cb_4_6_io_eo[49] ,
    \cb_4_6_io_eo[48] ,
    \cb_4_6_io_eo[47] ,
    \cb_4_6_io_eo[46] ,
    \cb_4_6_io_eo[45] ,
    \cb_4_6_io_eo[44] ,
    \cb_4_6_io_eo[43] ,
    \cb_4_6_io_eo[42] ,
    \cb_4_6_io_eo[41] ,
    \cb_4_6_io_eo[40] ,
    \cb_4_6_io_eo[39] ,
    \cb_4_6_io_eo[38] ,
    \cb_4_6_io_eo[37] ,
    \cb_4_6_io_eo[36] ,
    \cb_4_6_io_eo[35] ,
    \cb_4_6_io_eo[34] ,
    \cb_4_6_io_eo[33] ,
    \cb_4_6_io_eo[32] ,
    \cb_4_6_io_eo[31] ,
    \cb_4_6_io_eo[30] ,
    \cb_4_6_io_eo[29] ,
    \cb_4_6_io_eo[28] ,
    \cb_4_6_io_eo[27] ,
    \cb_4_6_io_eo[26] ,
    \cb_4_6_io_eo[25] ,
    \cb_4_6_io_eo[24] ,
    \cb_4_6_io_eo[23] ,
    \cb_4_6_io_eo[22] ,
    \cb_4_6_io_eo[21] ,
    \cb_4_6_io_eo[20] ,
    \cb_4_6_io_eo[19] ,
    \cb_4_6_io_eo[18] ,
    \cb_4_6_io_eo[17] ,
    \cb_4_6_io_eo[16] ,
    \cb_4_6_io_eo[15] ,
    \cb_4_6_io_eo[14] ,
    \cb_4_6_io_eo[13] ,
    \cb_4_6_io_eo[12] ,
    \cb_4_6_io_eo[11] ,
    \cb_4_6_io_eo[10] ,
    \cb_4_6_io_eo[9] ,
    \cb_4_6_io_eo[8] ,
    \cb_4_6_io_eo[7] ,
    \cb_4_6_io_eo[6] ,
    \cb_4_6_io_eo[5] ,
    \cb_4_6_io_eo[4] ,
    \cb_4_6_io_eo[3] ,
    \cb_4_6_io_eo[2] ,
    \cb_4_6_io_eo[1] ,
    \cb_4_6_io_eo[0] }),
    .io_i_0_in1({\cb_4_5_io_o_0_out[7] ,
    \cb_4_5_io_o_0_out[6] ,
    \cb_4_5_io_o_0_out[5] ,
    \cb_4_5_io_o_0_out[4] ,
    \cb_4_5_io_o_0_out[3] ,
    \cb_4_5_io_o_0_out[2] ,
    \cb_4_5_io_o_0_out[1] ,
    \cb_4_5_io_o_0_out[0] }),
    .io_i_1_in1({\cb_4_5_io_o_1_out[7] ,
    \cb_4_5_io_o_1_out[6] ,
    \cb_4_5_io_o_1_out[5] ,
    \cb_4_5_io_o_1_out[4] ,
    \cb_4_5_io_o_1_out[3] ,
    \cb_4_5_io_o_1_out[2] ,
    \cb_4_5_io_o_1_out[1] ,
    \cb_4_5_io_o_1_out[0] }),
    .io_i_2_in1({\cb_4_5_io_o_2_out[7] ,
    \cb_4_5_io_o_2_out[6] ,
    \cb_4_5_io_o_2_out[5] ,
    \cb_4_5_io_o_2_out[4] ,
    \cb_4_5_io_o_2_out[3] ,
    \cb_4_5_io_o_2_out[2] ,
    \cb_4_5_io_o_2_out[1] ,
    \cb_4_5_io_o_2_out[0] }),
    .io_i_3_in1({\cb_4_5_io_o_3_out[7] ,
    \cb_4_5_io_o_3_out[6] ,
    \cb_4_5_io_o_3_out[5] ,
    \cb_4_5_io_o_3_out[4] ,
    \cb_4_5_io_o_3_out[3] ,
    \cb_4_5_io_o_3_out[2] ,
    \cb_4_5_io_o_3_out[1] ,
    \cb_4_5_io_o_3_out[0] }),
    .io_i_4_in1({\cb_4_5_io_o_4_out[7] ,
    \cb_4_5_io_o_4_out[6] ,
    \cb_4_5_io_o_4_out[5] ,
    \cb_4_5_io_o_4_out[4] ,
    \cb_4_5_io_o_4_out[3] ,
    \cb_4_5_io_o_4_out[2] ,
    \cb_4_5_io_o_4_out[1] ,
    \cb_4_5_io_o_4_out[0] }),
    .io_i_5_in1({\cb_4_5_io_o_5_out[7] ,
    \cb_4_5_io_o_5_out[6] ,
    \cb_4_5_io_o_5_out[5] ,
    \cb_4_5_io_o_5_out[4] ,
    \cb_4_5_io_o_5_out[3] ,
    \cb_4_5_io_o_5_out[2] ,
    \cb_4_5_io_o_5_out[1] ,
    \cb_4_5_io_o_5_out[0] }),
    .io_i_6_in1({\cb_4_5_io_o_6_out[7] ,
    \cb_4_5_io_o_6_out[6] ,
    \cb_4_5_io_o_6_out[5] ,
    \cb_4_5_io_o_6_out[4] ,
    \cb_4_5_io_o_6_out[3] ,
    \cb_4_5_io_o_6_out[2] ,
    \cb_4_5_io_o_6_out[1] ,
    \cb_4_5_io_o_6_out[0] }),
    .io_i_7_in1({\cb_4_5_io_o_7_out[7] ,
    \cb_4_5_io_o_7_out[6] ,
    \cb_4_5_io_o_7_out[5] ,
    \cb_4_5_io_o_7_out[4] ,
    \cb_4_5_io_o_7_out[3] ,
    \cb_4_5_io_o_7_out[2] ,
    \cb_4_5_io_o_7_out[1] ,
    \cb_4_5_io_o_7_out[0] }),
    .io_o_0_out({\cb_4_6_io_o_0_out[7] ,
    \cb_4_6_io_o_0_out[6] ,
    \cb_4_6_io_o_0_out[5] ,
    \cb_4_6_io_o_0_out[4] ,
    \cb_4_6_io_o_0_out[3] ,
    \cb_4_6_io_o_0_out[2] ,
    \cb_4_6_io_o_0_out[1] ,
    \cb_4_6_io_o_0_out[0] }),
    .io_o_1_out({\cb_4_6_io_o_1_out[7] ,
    \cb_4_6_io_o_1_out[6] ,
    \cb_4_6_io_o_1_out[5] ,
    \cb_4_6_io_o_1_out[4] ,
    \cb_4_6_io_o_1_out[3] ,
    \cb_4_6_io_o_1_out[2] ,
    \cb_4_6_io_o_1_out[1] ,
    \cb_4_6_io_o_1_out[0] }),
    .io_o_2_out({\cb_4_6_io_o_2_out[7] ,
    \cb_4_6_io_o_2_out[6] ,
    \cb_4_6_io_o_2_out[5] ,
    \cb_4_6_io_o_2_out[4] ,
    \cb_4_6_io_o_2_out[3] ,
    \cb_4_6_io_o_2_out[2] ,
    \cb_4_6_io_o_2_out[1] ,
    \cb_4_6_io_o_2_out[0] }),
    .io_o_3_out({\cb_4_6_io_o_3_out[7] ,
    \cb_4_6_io_o_3_out[6] ,
    \cb_4_6_io_o_3_out[5] ,
    \cb_4_6_io_o_3_out[4] ,
    \cb_4_6_io_o_3_out[3] ,
    \cb_4_6_io_o_3_out[2] ,
    \cb_4_6_io_o_3_out[1] ,
    \cb_4_6_io_o_3_out[0] }),
    .io_o_4_out({\cb_4_6_io_o_4_out[7] ,
    \cb_4_6_io_o_4_out[6] ,
    \cb_4_6_io_o_4_out[5] ,
    \cb_4_6_io_o_4_out[4] ,
    \cb_4_6_io_o_4_out[3] ,
    \cb_4_6_io_o_4_out[2] ,
    \cb_4_6_io_o_4_out[1] ,
    \cb_4_6_io_o_4_out[0] }),
    .io_o_5_out({\cb_4_6_io_o_5_out[7] ,
    \cb_4_6_io_o_5_out[6] ,
    \cb_4_6_io_o_5_out[5] ,
    \cb_4_6_io_o_5_out[4] ,
    \cb_4_6_io_o_5_out[3] ,
    \cb_4_6_io_o_5_out[2] ,
    \cb_4_6_io_o_5_out[1] ,
    \cb_4_6_io_o_5_out[0] }),
    .io_o_6_out({\cb_4_6_io_o_6_out[7] ,
    \cb_4_6_io_o_6_out[6] ,
    \cb_4_6_io_o_6_out[5] ,
    \cb_4_6_io_o_6_out[4] ,
    \cb_4_6_io_o_6_out[3] ,
    \cb_4_6_io_o_6_out[2] ,
    \cb_4_6_io_o_6_out[1] ,
    \cb_4_6_io_o_6_out[0] }),
    .io_o_7_out({\cb_4_6_io_o_7_out[7] ,
    \cb_4_6_io_o_7_out[6] ,
    \cb_4_6_io_o_7_out[5] ,
    \cb_4_6_io_o_7_out[4] ,
    \cb_4_6_io_o_7_out[3] ,
    \cb_4_6_io_o_7_out[2] ,
    \cb_4_6_io_o_7_out[1] ,
    \cb_4_6_io_o_7_out[0] }),
    .io_wo({\cb_4_5_io_eo[63] ,
    \cb_4_5_io_eo[62] ,
    \cb_4_5_io_eo[61] ,
    \cb_4_5_io_eo[60] ,
    \cb_4_5_io_eo[59] ,
    \cb_4_5_io_eo[58] ,
    \cb_4_5_io_eo[57] ,
    \cb_4_5_io_eo[56] ,
    \cb_4_5_io_eo[55] ,
    \cb_4_5_io_eo[54] ,
    \cb_4_5_io_eo[53] ,
    \cb_4_5_io_eo[52] ,
    \cb_4_5_io_eo[51] ,
    \cb_4_5_io_eo[50] ,
    \cb_4_5_io_eo[49] ,
    \cb_4_5_io_eo[48] ,
    \cb_4_5_io_eo[47] ,
    \cb_4_5_io_eo[46] ,
    \cb_4_5_io_eo[45] ,
    \cb_4_5_io_eo[44] ,
    \cb_4_5_io_eo[43] ,
    \cb_4_5_io_eo[42] ,
    \cb_4_5_io_eo[41] ,
    \cb_4_5_io_eo[40] ,
    \cb_4_5_io_eo[39] ,
    \cb_4_5_io_eo[38] ,
    \cb_4_5_io_eo[37] ,
    \cb_4_5_io_eo[36] ,
    \cb_4_5_io_eo[35] ,
    \cb_4_5_io_eo[34] ,
    \cb_4_5_io_eo[33] ,
    \cb_4_5_io_eo[32] ,
    \cb_4_5_io_eo[31] ,
    \cb_4_5_io_eo[30] ,
    \cb_4_5_io_eo[29] ,
    \cb_4_5_io_eo[28] ,
    \cb_4_5_io_eo[27] ,
    \cb_4_5_io_eo[26] ,
    \cb_4_5_io_eo[25] ,
    \cb_4_5_io_eo[24] ,
    \cb_4_5_io_eo[23] ,
    \cb_4_5_io_eo[22] ,
    \cb_4_5_io_eo[21] ,
    \cb_4_5_io_eo[20] ,
    \cb_4_5_io_eo[19] ,
    \cb_4_5_io_eo[18] ,
    \cb_4_5_io_eo[17] ,
    \cb_4_5_io_eo[16] ,
    \cb_4_5_io_eo[15] ,
    \cb_4_5_io_eo[14] ,
    \cb_4_5_io_eo[13] ,
    \cb_4_5_io_eo[12] ,
    \cb_4_5_io_eo[11] ,
    \cb_4_5_io_eo[10] ,
    \cb_4_5_io_eo[9] ,
    \cb_4_5_io_eo[8] ,
    \cb_4_5_io_eo[7] ,
    \cb_4_5_io_eo[6] ,
    \cb_4_5_io_eo[5] ,
    \cb_4_5_io_eo[4] ,
    \cb_4_5_io_eo[3] ,
    \cb_4_5_io_eo[2] ,
    \cb_4_5_io_eo[1] ,
    \cb_4_5_io_eo[0] }));
 cic_block cb_4_7 (.io_cs_i(cb_4_7_io_cs_i),
    .io_i_0_ci(cb_4_6_io_o_0_co),
    .io_i_1_ci(cb_4_6_io_o_1_co),
    .io_i_2_ci(cb_4_6_io_o_2_co),
    .io_i_3_ci(cb_4_6_io_o_3_co),
    .io_i_4_ci(cb_4_6_io_o_4_co),
    .io_i_5_ci(cb_4_6_io_o_5_co),
    .io_i_6_ci(cb_4_6_io_o_6_co),
    .io_i_7_ci(cb_4_6_io_o_7_co),
    .io_o_0_co(cb_4_7_io_o_0_co),
    .io_o_1_co(cb_4_7_io_o_1_co),
    .io_o_2_co(cb_4_7_io_o_2_co),
    .io_o_3_co(cb_4_7_io_o_3_co),
    .io_o_4_co(cb_4_7_io_o_4_co),
    .io_o_5_co(cb_4_7_io_o_5_co),
    .io_o_6_co(cb_4_7_io_o_6_co),
    .io_o_7_co(cb_4_7_io_o_7_co),
    .io_vci(cb_4_6_io_vco),
    .io_vco(cb_4_7_io_vco),
    .io_vi(cb_4_7_io_vi),
    .io_we_i(cb_4_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_4_0_io_adr_i[1] ,
    \cb_4_0_io_adr_i[0] }),
    .io_dat_i({\cb_4_0_io_dat_i[15] ,
    \cb_4_0_io_dat_i[14] ,
    \cb_4_0_io_dat_i[13] ,
    \cb_4_0_io_dat_i[12] ,
    \cb_4_0_io_dat_i[11] ,
    \cb_4_0_io_dat_i[10] ,
    \cb_4_0_io_dat_i[9] ,
    \cb_4_0_io_dat_i[8] ,
    \cb_4_0_io_dat_i[7] ,
    \cb_4_0_io_dat_i[6] ,
    \cb_4_0_io_dat_i[5] ,
    \cb_4_0_io_dat_i[4] ,
    \cb_4_0_io_dat_i[3] ,
    \cb_4_0_io_dat_i[2] ,
    \cb_4_0_io_dat_i[1] ,
    \cb_4_0_io_dat_i[0] }),
    .io_dat_o({\cb_4_7_io_dat_o[15] ,
    \cb_4_7_io_dat_o[14] ,
    \cb_4_7_io_dat_o[13] ,
    \cb_4_7_io_dat_o[12] ,
    \cb_4_7_io_dat_o[11] ,
    \cb_4_7_io_dat_o[10] ,
    \cb_4_7_io_dat_o[9] ,
    \cb_4_7_io_dat_o[8] ,
    \cb_4_7_io_dat_o[7] ,
    \cb_4_7_io_dat_o[6] ,
    \cb_4_7_io_dat_o[5] ,
    \cb_4_7_io_dat_o[4] ,
    \cb_4_7_io_dat_o[3] ,
    \cb_4_7_io_dat_o[2] ,
    \cb_4_7_io_dat_o[1] ,
    \cb_4_7_io_dat_o[0] }),
    .io_eo({\cb_4_7_io_eo[63] ,
    \cb_4_7_io_eo[62] ,
    \cb_4_7_io_eo[61] ,
    \cb_4_7_io_eo[60] ,
    \cb_4_7_io_eo[59] ,
    \cb_4_7_io_eo[58] ,
    \cb_4_7_io_eo[57] ,
    \cb_4_7_io_eo[56] ,
    \cb_4_7_io_eo[55] ,
    \cb_4_7_io_eo[54] ,
    \cb_4_7_io_eo[53] ,
    \cb_4_7_io_eo[52] ,
    \cb_4_7_io_eo[51] ,
    \cb_4_7_io_eo[50] ,
    \cb_4_7_io_eo[49] ,
    \cb_4_7_io_eo[48] ,
    \cb_4_7_io_eo[47] ,
    \cb_4_7_io_eo[46] ,
    \cb_4_7_io_eo[45] ,
    \cb_4_7_io_eo[44] ,
    \cb_4_7_io_eo[43] ,
    \cb_4_7_io_eo[42] ,
    \cb_4_7_io_eo[41] ,
    \cb_4_7_io_eo[40] ,
    \cb_4_7_io_eo[39] ,
    \cb_4_7_io_eo[38] ,
    \cb_4_7_io_eo[37] ,
    \cb_4_7_io_eo[36] ,
    \cb_4_7_io_eo[35] ,
    \cb_4_7_io_eo[34] ,
    \cb_4_7_io_eo[33] ,
    \cb_4_7_io_eo[32] ,
    \cb_4_7_io_eo[31] ,
    \cb_4_7_io_eo[30] ,
    \cb_4_7_io_eo[29] ,
    \cb_4_7_io_eo[28] ,
    \cb_4_7_io_eo[27] ,
    \cb_4_7_io_eo[26] ,
    \cb_4_7_io_eo[25] ,
    \cb_4_7_io_eo[24] ,
    \cb_4_7_io_eo[23] ,
    \cb_4_7_io_eo[22] ,
    \cb_4_7_io_eo[21] ,
    \cb_4_7_io_eo[20] ,
    \cb_4_7_io_eo[19] ,
    \cb_4_7_io_eo[18] ,
    \cb_4_7_io_eo[17] ,
    \cb_4_7_io_eo[16] ,
    \cb_4_7_io_eo[15] ,
    \cb_4_7_io_eo[14] ,
    \cb_4_7_io_eo[13] ,
    \cb_4_7_io_eo[12] ,
    \cb_4_7_io_eo[11] ,
    \cb_4_7_io_eo[10] ,
    \cb_4_7_io_eo[9] ,
    \cb_4_7_io_eo[8] ,
    \cb_4_7_io_eo[7] ,
    \cb_4_7_io_eo[6] ,
    \cb_4_7_io_eo[5] ,
    \cb_4_7_io_eo[4] ,
    \cb_4_7_io_eo[3] ,
    \cb_4_7_io_eo[2] ,
    \cb_4_7_io_eo[1] ,
    \cb_4_7_io_eo[0] }),
    .io_i_0_in1({\cb_4_6_io_o_0_out[7] ,
    \cb_4_6_io_o_0_out[6] ,
    \cb_4_6_io_o_0_out[5] ,
    \cb_4_6_io_o_0_out[4] ,
    \cb_4_6_io_o_0_out[3] ,
    \cb_4_6_io_o_0_out[2] ,
    \cb_4_6_io_o_0_out[1] ,
    \cb_4_6_io_o_0_out[0] }),
    .io_i_1_in1({\cb_4_6_io_o_1_out[7] ,
    \cb_4_6_io_o_1_out[6] ,
    \cb_4_6_io_o_1_out[5] ,
    \cb_4_6_io_o_1_out[4] ,
    \cb_4_6_io_o_1_out[3] ,
    \cb_4_6_io_o_1_out[2] ,
    \cb_4_6_io_o_1_out[1] ,
    \cb_4_6_io_o_1_out[0] }),
    .io_i_2_in1({\cb_4_6_io_o_2_out[7] ,
    \cb_4_6_io_o_2_out[6] ,
    \cb_4_6_io_o_2_out[5] ,
    \cb_4_6_io_o_2_out[4] ,
    \cb_4_6_io_o_2_out[3] ,
    \cb_4_6_io_o_2_out[2] ,
    \cb_4_6_io_o_2_out[1] ,
    \cb_4_6_io_o_2_out[0] }),
    .io_i_3_in1({\cb_4_6_io_o_3_out[7] ,
    \cb_4_6_io_o_3_out[6] ,
    \cb_4_6_io_o_3_out[5] ,
    \cb_4_6_io_o_3_out[4] ,
    \cb_4_6_io_o_3_out[3] ,
    \cb_4_6_io_o_3_out[2] ,
    \cb_4_6_io_o_3_out[1] ,
    \cb_4_6_io_o_3_out[0] }),
    .io_i_4_in1({\cb_4_6_io_o_4_out[7] ,
    \cb_4_6_io_o_4_out[6] ,
    \cb_4_6_io_o_4_out[5] ,
    \cb_4_6_io_o_4_out[4] ,
    \cb_4_6_io_o_4_out[3] ,
    \cb_4_6_io_o_4_out[2] ,
    \cb_4_6_io_o_4_out[1] ,
    \cb_4_6_io_o_4_out[0] }),
    .io_i_5_in1({\cb_4_6_io_o_5_out[7] ,
    \cb_4_6_io_o_5_out[6] ,
    \cb_4_6_io_o_5_out[5] ,
    \cb_4_6_io_o_5_out[4] ,
    \cb_4_6_io_o_5_out[3] ,
    \cb_4_6_io_o_5_out[2] ,
    \cb_4_6_io_o_5_out[1] ,
    \cb_4_6_io_o_5_out[0] }),
    .io_i_6_in1({\cb_4_6_io_o_6_out[7] ,
    \cb_4_6_io_o_6_out[6] ,
    \cb_4_6_io_o_6_out[5] ,
    \cb_4_6_io_o_6_out[4] ,
    \cb_4_6_io_o_6_out[3] ,
    \cb_4_6_io_o_6_out[2] ,
    \cb_4_6_io_o_6_out[1] ,
    \cb_4_6_io_o_6_out[0] }),
    .io_i_7_in1({\cb_4_6_io_o_7_out[7] ,
    \cb_4_6_io_o_7_out[6] ,
    \cb_4_6_io_o_7_out[5] ,
    \cb_4_6_io_o_7_out[4] ,
    \cb_4_6_io_o_7_out[3] ,
    \cb_4_6_io_o_7_out[2] ,
    \cb_4_6_io_o_7_out[1] ,
    \cb_4_6_io_o_7_out[0] }),
    .io_o_0_out({\cb_4_7_io_o_0_out[7] ,
    \cb_4_7_io_o_0_out[6] ,
    \cb_4_7_io_o_0_out[5] ,
    \cb_4_7_io_o_0_out[4] ,
    \cb_4_7_io_o_0_out[3] ,
    \cb_4_7_io_o_0_out[2] ,
    \cb_4_7_io_o_0_out[1] ,
    \cb_4_7_io_o_0_out[0] }),
    .io_o_1_out({\cb_4_7_io_o_1_out[7] ,
    \cb_4_7_io_o_1_out[6] ,
    \cb_4_7_io_o_1_out[5] ,
    \cb_4_7_io_o_1_out[4] ,
    \cb_4_7_io_o_1_out[3] ,
    \cb_4_7_io_o_1_out[2] ,
    \cb_4_7_io_o_1_out[1] ,
    \cb_4_7_io_o_1_out[0] }),
    .io_o_2_out({\cb_4_7_io_o_2_out[7] ,
    \cb_4_7_io_o_2_out[6] ,
    \cb_4_7_io_o_2_out[5] ,
    \cb_4_7_io_o_2_out[4] ,
    \cb_4_7_io_o_2_out[3] ,
    \cb_4_7_io_o_2_out[2] ,
    \cb_4_7_io_o_2_out[1] ,
    \cb_4_7_io_o_2_out[0] }),
    .io_o_3_out({\cb_4_7_io_o_3_out[7] ,
    \cb_4_7_io_o_3_out[6] ,
    \cb_4_7_io_o_3_out[5] ,
    \cb_4_7_io_o_3_out[4] ,
    \cb_4_7_io_o_3_out[3] ,
    \cb_4_7_io_o_3_out[2] ,
    \cb_4_7_io_o_3_out[1] ,
    \cb_4_7_io_o_3_out[0] }),
    .io_o_4_out({\cb_4_7_io_o_4_out[7] ,
    \cb_4_7_io_o_4_out[6] ,
    \cb_4_7_io_o_4_out[5] ,
    \cb_4_7_io_o_4_out[4] ,
    \cb_4_7_io_o_4_out[3] ,
    \cb_4_7_io_o_4_out[2] ,
    \cb_4_7_io_o_4_out[1] ,
    \cb_4_7_io_o_4_out[0] }),
    .io_o_5_out({\cb_4_7_io_o_5_out[7] ,
    \cb_4_7_io_o_5_out[6] ,
    \cb_4_7_io_o_5_out[5] ,
    \cb_4_7_io_o_5_out[4] ,
    \cb_4_7_io_o_5_out[3] ,
    \cb_4_7_io_o_5_out[2] ,
    \cb_4_7_io_o_5_out[1] ,
    \cb_4_7_io_o_5_out[0] }),
    .io_o_6_out({\cb_4_7_io_o_6_out[7] ,
    \cb_4_7_io_o_6_out[6] ,
    \cb_4_7_io_o_6_out[5] ,
    \cb_4_7_io_o_6_out[4] ,
    \cb_4_7_io_o_6_out[3] ,
    \cb_4_7_io_o_6_out[2] ,
    \cb_4_7_io_o_6_out[1] ,
    \cb_4_7_io_o_6_out[0] }),
    .io_o_7_out({\cb_4_7_io_o_7_out[7] ,
    \cb_4_7_io_o_7_out[6] ,
    \cb_4_7_io_o_7_out[5] ,
    \cb_4_7_io_o_7_out[4] ,
    \cb_4_7_io_o_7_out[3] ,
    \cb_4_7_io_o_7_out[2] ,
    \cb_4_7_io_o_7_out[1] ,
    \cb_4_7_io_o_7_out[0] }),
    .io_wo({\cb_4_6_io_eo[63] ,
    \cb_4_6_io_eo[62] ,
    \cb_4_6_io_eo[61] ,
    \cb_4_6_io_eo[60] ,
    \cb_4_6_io_eo[59] ,
    \cb_4_6_io_eo[58] ,
    \cb_4_6_io_eo[57] ,
    \cb_4_6_io_eo[56] ,
    \cb_4_6_io_eo[55] ,
    \cb_4_6_io_eo[54] ,
    \cb_4_6_io_eo[53] ,
    \cb_4_6_io_eo[52] ,
    \cb_4_6_io_eo[51] ,
    \cb_4_6_io_eo[50] ,
    \cb_4_6_io_eo[49] ,
    \cb_4_6_io_eo[48] ,
    \cb_4_6_io_eo[47] ,
    \cb_4_6_io_eo[46] ,
    \cb_4_6_io_eo[45] ,
    \cb_4_6_io_eo[44] ,
    \cb_4_6_io_eo[43] ,
    \cb_4_6_io_eo[42] ,
    \cb_4_6_io_eo[41] ,
    \cb_4_6_io_eo[40] ,
    \cb_4_6_io_eo[39] ,
    \cb_4_6_io_eo[38] ,
    \cb_4_6_io_eo[37] ,
    \cb_4_6_io_eo[36] ,
    \cb_4_6_io_eo[35] ,
    \cb_4_6_io_eo[34] ,
    \cb_4_6_io_eo[33] ,
    \cb_4_6_io_eo[32] ,
    \cb_4_6_io_eo[31] ,
    \cb_4_6_io_eo[30] ,
    \cb_4_6_io_eo[29] ,
    \cb_4_6_io_eo[28] ,
    \cb_4_6_io_eo[27] ,
    \cb_4_6_io_eo[26] ,
    \cb_4_6_io_eo[25] ,
    \cb_4_6_io_eo[24] ,
    \cb_4_6_io_eo[23] ,
    \cb_4_6_io_eo[22] ,
    \cb_4_6_io_eo[21] ,
    \cb_4_6_io_eo[20] ,
    \cb_4_6_io_eo[19] ,
    \cb_4_6_io_eo[18] ,
    \cb_4_6_io_eo[17] ,
    \cb_4_6_io_eo[16] ,
    \cb_4_6_io_eo[15] ,
    \cb_4_6_io_eo[14] ,
    \cb_4_6_io_eo[13] ,
    \cb_4_6_io_eo[12] ,
    \cb_4_6_io_eo[11] ,
    \cb_4_6_io_eo[10] ,
    \cb_4_6_io_eo[9] ,
    \cb_4_6_io_eo[8] ,
    \cb_4_6_io_eo[7] ,
    \cb_4_6_io_eo[6] ,
    \cb_4_6_io_eo[5] ,
    \cb_4_6_io_eo[4] ,
    \cb_4_6_io_eo[3] ,
    \cb_4_6_io_eo[2] ,
    \cb_4_6_io_eo[1] ,
    \cb_4_6_io_eo[0] }));
 cic_block cb_4_8 (.io_cs_i(cb_4_8_io_cs_i),
    .io_i_0_ci(cb_4_7_io_o_0_co),
    .io_i_1_ci(cb_4_7_io_o_1_co),
    .io_i_2_ci(cb_4_7_io_o_2_co),
    .io_i_3_ci(cb_4_7_io_o_3_co),
    .io_i_4_ci(cb_4_7_io_o_4_co),
    .io_i_5_ci(cb_4_7_io_o_5_co),
    .io_i_6_ci(cb_4_7_io_o_6_co),
    .io_i_7_ci(cb_4_7_io_o_7_co),
    .io_o_0_co(cb_4_8_io_o_0_co),
    .io_o_1_co(cb_4_8_io_o_1_co),
    .io_o_2_co(cb_4_8_io_o_2_co),
    .io_o_3_co(cb_4_8_io_o_3_co),
    .io_o_4_co(cb_4_8_io_o_4_co),
    .io_o_5_co(cb_4_8_io_o_5_co),
    .io_o_6_co(cb_4_8_io_o_6_co),
    .io_o_7_co(cb_4_8_io_o_7_co),
    .io_vci(cb_4_7_io_vco),
    .io_vco(cb_4_8_io_vco),
    .io_vi(cb_4_8_io_vi),
    .io_we_i(cb_4_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_4_0_io_adr_i[1] ,
    \cb_4_0_io_adr_i[0] }),
    .io_dat_i({\cb_4_0_io_dat_i[15] ,
    \cb_4_0_io_dat_i[14] ,
    \cb_4_0_io_dat_i[13] ,
    \cb_4_0_io_dat_i[12] ,
    \cb_4_0_io_dat_i[11] ,
    \cb_4_0_io_dat_i[10] ,
    \cb_4_0_io_dat_i[9] ,
    \cb_4_0_io_dat_i[8] ,
    \cb_4_0_io_dat_i[7] ,
    \cb_4_0_io_dat_i[6] ,
    \cb_4_0_io_dat_i[5] ,
    \cb_4_0_io_dat_i[4] ,
    \cb_4_0_io_dat_i[3] ,
    \cb_4_0_io_dat_i[2] ,
    \cb_4_0_io_dat_i[1] ,
    \cb_4_0_io_dat_i[0] }),
    .io_dat_o({\cb_4_8_io_dat_o[15] ,
    \cb_4_8_io_dat_o[14] ,
    \cb_4_8_io_dat_o[13] ,
    \cb_4_8_io_dat_o[12] ,
    \cb_4_8_io_dat_o[11] ,
    \cb_4_8_io_dat_o[10] ,
    \cb_4_8_io_dat_o[9] ,
    \cb_4_8_io_dat_o[8] ,
    \cb_4_8_io_dat_o[7] ,
    \cb_4_8_io_dat_o[6] ,
    \cb_4_8_io_dat_o[5] ,
    \cb_4_8_io_dat_o[4] ,
    \cb_4_8_io_dat_o[3] ,
    \cb_4_8_io_dat_o[2] ,
    \cb_4_8_io_dat_o[1] ,
    \cb_4_8_io_dat_o[0] }),
    .io_eo({\cb_4_8_io_eo[63] ,
    \cb_4_8_io_eo[62] ,
    \cb_4_8_io_eo[61] ,
    \cb_4_8_io_eo[60] ,
    \cb_4_8_io_eo[59] ,
    \cb_4_8_io_eo[58] ,
    \cb_4_8_io_eo[57] ,
    \cb_4_8_io_eo[56] ,
    \cb_4_8_io_eo[55] ,
    \cb_4_8_io_eo[54] ,
    \cb_4_8_io_eo[53] ,
    \cb_4_8_io_eo[52] ,
    \cb_4_8_io_eo[51] ,
    \cb_4_8_io_eo[50] ,
    \cb_4_8_io_eo[49] ,
    \cb_4_8_io_eo[48] ,
    \cb_4_8_io_eo[47] ,
    \cb_4_8_io_eo[46] ,
    \cb_4_8_io_eo[45] ,
    \cb_4_8_io_eo[44] ,
    \cb_4_8_io_eo[43] ,
    \cb_4_8_io_eo[42] ,
    \cb_4_8_io_eo[41] ,
    \cb_4_8_io_eo[40] ,
    \cb_4_8_io_eo[39] ,
    \cb_4_8_io_eo[38] ,
    \cb_4_8_io_eo[37] ,
    \cb_4_8_io_eo[36] ,
    \cb_4_8_io_eo[35] ,
    \cb_4_8_io_eo[34] ,
    \cb_4_8_io_eo[33] ,
    \cb_4_8_io_eo[32] ,
    \cb_4_8_io_eo[31] ,
    \cb_4_8_io_eo[30] ,
    \cb_4_8_io_eo[29] ,
    \cb_4_8_io_eo[28] ,
    \cb_4_8_io_eo[27] ,
    \cb_4_8_io_eo[26] ,
    \cb_4_8_io_eo[25] ,
    \cb_4_8_io_eo[24] ,
    \cb_4_8_io_eo[23] ,
    \cb_4_8_io_eo[22] ,
    \cb_4_8_io_eo[21] ,
    \cb_4_8_io_eo[20] ,
    \cb_4_8_io_eo[19] ,
    \cb_4_8_io_eo[18] ,
    \cb_4_8_io_eo[17] ,
    \cb_4_8_io_eo[16] ,
    \cb_4_8_io_eo[15] ,
    \cb_4_8_io_eo[14] ,
    \cb_4_8_io_eo[13] ,
    \cb_4_8_io_eo[12] ,
    \cb_4_8_io_eo[11] ,
    \cb_4_8_io_eo[10] ,
    \cb_4_8_io_eo[9] ,
    \cb_4_8_io_eo[8] ,
    \cb_4_8_io_eo[7] ,
    \cb_4_8_io_eo[6] ,
    \cb_4_8_io_eo[5] ,
    \cb_4_8_io_eo[4] ,
    \cb_4_8_io_eo[3] ,
    \cb_4_8_io_eo[2] ,
    \cb_4_8_io_eo[1] ,
    \cb_4_8_io_eo[0] }),
    .io_i_0_in1({\cb_4_7_io_o_0_out[7] ,
    \cb_4_7_io_o_0_out[6] ,
    \cb_4_7_io_o_0_out[5] ,
    \cb_4_7_io_o_0_out[4] ,
    \cb_4_7_io_o_0_out[3] ,
    \cb_4_7_io_o_0_out[2] ,
    \cb_4_7_io_o_0_out[1] ,
    \cb_4_7_io_o_0_out[0] }),
    .io_i_1_in1({\cb_4_7_io_o_1_out[7] ,
    \cb_4_7_io_o_1_out[6] ,
    \cb_4_7_io_o_1_out[5] ,
    \cb_4_7_io_o_1_out[4] ,
    \cb_4_7_io_o_1_out[3] ,
    \cb_4_7_io_o_1_out[2] ,
    \cb_4_7_io_o_1_out[1] ,
    \cb_4_7_io_o_1_out[0] }),
    .io_i_2_in1({\cb_4_7_io_o_2_out[7] ,
    \cb_4_7_io_o_2_out[6] ,
    \cb_4_7_io_o_2_out[5] ,
    \cb_4_7_io_o_2_out[4] ,
    \cb_4_7_io_o_2_out[3] ,
    \cb_4_7_io_o_2_out[2] ,
    \cb_4_7_io_o_2_out[1] ,
    \cb_4_7_io_o_2_out[0] }),
    .io_i_3_in1({\cb_4_7_io_o_3_out[7] ,
    \cb_4_7_io_o_3_out[6] ,
    \cb_4_7_io_o_3_out[5] ,
    \cb_4_7_io_o_3_out[4] ,
    \cb_4_7_io_o_3_out[3] ,
    \cb_4_7_io_o_3_out[2] ,
    \cb_4_7_io_o_3_out[1] ,
    \cb_4_7_io_o_3_out[0] }),
    .io_i_4_in1({\cb_4_7_io_o_4_out[7] ,
    \cb_4_7_io_o_4_out[6] ,
    \cb_4_7_io_o_4_out[5] ,
    \cb_4_7_io_o_4_out[4] ,
    \cb_4_7_io_o_4_out[3] ,
    \cb_4_7_io_o_4_out[2] ,
    \cb_4_7_io_o_4_out[1] ,
    \cb_4_7_io_o_4_out[0] }),
    .io_i_5_in1({\cb_4_7_io_o_5_out[7] ,
    \cb_4_7_io_o_5_out[6] ,
    \cb_4_7_io_o_5_out[5] ,
    \cb_4_7_io_o_5_out[4] ,
    \cb_4_7_io_o_5_out[3] ,
    \cb_4_7_io_o_5_out[2] ,
    \cb_4_7_io_o_5_out[1] ,
    \cb_4_7_io_o_5_out[0] }),
    .io_i_6_in1({\cb_4_7_io_o_6_out[7] ,
    \cb_4_7_io_o_6_out[6] ,
    \cb_4_7_io_o_6_out[5] ,
    \cb_4_7_io_o_6_out[4] ,
    \cb_4_7_io_o_6_out[3] ,
    \cb_4_7_io_o_6_out[2] ,
    \cb_4_7_io_o_6_out[1] ,
    \cb_4_7_io_o_6_out[0] }),
    .io_i_7_in1({\cb_4_7_io_o_7_out[7] ,
    \cb_4_7_io_o_7_out[6] ,
    \cb_4_7_io_o_7_out[5] ,
    \cb_4_7_io_o_7_out[4] ,
    \cb_4_7_io_o_7_out[3] ,
    \cb_4_7_io_o_7_out[2] ,
    \cb_4_7_io_o_7_out[1] ,
    \cb_4_7_io_o_7_out[0] }),
    .io_o_0_out({\cb_4_8_io_o_0_out[7] ,
    \cb_4_8_io_o_0_out[6] ,
    \cb_4_8_io_o_0_out[5] ,
    \cb_4_8_io_o_0_out[4] ,
    \cb_4_8_io_o_0_out[3] ,
    \cb_4_8_io_o_0_out[2] ,
    \cb_4_8_io_o_0_out[1] ,
    \cb_4_8_io_o_0_out[0] }),
    .io_o_1_out({\cb_4_8_io_o_1_out[7] ,
    \cb_4_8_io_o_1_out[6] ,
    \cb_4_8_io_o_1_out[5] ,
    \cb_4_8_io_o_1_out[4] ,
    \cb_4_8_io_o_1_out[3] ,
    \cb_4_8_io_o_1_out[2] ,
    \cb_4_8_io_o_1_out[1] ,
    \cb_4_8_io_o_1_out[0] }),
    .io_o_2_out({\cb_4_8_io_o_2_out[7] ,
    \cb_4_8_io_o_2_out[6] ,
    \cb_4_8_io_o_2_out[5] ,
    \cb_4_8_io_o_2_out[4] ,
    \cb_4_8_io_o_2_out[3] ,
    \cb_4_8_io_o_2_out[2] ,
    \cb_4_8_io_o_2_out[1] ,
    \cb_4_8_io_o_2_out[0] }),
    .io_o_3_out({\cb_4_8_io_o_3_out[7] ,
    \cb_4_8_io_o_3_out[6] ,
    \cb_4_8_io_o_3_out[5] ,
    \cb_4_8_io_o_3_out[4] ,
    \cb_4_8_io_o_3_out[3] ,
    \cb_4_8_io_o_3_out[2] ,
    \cb_4_8_io_o_3_out[1] ,
    \cb_4_8_io_o_3_out[0] }),
    .io_o_4_out({\cb_4_8_io_o_4_out[7] ,
    \cb_4_8_io_o_4_out[6] ,
    \cb_4_8_io_o_4_out[5] ,
    \cb_4_8_io_o_4_out[4] ,
    \cb_4_8_io_o_4_out[3] ,
    \cb_4_8_io_o_4_out[2] ,
    \cb_4_8_io_o_4_out[1] ,
    \cb_4_8_io_o_4_out[0] }),
    .io_o_5_out({\cb_4_8_io_o_5_out[7] ,
    \cb_4_8_io_o_5_out[6] ,
    \cb_4_8_io_o_5_out[5] ,
    \cb_4_8_io_o_5_out[4] ,
    \cb_4_8_io_o_5_out[3] ,
    \cb_4_8_io_o_5_out[2] ,
    \cb_4_8_io_o_5_out[1] ,
    \cb_4_8_io_o_5_out[0] }),
    .io_o_6_out({\cb_4_8_io_o_6_out[7] ,
    \cb_4_8_io_o_6_out[6] ,
    \cb_4_8_io_o_6_out[5] ,
    \cb_4_8_io_o_6_out[4] ,
    \cb_4_8_io_o_6_out[3] ,
    \cb_4_8_io_o_6_out[2] ,
    \cb_4_8_io_o_6_out[1] ,
    \cb_4_8_io_o_6_out[0] }),
    .io_o_7_out({\cb_4_8_io_o_7_out[7] ,
    \cb_4_8_io_o_7_out[6] ,
    \cb_4_8_io_o_7_out[5] ,
    \cb_4_8_io_o_7_out[4] ,
    \cb_4_8_io_o_7_out[3] ,
    \cb_4_8_io_o_7_out[2] ,
    \cb_4_8_io_o_7_out[1] ,
    \cb_4_8_io_o_7_out[0] }),
    .io_wo({\cb_4_7_io_eo[63] ,
    \cb_4_7_io_eo[62] ,
    \cb_4_7_io_eo[61] ,
    \cb_4_7_io_eo[60] ,
    \cb_4_7_io_eo[59] ,
    \cb_4_7_io_eo[58] ,
    \cb_4_7_io_eo[57] ,
    \cb_4_7_io_eo[56] ,
    \cb_4_7_io_eo[55] ,
    \cb_4_7_io_eo[54] ,
    \cb_4_7_io_eo[53] ,
    \cb_4_7_io_eo[52] ,
    \cb_4_7_io_eo[51] ,
    \cb_4_7_io_eo[50] ,
    \cb_4_7_io_eo[49] ,
    \cb_4_7_io_eo[48] ,
    \cb_4_7_io_eo[47] ,
    \cb_4_7_io_eo[46] ,
    \cb_4_7_io_eo[45] ,
    \cb_4_7_io_eo[44] ,
    \cb_4_7_io_eo[43] ,
    \cb_4_7_io_eo[42] ,
    \cb_4_7_io_eo[41] ,
    \cb_4_7_io_eo[40] ,
    \cb_4_7_io_eo[39] ,
    \cb_4_7_io_eo[38] ,
    \cb_4_7_io_eo[37] ,
    \cb_4_7_io_eo[36] ,
    \cb_4_7_io_eo[35] ,
    \cb_4_7_io_eo[34] ,
    \cb_4_7_io_eo[33] ,
    \cb_4_7_io_eo[32] ,
    \cb_4_7_io_eo[31] ,
    \cb_4_7_io_eo[30] ,
    \cb_4_7_io_eo[29] ,
    \cb_4_7_io_eo[28] ,
    \cb_4_7_io_eo[27] ,
    \cb_4_7_io_eo[26] ,
    \cb_4_7_io_eo[25] ,
    \cb_4_7_io_eo[24] ,
    \cb_4_7_io_eo[23] ,
    \cb_4_7_io_eo[22] ,
    \cb_4_7_io_eo[21] ,
    \cb_4_7_io_eo[20] ,
    \cb_4_7_io_eo[19] ,
    \cb_4_7_io_eo[18] ,
    \cb_4_7_io_eo[17] ,
    \cb_4_7_io_eo[16] ,
    \cb_4_7_io_eo[15] ,
    \cb_4_7_io_eo[14] ,
    \cb_4_7_io_eo[13] ,
    \cb_4_7_io_eo[12] ,
    \cb_4_7_io_eo[11] ,
    \cb_4_7_io_eo[10] ,
    \cb_4_7_io_eo[9] ,
    \cb_4_7_io_eo[8] ,
    \cb_4_7_io_eo[7] ,
    \cb_4_7_io_eo[6] ,
    \cb_4_7_io_eo[5] ,
    \cb_4_7_io_eo[4] ,
    \cb_4_7_io_eo[3] ,
    \cb_4_7_io_eo[2] ,
    \cb_4_7_io_eo[1] ,
    \cb_4_7_io_eo[0] }));
 cic_block cb_4_9 (.io_cs_i(cb_4_9_io_cs_i),
    .io_i_0_ci(cb_4_8_io_o_0_co),
    .io_i_1_ci(cb_4_8_io_o_1_co),
    .io_i_2_ci(cb_4_8_io_o_2_co),
    .io_i_3_ci(cb_4_8_io_o_3_co),
    .io_i_4_ci(cb_4_8_io_o_4_co),
    .io_i_5_ci(cb_4_8_io_o_5_co),
    .io_i_6_ci(cb_4_8_io_o_6_co),
    .io_i_7_ci(cb_4_8_io_o_7_co),
    .io_o_0_co(cb_4_10_io_i_0_ci),
    .io_o_1_co(cb_4_10_io_i_1_ci),
    .io_o_2_co(cb_4_10_io_i_2_ci),
    .io_o_3_co(cb_4_10_io_i_3_ci),
    .io_o_4_co(cb_4_10_io_i_4_ci),
    .io_o_5_co(cb_4_10_io_i_5_ci),
    .io_o_6_co(cb_4_10_io_i_6_ci),
    .io_o_7_co(cb_4_10_io_i_7_ci),
    .io_vci(cb_4_8_io_vco),
    .io_vco(cb_4_10_io_vci),
    .io_vi(cb_4_9_io_vi),
    .io_we_i(cb_4_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_4_0_io_adr_i[1] ,
    \cb_4_0_io_adr_i[0] }),
    .io_dat_i({\cb_4_0_io_dat_i[15] ,
    \cb_4_0_io_dat_i[14] ,
    \cb_4_0_io_dat_i[13] ,
    \cb_4_0_io_dat_i[12] ,
    \cb_4_0_io_dat_i[11] ,
    \cb_4_0_io_dat_i[10] ,
    \cb_4_0_io_dat_i[9] ,
    \cb_4_0_io_dat_i[8] ,
    \cb_4_0_io_dat_i[7] ,
    \cb_4_0_io_dat_i[6] ,
    \cb_4_0_io_dat_i[5] ,
    \cb_4_0_io_dat_i[4] ,
    \cb_4_0_io_dat_i[3] ,
    \cb_4_0_io_dat_i[2] ,
    \cb_4_0_io_dat_i[1] ,
    \cb_4_0_io_dat_i[0] }),
    .io_dat_o({\cb_4_9_io_dat_o[15] ,
    \cb_4_9_io_dat_o[14] ,
    \cb_4_9_io_dat_o[13] ,
    \cb_4_9_io_dat_o[12] ,
    \cb_4_9_io_dat_o[11] ,
    \cb_4_9_io_dat_o[10] ,
    \cb_4_9_io_dat_o[9] ,
    \cb_4_9_io_dat_o[8] ,
    \cb_4_9_io_dat_o[7] ,
    \cb_4_9_io_dat_o[6] ,
    \cb_4_9_io_dat_o[5] ,
    \cb_4_9_io_dat_o[4] ,
    \cb_4_9_io_dat_o[3] ,
    \cb_4_9_io_dat_o[2] ,
    \cb_4_9_io_dat_o[1] ,
    \cb_4_9_io_dat_o[0] }),
    .io_eo({\cb_4_10_io_wo[63] ,
    \cb_4_10_io_wo[62] ,
    \cb_4_10_io_wo[61] ,
    \cb_4_10_io_wo[60] ,
    \cb_4_10_io_wo[59] ,
    \cb_4_10_io_wo[58] ,
    \cb_4_10_io_wo[57] ,
    \cb_4_10_io_wo[56] ,
    \cb_4_10_io_wo[55] ,
    \cb_4_10_io_wo[54] ,
    \cb_4_10_io_wo[53] ,
    \cb_4_10_io_wo[52] ,
    \cb_4_10_io_wo[51] ,
    \cb_4_10_io_wo[50] ,
    \cb_4_10_io_wo[49] ,
    \cb_4_10_io_wo[48] ,
    \cb_4_10_io_wo[47] ,
    \cb_4_10_io_wo[46] ,
    \cb_4_10_io_wo[45] ,
    \cb_4_10_io_wo[44] ,
    \cb_4_10_io_wo[43] ,
    \cb_4_10_io_wo[42] ,
    \cb_4_10_io_wo[41] ,
    \cb_4_10_io_wo[40] ,
    \cb_4_10_io_wo[39] ,
    \cb_4_10_io_wo[38] ,
    \cb_4_10_io_wo[37] ,
    \cb_4_10_io_wo[36] ,
    \cb_4_10_io_wo[35] ,
    \cb_4_10_io_wo[34] ,
    \cb_4_10_io_wo[33] ,
    \cb_4_10_io_wo[32] ,
    \cb_4_10_io_wo[31] ,
    \cb_4_10_io_wo[30] ,
    \cb_4_10_io_wo[29] ,
    \cb_4_10_io_wo[28] ,
    \cb_4_10_io_wo[27] ,
    \cb_4_10_io_wo[26] ,
    \cb_4_10_io_wo[25] ,
    \cb_4_10_io_wo[24] ,
    \cb_4_10_io_wo[23] ,
    \cb_4_10_io_wo[22] ,
    \cb_4_10_io_wo[21] ,
    \cb_4_10_io_wo[20] ,
    \cb_4_10_io_wo[19] ,
    \cb_4_10_io_wo[18] ,
    \cb_4_10_io_wo[17] ,
    \cb_4_10_io_wo[16] ,
    \cb_4_10_io_wo[15] ,
    \cb_4_10_io_wo[14] ,
    \cb_4_10_io_wo[13] ,
    \cb_4_10_io_wo[12] ,
    \cb_4_10_io_wo[11] ,
    \cb_4_10_io_wo[10] ,
    \cb_4_10_io_wo[9] ,
    \cb_4_10_io_wo[8] ,
    \cb_4_10_io_wo[7] ,
    \cb_4_10_io_wo[6] ,
    \cb_4_10_io_wo[5] ,
    \cb_4_10_io_wo[4] ,
    \cb_4_10_io_wo[3] ,
    \cb_4_10_io_wo[2] ,
    \cb_4_10_io_wo[1] ,
    \cb_4_10_io_wo[0] }),
    .io_i_0_in1({\cb_4_8_io_o_0_out[7] ,
    \cb_4_8_io_o_0_out[6] ,
    \cb_4_8_io_o_0_out[5] ,
    \cb_4_8_io_o_0_out[4] ,
    \cb_4_8_io_o_0_out[3] ,
    \cb_4_8_io_o_0_out[2] ,
    \cb_4_8_io_o_0_out[1] ,
    \cb_4_8_io_o_0_out[0] }),
    .io_i_1_in1({\cb_4_8_io_o_1_out[7] ,
    \cb_4_8_io_o_1_out[6] ,
    \cb_4_8_io_o_1_out[5] ,
    \cb_4_8_io_o_1_out[4] ,
    \cb_4_8_io_o_1_out[3] ,
    \cb_4_8_io_o_1_out[2] ,
    \cb_4_8_io_o_1_out[1] ,
    \cb_4_8_io_o_1_out[0] }),
    .io_i_2_in1({\cb_4_8_io_o_2_out[7] ,
    \cb_4_8_io_o_2_out[6] ,
    \cb_4_8_io_o_2_out[5] ,
    \cb_4_8_io_o_2_out[4] ,
    \cb_4_8_io_o_2_out[3] ,
    \cb_4_8_io_o_2_out[2] ,
    \cb_4_8_io_o_2_out[1] ,
    \cb_4_8_io_o_2_out[0] }),
    .io_i_3_in1({\cb_4_8_io_o_3_out[7] ,
    \cb_4_8_io_o_3_out[6] ,
    \cb_4_8_io_o_3_out[5] ,
    \cb_4_8_io_o_3_out[4] ,
    \cb_4_8_io_o_3_out[3] ,
    \cb_4_8_io_o_3_out[2] ,
    \cb_4_8_io_o_3_out[1] ,
    \cb_4_8_io_o_3_out[0] }),
    .io_i_4_in1({\cb_4_8_io_o_4_out[7] ,
    \cb_4_8_io_o_4_out[6] ,
    \cb_4_8_io_o_4_out[5] ,
    \cb_4_8_io_o_4_out[4] ,
    \cb_4_8_io_o_4_out[3] ,
    \cb_4_8_io_o_4_out[2] ,
    \cb_4_8_io_o_4_out[1] ,
    \cb_4_8_io_o_4_out[0] }),
    .io_i_5_in1({\cb_4_8_io_o_5_out[7] ,
    \cb_4_8_io_o_5_out[6] ,
    \cb_4_8_io_o_5_out[5] ,
    \cb_4_8_io_o_5_out[4] ,
    \cb_4_8_io_o_5_out[3] ,
    \cb_4_8_io_o_5_out[2] ,
    \cb_4_8_io_o_5_out[1] ,
    \cb_4_8_io_o_5_out[0] }),
    .io_i_6_in1({\cb_4_8_io_o_6_out[7] ,
    \cb_4_8_io_o_6_out[6] ,
    \cb_4_8_io_o_6_out[5] ,
    \cb_4_8_io_o_6_out[4] ,
    \cb_4_8_io_o_6_out[3] ,
    \cb_4_8_io_o_6_out[2] ,
    \cb_4_8_io_o_6_out[1] ,
    \cb_4_8_io_o_6_out[0] }),
    .io_i_7_in1({\cb_4_8_io_o_7_out[7] ,
    \cb_4_8_io_o_7_out[6] ,
    \cb_4_8_io_o_7_out[5] ,
    \cb_4_8_io_o_7_out[4] ,
    \cb_4_8_io_o_7_out[3] ,
    \cb_4_8_io_o_7_out[2] ,
    \cb_4_8_io_o_7_out[1] ,
    \cb_4_8_io_o_7_out[0] }),
    .io_o_0_out({\cb_4_10_io_i_0_in1[7] ,
    \cb_4_10_io_i_0_in1[6] ,
    \cb_4_10_io_i_0_in1[5] ,
    \cb_4_10_io_i_0_in1[4] ,
    \cb_4_10_io_i_0_in1[3] ,
    \cb_4_10_io_i_0_in1[2] ,
    \cb_4_10_io_i_0_in1[1] ,
    \cb_4_10_io_i_0_in1[0] }),
    .io_o_1_out({\cb_4_10_io_i_1_in1[7] ,
    \cb_4_10_io_i_1_in1[6] ,
    \cb_4_10_io_i_1_in1[5] ,
    \cb_4_10_io_i_1_in1[4] ,
    \cb_4_10_io_i_1_in1[3] ,
    \cb_4_10_io_i_1_in1[2] ,
    \cb_4_10_io_i_1_in1[1] ,
    \cb_4_10_io_i_1_in1[0] }),
    .io_o_2_out({\cb_4_10_io_i_2_in1[7] ,
    \cb_4_10_io_i_2_in1[6] ,
    \cb_4_10_io_i_2_in1[5] ,
    \cb_4_10_io_i_2_in1[4] ,
    \cb_4_10_io_i_2_in1[3] ,
    \cb_4_10_io_i_2_in1[2] ,
    \cb_4_10_io_i_2_in1[1] ,
    \cb_4_10_io_i_2_in1[0] }),
    .io_o_3_out({\cb_4_10_io_i_3_in1[7] ,
    \cb_4_10_io_i_3_in1[6] ,
    \cb_4_10_io_i_3_in1[5] ,
    \cb_4_10_io_i_3_in1[4] ,
    \cb_4_10_io_i_3_in1[3] ,
    \cb_4_10_io_i_3_in1[2] ,
    \cb_4_10_io_i_3_in1[1] ,
    \cb_4_10_io_i_3_in1[0] }),
    .io_o_4_out({\cb_4_10_io_i_4_in1[7] ,
    \cb_4_10_io_i_4_in1[6] ,
    \cb_4_10_io_i_4_in1[5] ,
    \cb_4_10_io_i_4_in1[4] ,
    \cb_4_10_io_i_4_in1[3] ,
    \cb_4_10_io_i_4_in1[2] ,
    \cb_4_10_io_i_4_in1[1] ,
    \cb_4_10_io_i_4_in1[0] }),
    .io_o_5_out({\cb_4_10_io_i_5_in1[7] ,
    \cb_4_10_io_i_5_in1[6] ,
    \cb_4_10_io_i_5_in1[5] ,
    \cb_4_10_io_i_5_in1[4] ,
    \cb_4_10_io_i_5_in1[3] ,
    \cb_4_10_io_i_5_in1[2] ,
    \cb_4_10_io_i_5_in1[1] ,
    \cb_4_10_io_i_5_in1[0] }),
    .io_o_6_out({\cb_4_10_io_i_6_in1[7] ,
    \cb_4_10_io_i_6_in1[6] ,
    \cb_4_10_io_i_6_in1[5] ,
    \cb_4_10_io_i_6_in1[4] ,
    \cb_4_10_io_i_6_in1[3] ,
    \cb_4_10_io_i_6_in1[2] ,
    \cb_4_10_io_i_6_in1[1] ,
    \cb_4_10_io_i_6_in1[0] }),
    .io_o_7_out({\cb_4_10_io_i_7_in1[7] ,
    \cb_4_10_io_i_7_in1[6] ,
    \cb_4_10_io_i_7_in1[5] ,
    \cb_4_10_io_i_7_in1[4] ,
    \cb_4_10_io_i_7_in1[3] ,
    \cb_4_10_io_i_7_in1[2] ,
    \cb_4_10_io_i_7_in1[1] ,
    \cb_4_10_io_i_7_in1[0] }),
    .io_wo({\cb_4_8_io_eo[63] ,
    \cb_4_8_io_eo[62] ,
    \cb_4_8_io_eo[61] ,
    \cb_4_8_io_eo[60] ,
    \cb_4_8_io_eo[59] ,
    \cb_4_8_io_eo[58] ,
    \cb_4_8_io_eo[57] ,
    \cb_4_8_io_eo[56] ,
    \cb_4_8_io_eo[55] ,
    \cb_4_8_io_eo[54] ,
    \cb_4_8_io_eo[53] ,
    \cb_4_8_io_eo[52] ,
    \cb_4_8_io_eo[51] ,
    \cb_4_8_io_eo[50] ,
    \cb_4_8_io_eo[49] ,
    \cb_4_8_io_eo[48] ,
    \cb_4_8_io_eo[47] ,
    \cb_4_8_io_eo[46] ,
    \cb_4_8_io_eo[45] ,
    \cb_4_8_io_eo[44] ,
    \cb_4_8_io_eo[43] ,
    \cb_4_8_io_eo[42] ,
    \cb_4_8_io_eo[41] ,
    \cb_4_8_io_eo[40] ,
    \cb_4_8_io_eo[39] ,
    \cb_4_8_io_eo[38] ,
    \cb_4_8_io_eo[37] ,
    \cb_4_8_io_eo[36] ,
    \cb_4_8_io_eo[35] ,
    \cb_4_8_io_eo[34] ,
    \cb_4_8_io_eo[33] ,
    \cb_4_8_io_eo[32] ,
    \cb_4_8_io_eo[31] ,
    \cb_4_8_io_eo[30] ,
    \cb_4_8_io_eo[29] ,
    \cb_4_8_io_eo[28] ,
    \cb_4_8_io_eo[27] ,
    \cb_4_8_io_eo[26] ,
    \cb_4_8_io_eo[25] ,
    \cb_4_8_io_eo[24] ,
    \cb_4_8_io_eo[23] ,
    \cb_4_8_io_eo[22] ,
    \cb_4_8_io_eo[21] ,
    \cb_4_8_io_eo[20] ,
    \cb_4_8_io_eo[19] ,
    \cb_4_8_io_eo[18] ,
    \cb_4_8_io_eo[17] ,
    \cb_4_8_io_eo[16] ,
    \cb_4_8_io_eo[15] ,
    \cb_4_8_io_eo[14] ,
    \cb_4_8_io_eo[13] ,
    \cb_4_8_io_eo[12] ,
    \cb_4_8_io_eo[11] ,
    \cb_4_8_io_eo[10] ,
    \cb_4_8_io_eo[9] ,
    \cb_4_8_io_eo[8] ,
    \cb_4_8_io_eo[7] ,
    \cb_4_8_io_eo[6] ,
    \cb_4_8_io_eo[5] ,
    \cb_4_8_io_eo[4] ,
    \cb_4_8_io_eo[3] ,
    \cb_4_8_io_eo[2] ,
    \cb_4_8_io_eo[1] ,
    \cb_4_8_io_eo[0] }));
 cic_block cb_5_0 (.io_cs_i(cb_5_0_io_cs_i),
    .io_i_0_ci(cb_5_0_io_i_0_ci),
    .io_o_0_co(cb_5_0_io_o_0_co),
    .io_o_1_co(cb_5_0_io_o_1_co),
    .io_o_2_co(cb_5_0_io_o_2_co),
    .io_o_3_co(cb_5_0_io_o_3_co),
    .io_o_4_co(cb_5_0_io_o_4_co),
    .io_o_5_co(cb_5_0_io_o_5_co),
    .io_o_6_co(cb_5_0_io_o_6_co),
    .io_o_7_co(cb_5_0_io_o_7_co),
    .io_vco(cb_5_0_io_vco),
    .io_vi(cb_5_0_io_vi),
    .io_we_i(cb_5_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_5_0_io_adr_i[1] ,
    \cb_5_0_io_adr_i[0] }),
    .io_dat_i({\cb_5_0_io_dat_i[15] ,
    \cb_5_0_io_dat_i[14] ,
    \cb_5_0_io_dat_i[13] ,
    \cb_5_0_io_dat_i[12] ,
    \cb_5_0_io_dat_i[11] ,
    \cb_5_0_io_dat_i[10] ,
    \cb_5_0_io_dat_i[9] ,
    \cb_5_0_io_dat_i[8] ,
    \cb_5_0_io_dat_i[7] ,
    \cb_5_0_io_dat_i[6] ,
    \cb_5_0_io_dat_i[5] ,
    \cb_5_0_io_dat_i[4] ,
    \cb_5_0_io_dat_i[3] ,
    \cb_5_0_io_dat_i[2] ,
    \cb_5_0_io_dat_i[1] ,
    \cb_5_0_io_dat_i[0] }),
    .io_dat_o({\cb_5_0_io_dat_o[15] ,
    \cb_5_0_io_dat_o[14] ,
    \cb_5_0_io_dat_o[13] ,
    \cb_5_0_io_dat_o[12] ,
    \cb_5_0_io_dat_o[11] ,
    \cb_5_0_io_dat_o[10] ,
    \cb_5_0_io_dat_o[9] ,
    \cb_5_0_io_dat_o[8] ,
    \cb_5_0_io_dat_o[7] ,
    \cb_5_0_io_dat_o[6] ,
    \cb_5_0_io_dat_o[5] ,
    \cb_5_0_io_dat_o[4] ,
    \cb_5_0_io_dat_o[3] ,
    \cb_5_0_io_dat_o[2] ,
    \cb_5_0_io_dat_o[1] ,
    \cb_5_0_io_dat_o[0] }),
    .io_eo({\cb_5_0_io_eo[63] ,
    \cb_5_0_io_eo[62] ,
    \cb_5_0_io_eo[61] ,
    \cb_5_0_io_eo[60] ,
    \cb_5_0_io_eo[59] ,
    \cb_5_0_io_eo[58] ,
    \cb_5_0_io_eo[57] ,
    \cb_5_0_io_eo[56] ,
    \cb_5_0_io_eo[55] ,
    \cb_5_0_io_eo[54] ,
    \cb_5_0_io_eo[53] ,
    \cb_5_0_io_eo[52] ,
    \cb_5_0_io_eo[51] ,
    \cb_5_0_io_eo[50] ,
    \cb_5_0_io_eo[49] ,
    \cb_5_0_io_eo[48] ,
    \cb_5_0_io_eo[47] ,
    \cb_5_0_io_eo[46] ,
    \cb_5_0_io_eo[45] ,
    \cb_5_0_io_eo[44] ,
    \cb_5_0_io_eo[43] ,
    \cb_5_0_io_eo[42] ,
    \cb_5_0_io_eo[41] ,
    \cb_5_0_io_eo[40] ,
    \cb_5_0_io_eo[39] ,
    \cb_5_0_io_eo[38] ,
    \cb_5_0_io_eo[37] ,
    \cb_5_0_io_eo[36] ,
    \cb_5_0_io_eo[35] ,
    \cb_5_0_io_eo[34] ,
    \cb_5_0_io_eo[33] ,
    \cb_5_0_io_eo[32] ,
    \cb_5_0_io_eo[31] ,
    \cb_5_0_io_eo[30] ,
    \cb_5_0_io_eo[29] ,
    \cb_5_0_io_eo[28] ,
    \cb_5_0_io_eo[27] ,
    \cb_5_0_io_eo[26] ,
    \cb_5_0_io_eo[25] ,
    \cb_5_0_io_eo[24] ,
    \cb_5_0_io_eo[23] ,
    \cb_5_0_io_eo[22] ,
    \cb_5_0_io_eo[21] ,
    \cb_5_0_io_eo[20] ,
    \cb_5_0_io_eo[19] ,
    \cb_5_0_io_eo[18] ,
    \cb_5_0_io_eo[17] ,
    \cb_5_0_io_eo[16] ,
    \cb_5_0_io_eo[15] ,
    \cb_5_0_io_eo[14] ,
    \cb_5_0_io_eo[13] ,
    \cb_5_0_io_eo[12] ,
    \cb_5_0_io_eo[11] ,
    \cb_5_0_io_eo[10] ,
    \cb_5_0_io_eo[9] ,
    \cb_5_0_io_eo[8] ,
    \cb_5_0_io_eo[7] ,
    \cb_5_0_io_eo[6] ,
    \cb_5_0_io_eo[5] ,
    \cb_5_0_io_eo[4] ,
    \cb_5_0_io_eo[3] ,
    \cb_5_0_io_eo[2] ,
    \cb_5_0_io_eo[1] ,
    \cb_5_0_io_eo[0] }),
    .io_i_0_in1({_NC321,
    _NC322,
    _NC323,
    _NC324,
    _NC325,
    _NC326,
    _NC327,
    _NC328}),
    .io_i_1_in1({_NC329,
    _NC330,
    _NC331,
    _NC332,
    _NC333,
    _NC334,
    _NC335,
    _NC336}),
    .io_i_2_in1({_NC337,
    _NC338,
    _NC339,
    _NC340,
    _NC341,
    _NC342,
    _NC343,
    _NC344}),
    .io_i_3_in1({_NC345,
    _NC346,
    _NC347,
    _NC348,
    _NC349,
    _NC350,
    _NC351,
    _NC352}),
    .io_i_4_in1({_NC353,
    _NC354,
    _NC355,
    _NC356,
    _NC357,
    _NC358,
    _NC359,
    _NC360}),
    .io_i_5_in1({_NC361,
    _NC362,
    _NC363,
    _NC364,
    _NC365,
    _NC366,
    _NC367,
    _NC368}),
    .io_i_6_in1({_NC369,
    _NC370,
    _NC371,
    _NC372,
    _NC373,
    _NC374,
    _NC375,
    _NC376}),
    .io_i_7_in1({_NC377,
    _NC378,
    _NC379,
    _NC380,
    _NC381,
    _NC382,
    _NC383,
    _NC384}),
    .io_o_0_out({\cb_5_0_io_o_0_out[7] ,
    \cb_5_0_io_o_0_out[6] ,
    \cb_5_0_io_o_0_out[5] ,
    \cb_5_0_io_o_0_out[4] ,
    \cb_5_0_io_o_0_out[3] ,
    \cb_5_0_io_o_0_out[2] ,
    \cb_5_0_io_o_0_out[1] ,
    \cb_5_0_io_o_0_out[0] }),
    .io_o_1_out({\cb_5_0_io_o_1_out[7] ,
    \cb_5_0_io_o_1_out[6] ,
    \cb_5_0_io_o_1_out[5] ,
    \cb_5_0_io_o_1_out[4] ,
    \cb_5_0_io_o_1_out[3] ,
    \cb_5_0_io_o_1_out[2] ,
    \cb_5_0_io_o_1_out[1] ,
    \cb_5_0_io_o_1_out[0] }),
    .io_o_2_out({\cb_5_0_io_o_2_out[7] ,
    \cb_5_0_io_o_2_out[6] ,
    \cb_5_0_io_o_2_out[5] ,
    \cb_5_0_io_o_2_out[4] ,
    \cb_5_0_io_o_2_out[3] ,
    \cb_5_0_io_o_2_out[2] ,
    \cb_5_0_io_o_2_out[1] ,
    \cb_5_0_io_o_2_out[0] }),
    .io_o_3_out({\cb_5_0_io_o_3_out[7] ,
    \cb_5_0_io_o_3_out[6] ,
    \cb_5_0_io_o_3_out[5] ,
    \cb_5_0_io_o_3_out[4] ,
    \cb_5_0_io_o_3_out[3] ,
    \cb_5_0_io_o_3_out[2] ,
    \cb_5_0_io_o_3_out[1] ,
    \cb_5_0_io_o_3_out[0] }),
    .io_o_4_out({\cb_5_0_io_o_4_out[7] ,
    \cb_5_0_io_o_4_out[6] ,
    \cb_5_0_io_o_4_out[5] ,
    \cb_5_0_io_o_4_out[4] ,
    \cb_5_0_io_o_4_out[3] ,
    \cb_5_0_io_o_4_out[2] ,
    \cb_5_0_io_o_4_out[1] ,
    \cb_5_0_io_o_4_out[0] }),
    .io_o_5_out({\cb_5_0_io_o_5_out[7] ,
    \cb_5_0_io_o_5_out[6] ,
    \cb_5_0_io_o_5_out[5] ,
    \cb_5_0_io_o_5_out[4] ,
    \cb_5_0_io_o_5_out[3] ,
    \cb_5_0_io_o_5_out[2] ,
    \cb_5_0_io_o_5_out[1] ,
    \cb_5_0_io_o_5_out[0] }),
    .io_o_6_out({\cb_5_0_io_o_6_out[7] ,
    \cb_5_0_io_o_6_out[6] ,
    \cb_5_0_io_o_6_out[5] ,
    \cb_5_0_io_o_6_out[4] ,
    \cb_5_0_io_o_6_out[3] ,
    \cb_5_0_io_o_6_out[2] ,
    \cb_5_0_io_o_6_out[1] ,
    \cb_5_0_io_o_6_out[0] }),
    .io_o_7_out({\cb_5_0_io_o_7_out[7] ,
    \cb_5_0_io_o_7_out[6] ,
    \cb_5_0_io_o_7_out[5] ,
    \cb_5_0_io_o_7_out[4] ,
    \cb_5_0_io_o_7_out[3] ,
    \cb_5_0_io_o_7_out[2] ,
    \cb_5_0_io_o_7_out[1] ,
    \cb_5_0_io_o_7_out[0] }),
    .io_wo({\cb_5_0_io_wo[63] ,
    \cb_5_0_io_wo[62] ,
    \cb_5_0_io_wo[61] ,
    \cb_5_0_io_wo[60] ,
    \cb_5_0_io_wo[59] ,
    \cb_5_0_io_wo[58] ,
    \cb_5_0_io_wo[57] ,
    \cb_5_0_io_wo[56] ,
    \cb_5_0_io_wo[55] ,
    \cb_5_0_io_wo[54] ,
    \cb_5_0_io_wo[53] ,
    \cb_5_0_io_wo[52] ,
    \cb_5_0_io_wo[51] ,
    \cb_5_0_io_wo[50] ,
    \cb_5_0_io_wo[49] ,
    \cb_5_0_io_wo[48] ,
    \cb_5_0_io_wo[47] ,
    \cb_5_0_io_wo[46] ,
    \cb_5_0_io_wo[45] ,
    \cb_5_0_io_wo[44] ,
    \cb_5_0_io_wo[43] ,
    \cb_5_0_io_wo[42] ,
    \cb_5_0_io_wo[41] ,
    \cb_5_0_io_wo[40] ,
    \cb_5_0_io_wo[39] ,
    \cb_5_0_io_wo[38] ,
    \cb_5_0_io_wo[37] ,
    \cb_5_0_io_wo[36] ,
    \cb_5_0_io_wo[35] ,
    \cb_5_0_io_wo[34] ,
    \cb_5_0_io_wo[33] ,
    \cb_5_0_io_wo[32] ,
    \cb_5_0_io_wo[31] ,
    \cb_5_0_io_wo[30] ,
    \cb_5_0_io_wo[29] ,
    \cb_5_0_io_wo[28] ,
    \cb_5_0_io_wo[27] ,
    \cb_5_0_io_wo[26] ,
    \cb_5_0_io_wo[25] ,
    \cb_5_0_io_wo[24] ,
    \cb_5_0_io_wo[23] ,
    \cb_5_0_io_wo[22] ,
    \cb_5_0_io_wo[21] ,
    \cb_5_0_io_wo[20] ,
    \cb_5_0_io_wo[19] ,
    \cb_5_0_io_wo[18] ,
    \cb_5_0_io_wo[17] ,
    \cb_5_0_io_wo[16] ,
    \cb_5_0_io_wo[15] ,
    \cb_5_0_io_wo[14] ,
    \cb_5_0_io_wo[13] ,
    \cb_5_0_io_wo[12] ,
    \cb_5_0_io_wo[11] ,
    \cb_5_0_io_wo[10] ,
    \cb_5_0_io_wo[9] ,
    \cb_5_0_io_wo[8] ,
    \cb_5_0_io_wo[7] ,
    \cb_5_0_io_wo[6] ,
    \cb_5_0_io_wo[5] ,
    \cb_5_0_io_wo[4] ,
    \cb_5_0_io_wo[3] ,
    \cb_5_0_io_wo[2] ,
    \cb_5_0_io_wo[1] ,
    \cb_5_0_io_wo[0] }));
 cic_block cb_5_1 (.io_cs_i(cb_5_1_io_cs_i),
    .io_i_0_ci(cb_5_0_io_o_0_co),
    .io_i_1_ci(cb_5_0_io_o_1_co),
    .io_i_2_ci(cb_5_0_io_o_2_co),
    .io_i_3_ci(cb_5_0_io_o_3_co),
    .io_i_4_ci(cb_5_0_io_o_4_co),
    .io_i_5_ci(cb_5_0_io_o_5_co),
    .io_i_6_ci(cb_5_0_io_o_6_co),
    .io_i_7_ci(cb_5_0_io_o_7_co),
    .io_o_0_co(cb_5_1_io_o_0_co),
    .io_o_1_co(cb_5_1_io_o_1_co),
    .io_o_2_co(cb_5_1_io_o_2_co),
    .io_o_3_co(cb_5_1_io_o_3_co),
    .io_o_4_co(cb_5_1_io_o_4_co),
    .io_o_5_co(cb_5_1_io_o_5_co),
    .io_o_6_co(cb_5_1_io_o_6_co),
    .io_o_7_co(cb_5_1_io_o_7_co),
    .io_vci(cb_5_0_io_vco),
    .io_vco(cb_5_1_io_vco),
    .io_vi(cb_5_1_io_vi),
    .io_we_i(cb_5_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_5_0_io_adr_i[1] ,
    \cb_5_0_io_adr_i[0] }),
    .io_dat_i({\cb_5_0_io_dat_i[15] ,
    \cb_5_0_io_dat_i[14] ,
    \cb_5_0_io_dat_i[13] ,
    \cb_5_0_io_dat_i[12] ,
    \cb_5_0_io_dat_i[11] ,
    \cb_5_0_io_dat_i[10] ,
    \cb_5_0_io_dat_i[9] ,
    \cb_5_0_io_dat_i[8] ,
    \cb_5_0_io_dat_i[7] ,
    \cb_5_0_io_dat_i[6] ,
    \cb_5_0_io_dat_i[5] ,
    \cb_5_0_io_dat_i[4] ,
    \cb_5_0_io_dat_i[3] ,
    \cb_5_0_io_dat_i[2] ,
    \cb_5_0_io_dat_i[1] ,
    \cb_5_0_io_dat_i[0] }),
    .io_dat_o({\cb_5_1_io_dat_o[15] ,
    \cb_5_1_io_dat_o[14] ,
    \cb_5_1_io_dat_o[13] ,
    \cb_5_1_io_dat_o[12] ,
    \cb_5_1_io_dat_o[11] ,
    \cb_5_1_io_dat_o[10] ,
    \cb_5_1_io_dat_o[9] ,
    \cb_5_1_io_dat_o[8] ,
    \cb_5_1_io_dat_o[7] ,
    \cb_5_1_io_dat_o[6] ,
    \cb_5_1_io_dat_o[5] ,
    \cb_5_1_io_dat_o[4] ,
    \cb_5_1_io_dat_o[3] ,
    \cb_5_1_io_dat_o[2] ,
    \cb_5_1_io_dat_o[1] ,
    \cb_5_1_io_dat_o[0] }),
    .io_eo({\cb_5_1_io_eo[63] ,
    \cb_5_1_io_eo[62] ,
    \cb_5_1_io_eo[61] ,
    \cb_5_1_io_eo[60] ,
    \cb_5_1_io_eo[59] ,
    \cb_5_1_io_eo[58] ,
    \cb_5_1_io_eo[57] ,
    \cb_5_1_io_eo[56] ,
    \cb_5_1_io_eo[55] ,
    \cb_5_1_io_eo[54] ,
    \cb_5_1_io_eo[53] ,
    \cb_5_1_io_eo[52] ,
    \cb_5_1_io_eo[51] ,
    \cb_5_1_io_eo[50] ,
    \cb_5_1_io_eo[49] ,
    \cb_5_1_io_eo[48] ,
    \cb_5_1_io_eo[47] ,
    \cb_5_1_io_eo[46] ,
    \cb_5_1_io_eo[45] ,
    \cb_5_1_io_eo[44] ,
    \cb_5_1_io_eo[43] ,
    \cb_5_1_io_eo[42] ,
    \cb_5_1_io_eo[41] ,
    \cb_5_1_io_eo[40] ,
    \cb_5_1_io_eo[39] ,
    \cb_5_1_io_eo[38] ,
    \cb_5_1_io_eo[37] ,
    \cb_5_1_io_eo[36] ,
    \cb_5_1_io_eo[35] ,
    \cb_5_1_io_eo[34] ,
    \cb_5_1_io_eo[33] ,
    \cb_5_1_io_eo[32] ,
    \cb_5_1_io_eo[31] ,
    \cb_5_1_io_eo[30] ,
    \cb_5_1_io_eo[29] ,
    \cb_5_1_io_eo[28] ,
    \cb_5_1_io_eo[27] ,
    \cb_5_1_io_eo[26] ,
    \cb_5_1_io_eo[25] ,
    \cb_5_1_io_eo[24] ,
    \cb_5_1_io_eo[23] ,
    \cb_5_1_io_eo[22] ,
    \cb_5_1_io_eo[21] ,
    \cb_5_1_io_eo[20] ,
    \cb_5_1_io_eo[19] ,
    \cb_5_1_io_eo[18] ,
    \cb_5_1_io_eo[17] ,
    \cb_5_1_io_eo[16] ,
    \cb_5_1_io_eo[15] ,
    \cb_5_1_io_eo[14] ,
    \cb_5_1_io_eo[13] ,
    \cb_5_1_io_eo[12] ,
    \cb_5_1_io_eo[11] ,
    \cb_5_1_io_eo[10] ,
    \cb_5_1_io_eo[9] ,
    \cb_5_1_io_eo[8] ,
    \cb_5_1_io_eo[7] ,
    \cb_5_1_io_eo[6] ,
    \cb_5_1_io_eo[5] ,
    \cb_5_1_io_eo[4] ,
    \cb_5_1_io_eo[3] ,
    \cb_5_1_io_eo[2] ,
    \cb_5_1_io_eo[1] ,
    \cb_5_1_io_eo[0] }),
    .io_i_0_in1({\cb_5_0_io_o_0_out[7] ,
    \cb_5_0_io_o_0_out[6] ,
    \cb_5_0_io_o_0_out[5] ,
    \cb_5_0_io_o_0_out[4] ,
    \cb_5_0_io_o_0_out[3] ,
    \cb_5_0_io_o_0_out[2] ,
    \cb_5_0_io_o_0_out[1] ,
    \cb_5_0_io_o_0_out[0] }),
    .io_i_1_in1({\cb_5_0_io_o_1_out[7] ,
    \cb_5_0_io_o_1_out[6] ,
    \cb_5_0_io_o_1_out[5] ,
    \cb_5_0_io_o_1_out[4] ,
    \cb_5_0_io_o_1_out[3] ,
    \cb_5_0_io_o_1_out[2] ,
    \cb_5_0_io_o_1_out[1] ,
    \cb_5_0_io_o_1_out[0] }),
    .io_i_2_in1({\cb_5_0_io_o_2_out[7] ,
    \cb_5_0_io_o_2_out[6] ,
    \cb_5_0_io_o_2_out[5] ,
    \cb_5_0_io_o_2_out[4] ,
    \cb_5_0_io_o_2_out[3] ,
    \cb_5_0_io_o_2_out[2] ,
    \cb_5_0_io_o_2_out[1] ,
    \cb_5_0_io_o_2_out[0] }),
    .io_i_3_in1({\cb_5_0_io_o_3_out[7] ,
    \cb_5_0_io_o_3_out[6] ,
    \cb_5_0_io_o_3_out[5] ,
    \cb_5_0_io_o_3_out[4] ,
    \cb_5_0_io_o_3_out[3] ,
    \cb_5_0_io_o_3_out[2] ,
    \cb_5_0_io_o_3_out[1] ,
    \cb_5_0_io_o_3_out[0] }),
    .io_i_4_in1({\cb_5_0_io_o_4_out[7] ,
    \cb_5_0_io_o_4_out[6] ,
    \cb_5_0_io_o_4_out[5] ,
    \cb_5_0_io_o_4_out[4] ,
    \cb_5_0_io_o_4_out[3] ,
    \cb_5_0_io_o_4_out[2] ,
    \cb_5_0_io_o_4_out[1] ,
    \cb_5_0_io_o_4_out[0] }),
    .io_i_5_in1({\cb_5_0_io_o_5_out[7] ,
    \cb_5_0_io_o_5_out[6] ,
    \cb_5_0_io_o_5_out[5] ,
    \cb_5_0_io_o_5_out[4] ,
    \cb_5_0_io_o_5_out[3] ,
    \cb_5_0_io_o_5_out[2] ,
    \cb_5_0_io_o_5_out[1] ,
    \cb_5_0_io_o_5_out[0] }),
    .io_i_6_in1({\cb_5_0_io_o_6_out[7] ,
    \cb_5_0_io_o_6_out[6] ,
    \cb_5_0_io_o_6_out[5] ,
    \cb_5_0_io_o_6_out[4] ,
    \cb_5_0_io_o_6_out[3] ,
    \cb_5_0_io_o_6_out[2] ,
    \cb_5_0_io_o_6_out[1] ,
    \cb_5_0_io_o_6_out[0] }),
    .io_i_7_in1({\cb_5_0_io_o_7_out[7] ,
    \cb_5_0_io_o_7_out[6] ,
    \cb_5_0_io_o_7_out[5] ,
    \cb_5_0_io_o_7_out[4] ,
    \cb_5_0_io_o_7_out[3] ,
    \cb_5_0_io_o_7_out[2] ,
    \cb_5_0_io_o_7_out[1] ,
    \cb_5_0_io_o_7_out[0] }),
    .io_o_0_out({\cb_5_1_io_o_0_out[7] ,
    \cb_5_1_io_o_0_out[6] ,
    \cb_5_1_io_o_0_out[5] ,
    \cb_5_1_io_o_0_out[4] ,
    \cb_5_1_io_o_0_out[3] ,
    \cb_5_1_io_o_0_out[2] ,
    \cb_5_1_io_o_0_out[1] ,
    \cb_5_1_io_o_0_out[0] }),
    .io_o_1_out({\cb_5_1_io_o_1_out[7] ,
    \cb_5_1_io_o_1_out[6] ,
    \cb_5_1_io_o_1_out[5] ,
    \cb_5_1_io_o_1_out[4] ,
    \cb_5_1_io_o_1_out[3] ,
    \cb_5_1_io_o_1_out[2] ,
    \cb_5_1_io_o_1_out[1] ,
    \cb_5_1_io_o_1_out[0] }),
    .io_o_2_out({\cb_5_1_io_o_2_out[7] ,
    \cb_5_1_io_o_2_out[6] ,
    \cb_5_1_io_o_2_out[5] ,
    \cb_5_1_io_o_2_out[4] ,
    \cb_5_1_io_o_2_out[3] ,
    \cb_5_1_io_o_2_out[2] ,
    \cb_5_1_io_o_2_out[1] ,
    \cb_5_1_io_o_2_out[0] }),
    .io_o_3_out({\cb_5_1_io_o_3_out[7] ,
    \cb_5_1_io_o_3_out[6] ,
    \cb_5_1_io_o_3_out[5] ,
    \cb_5_1_io_o_3_out[4] ,
    \cb_5_1_io_o_3_out[3] ,
    \cb_5_1_io_o_3_out[2] ,
    \cb_5_1_io_o_3_out[1] ,
    \cb_5_1_io_o_3_out[0] }),
    .io_o_4_out({\cb_5_1_io_o_4_out[7] ,
    \cb_5_1_io_o_4_out[6] ,
    \cb_5_1_io_o_4_out[5] ,
    \cb_5_1_io_o_4_out[4] ,
    \cb_5_1_io_o_4_out[3] ,
    \cb_5_1_io_o_4_out[2] ,
    \cb_5_1_io_o_4_out[1] ,
    \cb_5_1_io_o_4_out[0] }),
    .io_o_5_out({\cb_5_1_io_o_5_out[7] ,
    \cb_5_1_io_o_5_out[6] ,
    \cb_5_1_io_o_5_out[5] ,
    \cb_5_1_io_o_5_out[4] ,
    \cb_5_1_io_o_5_out[3] ,
    \cb_5_1_io_o_5_out[2] ,
    \cb_5_1_io_o_5_out[1] ,
    \cb_5_1_io_o_5_out[0] }),
    .io_o_6_out({\cb_5_1_io_o_6_out[7] ,
    \cb_5_1_io_o_6_out[6] ,
    \cb_5_1_io_o_6_out[5] ,
    \cb_5_1_io_o_6_out[4] ,
    \cb_5_1_io_o_6_out[3] ,
    \cb_5_1_io_o_6_out[2] ,
    \cb_5_1_io_o_6_out[1] ,
    \cb_5_1_io_o_6_out[0] }),
    .io_o_7_out({\cb_5_1_io_o_7_out[7] ,
    \cb_5_1_io_o_7_out[6] ,
    \cb_5_1_io_o_7_out[5] ,
    \cb_5_1_io_o_7_out[4] ,
    \cb_5_1_io_o_7_out[3] ,
    \cb_5_1_io_o_7_out[2] ,
    \cb_5_1_io_o_7_out[1] ,
    \cb_5_1_io_o_7_out[0] }),
    .io_wo({\cb_5_0_io_eo[63] ,
    \cb_5_0_io_eo[62] ,
    \cb_5_0_io_eo[61] ,
    \cb_5_0_io_eo[60] ,
    \cb_5_0_io_eo[59] ,
    \cb_5_0_io_eo[58] ,
    \cb_5_0_io_eo[57] ,
    \cb_5_0_io_eo[56] ,
    \cb_5_0_io_eo[55] ,
    \cb_5_0_io_eo[54] ,
    \cb_5_0_io_eo[53] ,
    \cb_5_0_io_eo[52] ,
    \cb_5_0_io_eo[51] ,
    \cb_5_0_io_eo[50] ,
    \cb_5_0_io_eo[49] ,
    \cb_5_0_io_eo[48] ,
    \cb_5_0_io_eo[47] ,
    \cb_5_0_io_eo[46] ,
    \cb_5_0_io_eo[45] ,
    \cb_5_0_io_eo[44] ,
    \cb_5_0_io_eo[43] ,
    \cb_5_0_io_eo[42] ,
    \cb_5_0_io_eo[41] ,
    \cb_5_0_io_eo[40] ,
    \cb_5_0_io_eo[39] ,
    \cb_5_0_io_eo[38] ,
    \cb_5_0_io_eo[37] ,
    \cb_5_0_io_eo[36] ,
    \cb_5_0_io_eo[35] ,
    \cb_5_0_io_eo[34] ,
    \cb_5_0_io_eo[33] ,
    \cb_5_0_io_eo[32] ,
    \cb_5_0_io_eo[31] ,
    \cb_5_0_io_eo[30] ,
    \cb_5_0_io_eo[29] ,
    \cb_5_0_io_eo[28] ,
    \cb_5_0_io_eo[27] ,
    \cb_5_0_io_eo[26] ,
    \cb_5_0_io_eo[25] ,
    \cb_5_0_io_eo[24] ,
    \cb_5_0_io_eo[23] ,
    \cb_5_0_io_eo[22] ,
    \cb_5_0_io_eo[21] ,
    \cb_5_0_io_eo[20] ,
    \cb_5_0_io_eo[19] ,
    \cb_5_0_io_eo[18] ,
    \cb_5_0_io_eo[17] ,
    \cb_5_0_io_eo[16] ,
    \cb_5_0_io_eo[15] ,
    \cb_5_0_io_eo[14] ,
    \cb_5_0_io_eo[13] ,
    \cb_5_0_io_eo[12] ,
    \cb_5_0_io_eo[11] ,
    \cb_5_0_io_eo[10] ,
    \cb_5_0_io_eo[9] ,
    \cb_5_0_io_eo[8] ,
    \cb_5_0_io_eo[7] ,
    \cb_5_0_io_eo[6] ,
    \cb_5_0_io_eo[5] ,
    \cb_5_0_io_eo[4] ,
    \cb_5_0_io_eo[3] ,
    \cb_5_0_io_eo[2] ,
    \cb_5_0_io_eo[1] ,
    \cb_5_0_io_eo[0] }));
 cic_block cb_5_10 (.io_cs_i(cb_5_10_io_cs_i),
    .io_i_0_ci(cb_5_10_io_i_0_ci),
    .io_i_1_ci(cb_5_10_io_i_1_ci),
    .io_i_2_ci(cb_5_10_io_i_2_ci),
    .io_i_3_ci(cb_5_10_io_i_3_ci),
    .io_i_4_ci(cb_5_10_io_i_4_ci),
    .io_i_5_ci(cb_5_10_io_i_5_ci),
    .io_i_6_ci(cb_5_10_io_i_6_ci),
    .io_i_7_ci(cb_5_10_io_i_7_ci),
    .io_o_0_co(cb_5_10_io_o_0_co),
    .io_o_1_co(cb_5_10_io_o_1_co),
    .io_o_2_co(cb_5_10_io_o_2_co),
    .io_o_3_co(cb_5_10_io_o_3_co),
    .io_o_4_co(cb_5_10_io_o_4_co),
    .io_o_5_co(cb_5_10_io_o_5_co),
    .io_o_6_co(cb_5_10_io_o_6_co),
    .io_o_7_co(cb_5_10_io_o_7_co),
    .io_vci(cb_5_10_io_vci),
    .io_vco(cb_5_10_io_vco),
    .io_vi(cb_5_10_io_vi),
    .io_we_i(cb_5_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_5_0_io_adr_i[1] ,
    \cb_5_0_io_adr_i[0] }),
    .io_dat_i({\cb_5_0_io_dat_i[15] ,
    \cb_5_0_io_dat_i[14] ,
    \cb_5_0_io_dat_i[13] ,
    \cb_5_0_io_dat_i[12] ,
    \cb_5_0_io_dat_i[11] ,
    \cb_5_0_io_dat_i[10] ,
    \cb_5_0_io_dat_i[9] ,
    \cb_5_0_io_dat_i[8] ,
    \cb_5_0_io_dat_i[7] ,
    \cb_5_0_io_dat_i[6] ,
    \cb_5_0_io_dat_i[5] ,
    \cb_5_0_io_dat_i[4] ,
    \cb_5_0_io_dat_i[3] ,
    \cb_5_0_io_dat_i[2] ,
    \cb_5_0_io_dat_i[1] ,
    \cb_5_0_io_dat_i[0] }),
    .io_dat_o({\cb_5_10_io_dat_o[15] ,
    \cb_5_10_io_dat_o[14] ,
    \cb_5_10_io_dat_o[13] ,
    \cb_5_10_io_dat_o[12] ,
    \cb_5_10_io_dat_o[11] ,
    \cb_5_10_io_dat_o[10] ,
    \cb_5_10_io_dat_o[9] ,
    \cb_5_10_io_dat_o[8] ,
    \cb_5_10_io_dat_o[7] ,
    \cb_5_10_io_dat_o[6] ,
    \cb_5_10_io_dat_o[5] ,
    \cb_5_10_io_dat_o[4] ,
    \cb_5_10_io_dat_o[3] ,
    \cb_5_10_io_dat_o[2] ,
    \cb_5_10_io_dat_o[1] ,
    \cb_5_10_io_dat_o[0] }),
    .io_eo({\_T_123[31] ,
    \_T_123[30] ,
    \_T_123[29] ,
    \_T_123[28] ,
    \_T_123[27] ,
    \_T_123[26] ,
    \_T_123[25] ,
    \_T_123[24] ,
    \_T_123[23] ,
    \_T_123[22] ,
    \_T_123[21] ,
    \_T_123[20] ,
    \_T_123[19] ,
    \_T_123[18] ,
    \_T_123[17] ,
    \_T_123[16] ,
    \_T_123[15] ,
    \_T_123[14] ,
    \_T_123[13] ,
    \_T_123[12] ,
    \_T_123[11] ,
    \_T_123[10] ,
    \_T_123[9] ,
    \_T_123[8] ,
    \_T_123[7] ,
    \_T_123[6] ,
    \_T_123[5] ,
    \_T_123[4] ,
    \_T_123[3] ,
    \_T_123[2] ,
    \_T_123[1] ,
    \_T_123[0] ,
    \_T_120[31] ,
    \_T_120[30] ,
    \_T_120[29] ,
    \_T_120[28] ,
    \_T_120[27] ,
    \_T_120[26] ,
    \_T_120[25] ,
    \_T_120[24] ,
    \_T_120[23] ,
    \_T_120[22] ,
    \_T_120[21] ,
    \_T_120[20] ,
    \_T_120[19] ,
    \_T_120[18] ,
    \_T_120[17] ,
    \_T_120[16] ,
    \_T_120[15] ,
    \_T_120[14] ,
    \_T_120[13] ,
    \_T_120[12] ,
    \_T_120[11] ,
    \_T_120[10] ,
    \_T_120[9] ,
    \_T_120[8] ,
    \_T_120[7] ,
    \_T_120[6] ,
    \_T_120[5] ,
    \_T_120[4] ,
    \_T_120[3] ,
    \_T_120[2] ,
    \_T_120[1] ,
    \_T_120[0] }),
    .io_i_0_in1({\cb_5_10_io_i_0_in1[7] ,
    \cb_5_10_io_i_0_in1[6] ,
    \cb_5_10_io_i_0_in1[5] ,
    \cb_5_10_io_i_0_in1[4] ,
    \cb_5_10_io_i_0_in1[3] ,
    \cb_5_10_io_i_0_in1[2] ,
    \cb_5_10_io_i_0_in1[1] ,
    \cb_5_10_io_i_0_in1[0] }),
    .io_i_1_in1({\cb_5_10_io_i_1_in1[7] ,
    \cb_5_10_io_i_1_in1[6] ,
    \cb_5_10_io_i_1_in1[5] ,
    \cb_5_10_io_i_1_in1[4] ,
    \cb_5_10_io_i_1_in1[3] ,
    \cb_5_10_io_i_1_in1[2] ,
    \cb_5_10_io_i_1_in1[1] ,
    \cb_5_10_io_i_1_in1[0] }),
    .io_i_2_in1({\cb_5_10_io_i_2_in1[7] ,
    \cb_5_10_io_i_2_in1[6] ,
    \cb_5_10_io_i_2_in1[5] ,
    \cb_5_10_io_i_2_in1[4] ,
    \cb_5_10_io_i_2_in1[3] ,
    \cb_5_10_io_i_2_in1[2] ,
    \cb_5_10_io_i_2_in1[1] ,
    \cb_5_10_io_i_2_in1[0] }),
    .io_i_3_in1({\cb_5_10_io_i_3_in1[7] ,
    \cb_5_10_io_i_3_in1[6] ,
    \cb_5_10_io_i_3_in1[5] ,
    \cb_5_10_io_i_3_in1[4] ,
    \cb_5_10_io_i_3_in1[3] ,
    \cb_5_10_io_i_3_in1[2] ,
    \cb_5_10_io_i_3_in1[1] ,
    \cb_5_10_io_i_3_in1[0] }),
    .io_i_4_in1({\cb_5_10_io_i_4_in1[7] ,
    \cb_5_10_io_i_4_in1[6] ,
    \cb_5_10_io_i_4_in1[5] ,
    \cb_5_10_io_i_4_in1[4] ,
    \cb_5_10_io_i_4_in1[3] ,
    \cb_5_10_io_i_4_in1[2] ,
    \cb_5_10_io_i_4_in1[1] ,
    \cb_5_10_io_i_4_in1[0] }),
    .io_i_5_in1({\cb_5_10_io_i_5_in1[7] ,
    \cb_5_10_io_i_5_in1[6] ,
    \cb_5_10_io_i_5_in1[5] ,
    \cb_5_10_io_i_5_in1[4] ,
    \cb_5_10_io_i_5_in1[3] ,
    \cb_5_10_io_i_5_in1[2] ,
    \cb_5_10_io_i_5_in1[1] ,
    \cb_5_10_io_i_5_in1[0] }),
    .io_i_6_in1({\cb_5_10_io_i_6_in1[7] ,
    \cb_5_10_io_i_6_in1[6] ,
    \cb_5_10_io_i_6_in1[5] ,
    \cb_5_10_io_i_6_in1[4] ,
    \cb_5_10_io_i_6_in1[3] ,
    \cb_5_10_io_i_6_in1[2] ,
    \cb_5_10_io_i_6_in1[1] ,
    \cb_5_10_io_i_6_in1[0] }),
    .io_i_7_in1({\cb_5_10_io_i_7_in1[7] ,
    \cb_5_10_io_i_7_in1[6] ,
    \cb_5_10_io_i_7_in1[5] ,
    \cb_5_10_io_i_7_in1[4] ,
    \cb_5_10_io_i_7_in1[3] ,
    \cb_5_10_io_i_7_in1[2] ,
    \cb_5_10_io_i_7_in1[1] ,
    \cb_5_10_io_i_7_in1[0] }),
    .io_o_0_out({\_T_120[7] ,
    \_T_120[6] ,
    \_T_120[5] ,
    \_T_120[4] ,
    \_T_120[3] ,
    \_T_120[2] ,
    \_T_120[1] ,
    \_T_120[0] }),
    .io_o_1_out({\_T_120[15] ,
    \_T_120[14] ,
    \_T_120[13] ,
    \_T_120[12] ,
    \_T_120[11] ,
    \_T_120[10] ,
    \_T_120[9] ,
    \_T_120[8] }),
    .io_o_2_out({\_T_120[23] ,
    \_T_120[22] ,
    \_T_120[21] ,
    \_T_120[20] ,
    \_T_120[19] ,
    \_T_120[18] ,
    \_T_120[17] ,
    \_T_120[16] }),
    .io_o_3_out({\_T_120[31] ,
    \_T_120[30] ,
    \_T_120[29] ,
    \_T_120[28] ,
    \_T_120[27] ,
    \_T_120[26] ,
    \_T_120[25] ,
    \_T_120[24] }),
    .io_o_4_out({\_T_123[7] ,
    \_T_123[6] ,
    \_T_123[5] ,
    \_T_123[4] ,
    \_T_123[3] ,
    \_T_123[2] ,
    \_T_123[1] ,
    \_T_123[0] }),
    .io_o_5_out({\_T_123[15] ,
    \_T_123[14] ,
    \_T_123[13] ,
    \_T_123[12] ,
    \_T_123[11] ,
    \_T_123[10] ,
    \_T_123[9] ,
    \_T_123[8] }),
    .io_o_6_out({\_T_123[23] ,
    \_T_123[22] ,
    \_T_123[21] ,
    \_T_123[20] ,
    \_T_123[19] ,
    \_T_123[18] ,
    \_T_123[17] ,
    \_T_123[16] }),
    .io_o_7_out({\_T_123[31] ,
    \_T_123[30] ,
    \_T_123[29] ,
    \_T_123[28] ,
    \_T_123[27] ,
    \_T_123[26] ,
    \_T_123[25] ,
    \_T_123[24] }),
    .io_wo({\cb_5_10_io_wo[63] ,
    \cb_5_10_io_wo[62] ,
    \cb_5_10_io_wo[61] ,
    \cb_5_10_io_wo[60] ,
    \cb_5_10_io_wo[59] ,
    \cb_5_10_io_wo[58] ,
    \cb_5_10_io_wo[57] ,
    \cb_5_10_io_wo[56] ,
    \cb_5_10_io_wo[55] ,
    \cb_5_10_io_wo[54] ,
    \cb_5_10_io_wo[53] ,
    \cb_5_10_io_wo[52] ,
    \cb_5_10_io_wo[51] ,
    \cb_5_10_io_wo[50] ,
    \cb_5_10_io_wo[49] ,
    \cb_5_10_io_wo[48] ,
    \cb_5_10_io_wo[47] ,
    \cb_5_10_io_wo[46] ,
    \cb_5_10_io_wo[45] ,
    \cb_5_10_io_wo[44] ,
    \cb_5_10_io_wo[43] ,
    \cb_5_10_io_wo[42] ,
    \cb_5_10_io_wo[41] ,
    \cb_5_10_io_wo[40] ,
    \cb_5_10_io_wo[39] ,
    \cb_5_10_io_wo[38] ,
    \cb_5_10_io_wo[37] ,
    \cb_5_10_io_wo[36] ,
    \cb_5_10_io_wo[35] ,
    \cb_5_10_io_wo[34] ,
    \cb_5_10_io_wo[33] ,
    \cb_5_10_io_wo[32] ,
    \cb_5_10_io_wo[31] ,
    \cb_5_10_io_wo[30] ,
    \cb_5_10_io_wo[29] ,
    \cb_5_10_io_wo[28] ,
    \cb_5_10_io_wo[27] ,
    \cb_5_10_io_wo[26] ,
    \cb_5_10_io_wo[25] ,
    \cb_5_10_io_wo[24] ,
    \cb_5_10_io_wo[23] ,
    \cb_5_10_io_wo[22] ,
    \cb_5_10_io_wo[21] ,
    \cb_5_10_io_wo[20] ,
    \cb_5_10_io_wo[19] ,
    \cb_5_10_io_wo[18] ,
    \cb_5_10_io_wo[17] ,
    \cb_5_10_io_wo[16] ,
    \cb_5_10_io_wo[15] ,
    \cb_5_10_io_wo[14] ,
    \cb_5_10_io_wo[13] ,
    \cb_5_10_io_wo[12] ,
    \cb_5_10_io_wo[11] ,
    \cb_5_10_io_wo[10] ,
    \cb_5_10_io_wo[9] ,
    \cb_5_10_io_wo[8] ,
    \cb_5_10_io_wo[7] ,
    \cb_5_10_io_wo[6] ,
    \cb_5_10_io_wo[5] ,
    \cb_5_10_io_wo[4] ,
    \cb_5_10_io_wo[3] ,
    \cb_5_10_io_wo[2] ,
    \cb_5_10_io_wo[1] ,
    \cb_5_10_io_wo[0] }));
 cic_block cb_5_2 (.io_cs_i(cb_5_2_io_cs_i),
    .io_i_0_ci(cb_5_1_io_o_0_co),
    .io_i_1_ci(cb_5_1_io_o_1_co),
    .io_i_2_ci(cb_5_1_io_o_2_co),
    .io_i_3_ci(cb_5_1_io_o_3_co),
    .io_i_4_ci(cb_5_1_io_o_4_co),
    .io_i_5_ci(cb_5_1_io_o_5_co),
    .io_i_6_ci(cb_5_1_io_o_6_co),
    .io_i_7_ci(cb_5_1_io_o_7_co),
    .io_o_0_co(cb_5_2_io_o_0_co),
    .io_o_1_co(cb_5_2_io_o_1_co),
    .io_o_2_co(cb_5_2_io_o_2_co),
    .io_o_3_co(cb_5_2_io_o_3_co),
    .io_o_4_co(cb_5_2_io_o_4_co),
    .io_o_5_co(cb_5_2_io_o_5_co),
    .io_o_6_co(cb_5_2_io_o_6_co),
    .io_o_7_co(cb_5_2_io_o_7_co),
    .io_vci(cb_5_1_io_vco),
    .io_vco(cb_5_2_io_vco),
    .io_vi(cb_5_2_io_vi),
    .io_we_i(cb_5_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_5_0_io_adr_i[1] ,
    \cb_5_0_io_adr_i[0] }),
    .io_dat_i({\cb_5_0_io_dat_i[15] ,
    \cb_5_0_io_dat_i[14] ,
    \cb_5_0_io_dat_i[13] ,
    \cb_5_0_io_dat_i[12] ,
    \cb_5_0_io_dat_i[11] ,
    \cb_5_0_io_dat_i[10] ,
    \cb_5_0_io_dat_i[9] ,
    \cb_5_0_io_dat_i[8] ,
    \cb_5_0_io_dat_i[7] ,
    \cb_5_0_io_dat_i[6] ,
    \cb_5_0_io_dat_i[5] ,
    \cb_5_0_io_dat_i[4] ,
    \cb_5_0_io_dat_i[3] ,
    \cb_5_0_io_dat_i[2] ,
    \cb_5_0_io_dat_i[1] ,
    \cb_5_0_io_dat_i[0] }),
    .io_dat_o({\cb_5_2_io_dat_o[15] ,
    \cb_5_2_io_dat_o[14] ,
    \cb_5_2_io_dat_o[13] ,
    \cb_5_2_io_dat_o[12] ,
    \cb_5_2_io_dat_o[11] ,
    \cb_5_2_io_dat_o[10] ,
    \cb_5_2_io_dat_o[9] ,
    \cb_5_2_io_dat_o[8] ,
    \cb_5_2_io_dat_o[7] ,
    \cb_5_2_io_dat_o[6] ,
    \cb_5_2_io_dat_o[5] ,
    \cb_5_2_io_dat_o[4] ,
    \cb_5_2_io_dat_o[3] ,
    \cb_5_2_io_dat_o[2] ,
    \cb_5_2_io_dat_o[1] ,
    \cb_5_2_io_dat_o[0] }),
    .io_eo({\cb_5_2_io_eo[63] ,
    \cb_5_2_io_eo[62] ,
    \cb_5_2_io_eo[61] ,
    \cb_5_2_io_eo[60] ,
    \cb_5_2_io_eo[59] ,
    \cb_5_2_io_eo[58] ,
    \cb_5_2_io_eo[57] ,
    \cb_5_2_io_eo[56] ,
    \cb_5_2_io_eo[55] ,
    \cb_5_2_io_eo[54] ,
    \cb_5_2_io_eo[53] ,
    \cb_5_2_io_eo[52] ,
    \cb_5_2_io_eo[51] ,
    \cb_5_2_io_eo[50] ,
    \cb_5_2_io_eo[49] ,
    \cb_5_2_io_eo[48] ,
    \cb_5_2_io_eo[47] ,
    \cb_5_2_io_eo[46] ,
    \cb_5_2_io_eo[45] ,
    \cb_5_2_io_eo[44] ,
    \cb_5_2_io_eo[43] ,
    \cb_5_2_io_eo[42] ,
    \cb_5_2_io_eo[41] ,
    \cb_5_2_io_eo[40] ,
    \cb_5_2_io_eo[39] ,
    \cb_5_2_io_eo[38] ,
    \cb_5_2_io_eo[37] ,
    \cb_5_2_io_eo[36] ,
    \cb_5_2_io_eo[35] ,
    \cb_5_2_io_eo[34] ,
    \cb_5_2_io_eo[33] ,
    \cb_5_2_io_eo[32] ,
    \cb_5_2_io_eo[31] ,
    \cb_5_2_io_eo[30] ,
    \cb_5_2_io_eo[29] ,
    \cb_5_2_io_eo[28] ,
    \cb_5_2_io_eo[27] ,
    \cb_5_2_io_eo[26] ,
    \cb_5_2_io_eo[25] ,
    \cb_5_2_io_eo[24] ,
    \cb_5_2_io_eo[23] ,
    \cb_5_2_io_eo[22] ,
    \cb_5_2_io_eo[21] ,
    \cb_5_2_io_eo[20] ,
    \cb_5_2_io_eo[19] ,
    \cb_5_2_io_eo[18] ,
    \cb_5_2_io_eo[17] ,
    \cb_5_2_io_eo[16] ,
    \cb_5_2_io_eo[15] ,
    \cb_5_2_io_eo[14] ,
    \cb_5_2_io_eo[13] ,
    \cb_5_2_io_eo[12] ,
    \cb_5_2_io_eo[11] ,
    \cb_5_2_io_eo[10] ,
    \cb_5_2_io_eo[9] ,
    \cb_5_2_io_eo[8] ,
    \cb_5_2_io_eo[7] ,
    \cb_5_2_io_eo[6] ,
    \cb_5_2_io_eo[5] ,
    \cb_5_2_io_eo[4] ,
    \cb_5_2_io_eo[3] ,
    \cb_5_2_io_eo[2] ,
    \cb_5_2_io_eo[1] ,
    \cb_5_2_io_eo[0] }),
    .io_i_0_in1({\cb_5_1_io_o_0_out[7] ,
    \cb_5_1_io_o_0_out[6] ,
    \cb_5_1_io_o_0_out[5] ,
    \cb_5_1_io_o_0_out[4] ,
    \cb_5_1_io_o_0_out[3] ,
    \cb_5_1_io_o_0_out[2] ,
    \cb_5_1_io_o_0_out[1] ,
    \cb_5_1_io_o_0_out[0] }),
    .io_i_1_in1({\cb_5_1_io_o_1_out[7] ,
    \cb_5_1_io_o_1_out[6] ,
    \cb_5_1_io_o_1_out[5] ,
    \cb_5_1_io_o_1_out[4] ,
    \cb_5_1_io_o_1_out[3] ,
    \cb_5_1_io_o_1_out[2] ,
    \cb_5_1_io_o_1_out[1] ,
    \cb_5_1_io_o_1_out[0] }),
    .io_i_2_in1({\cb_5_1_io_o_2_out[7] ,
    \cb_5_1_io_o_2_out[6] ,
    \cb_5_1_io_o_2_out[5] ,
    \cb_5_1_io_o_2_out[4] ,
    \cb_5_1_io_o_2_out[3] ,
    \cb_5_1_io_o_2_out[2] ,
    \cb_5_1_io_o_2_out[1] ,
    \cb_5_1_io_o_2_out[0] }),
    .io_i_3_in1({\cb_5_1_io_o_3_out[7] ,
    \cb_5_1_io_o_3_out[6] ,
    \cb_5_1_io_o_3_out[5] ,
    \cb_5_1_io_o_3_out[4] ,
    \cb_5_1_io_o_3_out[3] ,
    \cb_5_1_io_o_3_out[2] ,
    \cb_5_1_io_o_3_out[1] ,
    \cb_5_1_io_o_3_out[0] }),
    .io_i_4_in1({\cb_5_1_io_o_4_out[7] ,
    \cb_5_1_io_o_4_out[6] ,
    \cb_5_1_io_o_4_out[5] ,
    \cb_5_1_io_o_4_out[4] ,
    \cb_5_1_io_o_4_out[3] ,
    \cb_5_1_io_o_4_out[2] ,
    \cb_5_1_io_o_4_out[1] ,
    \cb_5_1_io_o_4_out[0] }),
    .io_i_5_in1({\cb_5_1_io_o_5_out[7] ,
    \cb_5_1_io_o_5_out[6] ,
    \cb_5_1_io_o_5_out[5] ,
    \cb_5_1_io_o_5_out[4] ,
    \cb_5_1_io_o_5_out[3] ,
    \cb_5_1_io_o_5_out[2] ,
    \cb_5_1_io_o_5_out[1] ,
    \cb_5_1_io_o_5_out[0] }),
    .io_i_6_in1({\cb_5_1_io_o_6_out[7] ,
    \cb_5_1_io_o_6_out[6] ,
    \cb_5_1_io_o_6_out[5] ,
    \cb_5_1_io_o_6_out[4] ,
    \cb_5_1_io_o_6_out[3] ,
    \cb_5_1_io_o_6_out[2] ,
    \cb_5_1_io_o_6_out[1] ,
    \cb_5_1_io_o_6_out[0] }),
    .io_i_7_in1({\cb_5_1_io_o_7_out[7] ,
    \cb_5_1_io_o_7_out[6] ,
    \cb_5_1_io_o_7_out[5] ,
    \cb_5_1_io_o_7_out[4] ,
    \cb_5_1_io_o_7_out[3] ,
    \cb_5_1_io_o_7_out[2] ,
    \cb_5_1_io_o_7_out[1] ,
    \cb_5_1_io_o_7_out[0] }),
    .io_o_0_out({\cb_5_2_io_o_0_out[7] ,
    \cb_5_2_io_o_0_out[6] ,
    \cb_5_2_io_o_0_out[5] ,
    \cb_5_2_io_o_0_out[4] ,
    \cb_5_2_io_o_0_out[3] ,
    \cb_5_2_io_o_0_out[2] ,
    \cb_5_2_io_o_0_out[1] ,
    \cb_5_2_io_o_0_out[0] }),
    .io_o_1_out({\cb_5_2_io_o_1_out[7] ,
    \cb_5_2_io_o_1_out[6] ,
    \cb_5_2_io_o_1_out[5] ,
    \cb_5_2_io_o_1_out[4] ,
    \cb_5_2_io_o_1_out[3] ,
    \cb_5_2_io_o_1_out[2] ,
    \cb_5_2_io_o_1_out[1] ,
    \cb_5_2_io_o_1_out[0] }),
    .io_o_2_out({\cb_5_2_io_o_2_out[7] ,
    \cb_5_2_io_o_2_out[6] ,
    \cb_5_2_io_o_2_out[5] ,
    \cb_5_2_io_o_2_out[4] ,
    \cb_5_2_io_o_2_out[3] ,
    \cb_5_2_io_o_2_out[2] ,
    \cb_5_2_io_o_2_out[1] ,
    \cb_5_2_io_o_2_out[0] }),
    .io_o_3_out({\cb_5_2_io_o_3_out[7] ,
    \cb_5_2_io_o_3_out[6] ,
    \cb_5_2_io_o_3_out[5] ,
    \cb_5_2_io_o_3_out[4] ,
    \cb_5_2_io_o_3_out[3] ,
    \cb_5_2_io_o_3_out[2] ,
    \cb_5_2_io_o_3_out[1] ,
    \cb_5_2_io_o_3_out[0] }),
    .io_o_4_out({\cb_5_2_io_o_4_out[7] ,
    \cb_5_2_io_o_4_out[6] ,
    \cb_5_2_io_o_4_out[5] ,
    \cb_5_2_io_o_4_out[4] ,
    \cb_5_2_io_o_4_out[3] ,
    \cb_5_2_io_o_4_out[2] ,
    \cb_5_2_io_o_4_out[1] ,
    \cb_5_2_io_o_4_out[0] }),
    .io_o_5_out({\cb_5_2_io_o_5_out[7] ,
    \cb_5_2_io_o_5_out[6] ,
    \cb_5_2_io_o_5_out[5] ,
    \cb_5_2_io_o_5_out[4] ,
    \cb_5_2_io_o_5_out[3] ,
    \cb_5_2_io_o_5_out[2] ,
    \cb_5_2_io_o_5_out[1] ,
    \cb_5_2_io_o_5_out[0] }),
    .io_o_6_out({\cb_5_2_io_o_6_out[7] ,
    \cb_5_2_io_o_6_out[6] ,
    \cb_5_2_io_o_6_out[5] ,
    \cb_5_2_io_o_6_out[4] ,
    \cb_5_2_io_o_6_out[3] ,
    \cb_5_2_io_o_6_out[2] ,
    \cb_5_2_io_o_6_out[1] ,
    \cb_5_2_io_o_6_out[0] }),
    .io_o_7_out({\cb_5_2_io_o_7_out[7] ,
    \cb_5_2_io_o_7_out[6] ,
    \cb_5_2_io_o_7_out[5] ,
    \cb_5_2_io_o_7_out[4] ,
    \cb_5_2_io_o_7_out[3] ,
    \cb_5_2_io_o_7_out[2] ,
    \cb_5_2_io_o_7_out[1] ,
    \cb_5_2_io_o_7_out[0] }),
    .io_wo({\cb_5_1_io_eo[63] ,
    \cb_5_1_io_eo[62] ,
    \cb_5_1_io_eo[61] ,
    \cb_5_1_io_eo[60] ,
    \cb_5_1_io_eo[59] ,
    \cb_5_1_io_eo[58] ,
    \cb_5_1_io_eo[57] ,
    \cb_5_1_io_eo[56] ,
    \cb_5_1_io_eo[55] ,
    \cb_5_1_io_eo[54] ,
    \cb_5_1_io_eo[53] ,
    \cb_5_1_io_eo[52] ,
    \cb_5_1_io_eo[51] ,
    \cb_5_1_io_eo[50] ,
    \cb_5_1_io_eo[49] ,
    \cb_5_1_io_eo[48] ,
    \cb_5_1_io_eo[47] ,
    \cb_5_1_io_eo[46] ,
    \cb_5_1_io_eo[45] ,
    \cb_5_1_io_eo[44] ,
    \cb_5_1_io_eo[43] ,
    \cb_5_1_io_eo[42] ,
    \cb_5_1_io_eo[41] ,
    \cb_5_1_io_eo[40] ,
    \cb_5_1_io_eo[39] ,
    \cb_5_1_io_eo[38] ,
    \cb_5_1_io_eo[37] ,
    \cb_5_1_io_eo[36] ,
    \cb_5_1_io_eo[35] ,
    \cb_5_1_io_eo[34] ,
    \cb_5_1_io_eo[33] ,
    \cb_5_1_io_eo[32] ,
    \cb_5_1_io_eo[31] ,
    \cb_5_1_io_eo[30] ,
    \cb_5_1_io_eo[29] ,
    \cb_5_1_io_eo[28] ,
    \cb_5_1_io_eo[27] ,
    \cb_5_1_io_eo[26] ,
    \cb_5_1_io_eo[25] ,
    \cb_5_1_io_eo[24] ,
    \cb_5_1_io_eo[23] ,
    \cb_5_1_io_eo[22] ,
    \cb_5_1_io_eo[21] ,
    \cb_5_1_io_eo[20] ,
    \cb_5_1_io_eo[19] ,
    \cb_5_1_io_eo[18] ,
    \cb_5_1_io_eo[17] ,
    \cb_5_1_io_eo[16] ,
    \cb_5_1_io_eo[15] ,
    \cb_5_1_io_eo[14] ,
    \cb_5_1_io_eo[13] ,
    \cb_5_1_io_eo[12] ,
    \cb_5_1_io_eo[11] ,
    \cb_5_1_io_eo[10] ,
    \cb_5_1_io_eo[9] ,
    \cb_5_1_io_eo[8] ,
    \cb_5_1_io_eo[7] ,
    \cb_5_1_io_eo[6] ,
    \cb_5_1_io_eo[5] ,
    \cb_5_1_io_eo[4] ,
    \cb_5_1_io_eo[3] ,
    \cb_5_1_io_eo[2] ,
    \cb_5_1_io_eo[1] ,
    \cb_5_1_io_eo[0] }));
 cic_block cb_5_3 (.io_cs_i(cb_5_3_io_cs_i),
    .io_i_0_ci(cb_5_2_io_o_0_co),
    .io_i_1_ci(cb_5_2_io_o_1_co),
    .io_i_2_ci(cb_5_2_io_o_2_co),
    .io_i_3_ci(cb_5_2_io_o_3_co),
    .io_i_4_ci(cb_5_2_io_o_4_co),
    .io_i_5_ci(cb_5_2_io_o_5_co),
    .io_i_6_ci(cb_5_2_io_o_6_co),
    .io_i_7_ci(cb_5_2_io_o_7_co),
    .io_o_0_co(cb_5_3_io_o_0_co),
    .io_o_1_co(cb_5_3_io_o_1_co),
    .io_o_2_co(cb_5_3_io_o_2_co),
    .io_o_3_co(cb_5_3_io_o_3_co),
    .io_o_4_co(cb_5_3_io_o_4_co),
    .io_o_5_co(cb_5_3_io_o_5_co),
    .io_o_6_co(cb_5_3_io_o_6_co),
    .io_o_7_co(cb_5_3_io_o_7_co),
    .io_vci(cb_5_2_io_vco),
    .io_vco(cb_5_3_io_vco),
    .io_vi(cb_5_3_io_vi),
    .io_we_i(cb_5_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_5_0_io_adr_i[1] ,
    \cb_5_0_io_adr_i[0] }),
    .io_dat_i({\cb_5_0_io_dat_i[15] ,
    \cb_5_0_io_dat_i[14] ,
    \cb_5_0_io_dat_i[13] ,
    \cb_5_0_io_dat_i[12] ,
    \cb_5_0_io_dat_i[11] ,
    \cb_5_0_io_dat_i[10] ,
    \cb_5_0_io_dat_i[9] ,
    \cb_5_0_io_dat_i[8] ,
    \cb_5_0_io_dat_i[7] ,
    \cb_5_0_io_dat_i[6] ,
    \cb_5_0_io_dat_i[5] ,
    \cb_5_0_io_dat_i[4] ,
    \cb_5_0_io_dat_i[3] ,
    \cb_5_0_io_dat_i[2] ,
    \cb_5_0_io_dat_i[1] ,
    \cb_5_0_io_dat_i[0] }),
    .io_dat_o({\cb_5_3_io_dat_o[15] ,
    \cb_5_3_io_dat_o[14] ,
    \cb_5_3_io_dat_o[13] ,
    \cb_5_3_io_dat_o[12] ,
    \cb_5_3_io_dat_o[11] ,
    \cb_5_3_io_dat_o[10] ,
    \cb_5_3_io_dat_o[9] ,
    \cb_5_3_io_dat_o[8] ,
    \cb_5_3_io_dat_o[7] ,
    \cb_5_3_io_dat_o[6] ,
    \cb_5_3_io_dat_o[5] ,
    \cb_5_3_io_dat_o[4] ,
    \cb_5_3_io_dat_o[3] ,
    \cb_5_3_io_dat_o[2] ,
    \cb_5_3_io_dat_o[1] ,
    \cb_5_3_io_dat_o[0] }),
    .io_eo({\cb_5_3_io_eo[63] ,
    \cb_5_3_io_eo[62] ,
    \cb_5_3_io_eo[61] ,
    \cb_5_3_io_eo[60] ,
    \cb_5_3_io_eo[59] ,
    \cb_5_3_io_eo[58] ,
    \cb_5_3_io_eo[57] ,
    \cb_5_3_io_eo[56] ,
    \cb_5_3_io_eo[55] ,
    \cb_5_3_io_eo[54] ,
    \cb_5_3_io_eo[53] ,
    \cb_5_3_io_eo[52] ,
    \cb_5_3_io_eo[51] ,
    \cb_5_3_io_eo[50] ,
    \cb_5_3_io_eo[49] ,
    \cb_5_3_io_eo[48] ,
    \cb_5_3_io_eo[47] ,
    \cb_5_3_io_eo[46] ,
    \cb_5_3_io_eo[45] ,
    \cb_5_3_io_eo[44] ,
    \cb_5_3_io_eo[43] ,
    \cb_5_3_io_eo[42] ,
    \cb_5_3_io_eo[41] ,
    \cb_5_3_io_eo[40] ,
    \cb_5_3_io_eo[39] ,
    \cb_5_3_io_eo[38] ,
    \cb_5_3_io_eo[37] ,
    \cb_5_3_io_eo[36] ,
    \cb_5_3_io_eo[35] ,
    \cb_5_3_io_eo[34] ,
    \cb_5_3_io_eo[33] ,
    \cb_5_3_io_eo[32] ,
    \cb_5_3_io_eo[31] ,
    \cb_5_3_io_eo[30] ,
    \cb_5_3_io_eo[29] ,
    \cb_5_3_io_eo[28] ,
    \cb_5_3_io_eo[27] ,
    \cb_5_3_io_eo[26] ,
    \cb_5_3_io_eo[25] ,
    \cb_5_3_io_eo[24] ,
    \cb_5_3_io_eo[23] ,
    \cb_5_3_io_eo[22] ,
    \cb_5_3_io_eo[21] ,
    \cb_5_3_io_eo[20] ,
    \cb_5_3_io_eo[19] ,
    \cb_5_3_io_eo[18] ,
    \cb_5_3_io_eo[17] ,
    \cb_5_3_io_eo[16] ,
    \cb_5_3_io_eo[15] ,
    \cb_5_3_io_eo[14] ,
    \cb_5_3_io_eo[13] ,
    \cb_5_3_io_eo[12] ,
    \cb_5_3_io_eo[11] ,
    \cb_5_3_io_eo[10] ,
    \cb_5_3_io_eo[9] ,
    \cb_5_3_io_eo[8] ,
    \cb_5_3_io_eo[7] ,
    \cb_5_3_io_eo[6] ,
    \cb_5_3_io_eo[5] ,
    \cb_5_3_io_eo[4] ,
    \cb_5_3_io_eo[3] ,
    \cb_5_3_io_eo[2] ,
    \cb_5_3_io_eo[1] ,
    \cb_5_3_io_eo[0] }),
    .io_i_0_in1({\cb_5_2_io_o_0_out[7] ,
    \cb_5_2_io_o_0_out[6] ,
    \cb_5_2_io_o_0_out[5] ,
    \cb_5_2_io_o_0_out[4] ,
    \cb_5_2_io_o_0_out[3] ,
    \cb_5_2_io_o_0_out[2] ,
    \cb_5_2_io_o_0_out[1] ,
    \cb_5_2_io_o_0_out[0] }),
    .io_i_1_in1({\cb_5_2_io_o_1_out[7] ,
    \cb_5_2_io_o_1_out[6] ,
    \cb_5_2_io_o_1_out[5] ,
    \cb_5_2_io_o_1_out[4] ,
    \cb_5_2_io_o_1_out[3] ,
    \cb_5_2_io_o_1_out[2] ,
    \cb_5_2_io_o_1_out[1] ,
    \cb_5_2_io_o_1_out[0] }),
    .io_i_2_in1({\cb_5_2_io_o_2_out[7] ,
    \cb_5_2_io_o_2_out[6] ,
    \cb_5_2_io_o_2_out[5] ,
    \cb_5_2_io_o_2_out[4] ,
    \cb_5_2_io_o_2_out[3] ,
    \cb_5_2_io_o_2_out[2] ,
    \cb_5_2_io_o_2_out[1] ,
    \cb_5_2_io_o_2_out[0] }),
    .io_i_3_in1({\cb_5_2_io_o_3_out[7] ,
    \cb_5_2_io_o_3_out[6] ,
    \cb_5_2_io_o_3_out[5] ,
    \cb_5_2_io_o_3_out[4] ,
    \cb_5_2_io_o_3_out[3] ,
    \cb_5_2_io_o_3_out[2] ,
    \cb_5_2_io_o_3_out[1] ,
    \cb_5_2_io_o_3_out[0] }),
    .io_i_4_in1({\cb_5_2_io_o_4_out[7] ,
    \cb_5_2_io_o_4_out[6] ,
    \cb_5_2_io_o_4_out[5] ,
    \cb_5_2_io_o_4_out[4] ,
    \cb_5_2_io_o_4_out[3] ,
    \cb_5_2_io_o_4_out[2] ,
    \cb_5_2_io_o_4_out[1] ,
    \cb_5_2_io_o_4_out[0] }),
    .io_i_5_in1({\cb_5_2_io_o_5_out[7] ,
    \cb_5_2_io_o_5_out[6] ,
    \cb_5_2_io_o_5_out[5] ,
    \cb_5_2_io_o_5_out[4] ,
    \cb_5_2_io_o_5_out[3] ,
    \cb_5_2_io_o_5_out[2] ,
    \cb_5_2_io_o_5_out[1] ,
    \cb_5_2_io_o_5_out[0] }),
    .io_i_6_in1({\cb_5_2_io_o_6_out[7] ,
    \cb_5_2_io_o_6_out[6] ,
    \cb_5_2_io_o_6_out[5] ,
    \cb_5_2_io_o_6_out[4] ,
    \cb_5_2_io_o_6_out[3] ,
    \cb_5_2_io_o_6_out[2] ,
    \cb_5_2_io_o_6_out[1] ,
    \cb_5_2_io_o_6_out[0] }),
    .io_i_7_in1({\cb_5_2_io_o_7_out[7] ,
    \cb_5_2_io_o_7_out[6] ,
    \cb_5_2_io_o_7_out[5] ,
    \cb_5_2_io_o_7_out[4] ,
    \cb_5_2_io_o_7_out[3] ,
    \cb_5_2_io_o_7_out[2] ,
    \cb_5_2_io_o_7_out[1] ,
    \cb_5_2_io_o_7_out[0] }),
    .io_o_0_out({\cb_5_3_io_o_0_out[7] ,
    \cb_5_3_io_o_0_out[6] ,
    \cb_5_3_io_o_0_out[5] ,
    \cb_5_3_io_o_0_out[4] ,
    \cb_5_3_io_o_0_out[3] ,
    \cb_5_3_io_o_0_out[2] ,
    \cb_5_3_io_o_0_out[1] ,
    \cb_5_3_io_o_0_out[0] }),
    .io_o_1_out({\cb_5_3_io_o_1_out[7] ,
    \cb_5_3_io_o_1_out[6] ,
    \cb_5_3_io_o_1_out[5] ,
    \cb_5_3_io_o_1_out[4] ,
    \cb_5_3_io_o_1_out[3] ,
    \cb_5_3_io_o_1_out[2] ,
    \cb_5_3_io_o_1_out[1] ,
    \cb_5_3_io_o_1_out[0] }),
    .io_o_2_out({\cb_5_3_io_o_2_out[7] ,
    \cb_5_3_io_o_2_out[6] ,
    \cb_5_3_io_o_2_out[5] ,
    \cb_5_3_io_o_2_out[4] ,
    \cb_5_3_io_o_2_out[3] ,
    \cb_5_3_io_o_2_out[2] ,
    \cb_5_3_io_o_2_out[1] ,
    \cb_5_3_io_o_2_out[0] }),
    .io_o_3_out({\cb_5_3_io_o_3_out[7] ,
    \cb_5_3_io_o_3_out[6] ,
    \cb_5_3_io_o_3_out[5] ,
    \cb_5_3_io_o_3_out[4] ,
    \cb_5_3_io_o_3_out[3] ,
    \cb_5_3_io_o_3_out[2] ,
    \cb_5_3_io_o_3_out[1] ,
    \cb_5_3_io_o_3_out[0] }),
    .io_o_4_out({\cb_5_3_io_o_4_out[7] ,
    \cb_5_3_io_o_4_out[6] ,
    \cb_5_3_io_o_4_out[5] ,
    \cb_5_3_io_o_4_out[4] ,
    \cb_5_3_io_o_4_out[3] ,
    \cb_5_3_io_o_4_out[2] ,
    \cb_5_3_io_o_4_out[1] ,
    \cb_5_3_io_o_4_out[0] }),
    .io_o_5_out({\cb_5_3_io_o_5_out[7] ,
    \cb_5_3_io_o_5_out[6] ,
    \cb_5_3_io_o_5_out[5] ,
    \cb_5_3_io_o_5_out[4] ,
    \cb_5_3_io_o_5_out[3] ,
    \cb_5_3_io_o_5_out[2] ,
    \cb_5_3_io_o_5_out[1] ,
    \cb_5_3_io_o_5_out[0] }),
    .io_o_6_out({\cb_5_3_io_o_6_out[7] ,
    \cb_5_3_io_o_6_out[6] ,
    \cb_5_3_io_o_6_out[5] ,
    \cb_5_3_io_o_6_out[4] ,
    \cb_5_3_io_o_6_out[3] ,
    \cb_5_3_io_o_6_out[2] ,
    \cb_5_3_io_o_6_out[1] ,
    \cb_5_3_io_o_6_out[0] }),
    .io_o_7_out({\cb_5_3_io_o_7_out[7] ,
    \cb_5_3_io_o_7_out[6] ,
    \cb_5_3_io_o_7_out[5] ,
    \cb_5_3_io_o_7_out[4] ,
    \cb_5_3_io_o_7_out[3] ,
    \cb_5_3_io_o_7_out[2] ,
    \cb_5_3_io_o_7_out[1] ,
    \cb_5_3_io_o_7_out[0] }),
    .io_wo({\cb_5_2_io_eo[63] ,
    \cb_5_2_io_eo[62] ,
    \cb_5_2_io_eo[61] ,
    \cb_5_2_io_eo[60] ,
    \cb_5_2_io_eo[59] ,
    \cb_5_2_io_eo[58] ,
    \cb_5_2_io_eo[57] ,
    \cb_5_2_io_eo[56] ,
    \cb_5_2_io_eo[55] ,
    \cb_5_2_io_eo[54] ,
    \cb_5_2_io_eo[53] ,
    \cb_5_2_io_eo[52] ,
    \cb_5_2_io_eo[51] ,
    \cb_5_2_io_eo[50] ,
    \cb_5_2_io_eo[49] ,
    \cb_5_2_io_eo[48] ,
    \cb_5_2_io_eo[47] ,
    \cb_5_2_io_eo[46] ,
    \cb_5_2_io_eo[45] ,
    \cb_5_2_io_eo[44] ,
    \cb_5_2_io_eo[43] ,
    \cb_5_2_io_eo[42] ,
    \cb_5_2_io_eo[41] ,
    \cb_5_2_io_eo[40] ,
    \cb_5_2_io_eo[39] ,
    \cb_5_2_io_eo[38] ,
    \cb_5_2_io_eo[37] ,
    \cb_5_2_io_eo[36] ,
    \cb_5_2_io_eo[35] ,
    \cb_5_2_io_eo[34] ,
    \cb_5_2_io_eo[33] ,
    \cb_5_2_io_eo[32] ,
    \cb_5_2_io_eo[31] ,
    \cb_5_2_io_eo[30] ,
    \cb_5_2_io_eo[29] ,
    \cb_5_2_io_eo[28] ,
    \cb_5_2_io_eo[27] ,
    \cb_5_2_io_eo[26] ,
    \cb_5_2_io_eo[25] ,
    \cb_5_2_io_eo[24] ,
    \cb_5_2_io_eo[23] ,
    \cb_5_2_io_eo[22] ,
    \cb_5_2_io_eo[21] ,
    \cb_5_2_io_eo[20] ,
    \cb_5_2_io_eo[19] ,
    \cb_5_2_io_eo[18] ,
    \cb_5_2_io_eo[17] ,
    \cb_5_2_io_eo[16] ,
    \cb_5_2_io_eo[15] ,
    \cb_5_2_io_eo[14] ,
    \cb_5_2_io_eo[13] ,
    \cb_5_2_io_eo[12] ,
    \cb_5_2_io_eo[11] ,
    \cb_5_2_io_eo[10] ,
    \cb_5_2_io_eo[9] ,
    \cb_5_2_io_eo[8] ,
    \cb_5_2_io_eo[7] ,
    \cb_5_2_io_eo[6] ,
    \cb_5_2_io_eo[5] ,
    \cb_5_2_io_eo[4] ,
    \cb_5_2_io_eo[3] ,
    \cb_5_2_io_eo[2] ,
    \cb_5_2_io_eo[1] ,
    \cb_5_2_io_eo[0] }));
 cic_block cb_5_4 (.io_cs_i(cb_5_4_io_cs_i),
    .io_i_0_ci(cb_5_3_io_o_0_co),
    .io_i_1_ci(cb_5_3_io_o_1_co),
    .io_i_2_ci(cb_5_3_io_o_2_co),
    .io_i_3_ci(cb_5_3_io_o_3_co),
    .io_i_4_ci(cb_5_3_io_o_4_co),
    .io_i_5_ci(cb_5_3_io_o_5_co),
    .io_i_6_ci(cb_5_3_io_o_6_co),
    .io_i_7_ci(cb_5_3_io_o_7_co),
    .io_o_0_co(cb_5_4_io_o_0_co),
    .io_o_1_co(cb_5_4_io_o_1_co),
    .io_o_2_co(cb_5_4_io_o_2_co),
    .io_o_3_co(cb_5_4_io_o_3_co),
    .io_o_4_co(cb_5_4_io_o_4_co),
    .io_o_5_co(cb_5_4_io_o_5_co),
    .io_o_6_co(cb_5_4_io_o_6_co),
    .io_o_7_co(cb_5_4_io_o_7_co),
    .io_vci(cb_5_3_io_vco),
    .io_vco(cb_5_4_io_vco),
    .io_vi(cb_5_4_io_vi),
    .io_we_i(cb_5_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_5_0_io_adr_i[1] ,
    \cb_5_0_io_adr_i[0] }),
    .io_dat_i({\cb_5_0_io_dat_i[15] ,
    \cb_5_0_io_dat_i[14] ,
    \cb_5_0_io_dat_i[13] ,
    \cb_5_0_io_dat_i[12] ,
    \cb_5_0_io_dat_i[11] ,
    \cb_5_0_io_dat_i[10] ,
    \cb_5_0_io_dat_i[9] ,
    \cb_5_0_io_dat_i[8] ,
    \cb_5_0_io_dat_i[7] ,
    \cb_5_0_io_dat_i[6] ,
    \cb_5_0_io_dat_i[5] ,
    \cb_5_0_io_dat_i[4] ,
    \cb_5_0_io_dat_i[3] ,
    \cb_5_0_io_dat_i[2] ,
    \cb_5_0_io_dat_i[1] ,
    \cb_5_0_io_dat_i[0] }),
    .io_dat_o({\cb_5_4_io_dat_o[15] ,
    \cb_5_4_io_dat_o[14] ,
    \cb_5_4_io_dat_o[13] ,
    \cb_5_4_io_dat_o[12] ,
    \cb_5_4_io_dat_o[11] ,
    \cb_5_4_io_dat_o[10] ,
    \cb_5_4_io_dat_o[9] ,
    \cb_5_4_io_dat_o[8] ,
    \cb_5_4_io_dat_o[7] ,
    \cb_5_4_io_dat_o[6] ,
    \cb_5_4_io_dat_o[5] ,
    \cb_5_4_io_dat_o[4] ,
    \cb_5_4_io_dat_o[3] ,
    \cb_5_4_io_dat_o[2] ,
    \cb_5_4_io_dat_o[1] ,
    \cb_5_4_io_dat_o[0] }),
    .io_eo({\cb_5_4_io_eo[63] ,
    \cb_5_4_io_eo[62] ,
    \cb_5_4_io_eo[61] ,
    \cb_5_4_io_eo[60] ,
    \cb_5_4_io_eo[59] ,
    \cb_5_4_io_eo[58] ,
    \cb_5_4_io_eo[57] ,
    \cb_5_4_io_eo[56] ,
    \cb_5_4_io_eo[55] ,
    \cb_5_4_io_eo[54] ,
    \cb_5_4_io_eo[53] ,
    \cb_5_4_io_eo[52] ,
    \cb_5_4_io_eo[51] ,
    \cb_5_4_io_eo[50] ,
    \cb_5_4_io_eo[49] ,
    \cb_5_4_io_eo[48] ,
    \cb_5_4_io_eo[47] ,
    \cb_5_4_io_eo[46] ,
    \cb_5_4_io_eo[45] ,
    \cb_5_4_io_eo[44] ,
    \cb_5_4_io_eo[43] ,
    \cb_5_4_io_eo[42] ,
    \cb_5_4_io_eo[41] ,
    \cb_5_4_io_eo[40] ,
    \cb_5_4_io_eo[39] ,
    \cb_5_4_io_eo[38] ,
    \cb_5_4_io_eo[37] ,
    \cb_5_4_io_eo[36] ,
    \cb_5_4_io_eo[35] ,
    \cb_5_4_io_eo[34] ,
    \cb_5_4_io_eo[33] ,
    \cb_5_4_io_eo[32] ,
    \cb_5_4_io_eo[31] ,
    \cb_5_4_io_eo[30] ,
    \cb_5_4_io_eo[29] ,
    \cb_5_4_io_eo[28] ,
    \cb_5_4_io_eo[27] ,
    \cb_5_4_io_eo[26] ,
    \cb_5_4_io_eo[25] ,
    \cb_5_4_io_eo[24] ,
    \cb_5_4_io_eo[23] ,
    \cb_5_4_io_eo[22] ,
    \cb_5_4_io_eo[21] ,
    \cb_5_4_io_eo[20] ,
    \cb_5_4_io_eo[19] ,
    \cb_5_4_io_eo[18] ,
    \cb_5_4_io_eo[17] ,
    \cb_5_4_io_eo[16] ,
    \cb_5_4_io_eo[15] ,
    \cb_5_4_io_eo[14] ,
    \cb_5_4_io_eo[13] ,
    \cb_5_4_io_eo[12] ,
    \cb_5_4_io_eo[11] ,
    \cb_5_4_io_eo[10] ,
    \cb_5_4_io_eo[9] ,
    \cb_5_4_io_eo[8] ,
    \cb_5_4_io_eo[7] ,
    \cb_5_4_io_eo[6] ,
    \cb_5_4_io_eo[5] ,
    \cb_5_4_io_eo[4] ,
    \cb_5_4_io_eo[3] ,
    \cb_5_4_io_eo[2] ,
    \cb_5_4_io_eo[1] ,
    \cb_5_4_io_eo[0] }),
    .io_i_0_in1({\cb_5_3_io_o_0_out[7] ,
    \cb_5_3_io_o_0_out[6] ,
    \cb_5_3_io_o_0_out[5] ,
    \cb_5_3_io_o_0_out[4] ,
    \cb_5_3_io_o_0_out[3] ,
    \cb_5_3_io_o_0_out[2] ,
    \cb_5_3_io_o_0_out[1] ,
    \cb_5_3_io_o_0_out[0] }),
    .io_i_1_in1({\cb_5_3_io_o_1_out[7] ,
    \cb_5_3_io_o_1_out[6] ,
    \cb_5_3_io_o_1_out[5] ,
    \cb_5_3_io_o_1_out[4] ,
    \cb_5_3_io_o_1_out[3] ,
    \cb_5_3_io_o_1_out[2] ,
    \cb_5_3_io_o_1_out[1] ,
    \cb_5_3_io_o_1_out[0] }),
    .io_i_2_in1({\cb_5_3_io_o_2_out[7] ,
    \cb_5_3_io_o_2_out[6] ,
    \cb_5_3_io_o_2_out[5] ,
    \cb_5_3_io_o_2_out[4] ,
    \cb_5_3_io_o_2_out[3] ,
    \cb_5_3_io_o_2_out[2] ,
    \cb_5_3_io_o_2_out[1] ,
    \cb_5_3_io_o_2_out[0] }),
    .io_i_3_in1({\cb_5_3_io_o_3_out[7] ,
    \cb_5_3_io_o_3_out[6] ,
    \cb_5_3_io_o_3_out[5] ,
    \cb_5_3_io_o_3_out[4] ,
    \cb_5_3_io_o_3_out[3] ,
    \cb_5_3_io_o_3_out[2] ,
    \cb_5_3_io_o_3_out[1] ,
    \cb_5_3_io_o_3_out[0] }),
    .io_i_4_in1({\cb_5_3_io_o_4_out[7] ,
    \cb_5_3_io_o_4_out[6] ,
    \cb_5_3_io_o_4_out[5] ,
    \cb_5_3_io_o_4_out[4] ,
    \cb_5_3_io_o_4_out[3] ,
    \cb_5_3_io_o_4_out[2] ,
    \cb_5_3_io_o_4_out[1] ,
    \cb_5_3_io_o_4_out[0] }),
    .io_i_5_in1({\cb_5_3_io_o_5_out[7] ,
    \cb_5_3_io_o_5_out[6] ,
    \cb_5_3_io_o_5_out[5] ,
    \cb_5_3_io_o_5_out[4] ,
    \cb_5_3_io_o_5_out[3] ,
    \cb_5_3_io_o_5_out[2] ,
    \cb_5_3_io_o_5_out[1] ,
    \cb_5_3_io_o_5_out[0] }),
    .io_i_6_in1({\cb_5_3_io_o_6_out[7] ,
    \cb_5_3_io_o_6_out[6] ,
    \cb_5_3_io_o_6_out[5] ,
    \cb_5_3_io_o_6_out[4] ,
    \cb_5_3_io_o_6_out[3] ,
    \cb_5_3_io_o_6_out[2] ,
    \cb_5_3_io_o_6_out[1] ,
    \cb_5_3_io_o_6_out[0] }),
    .io_i_7_in1({\cb_5_3_io_o_7_out[7] ,
    \cb_5_3_io_o_7_out[6] ,
    \cb_5_3_io_o_7_out[5] ,
    \cb_5_3_io_o_7_out[4] ,
    \cb_5_3_io_o_7_out[3] ,
    \cb_5_3_io_o_7_out[2] ,
    \cb_5_3_io_o_7_out[1] ,
    \cb_5_3_io_o_7_out[0] }),
    .io_o_0_out({\cb_5_4_io_o_0_out[7] ,
    \cb_5_4_io_o_0_out[6] ,
    \cb_5_4_io_o_0_out[5] ,
    \cb_5_4_io_o_0_out[4] ,
    \cb_5_4_io_o_0_out[3] ,
    \cb_5_4_io_o_0_out[2] ,
    \cb_5_4_io_o_0_out[1] ,
    \cb_5_4_io_o_0_out[0] }),
    .io_o_1_out({\cb_5_4_io_o_1_out[7] ,
    \cb_5_4_io_o_1_out[6] ,
    \cb_5_4_io_o_1_out[5] ,
    \cb_5_4_io_o_1_out[4] ,
    \cb_5_4_io_o_1_out[3] ,
    \cb_5_4_io_o_1_out[2] ,
    \cb_5_4_io_o_1_out[1] ,
    \cb_5_4_io_o_1_out[0] }),
    .io_o_2_out({\cb_5_4_io_o_2_out[7] ,
    \cb_5_4_io_o_2_out[6] ,
    \cb_5_4_io_o_2_out[5] ,
    \cb_5_4_io_o_2_out[4] ,
    \cb_5_4_io_o_2_out[3] ,
    \cb_5_4_io_o_2_out[2] ,
    \cb_5_4_io_o_2_out[1] ,
    \cb_5_4_io_o_2_out[0] }),
    .io_o_3_out({\cb_5_4_io_o_3_out[7] ,
    \cb_5_4_io_o_3_out[6] ,
    \cb_5_4_io_o_3_out[5] ,
    \cb_5_4_io_o_3_out[4] ,
    \cb_5_4_io_o_3_out[3] ,
    \cb_5_4_io_o_3_out[2] ,
    \cb_5_4_io_o_3_out[1] ,
    \cb_5_4_io_o_3_out[0] }),
    .io_o_4_out({\cb_5_4_io_o_4_out[7] ,
    \cb_5_4_io_o_4_out[6] ,
    \cb_5_4_io_o_4_out[5] ,
    \cb_5_4_io_o_4_out[4] ,
    \cb_5_4_io_o_4_out[3] ,
    \cb_5_4_io_o_4_out[2] ,
    \cb_5_4_io_o_4_out[1] ,
    \cb_5_4_io_o_4_out[0] }),
    .io_o_5_out({\cb_5_4_io_o_5_out[7] ,
    \cb_5_4_io_o_5_out[6] ,
    \cb_5_4_io_o_5_out[5] ,
    \cb_5_4_io_o_5_out[4] ,
    \cb_5_4_io_o_5_out[3] ,
    \cb_5_4_io_o_5_out[2] ,
    \cb_5_4_io_o_5_out[1] ,
    \cb_5_4_io_o_5_out[0] }),
    .io_o_6_out({\cb_5_4_io_o_6_out[7] ,
    \cb_5_4_io_o_6_out[6] ,
    \cb_5_4_io_o_6_out[5] ,
    \cb_5_4_io_o_6_out[4] ,
    \cb_5_4_io_o_6_out[3] ,
    \cb_5_4_io_o_6_out[2] ,
    \cb_5_4_io_o_6_out[1] ,
    \cb_5_4_io_o_6_out[0] }),
    .io_o_7_out({\cb_5_4_io_o_7_out[7] ,
    \cb_5_4_io_o_7_out[6] ,
    \cb_5_4_io_o_7_out[5] ,
    \cb_5_4_io_o_7_out[4] ,
    \cb_5_4_io_o_7_out[3] ,
    \cb_5_4_io_o_7_out[2] ,
    \cb_5_4_io_o_7_out[1] ,
    \cb_5_4_io_o_7_out[0] }),
    .io_wo({\cb_5_3_io_eo[63] ,
    \cb_5_3_io_eo[62] ,
    \cb_5_3_io_eo[61] ,
    \cb_5_3_io_eo[60] ,
    \cb_5_3_io_eo[59] ,
    \cb_5_3_io_eo[58] ,
    \cb_5_3_io_eo[57] ,
    \cb_5_3_io_eo[56] ,
    \cb_5_3_io_eo[55] ,
    \cb_5_3_io_eo[54] ,
    \cb_5_3_io_eo[53] ,
    \cb_5_3_io_eo[52] ,
    \cb_5_3_io_eo[51] ,
    \cb_5_3_io_eo[50] ,
    \cb_5_3_io_eo[49] ,
    \cb_5_3_io_eo[48] ,
    \cb_5_3_io_eo[47] ,
    \cb_5_3_io_eo[46] ,
    \cb_5_3_io_eo[45] ,
    \cb_5_3_io_eo[44] ,
    \cb_5_3_io_eo[43] ,
    \cb_5_3_io_eo[42] ,
    \cb_5_3_io_eo[41] ,
    \cb_5_3_io_eo[40] ,
    \cb_5_3_io_eo[39] ,
    \cb_5_3_io_eo[38] ,
    \cb_5_3_io_eo[37] ,
    \cb_5_3_io_eo[36] ,
    \cb_5_3_io_eo[35] ,
    \cb_5_3_io_eo[34] ,
    \cb_5_3_io_eo[33] ,
    \cb_5_3_io_eo[32] ,
    \cb_5_3_io_eo[31] ,
    \cb_5_3_io_eo[30] ,
    \cb_5_3_io_eo[29] ,
    \cb_5_3_io_eo[28] ,
    \cb_5_3_io_eo[27] ,
    \cb_5_3_io_eo[26] ,
    \cb_5_3_io_eo[25] ,
    \cb_5_3_io_eo[24] ,
    \cb_5_3_io_eo[23] ,
    \cb_5_3_io_eo[22] ,
    \cb_5_3_io_eo[21] ,
    \cb_5_3_io_eo[20] ,
    \cb_5_3_io_eo[19] ,
    \cb_5_3_io_eo[18] ,
    \cb_5_3_io_eo[17] ,
    \cb_5_3_io_eo[16] ,
    \cb_5_3_io_eo[15] ,
    \cb_5_3_io_eo[14] ,
    \cb_5_3_io_eo[13] ,
    \cb_5_3_io_eo[12] ,
    \cb_5_3_io_eo[11] ,
    \cb_5_3_io_eo[10] ,
    \cb_5_3_io_eo[9] ,
    \cb_5_3_io_eo[8] ,
    \cb_5_3_io_eo[7] ,
    \cb_5_3_io_eo[6] ,
    \cb_5_3_io_eo[5] ,
    \cb_5_3_io_eo[4] ,
    \cb_5_3_io_eo[3] ,
    \cb_5_3_io_eo[2] ,
    \cb_5_3_io_eo[1] ,
    \cb_5_3_io_eo[0] }));
 cic_block cb_5_5 (.io_cs_i(cb_5_5_io_cs_i),
    .io_i_0_ci(cb_5_4_io_o_0_co),
    .io_i_1_ci(cb_5_4_io_o_1_co),
    .io_i_2_ci(cb_5_4_io_o_2_co),
    .io_i_3_ci(cb_5_4_io_o_3_co),
    .io_i_4_ci(cb_5_4_io_o_4_co),
    .io_i_5_ci(cb_5_4_io_o_5_co),
    .io_i_6_ci(cb_5_4_io_o_6_co),
    .io_i_7_ci(cb_5_4_io_o_7_co),
    .io_o_0_co(cb_5_5_io_o_0_co),
    .io_o_1_co(cb_5_5_io_o_1_co),
    .io_o_2_co(cb_5_5_io_o_2_co),
    .io_o_3_co(cb_5_5_io_o_3_co),
    .io_o_4_co(cb_5_5_io_o_4_co),
    .io_o_5_co(cb_5_5_io_o_5_co),
    .io_o_6_co(cb_5_5_io_o_6_co),
    .io_o_7_co(cb_5_5_io_o_7_co),
    .io_vci(cb_5_4_io_vco),
    .io_vco(cb_5_5_io_vco),
    .io_vi(cb_5_5_io_vi),
    .io_we_i(cb_5_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_5_0_io_adr_i[1] ,
    \cb_5_0_io_adr_i[0] }),
    .io_dat_i({\cb_5_0_io_dat_i[15] ,
    \cb_5_0_io_dat_i[14] ,
    \cb_5_0_io_dat_i[13] ,
    \cb_5_0_io_dat_i[12] ,
    \cb_5_0_io_dat_i[11] ,
    \cb_5_0_io_dat_i[10] ,
    \cb_5_0_io_dat_i[9] ,
    \cb_5_0_io_dat_i[8] ,
    \cb_5_0_io_dat_i[7] ,
    \cb_5_0_io_dat_i[6] ,
    \cb_5_0_io_dat_i[5] ,
    \cb_5_0_io_dat_i[4] ,
    \cb_5_0_io_dat_i[3] ,
    \cb_5_0_io_dat_i[2] ,
    \cb_5_0_io_dat_i[1] ,
    \cb_5_0_io_dat_i[0] }),
    .io_dat_o({\cb_5_5_io_dat_o[15] ,
    \cb_5_5_io_dat_o[14] ,
    \cb_5_5_io_dat_o[13] ,
    \cb_5_5_io_dat_o[12] ,
    \cb_5_5_io_dat_o[11] ,
    \cb_5_5_io_dat_o[10] ,
    \cb_5_5_io_dat_o[9] ,
    \cb_5_5_io_dat_o[8] ,
    \cb_5_5_io_dat_o[7] ,
    \cb_5_5_io_dat_o[6] ,
    \cb_5_5_io_dat_o[5] ,
    \cb_5_5_io_dat_o[4] ,
    \cb_5_5_io_dat_o[3] ,
    \cb_5_5_io_dat_o[2] ,
    \cb_5_5_io_dat_o[1] ,
    \cb_5_5_io_dat_o[0] }),
    .io_eo({\cb_5_5_io_eo[63] ,
    \cb_5_5_io_eo[62] ,
    \cb_5_5_io_eo[61] ,
    \cb_5_5_io_eo[60] ,
    \cb_5_5_io_eo[59] ,
    \cb_5_5_io_eo[58] ,
    \cb_5_5_io_eo[57] ,
    \cb_5_5_io_eo[56] ,
    \cb_5_5_io_eo[55] ,
    \cb_5_5_io_eo[54] ,
    \cb_5_5_io_eo[53] ,
    \cb_5_5_io_eo[52] ,
    \cb_5_5_io_eo[51] ,
    \cb_5_5_io_eo[50] ,
    \cb_5_5_io_eo[49] ,
    \cb_5_5_io_eo[48] ,
    \cb_5_5_io_eo[47] ,
    \cb_5_5_io_eo[46] ,
    \cb_5_5_io_eo[45] ,
    \cb_5_5_io_eo[44] ,
    \cb_5_5_io_eo[43] ,
    \cb_5_5_io_eo[42] ,
    \cb_5_5_io_eo[41] ,
    \cb_5_5_io_eo[40] ,
    \cb_5_5_io_eo[39] ,
    \cb_5_5_io_eo[38] ,
    \cb_5_5_io_eo[37] ,
    \cb_5_5_io_eo[36] ,
    \cb_5_5_io_eo[35] ,
    \cb_5_5_io_eo[34] ,
    \cb_5_5_io_eo[33] ,
    \cb_5_5_io_eo[32] ,
    \cb_5_5_io_eo[31] ,
    \cb_5_5_io_eo[30] ,
    \cb_5_5_io_eo[29] ,
    \cb_5_5_io_eo[28] ,
    \cb_5_5_io_eo[27] ,
    \cb_5_5_io_eo[26] ,
    \cb_5_5_io_eo[25] ,
    \cb_5_5_io_eo[24] ,
    \cb_5_5_io_eo[23] ,
    \cb_5_5_io_eo[22] ,
    \cb_5_5_io_eo[21] ,
    \cb_5_5_io_eo[20] ,
    \cb_5_5_io_eo[19] ,
    \cb_5_5_io_eo[18] ,
    \cb_5_5_io_eo[17] ,
    \cb_5_5_io_eo[16] ,
    \cb_5_5_io_eo[15] ,
    \cb_5_5_io_eo[14] ,
    \cb_5_5_io_eo[13] ,
    \cb_5_5_io_eo[12] ,
    \cb_5_5_io_eo[11] ,
    \cb_5_5_io_eo[10] ,
    \cb_5_5_io_eo[9] ,
    \cb_5_5_io_eo[8] ,
    \cb_5_5_io_eo[7] ,
    \cb_5_5_io_eo[6] ,
    \cb_5_5_io_eo[5] ,
    \cb_5_5_io_eo[4] ,
    \cb_5_5_io_eo[3] ,
    \cb_5_5_io_eo[2] ,
    \cb_5_5_io_eo[1] ,
    \cb_5_5_io_eo[0] }),
    .io_i_0_in1({\cb_5_4_io_o_0_out[7] ,
    \cb_5_4_io_o_0_out[6] ,
    \cb_5_4_io_o_0_out[5] ,
    \cb_5_4_io_o_0_out[4] ,
    \cb_5_4_io_o_0_out[3] ,
    \cb_5_4_io_o_0_out[2] ,
    \cb_5_4_io_o_0_out[1] ,
    \cb_5_4_io_o_0_out[0] }),
    .io_i_1_in1({\cb_5_4_io_o_1_out[7] ,
    \cb_5_4_io_o_1_out[6] ,
    \cb_5_4_io_o_1_out[5] ,
    \cb_5_4_io_o_1_out[4] ,
    \cb_5_4_io_o_1_out[3] ,
    \cb_5_4_io_o_1_out[2] ,
    \cb_5_4_io_o_1_out[1] ,
    \cb_5_4_io_o_1_out[0] }),
    .io_i_2_in1({\cb_5_4_io_o_2_out[7] ,
    \cb_5_4_io_o_2_out[6] ,
    \cb_5_4_io_o_2_out[5] ,
    \cb_5_4_io_o_2_out[4] ,
    \cb_5_4_io_o_2_out[3] ,
    \cb_5_4_io_o_2_out[2] ,
    \cb_5_4_io_o_2_out[1] ,
    \cb_5_4_io_o_2_out[0] }),
    .io_i_3_in1({\cb_5_4_io_o_3_out[7] ,
    \cb_5_4_io_o_3_out[6] ,
    \cb_5_4_io_o_3_out[5] ,
    \cb_5_4_io_o_3_out[4] ,
    \cb_5_4_io_o_3_out[3] ,
    \cb_5_4_io_o_3_out[2] ,
    \cb_5_4_io_o_3_out[1] ,
    \cb_5_4_io_o_3_out[0] }),
    .io_i_4_in1({\cb_5_4_io_o_4_out[7] ,
    \cb_5_4_io_o_4_out[6] ,
    \cb_5_4_io_o_4_out[5] ,
    \cb_5_4_io_o_4_out[4] ,
    \cb_5_4_io_o_4_out[3] ,
    \cb_5_4_io_o_4_out[2] ,
    \cb_5_4_io_o_4_out[1] ,
    \cb_5_4_io_o_4_out[0] }),
    .io_i_5_in1({\cb_5_4_io_o_5_out[7] ,
    \cb_5_4_io_o_5_out[6] ,
    \cb_5_4_io_o_5_out[5] ,
    \cb_5_4_io_o_5_out[4] ,
    \cb_5_4_io_o_5_out[3] ,
    \cb_5_4_io_o_5_out[2] ,
    \cb_5_4_io_o_5_out[1] ,
    \cb_5_4_io_o_5_out[0] }),
    .io_i_6_in1({\cb_5_4_io_o_6_out[7] ,
    \cb_5_4_io_o_6_out[6] ,
    \cb_5_4_io_o_6_out[5] ,
    \cb_5_4_io_o_6_out[4] ,
    \cb_5_4_io_o_6_out[3] ,
    \cb_5_4_io_o_6_out[2] ,
    \cb_5_4_io_o_6_out[1] ,
    \cb_5_4_io_o_6_out[0] }),
    .io_i_7_in1({\cb_5_4_io_o_7_out[7] ,
    \cb_5_4_io_o_7_out[6] ,
    \cb_5_4_io_o_7_out[5] ,
    \cb_5_4_io_o_7_out[4] ,
    \cb_5_4_io_o_7_out[3] ,
    \cb_5_4_io_o_7_out[2] ,
    \cb_5_4_io_o_7_out[1] ,
    \cb_5_4_io_o_7_out[0] }),
    .io_o_0_out({\cb_5_5_io_o_0_out[7] ,
    \cb_5_5_io_o_0_out[6] ,
    \cb_5_5_io_o_0_out[5] ,
    \cb_5_5_io_o_0_out[4] ,
    \cb_5_5_io_o_0_out[3] ,
    \cb_5_5_io_o_0_out[2] ,
    \cb_5_5_io_o_0_out[1] ,
    \cb_5_5_io_o_0_out[0] }),
    .io_o_1_out({\cb_5_5_io_o_1_out[7] ,
    \cb_5_5_io_o_1_out[6] ,
    \cb_5_5_io_o_1_out[5] ,
    \cb_5_5_io_o_1_out[4] ,
    \cb_5_5_io_o_1_out[3] ,
    \cb_5_5_io_o_1_out[2] ,
    \cb_5_5_io_o_1_out[1] ,
    \cb_5_5_io_o_1_out[0] }),
    .io_o_2_out({\cb_5_5_io_o_2_out[7] ,
    \cb_5_5_io_o_2_out[6] ,
    \cb_5_5_io_o_2_out[5] ,
    \cb_5_5_io_o_2_out[4] ,
    \cb_5_5_io_o_2_out[3] ,
    \cb_5_5_io_o_2_out[2] ,
    \cb_5_5_io_o_2_out[1] ,
    \cb_5_5_io_o_2_out[0] }),
    .io_o_3_out({\cb_5_5_io_o_3_out[7] ,
    \cb_5_5_io_o_3_out[6] ,
    \cb_5_5_io_o_3_out[5] ,
    \cb_5_5_io_o_3_out[4] ,
    \cb_5_5_io_o_3_out[3] ,
    \cb_5_5_io_o_3_out[2] ,
    \cb_5_5_io_o_3_out[1] ,
    \cb_5_5_io_o_3_out[0] }),
    .io_o_4_out({\cb_5_5_io_o_4_out[7] ,
    \cb_5_5_io_o_4_out[6] ,
    \cb_5_5_io_o_4_out[5] ,
    \cb_5_5_io_o_4_out[4] ,
    \cb_5_5_io_o_4_out[3] ,
    \cb_5_5_io_o_4_out[2] ,
    \cb_5_5_io_o_4_out[1] ,
    \cb_5_5_io_o_4_out[0] }),
    .io_o_5_out({\cb_5_5_io_o_5_out[7] ,
    \cb_5_5_io_o_5_out[6] ,
    \cb_5_5_io_o_5_out[5] ,
    \cb_5_5_io_o_5_out[4] ,
    \cb_5_5_io_o_5_out[3] ,
    \cb_5_5_io_o_5_out[2] ,
    \cb_5_5_io_o_5_out[1] ,
    \cb_5_5_io_o_5_out[0] }),
    .io_o_6_out({\cb_5_5_io_o_6_out[7] ,
    \cb_5_5_io_o_6_out[6] ,
    \cb_5_5_io_o_6_out[5] ,
    \cb_5_5_io_o_6_out[4] ,
    \cb_5_5_io_o_6_out[3] ,
    \cb_5_5_io_o_6_out[2] ,
    \cb_5_5_io_o_6_out[1] ,
    \cb_5_5_io_o_6_out[0] }),
    .io_o_7_out({\cb_5_5_io_o_7_out[7] ,
    \cb_5_5_io_o_7_out[6] ,
    \cb_5_5_io_o_7_out[5] ,
    \cb_5_5_io_o_7_out[4] ,
    \cb_5_5_io_o_7_out[3] ,
    \cb_5_5_io_o_7_out[2] ,
    \cb_5_5_io_o_7_out[1] ,
    \cb_5_5_io_o_7_out[0] }),
    .io_wo({\cb_5_4_io_eo[63] ,
    \cb_5_4_io_eo[62] ,
    \cb_5_4_io_eo[61] ,
    \cb_5_4_io_eo[60] ,
    \cb_5_4_io_eo[59] ,
    \cb_5_4_io_eo[58] ,
    \cb_5_4_io_eo[57] ,
    \cb_5_4_io_eo[56] ,
    \cb_5_4_io_eo[55] ,
    \cb_5_4_io_eo[54] ,
    \cb_5_4_io_eo[53] ,
    \cb_5_4_io_eo[52] ,
    \cb_5_4_io_eo[51] ,
    \cb_5_4_io_eo[50] ,
    \cb_5_4_io_eo[49] ,
    \cb_5_4_io_eo[48] ,
    \cb_5_4_io_eo[47] ,
    \cb_5_4_io_eo[46] ,
    \cb_5_4_io_eo[45] ,
    \cb_5_4_io_eo[44] ,
    \cb_5_4_io_eo[43] ,
    \cb_5_4_io_eo[42] ,
    \cb_5_4_io_eo[41] ,
    \cb_5_4_io_eo[40] ,
    \cb_5_4_io_eo[39] ,
    \cb_5_4_io_eo[38] ,
    \cb_5_4_io_eo[37] ,
    \cb_5_4_io_eo[36] ,
    \cb_5_4_io_eo[35] ,
    \cb_5_4_io_eo[34] ,
    \cb_5_4_io_eo[33] ,
    \cb_5_4_io_eo[32] ,
    \cb_5_4_io_eo[31] ,
    \cb_5_4_io_eo[30] ,
    \cb_5_4_io_eo[29] ,
    \cb_5_4_io_eo[28] ,
    \cb_5_4_io_eo[27] ,
    \cb_5_4_io_eo[26] ,
    \cb_5_4_io_eo[25] ,
    \cb_5_4_io_eo[24] ,
    \cb_5_4_io_eo[23] ,
    \cb_5_4_io_eo[22] ,
    \cb_5_4_io_eo[21] ,
    \cb_5_4_io_eo[20] ,
    \cb_5_4_io_eo[19] ,
    \cb_5_4_io_eo[18] ,
    \cb_5_4_io_eo[17] ,
    \cb_5_4_io_eo[16] ,
    \cb_5_4_io_eo[15] ,
    \cb_5_4_io_eo[14] ,
    \cb_5_4_io_eo[13] ,
    \cb_5_4_io_eo[12] ,
    \cb_5_4_io_eo[11] ,
    \cb_5_4_io_eo[10] ,
    \cb_5_4_io_eo[9] ,
    \cb_5_4_io_eo[8] ,
    \cb_5_4_io_eo[7] ,
    \cb_5_4_io_eo[6] ,
    \cb_5_4_io_eo[5] ,
    \cb_5_4_io_eo[4] ,
    \cb_5_4_io_eo[3] ,
    \cb_5_4_io_eo[2] ,
    \cb_5_4_io_eo[1] ,
    \cb_5_4_io_eo[0] }));
 cic_block cb_5_6 (.io_cs_i(cb_5_6_io_cs_i),
    .io_i_0_ci(cb_5_5_io_o_0_co),
    .io_i_1_ci(cb_5_5_io_o_1_co),
    .io_i_2_ci(cb_5_5_io_o_2_co),
    .io_i_3_ci(cb_5_5_io_o_3_co),
    .io_i_4_ci(cb_5_5_io_o_4_co),
    .io_i_5_ci(cb_5_5_io_o_5_co),
    .io_i_6_ci(cb_5_5_io_o_6_co),
    .io_i_7_ci(cb_5_5_io_o_7_co),
    .io_o_0_co(cb_5_6_io_o_0_co),
    .io_o_1_co(cb_5_6_io_o_1_co),
    .io_o_2_co(cb_5_6_io_o_2_co),
    .io_o_3_co(cb_5_6_io_o_3_co),
    .io_o_4_co(cb_5_6_io_o_4_co),
    .io_o_5_co(cb_5_6_io_o_5_co),
    .io_o_6_co(cb_5_6_io_o_6_co),
    .io_o_7_co(cb_5_6_io_o_7_co),
    .io_vci(cb_5_5_io_vco),
    .io_vco(cb_5_6_io_vco),
    .io_vi(cb_5_6_io_vi),
    .io_we_i(cb_5_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_5_0_io_adr_i[1] ,
    \cb_5_0_io_adr_i[0] }),
    .io_dat_i({\cb_5_0_io_dat_i[15] ,
    \cb_5_0_io_dat_i[14] ,
    \cb_5_0_io_dat_i[13] ,
    \cb_5_0_io_dat_i[12] ,
    \cb_5_0_io_dat_i[11] ,
    \cb_5_0_io_dat_i[10] ,
    \cb_5_0_io_dat_i[9] ,
    \cb_5_0_io_dat_i[8] ,
    \cb_5_0_io_dat_i[7] ,
    \cb_5_0_io_dat_i[6] ,
    \cb_5_0_io_dat_i[5] ,
    \cb_5_0_io_dat_i[4] ,
    \cb_5_0_io_dat_i[3] ,
    \cb_5_0_io_dat_i[2] ,
    \cb_5_0_io_dat_i[1] ,
    \cb_5_0_io_dat_i[0] }),
    .io_dat_o({\cb_5_6_io_dat_o[15] ,
    \cb_5_6_io_dat_o[14] ,
    \cb_5_6_io_dat_o[13] ,
    \cb_5_6_io_dat_o[12] ,
    \cb_5_6_io_dat_o[11] ,
    \cb_5_6_io_dat_o[10] ,
    \cb_5_6_io_dat_o[9] ,
    \cb_5_6_io_dat_o[8] ,
    \cb_5_6_io_dat_o[7] ,
    \cb_5_6_io_dat_o[6] ,
    \cb_5_6_io_dat_o[5] ,
    \cb_5_6_io_dat_o[4] ,
    \cb_5_6_io_dat_o[3] ,
    \cb_5_6_io_dat_o[2] ,
    \cb_5_6_io_dat_o[1] ,
    \cb_5_6_io_dat_o[0] }),
    .io_eo({\cb_5_6_io_eo[63] ,
    \cb_5_6_io_eo[62] ,
    \cb_5_6_io_eo[61] ,
    \cb_5_6_io_eo[60] ,
    \cb_5_6_io_eo[59] ,
    \cb_5_6_io_eo[58] ,
    \cb_5_6_io_eo[57] ,
    \cb_5_6_io_eo[56] ,
    \cb_5_6_io_eo[55] ,
    \cb_5_6_io_eo[54] ,
    \cb_5_6_io_eo[53] ,
    \cb_5_6_io_eo[52] ,
    \cb_5_6_io_eo[51] ,
    \cb_5_6_io_eo[50] ,
    \cb_5_6_io_eo[49] ,
    \cb_5_6_io_eo[48] ,
    \cb_5_6_io_eo[47] ,
    \cb_5_6_io_eo[46] ,
    \cb_5_6_io_eo[45] ,
    \cb_5_6_io_eo[44] ,
    \cb_5_6_io_eo[43] ,
    \cb_5_6_io_eo[42] ,
    \cb_5_6_io_eo[41] ,
    \cb_5_6_io_eo[40] ,
    \cb_5_6_io_eo[39] ,
    \cb_5_6_io_eo[38] ,
    \cb_5_6_io_eo[37] ,
    \cb_5_6_io_eo[36] ,
    \cb_5_6_io_eo[35] ,
    \cb_5_6_io_eo[34] ,
    \cb_5_6_io_eo[33] ,
    \cb_5_6_io_eo[32] ,
    \cb_5_6_io_eo[31] ,
    \cb_5_6_io_eo[30] ,
    \cb_5_6_io_eo[29] ,
    \cb_5_6_io_eo[28] ,
    \cb_5_6_io_eo[27] ,
    \cb_5_6_io_eo[26] ,
    \cb_5_6_io_eo[25] ,
    \cb_5_6_io_eo[24] ,
    \cb_5_6_io_eo[23] ,
    \cb_5_6_io_eo[22] ,
    \cb_5_6_io_eo[21] ,
    \cb_5_6_io_eo[20] ,
    \cb_5_6_io_eo[19] ,
    \cb_5_6_io_eo[18] ,
    \cb_5_6_io_eo[17] ,
    \cb_5_6_io_eo[16] ,
    \cb_5_6_io_eo[15] ,
    \cb_5_6_io_eo[14] ,
    \cb_5_6_io_eo[13] ,
    \cb_5_6_io_eo[12] ,
    \cb_5_6_io_eo[11] ,
    \cb_5_6_io_eo[10] ,
    \cb_5_6_io_eo[9] ,
    \cb_5_6_io_eo[8] ,
    \cb_5_6_io_eo[7] ,
    \cb_5_6_io_eo[6] ,
    \cb_5_6_io_eo[5] ,
    \cb_5_6_io_eo[4] ,
    \cb_5_6_io_eo[3] ,
    \cb_5_6_io_eo[2] ,
    \cb_5_6_io_eo[1] ,
    \cb_5_6_io_eo[0] }),
    .io_i_0_in1({\cb_5_5_io_o_0_out[7] ,
    \cb_5_5_io_o_0_out[6] ,
    \cb_5_5_io_o_0_out[5] ,
    \cb_5_5_io_o_0_out[4] ,
    \cb_5_5_io_o_0_out[3] ,
    \cb_5_5_io_o_0_out[2] ,
    \cb_5_5_io_o_0_out[1] ,
    \cb_5_5_io_o_0_out[0] }),
    .io_i_1_in1({\cb_5_5_io_o_1_out[7] ,
    \cb_5_5_io_o_1_out[6] ,
    \cb_5_5_io_o_1_out[5] ,
    \cb_5_5_io_o_1_out[4] ,
    \cb_5_5_io_o_1_out[3] ,
    \cb_5_5_io_o_1_out[2] ,
    \cb_5_5_io_o_1_out[1] ,
    \cb_5_5_io_o_1_out[0] }),
    .io_i_2_in1({\cb_5_5_io_o_2_out[7] ,
    \cb_5_5_io_o_2_out[6] ,
    \cb_5_5_io_o_2_out[5] ,
    \cb_5_5_io_o_2_out[4] ,
    \cb_5_5_io_o_2_out[3] ,
    \cb_5_5_io_o_2_out[2] ,
    \cb_5_5_io_o_2_out[1] ,
    \cb_5_5_io_o_2_out[0] }),
    .io_i_3_in1({\cb_5_5_io_o_3_out[7] ,
    \cb_5_5_io_o_3_out[6] ,
    \cb_5_5_io_o_3_out[5] ,
    \cb_5_5_io_o_3_out[4] ,
    \cb_5_5_io_o_3_out[3] ,
    \cb_5_5_io_o_3_out[2] ,
    \cb_5_5_io_o_3_out[1] ,
    \cb_5_5_io_o_3_out[0] }),
    .io_i_4_in1({\cb_5_5_io_o_4_out[7] ,
    \cb_5_5_io_o_4_out[6] ,
    \cb_5_5_io_o_4_out[5] ,
    \cb_5_5_io_o_4_out[4] ,
    \cb_5_5_io_o_4_out[3] ,
    \cb_5_5_io_o_4_out[2] ,
    \cb_5_5_io_o_4_out[1] ,
    \cb_5_5_io_o_4_out[0] }),
    .io_i_5_in1({\cb_5_5_io_o_5_out[7] ,
    \cb_5_5_io_o_5_out[6] ,
    \cb_5_5_io_o_5_out[5] ,
    \cb_5_5_io_o_5_out[4] ,
    \cb_5_5_io_o_5_out[3] ,
    \cb_5_5_io_o_5_out[2] ,
    \cb_5_5_io_o_5_out[1] ,
    \cb_5_5_io_o_5_out[0] }),
    .io_i_6_in1({\cb_5_5_io_o_6_out[7] ,
    \cb_5_5_io_o_6_out[6] ,
    \cb_5_5_io_o_6_out[5] ,
    \cb_5_5_io_o_6_out[4] ,
    \cb_5_5_io_o_6_out[3] ,
    \cb_5_5_io_o_6_out[2] ,
    \cb_5_5_io_o_6_out[1] ,
    \cb_5_5_io_o_6_out[0] }),
    .io_i_7_in1({\cb_5_5_io_o_7_out[7] ,
    \cb_5_5_io_o_7_out[6] ,
    \cb_5_5_io_o_7_out[5] ,
    \cb_5_5_io_o_7_out[4] ,
    \cb_5_5_io_o_7_out[3] ,
    \cb_5_5_io_o_7_out[2] ,
    \cb_5_5_io_o_7_out[1] ,
    \cb_5_5_io_o_7_out[0] }),
    .io_o_0_out({\cb_5_6_io_o_0_out[7] ,
    \cb_5_6_io_o_0_out[6] ,
    \cb_5_6_io_o_0_out[5] ,
    \cb_5_6_io_o_0_out[4] ,
    \cb_5_6_io_o_0_out[3] ,
    \cb_5_6_io_o_0_out[2] ,
    \cb_5_6_io_o_0_out[1] ,
    \cb_5_6_io_o_0_out[0] }),
    .io_o_1_out({\cb_5_6_io_o_1_out[7] ,
    \cb_5_6_io_o_1_out[6] ,
    \cb_5_6_io_o_1_out[5] ,
    \cb_5_6_io_o_1_out[4] ,
    \cb_5_6_io_o_1_out[3] ,
    \cb_5_6_io_o_1_out[2] ,
    \cb_5_6_io_o_1_out[1] ,
    \cb_5_6_io_o_1_out[0] }),
    .io_o_2_out({\cb_5_6_io_o_2_out[7] ,
    \cb_5_6_io_o_2_out[6] ,
    \cb_5_6_io_o_2_out[5] ,
    \cb_5_6_io_o_2_out[4] ,
    \cb_5_6_io_o_2_out[3] ,
    \cb_5_6_io_o_2_out[2] ,
    \cb_5_6_io_o_2_out[1] ,
    \cb_5_6_io_o_2_out[0] }),
    .io_o_3_out({\cb_5_6_io_o_3_out[7] ,
    \cb_5_6_io_o_3_out[6] ,
    \cb_5_6_io_o_3_out[5] ,
    \cb_5_6_io_o_3_out[4] ,
    \cb_5_6_io_o_3_out[3] ,
    \cb_5_6_io_o_3_out[2] ,
    \cb_5_6_io_o_3_out[1] ,
    \cb_5_6_io_o_3_out[0] }),
    .io_o_4_out({\cb_5_6_io_o_4_out[7] ,
    \cb_5_6_io_o_4_out[6] ,
    \cb_5_6_io_o_4_out[5] ,
    \cb_5_6_io_o_4_out[4] ,
    \cb_5_6_io_o_4_out[3] ,
    \cb_5_6_io_o_4_out[2] ,
    \cb_5_6_io_o_4_out[1] ,
    \cb_5_6_io_o_4_out[0] }),
    .io_o_5_out({\cb_5_6_io_o_5_out[7] ,
    \cb_5_6_io_o_5_out[6] ,
    \cb_5_6_io_o_5_out[5] ,
    \cb_5_6_io_o_5_out[4] ,
    \cb_5_6_io_o_5_out[3] ,
    \cb_5_6_io_o_5_out[2] ,
    \cb_5_6_io_o_5_out[1] ,
    \cb_5_6_io_o_5_out[0] }),
    .io_o_6_out({\cb_5_6_io_o_6_out[7] ,
    \cb_5_6_io_o_6_out[6] ,
    \cb_5_6_io_o_6_out[5] ,
    \cb_5_6_io_o_6_out[4] ,
    \cb_5_6_io_o_6_out[3] ,
    \cb_5_6_io_o_6_out[2] ,
    \cb_5_6_io_o_6_out[1] ,
    \cb_5_6_io_o_6_out[0] }),
    .io_o_7_out({\cb_5_6_io_o_7_out[7] ,
    \cb_5_6_io_o_7_out[6] ,
    \cb_5_6_io_o_7_out[5] ,
    \cb_5_6_io_o_7_out[4] ,
    \cb_5_6_io_o_7_out[3] ,
    \cb_5_6_io_o_7_out[2] ,
    \cb_5_6_io_o_7_out[1] ,
    \cb_5_6_io_o_7_out[0] }),
    .io_wo({\cb_5_5_io_eo[63] ,
    \cb_5_5_io_eo[62] ,
    \cb_5_5_io_eo[61] ,
    \cb_5_5_io_eo[60] ,
    \cb_5_5_io_eo[59] ,
    \cb_5_5_io_eo[58] ,
    \cb_5_5_io_eo[57] ,
    \cb_5_5_io_eo[56] ,
    \cb_5_5_io_eo[55] ,
    \cb_5_5_io_eo[54] ,
    \cb_5_5_io_eo[53] ,
    \cb_5_5_io_eo[52] ,
    \cb_5_5_io_eo[51] ,
    \cb_5_5_io_eo[50] ,
    \cb_5_5_io_eo[49] ,
    \cb_5_5_io_eo[48] ,
    \cb_5_5_io_eo[47] ,
    \cb_5_5_io_eo[46] ,
    \cb_5_5_io_eo[45] ,
    \cb_5_5_io_eo[44] ,
    \cb_5_5_io_eo[43] ,
    \cb_5_5_io_eo[42] ,
    \cb_5_5_io_eo[41] ,
    \cb_5_5_io_eo[40] ,
    \cb_5_5_io_eo[39] ,
    \cb_5_5_io_eo[38] ,
    \cb_5_5_io_eo[37] ,
    \cb_5_5_io_eo[36] ,
    \cb_5_5_io_eo[35] ,
    \cb_5_5_io_eo[34] ,
    \cb_5_5_io_eo[33] ,
    \cb_5_5_io_eo[32] ,
    \cb_5_5_io_eo[31] ,
    \cb_5_5_io_eo[30] ,
    \cb_5_5_io_eo[29] ,
    \cb_5_5_io_eo[28] ,
    \cb_5_5_io_eo[27] ,
    \cb_5_5_io_eo[26] ,
    \cb_5_5_io_eo[25] ,
    \cb_5_5_io_eo[24] ,
    \cb_5_5_io_eo[23] ,
    \cb_5_5_io_eo[22] ,
    \cb_5_5_io_eo[21] ,
    \cb_5_5_io_eo[20] ,
    \cb_5_5_io_eo[19] ,
    \cb_5_5_io_eo[18] ,
    \cb_5_5_io_eo[17] ,
    \cb_5_5_io_eo[16] ,
    \cb_5_5_io_eo[15] ,
    \cb_5_5_io_eo[14] ,
    \cb_5_5_io_eo[13] ,
    \cb_5_5_io_eo[12] ,
    \cb_5_5_io_eo[11] ,
    \cb_5_5_io_eo[10] ,
    \cb_5_5_io_eo[9] ,
    \cb_5_5_io_eo[8] ,
    \cb_5_5_io_eo[7] ,
    \cb_5_5_io_eo[6] ,
    \cb_5_5_io_eo[5] ,
    \cb_5_5_io_eo[4] ,
    \cb_5_5_io_eo[3] ,
    \cb_5_5_io_eo[2] ,
    \cb_5_5_io_eo[1] ,
    \cb_5_5_io_eo[0] }));
 cic_block cb_5_7 (.io_cs_i(cb_5_7_io_cs_i),
    .io_i_0_ci(cb_5_6_io_o_0_co),
    .io_i_1_ci(cb_5_6_io_o_1_co),
    .io_i_2_ci(cb_5_6_io_o_2_co),
    .io_i_3_ci(cb_5_6_io_o_3_co),
    .io_i_4_ci(cb_5_6_io_o_4_co),
    .io_i_5_ci(cb_5_6_io_o_5_co),
    .io_i_6_ci(cb_5_6_io_o_6_co),
    .io_i_7_ci(cb_5_6_io_o_7_co),
    .io_o_0_co(cb_5_7_io_o_0_co),
    .io_o_1_co(cb_5_7_io_o_1_co),
    .io_o_2_co(cb_5_7_io_o_2_co),
    .io_o_3_co(cb_5_7_io_o_3_co),
    .io_o_4_co(cb_5_7_io_o_4_co),
    .io_o_5_co(cb_5_7_io_o_5_co),
    .io_o_6_co(cb_5_7_io_o_6_co),
    .io_o_7_co(cb_5_7_io_o_7_co),
    .io_vci(cb_5_6_io_vco),
    .io_vco(cb_5_7_io_vco),
    .io_vi(cb_5_7_io_vi),
    .io_we_i(cb_5_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_5_0_io_adr_i[1] ,
    \cb_5_0_io_adr_i[0] }),
    .io_dat_i({\cb_5_0_io_dat_i[15] ,
    \cb_5_0_io_dat_i[14] ,
    \cb_5_0_io_dat_i[13] ,
    \cb_5_0_io_dat_i[12] ,
    \cb_5_0_io_dat_i[11] ,
    \cb_5_0_io_dat_i[10] ,
    \cb_5_0_io_dat_i[9] ,
    \cb_5_0_io_dat_i[8] ,
    \cb_5_0_io_dat_i[7] ,
    \cb_5_0_io_dat_i[6] ,
    \cb_5_0_io_dat_i[5] ,
    \cb_5_0_io_dat_i[4] ,
    \cb_5_0_io_dat_i[3] ,
    \cb_5_0_io_dat_i[2] ,
    \cb_5_0_io_dat_i[1] ,
    \cb_5_0_io_dat_i[0] }),
    .io_dat_o({\cb_5_7_io_dat_o[15] ,
    \cb_5_7_io_dat_o[14] ,
    \cb_5_7_io_dat_o[13] ,
    \cb_5_7_io_dat_o[12] ,
    \cb_5_7_io_dat_o[11] ,
    \cb_5_7_io_dat_o[10] ,
    \cb_5_7_io_dat_o[9] ,
    \cb_5_7_io_dat_o[8] ,
    \cb_5_7_io_dat_o[7] ,
    \cb_5_7_io_dat_o[6] ,
    \cb_5_7_io_dat_o[5] ,
    \cb_5_7_io_dat_o[4] ,
    \cb_5_7_io_dat_o[3] ,
    \cb_5_7_io_dat_o[2] ,
    \cb_5_7_io_dat_o[1] ,
    \cb_5_7_io_dat_o[0] }),
    .io_eo({\cb_5_7_io_eo[63] ,
    \cb_5_7_io_eo[62] ,
    \cb_5_7_io_eo[61] ,
    \cb_5_7_io_eo[60] ,
    \cb_5_7_io_eo[59] ,
    \cb_5_7_io_eo[58] ,
    \cb_5_7_io_eo[57] ,
    \cb_5_7_io_eo[56] ,
    \cb_5_7_io_eo[55] ,
    \cb_5_7_io_eo[54] ,
    \cb_5_7_io_eo[53] ,
    \cb_5_7_io_eo[52] ,
    \cb_5_7_io_eo[51] ,
    \cb_5_7_io_eo[50] ,
    \cb_5_7_io_eo[49] ,
    \cb_5_7_io_eo[48] ,
    \cb_5_7_io_eo[47] ,
    \cb_5_7_io_eo[46] ,
    \cb_5_7_io_eo[45] ,
    \cb_5_7_io_eo[44] ,
    \cb_5_7_io_eo[43] ,
    \cb_5_7_io_eo[42] ,
    \cb_5_7_io_eo[41] ,
    \cb_5_7_io_eo[40] ,
    \cb_5_7_io_eo[39] ,
    \cb_5_7_io_eo[38] ,
    \cb_5_7_io_eo[37] ,
    \cb_5_7_io_eo[36] ,
    \cb_5_7_io_eo[35] ,
    \cb_5_7_io_eo[34] ,
    \cb_5_7_io_eo[33] ,
    \cb_5_7_io_eo[32] ,
    \cb_5_7_io_eo[31] ,
    \cb_5_7_io_eo[30] ,
    \cb_5_7_io_eo[29] ,
    \cb_5_7_io_eo[28] ,
    \cb_5_7_io_eo[27] ,
    \cb_5_7_io_eo[26] ,
    \cb_5_7_io_eo[25] ,
    \cb_5_7_io_eo[24] ,
    \cb_5_7_io_eo[23] ,
    \cb_5_7_io_eo[22] ,
    \cb_5_7_io_eo[21] ,
    \cb_5_7_io_eo[20] ,
    \cb_5_7_io_eo[19] ,
    \cb_5_7_io_eo[18] ,
    \cb_5_7_io_eo[17] ,
    \cb_5_7_io_eo[16] ,
    \cb_5_7_io_eo[15] ,
    \cb_5_7_io_eo[14] ,
    \cb_5_7_io_eo[13] ,
    \cb_5_7_io_eo[12] ,
    \cb_5_7_io_eo[11] ,
    \cb_5_7_io_eo[10] ,
    \cb_5_7_io_eo[9] ,
    \cb_5_7_io_eo[8] ,
    \cb_5_7_io_eo[7] ,
    \cb_5_7_io_eo[6] ,
    \cb_5_7_io_eo[5] ,
    \cb_5_7_io_eo[4] ,
    \cb_5_7_io_eo[3] ,
    \cb_5_7_io_eo[2] ,
    \cb_5_7_io_eo[1] ,
    \cb_5_7_io_eo[0] }),
    .io_i_0_in1({\cb_5_6_io_o_0_out[7] ,
    \cb_5_6_io_o_0_out[6] ,
    \cb_5_6_io_o_0_out[5] ,
    \cb_5_6_io_o_0_out[4] ,
    \cb_5_6_io_o_0_out[3] ,
    \cb_5_6_io_o_0_out[2] ,
    \cb_5_6_io_o_0_out[1] ,
    \cb_5_6_io_o_0_out[0] }),
    .io_i_1_in1({\cb_5_6_io_o_1_out[7] ,
    \cb_5_6_io_o_1_out[6] ,
    \cb_5_6_io_o_1_out[5] ,
    \cb_5_6_io_o_1_out[4] ,
    \cb_5_6_io_o_1_out[3] ,
    \cb_5_6_io_o_1_out[2] ,
    \cb_5_6_io_o_1_out[1] ,
    \cb_5_6_io_o_1_out[0] }),
    .io_i_2_in1({\cb_5_6_io_o_2_out[7] ,
    \cb_5_6_io_o_2_out[6] ,
    \cb_5_6_io_o_2_out[5] ,
    \cb_5_6_io_o_2_out[4] ,
    \cb_5_6_io_o_2_out[3] ,
    \cb_5_6_io_o_2_out[2] ,
    \cb_5_6_io_o_2_out[1] ,
    \cb_5_6_io_o_2_out[0] }),
    .io_i_3_in1({\cb_5_6_io_o_3_out[7] ,
    \cb_5_6_io_o_3_out[6] ,
    \cb_5_6_io_o_3_out[5] ,
    \cb_5_6_io_o_3_out[4] ,
    \cb_5_6_io_o_3_out[3] ,
    \cb_5_6_io_o_3_out[2] ,
    \cb_5_6_io_o_3_out[1] ,
    \cb_5_6_io_o_3_out[0] }),
    .io_i_4_in1({\cb_5_6_io_o_4_out[7] ,
    \cb_5_6_io_o_4_out[6] ,
    \cb_5_6_io_o_4_out[5] ,
    \cb_5_6_io_o_4_out[4] ,
    \cb_5_6_io_o_4_out[3] ,
    \cb_5_6_io_o_4_out[2] ,
    \cb_5_6_io_o_4_out[1] ,
    \cb_5_6_io_o_4_out[0] }),
    .io_i_5_in1({\cb_5_6_io_o_5_out[7] ,
    \cb_5_6_io_o_5_out[6] ,
    \cb_5_6_io_o_5_out[5] ,
    \cb_5_6_io_o_5_out[4] ,
    \cb_5_6_io_o_5_out[3] ,
    \cb_5_6_io_o_5_out[2] ,
    \cb_5_6_io_o_5_out[1] ,
    \cb_5_6_io_o_5_out[0] }),
    .io_i_6_in1({\cb_5_6_io_o_6_out[7] ,
    \cb_5_6_io_o_6_out[6] ,
    \cb_5_6_io_o_6_out[5] ,
    \cb_5_6_io_o_6_out[4] ,
    \cb_5_6_io_o_6_out[3] ,
    \cb_5_6_io_o_6_out[2] ,
    \cb_5_6_io_o_6_out[1] ,
    \cb_5_6_io_o_6_out[0] }),
    .io_i_7_in1({\cb_5_6_io_o_7_out[7] ,
    \cb_5_6_io_o_7_out[6] ,
    \cb_5_6_io_o_7_out[5] ,
    \cb_5_6_io_o_7_out[4] ,
    \cb_5_6_io_o_7_out[3] ,
    \cb_5_6_io_o_7_out[2] ,
    \cb_5_6_io_o_7_out[1] ,
    \cb_5_6_io_o_7_out[0] }),
    .io_o_0_out({\cb_5_7_io_o_0_out[7] ,
    \cb_5_7_io_o_0_out[6] ,
    \cb_5_7_io_o_0_out[5] ,
    \cb_5_7_io_o_0_out[4] ,
    \cb_5_7_io_o_0_out[3] ,
    \cb_5_7_io_o_0_out[2] ,
    \cb_5_7_io_o_0_out[1] ,
    \cb_5_7_io_o_0_out[0] }),
    .io_o_1_out({\cb_5_7_io_o_1_out[7] ,
    \cb_5_7_io_o_1_out[6] ,
    \cb_5_7_io_o_1_out[5] ,
    \cb_5_7_io_o_1_out[4] ,
    \cb_5_7_io_o_1_out[3] ,
    \cb_5_7_io_o_1_out[2] ,
    \cb_5_7_io_o_1_out[1] ,
    \cb_5_7_io_o_1_out[0] }),
    .io_o_2_out({\cb_5_7_io_o_2_out[7] ,
    \cb_5_7_io_o_2_out[6] ,
    \cb_5_7_io_o_2_out[5] ,
    \cb_5_7_io_o_2_out[4] ,
    \cb_5_7_io_o_2_out[3] ,
    \cb_5_7_io_o_2_out[2] ,
    \cb_5_7_io_o_2_out[1] ,
    \cb_5_7_io_o_2_out[0] }),
    .io_o_3_out({\cb_5_7_io_o_3_out[7] ,
    \cb_5_7_io_o_3_out[6] ,
    \cb_5_7_io_o_3_out[5] ,
    \cb_5_7_io_o_3_out[4] ,
    \cb_5_7_io_o_3_out[3] ,
    \cb_5_7_io_o_3_out[2] ,
    \cb_5_7_io_o_3_out[1] ,
    \cb_5_7_io_o_3_out[0] }),
    .io_o_4_out({\cb_5_7_io_o_4_out[7] ,
    \cb_5_7_io_o_4_out[6] ,
    \cb_5_7_io_o_4_out[5] ,
    \cb_5_7_io_o_4_out[4] ,
    \cb_5_7_io_o_4_out[3] ,
    \cb_5_7_io_o_4_out[2] ,
    \cb_5_7_io_o_4_out[1] ,
    \cb_5_7_io_o_4_out[0] }),
    .io_o_5_out({\cb_5_7_io_o_5_out[7] ,
    \cb_5_7_io_o_5_out[6] ,
    \cb_5_7_io_o_5_out[5] ,
    \cb_5_7_io_o_5_out[4] ,
    \cb_5_7_io_o_5_out[3] ,
    \cb_5_7_io_o_5_out[2] ,
    \cb_5_7_io_o_5_out[1] ,
    \cb_5_7_io_o_5_out[0] }),
    .io_o_6_out({\cb_5_7_io_o_6_out[7] ,
    \cb_5_7_io_o_6_out[6] ,
    \cb_5_7_io_o_6_out[5] ,
    \cb_5_7_io_o_6_out[4] ,
    \cb_5_7_io_o_6_out[3] ,
    \cb_5_7_io_o_6_out[2] ,
    \cb_5_7_io_o_6_out[1] ,
    \cb_5_7_io_o_6_out[0] }),
    .io_o_7_out({\cb_5_7_io_o_7_out[7] ,
    \cb_5_7_io_o_7_out[6] ,
    \cb_5_7_io_o_7_out[5] ,
    \cb_5_7_io_o_7_out[4] ,
    \cb_5_7_io_o_7_out[3] ,
    \cb_5_7_io_o_7_out[2] ,
    \cb_5_7_io_o_7_out[1] ,
    \cb_5_7_io_o_7_out[0] }),
    .io_wo({\cb_5_6_io_eo[63] ,
    \cb_5_6_io_eo[62] ,
    \cb_5_6_io_eo[61] ,
    \cb_5_6_io_eo[60] ,
    \cb_5_6_io_eo[59] ,
    \cb_5_6_io_eo[58] ,
    \cb_5_6_io_eo[57] ,
    \cb_5_6_io_eo[56] ,
    \cb_5_6_io_eo[55] ,
    \cb_5_6_io_eo[54] ,
    \cb_5_6_io_eo[53] ,
    \cb_5_6_io_eo[52] ,
    \cb_5_6_io_eo[51] ,
    \cb_5_6_io_eo[50] ,
    \cb_5_6_io_eo[49] ,
    \cb_5_6_io_eo[48] ,
    \cb_5_6_io_eo[47] ,
    \cb_5_6_io_eo[46] ,
    \cb_5_6_io_eo[45] ,
    \cb_5_6_io_eo[44] ,
    \cb_5_6_io_eo[43] ,
    \cb_5_6_io_eo[42] ,
    \cb_5_6_io_eo[41] ,
    \cb_5_6_io_eo[40] ,
    \cb_5_6_io_eo[39] ,
    \cb_5_6_io_eo[38] ,
    \cb_5_6_io_eo[37] ,
    \cb_5_6_io_eo[36] ,
    \cb_5_6_io_eo[35] ,
    \cb_5_6_io_eo[34] ,
    \cb_5_6_io_eo[33] ,
    \cb_5_6_io_eo[32] ,
    \cb_5_6_io_eo[31] ,
    \cb_5_6_io_eo[30] ,
    \cb_5_6_io_eo[29] ,
    \cb_5_6_io_eo[28] ,
    \cb_5_6_io_eo[27] ,
    \cb_5_6_io_eo[26] ,
    \cb_5_6_io_eo[25] ,
    \cb_5_6_io_eo[24] ,
    \cb_5_6_io_eo[23] ,
    \cb_5_6_io_eo[22] ,
    \cb_5_6_io_eo[21] ,
    \cb_5_6_io_eo[20] ,
    \cb_5_6_io_eo[19] ,
    \cb_5_6_io_eo[18] ,
    \cb_5_6_io_eo[17] ,
    \cb_5_6_io_eo[16] ,
    \cb_5_6_io_eo[15] ,
    \cb_5_6_io_eo[14] ,
    \cb_5_6_io_eo[13] ,
    \cb_5_6_io_eo[12] ,
    \cb_5_6_io_eo[11] ,
    \cb_5_6_io_eo[10] ,
    \cb_5_6_io_eo[9] ,
    \cb_5_6_io_eo[8] ,
    \cb_5_6_io_eo[7] ,
    \cb_5_6_io_eo[6] ,
    \cb_5_6_io_eo[5] ,
    \cb_5_6_io_eo[4] ,
    \cb_5_6_io_eo[3] ,
    \cb_5_6_io_eo[2] ,
    \cb_5_6_io_eo[1] ,
    \cb_5_6_io_eo[0] }));
 cic_block cb_5_8 (.io_cs_i(cb_5_8_io_cs_i),
    .io_i_0_ci(cb_5_7_io_o_0_co),
    .io_i_1_ci(cb_5_7_io_o_1_co),
    .io_i_2_ci(cb_5_7_io_o_2_co),
    .io_i_3_ci(cb_5_7_io_o_3_co),
    .io_i_4_ci(cb_5_7_io_o_4_co),
    .io_i_5_ci(cb_5_7_io_o_5_co),
    .io_i_6_ci(cb_5_7_io_o_6_co),
    .io_i_7_ci(cb_5_7_io_o_7_co),
    .io_o_0_co(cb_5_8_io_o_0_co),
    .io_o_1_co(cb_5_8_io_o_1_co),
    .io_o_2_co(cb_5_8_io_o_2_co),
    .io_o_3_co(cb_5_8_io_o_3_co),
    .io_o_4_co(cb_5_8_io_o_4_co),
    .io_o_5_co(cb_5_8_io_o_5_co),
    .io_o_6_co(cb_5_8_io_o_6_co),
    .io_o_7_co(cb_5_8_io_o_7_co),
    .io_vci(cb_5_7_io_vco),
    .io_vco(cb_5_8_io_vco),
    .io_vi(cb_5_8_io_vi),
    .io_we_i(cb_5_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_5_0_io_adr_i[1] ,
    \cb_5_0_io_adr_i[0] }),
    .io_dat_i({\cb_5_0_io_dat_i[15] ,
    \cb_5_0_io_dat_i[14] ,
    \cb_5_0_io_dat_i[13] ,
    \cb_5_0_io_dat_i[12] ,
    \cb_5_0_io_dat_i[11] ,
    \cb_5_0_io_dat_i[10] ,
    \cb_5_0_io_dat_i[9] ,
    \cb_5_0_io_dat_i[8] ,
    \cb_5_0_io_dat_i[7] ,
    \cb_5_0_io_dat_i[6] ,
    \cb_5_0_io_dat_i[5] ,
    \cb_5_0_io_dat_i[4] ,
    \cb_5_0_io_dat_i[3] ,
    \cb_5_0_io_dat_i[2] ,
    \cb_5_0_io_dat_i[1] ,
    \cb_5_0_io_dat_i[0] }),
    .io_dat_o({\cb_5_8_io_dat_o[15] ,
    \cb_5_8_io_dat_o[14] ,
    \cb_5_8_io_dat_o[13] ,
    \cb_5_8_io_dat_o[12] ,
    \cb_5_8_io_dat_o[11] ,
    \cb_5_8_io_dat_o[10] ,
    \cb_5_8_io_dat_o[9] ,
    \cb_5_8_io_dat_o[8] ,
    \cb_5_8_io_dat_o[7] ,
    \cb_5_8_io_dat_o[6] ,
    \cb_5_8_io_dat_o[5] ,
    \cb_5_8_io_dat_o[4] ,
    \cb_5_8_io_dat_o[3] ,
    \cb_5_8_io_dat_o[2] ,
    \cb_5_8_io_dat_o[1] ,
    \cb_5_8_io_dat_o[0] }),
    .io_eo({\cb_5_8_io_eo[63] ,
    \cb_5_8_io_eo[62] ,
    \cb_5_8_io_eo[61] ,
    \cb_5_8_io_eo[60] ,
    \cb_5_8_io_eo[59] ,
    \cb_5_8_io_eo[58] ,
    \cb_5_8_io_eo[57] ,
    \cb_5_8_io_eo[56] ,
    \cb_5_8_io_eo[55] ,
    \cb_5_8_io_eo[54] ,
    \cb_5_8_io_eo[53] ,
    \cb_5_8_io_eo[52] ,
    \cb_5_8_io_eo[51] ,
    \cb_5_8_io_eo[50] ,
    \cb_5_8_io_eo[49] ,
    \cb_5_8_io_eo[48] ,
    \cb_5_8_io_eo[47] ,
    \cb_5_8_io_eo[46] ,
    \cb_5_8_io_eo[45] ,
    \cb_5_8_io_eo[44] ,
    \cb_5_8_io_eo[43] ,
    \cb_5_8_io_eo[42] ,
    \cb_5_8_io_eo[41] ,
    \cb_5_8_io_eo[40] ,
    \cb_5_8_io_eo[39] ,
    \cb_5_8_io_eo[38] ,
    \cb_5_8_io_eo[37] ,
    \cb_5_8_io_eo[36] ,
    \cb_5_8_io_eo[35] ,
    \cb_5_8_io_eo[34] ,
    \cb_5_8_io_eo[33] ,
    \cb_5_8_io_eo[32] ,
    \cb_5_8_io_eo[31] ,
    \cb_5_8_io_eo[30] ,
    \cb_5_8_io_eo[29] ,
    \cb_5_8_io_eo[28] ,
    \cb_5_8_io_eo[27] ,
    \cb_5_8_io_eo[26] ,
    \cb_5_8_io_eo[25] ,
    \cb_5_8_io_eo[24] ,
    \cb_5_8_io_eo[23] ,
    \cb_5_8_io_eo[22] ,
    \cb_5_8_io_eo[21] ,
    \cb_5_8_io_eo[20] ,
    \cb_5_8_io_eo[19] ,
    \cb_5_8_io_eo[18] ,
    \cb_5_8_io_eo[17] ,
    \cb_5_8_io_eo[16] ,
    \cb_5_8_io_eo[15] ,
    \cb_5_8_io_eo[14] ,
    \cb_5_8_io_eo[13] ,
    \cb_5_8_io_eo[12] ,
    \cb_5_8_io_eo[11] ,
    \cb_5_8_io_eo[10] ,
    \cb_5_8_io_eo[9] ,
    \cb_5_8_io_eo[8] ,
    \cb_5_8_io_eo[7] ,
    \cb_5_8_io_eo[6] ,
    \cb_5_8_io_eo[5] ,
    \cb_5_8_io_eo[4] ,
    \cb_5_8_io_eo[3] ,
    \cb_5_8_io_eo[2] ,
    \cb_5_8_io_eo[1] ,
    \cb_5_8_io_eo[0] }),
    .io_i_0_in1({\cb_5_7_io_o_0_out[7] ,
    \cb_5_7_io_o_0_out[6] ,
    \cb_5_7_io_o_0_out[5] ,
    \cb_5_7_io_o_0_out[4] ,
    \cb_5_7_io_o_0_out[3] ,
    \cb_5_7_io_o_0_out[2] ,
    \cb_5_7_io_o_0_out[1] ,
    \cb_5_7_io_o_0_out[0] }),
    .io_i_1_in1({\cb_5_7_io_o_1_out[7] ,
    \cb_5_7_io_o_1_out[6] ,
    \cb_5_7_io_o_1_out[5] ,
    \cb_5_7_io_o_1_out[4] ,
    \cb_5_7_io_o_1_out[3] ,
    \cb_5_7_io_o_1_out[2] ,
    \cb_5_7_io_o_1_out[1] ,
    \cb_5_7_io_o_1_out[0] }),
    .io_i_2_in1({\cb_5_7_io_o_2_out[7] ,
    \cb_5_7_io_o_2_out[6] ,
    \cb_5_7_io_o_2_out[5] ,
    \cb_5_7_io_o_2_out[4] ,
    \cb_5_7_io_o_2_out[3] ,
    \cb_5_7_io_o_2_out[2] ,
    \cb_5_7_io_o_2_out[1] ,
    \cb_5_7_io_o_2_out[0] }),
    .io_i_3_in1({\cb_5_7_io_o_3_out[7] ,
    \cb_5_7_io_o_3_out[6] ,
    \cb_5_7_io_o_3_out[5] ,
    \cb_5_7_io_o_3_out[4] ,
    \cb_5_7_io_o_3_out[3] ,
    \cb_5_7_io_o_3_out[2] ,
    \cb_5_7_io_o_3_out[1] ,
    \cb_5_7_io_o_3_out[0] }),
    .io_i_4_in1({\cb_5_7_io_o_4_out[7] ,
    \cb_5_7_io_o_4_out[6] ,
    \cb_5_7_io_o_4_out[5] ,
    \cb_5_7_io_o_4_out[4] ,
    \cb_5_7_io_o_4_out[3] ,
    \cb_5_7_io_o_4_out[2] ,
    \cb_5_7_io_o_4_out[1] ,
    \cb_5_7_io_o_4_out[0] }),
    .io_i_5_in1({\cb_5_7_io_o_5_out[7] ,
    \cb_5_7_io_o_5_out[6] ,
    \cb_5_7_io_o_5_out[5] ,
    \cb_5_7_io_o_5_out[4] ,
    \cb_5_7_io_o_5_out[3] ,
    \cb_5_7_io_o_5_out[2] ,
    \cb_5_7_io_o_5_out[1] ,
    \cb_5_7_io_o_5_out[0] }),
    .io_i_6_in1({\cb_5_7_io_o_6_out[7] ,
    \cb_5_7_io_o_6_out[6] ,
    \cb_5_7_io_o_6_out[5] ,
    \cb_5_7_io_o_6_out[4] ,
    \cb_5_7_io_o_6_out[3] ,
    \cb_5_7_io_o_6_out[2] ,
    \cb_5_7_io_o_6_out[1] ,
    \cb_5_7_io_o_6_out[0] }),
    .io_i_7_in1({\cb_5_7_io_o_7_out[7] ,
    \cb_5_7_io_o_7_out[6] ,
    \cb_5_7_io_o_7_out[5] ,
    \cb_5_7_io_o_7_out[4] ,
    \cb_5_7_io_o_7_out[3] ,
    \cb_5_7_io_o_7_out[2] ,
    \cb_5_7_io_o_7_out[1] ,
    \cb_5_7_io_o_7_out[0] }),
    .io_o_0_out({\cb_5_8_io_o_0_out[7] ,
    \cb_5_8_io_o_0_out[6] ,
    \cb_5_8_io_o_0_out[5] ,
    \cb_5_8_io_o_0_out[4] ,
    \cb_5_8_io_o_0_out[3] ,
    \cb_5_8_io_o_0_out[2] ,
    \cb_5_8_io_o_0_out[1] ,
    \cb_5_8_io_o_0_out[0] }),
    .io_o_1_out({\cb_5_8_io_o_1_out[7] ,
    \cb_5_8_io_o_1_out[6] ,
    \cb_5_8_io_o_1_out[5] ,
    \cb_5_8_io_o_1_out[4] ,
    \cb_5_8_io_o_1_out[3] ,
    \cb_5_8_io_o_1_out[2] ,
    \cb_5_8_io_o_1_out[1] ,
    \cb_5_8_io_o_1_out[0] }),
    .io_o_2_out({\cb_5_8_io_o_2_out[7] ,
    \cb_5_8_io_o_2_out[6] ,
    \cb_5_8_io_o_2_out[5] ,
    \cb_5_8_io_o_2_out[4] ,
    \cb_5_8_io_o_2_out[3] ,
    \cb_5_8_io_o_2_out[2] ,
    \cb_5_8_io_o_2_out[1] ,
    \cb_5_8_io_o_2_out[0] }),
    .io_o_3_out({\cb_5_8_io_o_3_out[7] ,
    \cb_5_8_io_o_3_out[6] ,
    \cb_5_8_io_o_3_out[5] ,
    \cb_5_8_io_o_3_out[4] ,
    \cb_5_8_io_o_3_out[3] ,
    \cb_5_8_io_o_3_out[2] ,
    \cb_5_8_io_o_3_out[1] ,
    \cb_5_8_io_o_3_out[0] }),
    .io_o_4_out({\cb_5_8_io_o_4_out[7] ,
    \cb_5_8_io_o_4_out[6] ,
    \cb_5_8_io_o_4_out[5] ,
    \cb_5_8_io_o_4_out[4] ,
    \cb_5_8_io_o_4_out[3] ,
    \cb_5_8_io_o_4_out[2] ,
    \cb_5_8_io_o_4_out[1] ,
    \cb_5_8_io_o_4_out[0] }),
    .io_o_5_out({\cb_5_8_io_o_5_out[7] ,
    \cb_5_8_io_o_5_out[6] ,
    \cb_5_8_io_o_5_out[5] ,
    \cb_5_8_io_o_5_out[4] ,
    \cb_5_8_io_o_5_out[3] ,
    \cb_5_8_io_o_5_out[2] ,
    \cb_5_8_io_o_5_out[1] ,
    \cb_5_8_io_o_5_out[0] }),
    .io_o_6_out({\cb_5_8_io_o_6_out[7] ,
    \cb_5_8_io_o_6_out[6] ,
    \cb_5_8_io_o_6_out[5] ,
    \cb_5_8_io_o_6_out[4] ,
    \cb_5_8_io_o_6_out[3] ,
    \cb_5_8_io_o_6_out[2] ,
    \cb_5_8_io_o_6_out[1] ,
    \cb_5_8_io_o_6_out[0] }),
    .io_o_7_out({\cb_5_8_io_o_7_out[7] ,
    \cb_5_8_io_o_7_out[6] ,
    \cb_5_8_io_o_7_out[5] ,
    \cb_5_8_io_o_7_out[4] ,
    \cb_5_8_io_o_7_out[3] ,
    \cb_5_8_io_o_7_out[2] ,
    \cb_5_8_io_o_7_out[1] ,
    \cb_5_8_io_o_7_out[0] }),
    .io_wo({\cb_5_7_io_eo[63] ,
    \cb_5_7_io_eo[62] ,
    \cb_5_7_io_eo[61] ,
    \cb_5_7_io_eo[60] ,
    \cb_5_7_io_eo[59] ,
    \cb_5_7_io_eo[58] ,
    \cb_5_7_io_eo[57] ,
    \cb_5_7_io_eo[56] ,
    \cb_5_7_io_eo[55] ,
    \cb_5_7_io_eo[54] ,
    \cb_5_7_io_eo[53] ,
    \cb_5_7_io_eo[52] ,
    \cb_5_7_io_eo[51] ,
    \cb_5_7_io_eo[50] ,
    \cb_5_7_io_eo[49] ,
    \cb_5_7_io_eo[48] ,
    \cb_5_7_io_eo[47] ,
    \cb_5_7_io_eo[46] ,
    \cb_5_7_io_eo[45] ,
    \cb_5_7_io_eo[44] ,
    \cb_5_7_io_eo[43] ,
    \cb_5_7_io_eo[42] ,
    \cb_5_7_io_eo[41] ,
    \cb_5_7_io_eo[40] ,
    \cb_5_7_io_eo[39] ,
    \cb_5_7_io_eo[38] ,
    \cb_5_7_io_eo[37] ,
    \cb_5_7_io_eo[36] ,
    \cb_5_7_io_eo[35] ,
    \cb_5_7_io_eo[34] ,
    \cb_5_7_io_eo[33] ,
    \cb_5_7_io_eo[32] ,
    \cb_5_7_io_eo[31] ,
    \cb_5_7_io_eo[30] ,
    \cb_5_7_io_eo[29] ,
    \cb_5_7_io_eo[28] ,
    \cb_5_7_io_eo[27] ,
    \cb_5_7_io_eo[26] ,
    \cb_5_7_io_eo[25] ,
    \cb_5_7_io_eo[24] ,
    \cb_5_7_io_eo[23] ,
    \cb_5_7_io_eo[22] ,
    \cb_5_7_io_eo[21] ,
    \cb_5_7_io_eo[20] ,
    \cb_5_7_io_eo[19] ,
    \cb_5_7_io_eo[18] ,
    \cb_5_7_io_eo[17] ,
    \cb_5_7_io_eo[16] ,
    \cb_5_7_io_eo[15] ,
    \cb_5_7_io_eo[14] ,
    \cb_5_7_io_eo[13] ,
    \cb_5_7_io_eo[12] ,
    \cb_5_7_io_eo[11] ,
    \cb_5_7_io_eo[10] ,
    \cb_5_7_io_eo[9] ,
    \cb_5_7_io_eo[8] ,
    \cb_5_7_io_eo[7] ,
    \cb_5_7_io_eo[6] ,
    \cb_5_7_io_eo[5] ,
    \cb_5_7_io_eo[4] ,
    \cb_5_7_io_eo[3] ,
    \cb_5_7_io_eo[2] ,
    \cb_5_7_io_eo[1] ,
    \cb_5_7_io_eo[0] }));
 cic_block cb_5_9 (.io_cs_i(cb_5_9_io_cs_i),
    .io_i_0_ci(cb_5_8_io_o_0_co),
    .io_i_1_ci(cb_5_8_io_o_1_co),
    .io_i_2_ci(cb_5_8_io_o_2_co),
    .io_i_3_ci(cb_5_8_io_o_3_co),
    .io_i_4_ci(cb_5_8_io_o_4_co),
    .io_i_5_ci(cb_5_8_io_o_5_co),
    .io_i_6_ci(cb_5_8_io_o_6_co),
    .io_i_7_ci(cb_5_8_io_o_7_co),
    .io_o_0_co(cb_5_10_io_i_0_ci),
    .io_o_1_co(cb_5_10_io_i_1_ci),
    .io_o_2_co(cb_5_10_io_i_2_ci),
    .io_o_3_co(cb_5_10_io_i_3_ci),
    .io_o_4_co(cb_5_10_io_i_4_ci),
    .io_o_5_co(cb_5_10_io_i_5_ci),
    .io_o_6_co(cb_5_10_io_i_6_ci),
    .io_o_7_co(cb_5_10_io_i_7_ci),
    .io_vci(cb_5_8_io_vco),
    .io_vco(cb_5_10_io_vci),
    .io_vi(cb_5_9_io_vi),
    .io_we_i(cb_5_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_5_0_io_adr_i[1] ,
    \cb_5_0_io_adr_i[0] }),
    .io_dat_i({\cb_5_0_io_dat_i[15] ,
    \cb_5_0_io_dat_i[14] ,
    \cb_5_0_io_dat_i[13] ,
    \cb_5_0_io_dat_i[12] ,
    \cb_5_0_io_dat_i[11] ,
    \cb_5_0_io_dat_i[10] ,
    \cb_5_0_io_dat_i[9] ,
    \cb_5_0_io_dat_i[8] ,
    \cb_5_0_io_dat_i[7] ,
    \cb_5_0_io_dat_i[6] ,
    \cb_5_0_io_dat_i[5] ,
    \cb_5_0_io_dat_i[4] ,
    \cb_5_0_io_dat_i[3] ,
    \cb_5_0_io_dat_i[2] ,
    \cb_5_0_io_dat_i[1] ,
    \cb_5_0_io_dat_i[0] }),
    .io_dat_o({\cb_5_9_io_dat_o[15] ,
    \cb_5_9_io_dat_o[14] ,
    \cb_5_9_io_dat_o[13] ,
    \cb_5_9_io_dat_o[12] ,
    \cb_5_9_io_dat_o[11] ,
    \cb_5_9_io_dat_o[10] ,
    \cb_5_9_io_dat_o[9] ,
    \cb_5_9_io_dat_o[8] ,
    \cb_5_9_io_dat_o[7] ,
    \cb_5_9_io_dat_o[6] ,
    \cb_5_9_io_dat_o[5] ,
    \cb_5_9_io_dat_o[4] ,
    \cb_5_9_io_dat_o[3] ,
    \cb_5_9_io_dat_o[2] ,
    \cb_5_9_io_dat_o[1] ,
    \cb_5_9_io_dat_o[0] }),
    .io_eo({\cb_5_10_io_wo[63] ,
    \cb_5_10_io_wo[62] ,
    \cb_5_10_io_wo[61] ,
    \cb_5_10_io_wo[60] ,
    \cb_5_10_io_wo[59] ,
    \cb_5_10_io_wo[58] ,
    \cb_5_10_io_wo[57] ,
    \cb_5_10_io_wo[56] ,
    \cb_5_10_io_wo[55] ,
    \cb_5_10_io_wo[54] ,
    \cb_5_10_io_wo[53] ,
    \cb_5_10_io_wo[52] ,
    \cb_5_10_io_wo[51] ,
    \cb_5_10_io_wo[50] ,
    \cb_5_10_io_wo[49] ,
    \cb_5_10_io_wo[48] ,
    \cb_5_10_io_wo[47] ,
    \cb_5_10_io_wo[46] ,
    \cb_5_10_io_wo[45] ,
    \cb_5_10_io_wo[44] ,
    \cb_5_10_io_wo[43] ,
    \cb_5_10_io_wo[42] ,
    \cb_5_10_io_wo[41] ,
    \cb_5_10_io_wo[40] ,
    \cb_5_10_io_wo[39] ,
    \cb_5_10_io_wo[38] ,
    \cb_5_10_io_wo[37] ,
    \cb_5_10_io_wo[36] ,
    \cb_5_10_io_wo[35] ,
    \cb_5_10_io_wo[34] ,
    \cb_5_10_io_wo[33] ,
    \cb_5_10_io_wo[32] ,
    \cb_5_10_io_wo[31] ,
    \cb_5_10_io_wo[30] ,
    \cb_5_10_io_wo[29] ,
    \cb_5_10_io_wo[28] ,
    \cb_5_10_io_wo[27] ,
    \cb_5_10_io_wo[26] ,
    \cb_5_10_io_wo[25] ,
    \cb_5_10_io_wo[24] ,
    \cb_5_10_io_wo[23] ,
    \cb_5_10_io_wo[22] ,
    \cb_5_10_io_wo[21] ,
    \cb_5_10_io_wo[20] ,
    \cb_5_10_io_wo[19] ,
    \cb_5_10_io_wo[18] ,
    \cb_5_10_io_wo[17] ,
    \cb_5_10_io_wo[16] ,
    \cb_5_10_io_wo[15] ,
    \cb_5_10_io_wo[14] ,
    \cb_5_10_io_wo[13] ,
    \cb_5_10_io_wo[12] ,
    \cb_5_10_io_wo[11] ,
    \cb_5_10_io_wo[10] ,
    \cb_5_10_io_wo[9] ,
    \cb_5_10_io_wo[8] ,
    \cb_5_10_io_wo[7] ,
    \cb_5_10_io_wo[6] ,
    \cb_5_10_io_wo[5] ,
    \cb_5_10_io_wo[4] ,
    \cb_5_10_io_wo[3] ,
    \cb_5_10_io_wo[2] ,
    \cb_5_10_io_wo[1] ,
    \cb_5_10_io_wo[0] }),
    .io_i_0_in1({\cb_5_8_io_o_0_out[7] ,
    \cb_5_8_io_o_0_out[6] ,
    \cb_5_8_io_o_0_out[5] ,
    \cb_5_8_io_o_0_out[4] ,
    \cb_5_8_io_o_0_out[3] ,
    \cb_5_8_io_o_0_out[2] ,
    \cb_5_8_io_o_0_out[1] ,
    \cb_5_8_io_o_0_out[0] }),
    .io_i_1_in1({\cb_5_8_io_o_1_out[7] ,
    \cb_5_8_io_o_1_out[6] ,
    \cb_5_8_io_o_1_out[5] ,
    \cb_5_8_io_o_1_out[4] ,
    \cb_5_8_io_o_1_out[3] ,
    \cb_5_8_io_o_1_out[2] ,
    \cb_5_8_io_o_1_out[1] ,
    \cb_5_8_io_o_1_out[0] }),
    .io_i_2_in1({\cb_5_8_io_o_2_out[7] ,
    \cb_5_8_io_o_2_out[6] ,
    \cb_5_8_io_o_2_out[5] ,
    \cb_5_8_io_o_2_out[4] ,
    \cb_5_8_io_o_2_out[3] ,
    \cb_5_8_io_o_2_out[2] ,
    \cb_5_8_io_o_2_out[1] ,
    \cb_5_8_io_o_2_out[0] }),
    .io_i_3_in1({\cb_5_8_io_o_3_out[7] ,
    \cb_5_8_io_o_3_out[6] ,
    \cb_5_8_io_o_3_out[5] ,
    \cb_5_8_io_o_3_out[4] ,
    \cb_5_8_io_o_3_out[3] ,
    \cb_5_8_io_o_3_out[2] ,
    \cb_5_8_io_o_3_out[1] ,
    \cb_5_8_io_o_3_out[0] }),
    .io_i_4_in1({\cb_5_8_io_o_4_out[7] ,
    \cb_5_8_io_o_4_out[6] ,
    \cb_5_8_io_o_4_out[5] ,
    \cb_5_8_io_o_4_out[4] ,
    \cb_5_8_io_o_4_out[3] ,
    \cb_5_8_io_o_4_out[2] ,
    \cb_5_8_io_o_4_out[1] ,
    \cb_5_8_io_o_4_out[0] }),
    .io_i_5_in1({\cb_5_8_io_o_5_out[7] ,
    \cb_5_8_io_o_5_out[6] ,
    \cb_5_8_io_o_5_out[5] ,
    \cb_5_8_io_o_5_out[4] ,
    \cb_5_8_io_o_5_out[3] ,
    \cb_5_8_io_o_5_out[2] ,
    \cb_5_8_io_o_5_out[1] ,
    \cb_5_8_io_o_5_out[0] }),
    .io_i_6_in1({\cb_5_8_io_o_6_out[7] ,
    \cb_5_8_io_o_6_out[6] ,
    \cb_5_8_io_o_6_out[5] ,
    \cb_5_8_io_o_6_out[4] ,
    \cb_5_8_io_o_6_out[3] ,
    \cb_5_8_io_o_6_out[2] ,
    \cb_5_8_io_o_6_out[1] ,
    \cb_5_8_io_o_6_out[0] }),
    .io_i_7_in1({\cb_5_8_io_o_7_out[7] ,
    \cb_5_8_io_o_7_out[6] ,
    \cb_5_8_io_o_7_out[5] ,
    \cb_5_8_io_o_7_out[4] ,
    \cb_5_8_io_o_7_out[3] ,
    \cb_5_8_io_o_7_out[2] ,
    \cb_5_8_io_o_7_out[1] ,
    \cb_5_8_io_o_7_out[0] }),
    .io_o_0_out({\cb_5_10_io_i_0_in1[7] ,
    \cb_5_10_io_i_0_in1[6] ,
    \cb_5_10_io_i_0_in1[5] ,
    \cb_5_10_io_i_0_in1[4] ,
    \cb_5_10_io_i_0_in1[3] ,
    \cb_5_10_io_i_0_in1[2] ,
    \cb_5_10_io_i_0_in1[1] ,
    \cb_5_10_io_i_0_in1[0] }),
    .io_o_1_out({\cb_5_10_io_i_1_in1[7] ,
    \cb_5_10_io_i_1_in1[6] ,
    \cb_5_10_io_i_1_in1[5] ,
    \cb_5_10_io_i_1_in1[4] ,
    \cb_5_10_io_i_1_in1[3] ,
    \cb_5_10_io_i_1_in1[2] ,
    \cb_5_10_io_i_1_in1[1] ,
    \cb_5_10_io_i_1_in1[0] }),
    .io_o_2_out({\cb_5_10_io_i_2_in1[7] ,
    \cb_5_10_io_i_2_in1[6] ,
    \cb_5_10_io_i_2_in1[5] ,
    \cb_5_10_io_i_2_in1[4] ,
    \cb_5_10_io_i_2_in1[3] ,
    \cb_5_10_io_i_2_in1[2] ,
    \cb_5_10_io_i_2_in1[1] ,
    \cb_5_10_io_i_2_in1[0] }),
    .io_o_3_out({\cb_5_10_io_i_3_in1[7] ,
    \cb_5_10_io_i_3_in1[6] ,
    \cb_5_10_io_i_3_in1[5] ,
    \cb_5_10_io_i_3_in1[4] ,
    \cb_5_10_io_i_3_in1[3] ,
    \cb_5_10_io_i_3_in1[2] ,
    \cb_5_10_io_i_3_in1[1] ,
    \cb_5_10_io_i_3_in1[0] }),
    .io_o_4_out({\cb_5_10_io_i_4_in1[7] ,
    \cb_5_10_io_i_4_in1[6] ,
    \cb_5_10_io_i_4_in1[5] ,
    \cb_5_10_io_i_4_in1[4] ,
    \cb_5_10_io_i_4_in1[3] ,
    \cb_5_10_io_i_4_in1[2] ,
    \cb_5_10_io_i_4_in1[1] ,
    \cb_5_10_io_i_4_in1[0] }),
    .io_o_5_out({\cb_5_10_io_i_5_in1[7] ,
    \cb_5_10_io_i_5_in1[6] ,
    \cb_5_10_io_i_5_in1[5] ,
    \cb_5_10_io_i_5_in1[4] ,
    \cb_5_10_io_i_5_in1[3] ,
    \cb_5_10_io_i_5_in1[2] ,
    \cb_5_10_io_i_5_in1[1] ,
    \cb_5_10_io_i_5_in1[0] }),
    .io_o_6_out({\cb_5_10_io_i_6_in1[7] ,
    \cb_5_10_io_i_6_in1[6] ,
    \cb_5_10_io_i_6_in1[5] ,
    \cb_5_10_io_i_6_in1[4] ,
    \cb_5_10_io_i_6_in1[3] ,
    \cb_5_10_io_i_6_in1[2] ,
    \cb_5_10_io_i_6_in1[1] ,
    \cb_5_10_io_i_6_in1[0] }),
    .io_o_7_out({\cb_5_10_io_i_7_in1[7] ,
    \cb_5_10_io_i_7_in1[6] ,
    \cb_5_10_io_i_7_in1[5] ,
    \cb_5_10_io_i_7_in1[4] ,
    \cb_5_10_io_i_7_in1[3] ,
    \cb_5_10_io_i_7_in1[2] ,
    \cb_5_10_io_i_7_in1[1] ,
    \cb_5_10_io_i_7_in1[0] }),
    .io_wo({\cb_5_8_io_eo[63] ,
    \cb_5_8_io_eo[62] ,
    \cb_5_8_io_eo[61] ,
    \cb_5_8_io_eo[60] ,
    \cb_5_8_io_eo[59] ,
    \cb_5_8_io_eo[58] ,
    \cb_5_8_io_eo[57] ,
    \cb_5_8_io_eo[56] ,
    \cb_5_8_io_eo[55] ,
    \cb_5_8_io_eo[54] ,
    \cb_5_8_io_eo[53] ,
    \cb_5_8_io_eo[52] ,
    \cb_5_8_io_eo[51] ,
    \cb_5_8_io_eo[50] ,
    \cb_5_8_io_eo[49] ,
    \cb_5_8_io_eo[48] ,
    \cb_5_8_io_eo[47] ,
    \cb_5_8_io_eo[46] ,
    \cb_5_8_io_eo[45] ,
    \cb_5_8_io_eo[44] ,
    \cb_5_8_io_eo[43] ,
    \cb_5_8_io_eo[42] ,
    \cb_5_8_io_eo[41] ,
    \cb_5_8_io_eo[40] ,
    \cb_5_8_io_eo[39] ,
    \cb_5_8_io_eo[38] ,
    \cb_5_8_io_eo[37] ,
    \cb_5_8_io_eo[36] ,
    \cb_5_8_io_eo[35] ,
    \cb_5_8_io_eo[34] ,
    \cb_5_8_io_eo[33] ,
    \cb_5_8_io_eo[32] ,
    \cb_5_8_io_eo[31] ,
    \cb_5_8_io_eo[30] ,
    \cb_5_8_io_eo[29] ,
    \cb_5_8_io_eo[28] ,
    \cb_5_8_io_eo[27] ,
    \cb_5_8_io_eo[26] ,
    \cb_5_8_io_eo[25] ,
    \cb_5_8_io_eo[24] ,
    \cb_5_8_io_eo[23] ,
    \cb_5_8_io_eo[22] ,
    \cb_5_8_io_eo[21] ,
    \cb_5_8_io_eo[20] ,
    \cb_5_8_io_eo[19] ,
    \cb_5_8_io_eo[18] ,
    \cb_5_8_io_eo[17] ,
    \cb_5_8_io_eo[16] ,
    \cb_5_8_io_eo[15] ,
    \cb_5_8_io_eo[14] ,
    \cb_5_8_io_eo[13] ,
    \cb_5_8_io_eo[12] ,
    \cb_5_8_io_eo[11] ,
    \cb_5_8_io_eo[10] ,
    \cb_5_8_io_eo[9] ,
    \cb_5_8_io_eo[8] ,
    \cb_5_8_io_eo[7] ,
    \cb_5_8_io_eo[6] ,
    \cb_5_8_io_eo[5] ,
    \cb_5_8_io_eo[4] ,
    \cb_5_8_io_eo[3] ,
    \cb_5_8_io_eo[2] ,
    \cb_5_8_io_eo[1] ,
    \cb_5_8_io_eo[0] }));
 cic_block cb_6_0 (.io_cs_i(cb_6_0_io_cs_i),
    .io_i_0_ci(cb_6_0_io_i_0_ci),
    .io_o_0_co(cb_6_0_io_o_0_co),
    .io_o_1_co(cb_6_0_io_o_1_co),
    .io_o_2_co(cb_6_0_io_o_2_co),
    .io_o_3_co(cb_6_0_io_o_3_co),
    .io_o_4_co(cb_6_0_io_o_4_co),
    .io_o_5_co(cb_6_0_io_o_5_co),
    .io_o_6_co(cb_6_0_io_o_6_co),
    .io_o_7_co(cb_6_0_io_o_7_co),
    .io_vco(cb_6_0_io_vco),
    .io_vi(cb_6_0_io_vi),
    .io_we_i(cb_6_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_6_0_io_adr_i[1] ,
    \cb_6_0_io_adr_i[0] }),
    .io_dat_i({\cb_6_0_io_dat_i[15] ,
    \cb_6_0_io_dat_i[14] ,
    \cb_6_0_io_dat_i[13] ,
    \cb_6_0_io_dat_i[12] ,
    \cb_6_0_io_dat_i[11] ,
    \cb_6_0_io_dat_i[10] ,
    \cb_6_0_io_dat_i[9] ,
    \cb_6_0_io_dat_i[8] ,
    \cb_6_0_io_dat_i[7] ,
    \cb_6_0_io_dat_i[6] ,
    \cb_6_0_io_dat_i[5] ,
    \cb_6_0_io_dat_i[4] ,
    \cb_6_0_io_dat_i[3] ,
    \cb_6_0_io_dat_i[2] ,
    \cb_6_0_io_dat_i[1] ,
    \cb_6_0_io_dat_i[0] }),
    .io_dat_o({\cb_6_0_io_dat_o[15] ,
    \cb_6_0_io_dat_o[14] ,
    \cb_6_0_io_dat_o[13] ,
    \cb_6_0_io_dat_o[12] ,
    \cb_6_0_io_dat_o[11] ,
    \cb_6_0_io_dat_o[10] ,
    \cb_6_0_io_dat_o[9] ,
    \cb_6_0_io_dat_o[8] ,
    \cb_6_0_io_dat_o[7] ,
    \cb_6_0_io_dat_o[6] ,
    \cb_6_0_io_dat_o[5] ,
    \cb_6_0_io_dat_o[4] ,
    \cb_6_0_io_dat_o[3] ,
    \cb_6_0_io_dat_o[2] ,
    \cb_6_0_io_dat_o[1] ,
    \cb_6_0_io_dat_o[0] }),
    .io_eo({\cb_6_0_io_eo[63] ,
    \cb_6_0_io_eo[62] ,
    \cb_6_0_io_eo[61] ,
    \cb_6_0_io_eo[60] ,
    \cb_6_0_io_eo[59] ,
    \cb_6_0_io_eo[58] ,
    \cb_6_0_io_eo[57] ,
    \cb_6_0_io_eo[56] ,
    \cb_6_0_io_eo[55] ,
    \cb_6_0_io_eo[54] ,
    \cb_6_0_io_eo[53] ,
    \cb_6_0_io_eo[52] ,
    \cb_6_0_io_eo[51] ,
    \cb_6_0_io_eo[50] ,
    \cb_6_0_io_eo[49] ,
    \cb_6_0_io_eo[48] ,
    \cb_6_0_io_eo[47] ,
    \cb_6_0_io_eo[46] ,
    \cb_6_0_io_eo[45] ,
    \cb_6_0_io_eo[44] ,
    \cb_6_0_io_eo[43] ,
    \cb_6_0_io_eo[42] ,
    \cb_6_0_io_eo[41] ,
    \cb_6_0_io_eo[40] ,
    \cb_6_0_io_eo[39] ,
    \cb_6_0_io_eo[38] ,
    \cb_6_0_io_eo[37] ,
    \cb_6_0_io_eo[36] ,
    \cb_6_0_io_eo[35] ,
    \cb_6_0_io_eo[34] ,
    \cb_6_0_io_eo[33] ,
    \cb_6_0_io_eo[32] ,
    \cb_6_0_io_eo[31] ,
    \cb_6_0_io_eo[30] ,
    \cb_6_0_io_eo[29] ,
    \cb_6_0_io_eo[28] ,
    \cb_6_0_io_eo[27] ,
    \cb_6_0_io_eo[26] ,
    \cb_6_0_io_eo[25] ,
    \cb_6_0_io_eo[24] ,
    \cb_6_0_io_eo[23] ,
    \cb_6_0_io_eo[22] ,
    \cb_6_0_io_eo[21] ,
    \cb_6_0_io_eo[20] ,
    \cb_6_0_io_eo[19] ,
    \cb_6_0_io_eo[18] ,
    \cb_6_0_io_eo[17] ,
    \cb_6_0_io_eo[16] ,
    \cb_6_0_io_eo[15] ,
    \cb_6_0_io_eo[14] ,
    \cb_6_0_io_eo[13] ,
    \cb_6_0_io_eo[12] ,
    \cb_6_0_io_eo[11] ,
    \cb_6_0_io_eo[10] ,
    \cb_6_0_io_eo[9] ,
    \cb_6_0_io_eo[8] ,
    \cb_6_0_io_eo[7] ,
    \cb_6_0_io_eo[6] ,
    \cb_6_0_io_eo[5] ,
    \cb_6_0_io_eo[4] ,
    \cb_6_0_io_eo[3] ,
    \cb_6_0_io_eo[2] ,
    \cb_6_0_io_eo[1] ,
    \cb_6_0_io_eo[0] }),
    .io_i_0_in1({_NC385,
    _NC386,
    _NC387,
    _NC388,
    _NC389,
    _NC390,
    _NC391,
    _NC392}),
    .io_i_1_in1({_NC393,
    _NC394,
    _NC395,
    _NC396,
    _NC397,
    _NC398,
    _NC399,
    _NC400}),
    .io_i_2_in1({_NC401,
    _NC402,
    _NC403,
    _NC404,
    _NC405,
    _NC406,
    _NC407,
    _NC408}),
    .io_i_3_in1({_NC409,
    _NC410,
    _NC411,
    _NC412,
    _NC413,
    _NC414,
    _NC415,
    _NC416}),
    .io_i_4_in1({_NC417,
    _NC418,
    _NC419,
    _NC420,
    _NC421,
    _NC422,
    _NC423,
    _NC424}),
    .io_i_5_in1({_NC425,
    _NC426,
    _NC427,
    _NC428,
    _NC429,
    _NC430,
    _NC431,
    _NC432}),
    .io_i_6_in1({_NC433,
    _NC434,
    _NC435,
    _NC436,
    _NC437,
    _NC438,
    _NC439,
    _NC440}),
    .io_i_7_in1({_NC441,
    _NC442,
    _NC443,
    _NC444,
    _NC445,
    _NC446,
    _NC447,
    _NC448}),
    .io_o_0_out({\cb_6_0_io_o_0_out[7] ,
    \cb_6_0_io_o_0_out[6] ,
    \cb_6_0_io_o_0_out[5] ,
    \cb_6_0_io_o_0_out[4] ,
    \cb_6_0_io_o_0_out[3] ,
    \cb_6_0_io_o_0_out[2] ,
    \cb_6_0_io_o_0_out[1] ,
    \cb_6_0_io_o_0_out[0] }),
    .io_o_1_out({\cb_6_0_io_o_1_out[7] ,
    \cb_6_0_io_o_1_out[6] ,
    \cb_6_0_io_o_1_out[5] ,
    \cb_6_0_io_o_1_out[4] ,
    \cb_6_0_io_o_1_out[3] ,
    \cb_6_0_io_o_1_out[2] ,
    \cb_6_0_io_o_1_out[1] ,
    \cb_6_0_io_o_1_out[0] }),
    .io_o_2_out({\cb_6_0_io_o_2_out[7] ,
    \cb_6_0_io_o_2_out[6] ,
    \cb_6_0_io_o_2_out[5] ,
    \cb_6_0_io_o_2_out[4] ,
    \cb_6_0_io_o_2_out[3] ,
    \cb_6_0_io_o_2_out[2] ,
    \cb_6_0_io_o_2_out[1] ,
    \cb_6_0_io_o_2_out[0] }),
    .io_o_3_out({\cb_6_0_io_o_3_out[7] ,
    \cb_6_0_io_o_3_out[6] ,
    \cb_6_0_io_o_3_out[5] ,
    \cb_6_0_io_o_3_out[4] ,
    \cb_6_0_io_o_3_out[3] ,
    \cb_6_0_io_o_3_out[2] ,
    \cb_6_0_io_o_3_out[1] ,
    \cb_6_0_io_o_3_out[0] }),
    .io_o_4_out({\cb_6_0_io_o_4_out[7] ,
    \cb_6_0_io_o_4_out[6] ,
    \cb_6_0_io_o_4_out[5] ,
    \cb_6_0_io_o_4_out[4] ,
    \cb_6_0_io_o_4_out[3] ,
    \cb_6_0_io_o_4_out[2] ,
    \cb_6_0_io_o_4_out[1] ,
    \cb_6_0_io_o_4_out[0] }),
    .io_o_5_out({\cb_6_0_io_o_5_out[7] ,
    \cb_6_0_io_o_5_out[6] ,
    \cb_6_0_io_o_5_out[5] ,
    \cb_6_0_io_o_5_out[4] ,
    \cb_6_0_io_o_5_out[3] ,
    \cb_6_0_io_o_5_out[2] ,
    \cb_6_0_io_o_5_out[1] ,
    \cb_6_0_io_o_5_out[0] }),
    .io_o_6_out({\cb_6_0_io_o_6_out[7] ,
    \cb_6_0_io_o_6_out[6] ,
    \cb_6_0_io_o_6_out[5] ,
    \cb_6_0_io_o_6_out[4] ,
    \cb_6_0_io_o_6_out[3] ,
    \cb_6_0_io_o_6_out[2] ,
    \cb_6_0_io_o_6_out[1] ,
    \cb_6_0_io_o_6_out[0] }),
    .io_o_7_out({\cb_6_0_io_o_7_out[7] ,
    \cb_6_0_io_o_7_out[6] ,
    \cb_6_0_io_o_7_out[5] ,
    \cb_6_0_io_o_7_out[4] ,
    \cb_6_0_io_o_7_out[3] ,
    \cb_6_0_io_o_7_out[2] ,
    \cb_6_0_io_o_7_out[1] ,
    \cb_6_0_io_o_7_out[0] }),
    .io_wo({\cb_6_0_io_wo[63] ,
    \cb_6_0_io_wo[62] ,
    \cb_6_0_io_wo[61] ,
    \cb_6_0_io_wo[60] ,
    \cb_6_0_io_wo[59] ,
    \cb_6_0_io_wo[58] ,
    \cb_6_0_io_wo[57] ,
    \cb_6_0_io_wo[56] ,
    \cb_6_0_io_wo[55] ,
    \cb_6_0_io_wo[54] ,
    \cb_6_0_io_wo[53] ,
    \cb_6_0_io_wo[52] ,
    \cb_6_0_io_wo[51] ,
    \cb_6_0_io_wo[50] ,
    \cb_6_0_io_wo[49] ,
    \cb_6_0_io_wo[48] ,
    \cb_6_0_io_wo[47] ,
    \cb_6_0_io_wo[46] ,
    \cb_6_0_io_wo[45] ,
    \cb_6_0_io_wo[44] ,
    \cb_6_0_io_wo[43] ,
    \cb_6_0_io_wo[42] ,
    \cb_6_0_io_wo[41] ,
    \cb_6_0_io_wo[40] ,
    \cb_6_0_io_wo[39] ,
    \cb_6_0_io_wo[38] ,
    \cb_6_0_io_wo[37] ,
    \cb_6_0_io_wo[36] ,
    \cb_6_0_io_wo[35] ,
    \cb_6_0_io_wo[34] ,
    \cb_6_0_io_wo[33] ,
    \cb_6_0_io_wo[32] ,
    \cb_6_0_io_wo[31] ,
    \cb_6_0_io_wo[30] ,
    \cb_6_0_io_wo[29] ,
    \cb_6_0_io_wo[28] ,
    \cb_6_0_io_wo[27] ,
    \cb_6_0_io_wo[26] ,
    \cb_6_0_io_wo[25] ,
    \cb_6_0_io_wo[24] ,
    \cb_6_0_io_wo[23] ,
    \cb_6_0_io_wo[22] ,
    \cb_6_0_io_wo[21] ,
    \cb_6_0_io_wo[20] ,
    \cb_6_0_io_wo[19] ,
    \cb_6_0_io_wo[18] ,
    \cb_6_0_io_wo[17] ,
    \cb_6_0_io_wo[16] ,
    \cb_6_0_io_wo[15] ,
    \cb_6_0_io_wo[14] ,
    \cb_6_0_io_wo[13] ,
    \cb_6_0_io_wo[12] ,
    \cb_6_0_io_wo[11] ,
    \cb_6_0_io_wo[10] ,
    \cb_6_0_io_wo[9] ,
    \cb_6_0_io_wo[8] ,
    \cb_6_0_io_wo[7] ,
    \cb_6_0_io_wo[6] ,
    \cb_6_0_io_wo[5] ,
    \cb_6_0_io_wo[4] ,
    \cb_6_0_io_wo[3] ,
    \cb_6_0_io_wo[2] ,
    \cb_6_0_io_wo[1] ,
    \cb_6_0_io_wo[0] }));
 cic_block cb_6_1 (.io_cs_i(cb_6_1_io_cs_i),
    .io_i_0_ci(cb_6_0_io_o_0_co),
    .io_i_1_ci(cb_6_0_io_o_1_co),
    .io_i_2_ci(cb_6_0_io_o_2_co),
    .io_i_3_ci(cb_6_0_io_o_3_co),
    .io_i_4_ci(cb_6_0_io_o_4_co),
    .io_i_5_ci(cb_6_0_io_o_5_co),
    .io_i_6_ci(cb_6_0_io_o_6_co),
    .io_i_7_ci(cb_6_0_io_o_7_co),
    .io_o_0_co(cb_6_1_io_o_0_co),
    .io_o_1_co(cb_6_1_io_o_1_co),
    .io_o_2_co(cb_6_1_io_o_2_co),
    .io_o_3_co(cb_6_1_io_o_3_co),
    .io_o_4_co(cb_6_1_io_o_4_co),
    .io_o_5_co(cb_6_1_io_o_5_co),
    .io_o_6_co(cb_6_1_io_o_6_co),
    .io_o_7_co(cb_6_1_io_o_7_co),
    .io_vci(cb_6_0_io_vco),
    .io_vco(cb_6_1_io_vco),
    .io_vi(cb_6_1_io_vi),
    .io_we_i(cb_6_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_6_0_io_adr_i[1] ,
    \cb_6_0_io_adr_i[0] }),
    .io_dat_i({\cb_6_0_io_dat_i[15] ,
    \cb_6_0_io_dat_i[14] ,
    \cb_6_0_io_dat_i[13] ,
    \cb_6_0_io_dat_i[12] ,
    \cb_6_0_io_dat_i[11] ,
    \cb_6_0_io_dat_i[10] ,
    \cb_6_0_io_dat_i[9] ,
    \cb_6_0_io_dat_i[8] ,
    \cb_6_0_io_dat_i[7] ,
    \cb_6_0_io_dat_i[6] ,
    \cb_6_0_io_dat_i[5] ,
    \cb_6_0_io_dat_i[4] ,
    \cb_6_0_io_dat_i[3] ,
    \cb_6_0_io_dat_i[2] ,
    \cb_6_0_io_dat_i[1] ,
    \cb_6_0_io_dat_i[0] }),
    .io_dat_o({\cb_6_1_io_dat_o[15] ,
    \cb_6_1_io_dat_o[14] ,
    \cb_6_1_io_dat_o[13] ,
    \cb_6_1_io_dat_o[12] ,
    \cb_6_1_io_dat_o[11] ,
    \cb_6_1_io_dat_o[10] ,
    \cb_6_1_io_dat_o[9] ,
    \cb_6_1_io_dat_o[8] ,
    \cb_6_1_io_dat_o[7] ,
    \cb_6_1_io_dat_o[6] ,
    \cb_6_1_io_dat_o[5] ,
    \cb_6_1_io_dat_o[4] ,
    \cb_6_1_io_dat_o[3] ,
    \cb_6_1_io_dat_o[2] ,
    \cb_6_1_io_dat_o[1] ,
    \cb_6_1_io_dat_o[0] }),
    .io_eo({\cb_6_1_io_eo[63] ,
    \cb_6_1_io_eo[62] ,
    \cb_6_1_io_eo[61] ,
    \cb_6_1_io_eo[60] ,
    \cb_6_1_io_eo[59] ,
    \cb_6_1_io_eo[58] ,
    \cb_6_1_io_eo[57] ,
    \cb_6_1_io_eo[56] ,
    \cb_6_1_io_eo[55] ,
    \cb_6_1_io_eo[54] ,
    \cb_6_1_io_eo[53] ,
    \cb_6_1_io_eo[52] ,
    \cb_6_1_io_eo[51] ,
    \cb_6_1_io_eo[50] ,
    \cb_6_1_io_eo[49] ,
    \cb_6_1_io_eo[48] ,
    \cb_6_1_io_eo[47] ,
    \cb_6_1_io_eo[46] ,
    \cb_6_1_io_eo[45] ,
    \cb_6_1_io_eo[44] ,
    \cb_6_1_io_eo[43] ,
    \cb_6_1_io_eo[42] ,
    \cb_6_1_io_eo[41] ,
    \cb_6_1_io_eo[40] ,
    \cb_6_1_io_eo[39] ,
    \cb_6_1_io_eo[38] ,
    \cb_6_1_io_eo[37] ,
    \cb_6_1_io_eo[36] ,
    \cb_6_1_io_eo[35] ,
    \cb_6_1_io_eo[34] ,
    \cb_6_1_io_eo[33] ,
    \cb_6_1_io_eo[32] ,
    \cb_6_1_io_eo[31] ,
    \cb_6_1_io_eo[30] ,
    \cb_6_1_io_eo[29] ,
    \cb_6_1_io_eo[28] ,
    \cb_6_1_io_eo[27] ,
    \cb_6_1_io_eo[26] ,
    \cb_6_1_io_eo[25] ,
    \cb_6_1_io_eo[24] ,
    \cb_6_1_io_eo[23] ,
    \cb_6_1_io_eo[22] ,
    \cb_6_1_io_eo[21] ,
    \cb_6_1_io_eo[20] ,
    \cb_6_1_io_eo[19] ,
    \cb_6_1_io_eo[18] ,
    \cb_6_1_io_eo[17] ,
    \cb_6_1_io_eo[16] ,
    \cb_6_1_io_eo[15] ,
    \cb_6_1_io_eo[14] ,
    \cb_6_1_io_eo[13] ,
    \cb_6_1_io_eo[12] ,
    \cb_6_1_io_eo[11] ,
    \cb_6_1_io_eo[10] ,
    \cb_6_1_io_eo[9] ,
    \cb_6_1_io_eo[8] ,
    \cb_6_1_io_eo[7] ,
    \cb_6_1_io_eo[6] ,
    \cb_6_1_io_eo[5] ,
    \cb_6_1_io_eo[4] ,
    \cb_6_1_io_eo[3] ,
    \cb_6_1_io_eo[2] ,
    \cb_6_1_io_eo[1] ,
    \cb_6_1_io_eo[0] }),
    .io_i_0_in1({\cb_6_0_io_o_0_out[7] ,
    \cb_6_0_io_o_0_out[6] ,
    \cb_6_0_io_o_0_out[5] ,
    \cb_6_0_io_o_0_out[4] ,
    \cb_6_0_io_o_0_out[3] ,
    \cb_6_0_io_o_0_out[2] ,
    \cb_6_0_io_o_0_out[1] ,
    \cb_6_0_io_o_0_out[0] }),
    .io_i_1_in1({\cb_6_0_io_o_1_out[7] ,
    \cb_6_0_io_o_1_out[6] ,
    \cb_6_0_io_o_1_out[5] ,
    \cb_6_0_io_o_1_out[4] ,
    \cb_6_0_io_o_1_out[3] ,
    \cb_6_0_io_o_1_out[2] ,
    \cb_6_0_io_o_1_out[1] ,
    \cb_6_0_io_o_1_out[0] }),
    .io_i_2_in1({\cb_6_0_io_o_2_out[7] ,
    \cb_6_0_io_o_2_out[6] ,
    \cb_6_0_io_o_2_out[5] ,
    \cb_6_0_io_o_2_out[4] ,
    \cb_6_0_io_o_2_out[3] ,
    \cb_6_0_io_o_2_out[2] ,
    \cb_6_0_io_o_2_out[1] ,
    \cb_6_0_io_o_2_out[0] }),
    .io_i_3_in1({\cb_6_0_io_o_3_out[7] ,
    \cb_6_0_io_o_3_out[6] ,
    \cb_6_0_io_o_3_out[5] ,
    \cb_6_0_io_o_3_out[4] ,
    \cb_6_0_io_o_3_out[3] ,
    \cb_6_0_io_o_3_out[2] ,
    \cb_6_0_io_o_3_out[1] ,
    \cb_6_0_io_o_3_out[0] }),
    .io_i_4_in1({\cb_6_0_io_o_4_out[7] ,
    \cb_6_0_io_o_4_out[6] ,
    \cb_6_0_io_o_4_out[5] ,
    \cb_6_0_io_o_4_out[4] ,
    \cb_6_0_io_o_4_out[3] ,
    \cb_6_0_io_o_4_out[2] ,
    \cb_6_0_io_o_4_out[1] ,
    \cb_6_0_io_o_4_out[0] }),
    .io_i_5_in1({\cb_6_0_io_o_5_out[7] ,
    \cb_6_0_io_o_5_out[6] ,
    \cb_6_0_io_o_5_out[5] ,
    \cb_6_0_io_o_5_out[4] ,
    \cb_6_0_io_o_5_out[3] ,
    \cb_6_0_io_o_5_out[2] ,
    \cb_6_0_io_o_5_out[1] ,
    \cb_6_0_io_o_5_out[0] }),
    .io_i_6_in1({\cb_6_0_io_o_6_out[7] ,
    \cb_6_0_io_o_6_out[6] ,
    \cb_6_0_io_o_6_out[5] ,
    \cb_6_0_io_o_6_out[4] ,
    \cb_6_0_io_o_6_out[3] ,
    \cb_6_0_io_o_6_out[2] ,
    \cb_6_0_io_o_6_out[1] ,
    \cb_6_0_io_o_6_out[0] }),
    .io_i_7_in1({\cb_6_0_io_o_7_out[7] ,
    \cb_6_0_io_o_7_out[6] ,
    \cb_6_0_io_o_7_out[5] ,
    \cb_6_0_io_o_7_out[4] ,
    \cb_6_0_io_o_7_out[3] ,
    \cb_6_0_io_o_7_out[2] ,
    \cb_6_0_io_o_7_out[1] ,
    \cb_6_0_io_o_7_out[0] }),
    .io_o_0_out({\cb_6_1_io_o_0_out[7] ,
    \cb_6_1_io_o_0_out[6] ,
    \cb_6_1_io_o_0_out[5] ,
    \cb_6_1_io_o_0_out[4] ,
    \cb_6_1_io_o_0_out[3] ,
    \cb_6_1_io_o_0_out[2] ,
    \cb_6_1_io_o_0_out[1] ,
    \cb_6_1_io_o_0_out[0] }),
    .io_o_1_out({\cb_6_1_io_o_1_out[7] ,
    \cb_6_1_io_o_1_out[6] ,
    \cb_6_1_io_o_1_out[5] ,
    \cb_6_1_io_o_1_out[4] ,
    \cb_6_1_io_o_1_out[3] ,
    \cb_6_1_io_o_1_out[2] ,
    \cb_6_1_io_o_1_out[1] ,
    \cb_6_1_io_o_1_out[0] }),
    .io_o_2_out({\cb_6_1_io_o_2_out[7] ,
    \cb_6_1_io_o_2_out[6] ,
    \cb_6_1_io_o_2_out[5] ,
    \cb_6_1_io_o_2_out[4] ,
    \cb_6_1_io_o_2_out[3] ,
    \cb_6_1_io_o_2_out[2] ,
    \cb_6_1_io_o_2_out[1] ,
    \cb_6_1_io_o_2_out[0] }),
    .io_o_3_out({\cb_6_1_io_o_3_out[7] ,
    \cb_6_1_io_o_3_out[6] ,
    \cb_6_1_io_o_3_out[5] ,
    \cb_6_1_io_o_3_out[4] ,
    \cb_6_1_io_o_3_out[3] ,
    \cb_6_1_io_o_3_out[2] ,
    \cb_6_1_io_o_3_out[1] ,
    \cb_6_1_io_o_3_out[0] }),
    .io_o_4_out({\cb_6_1_io_o_4_out[7] ,
    \cb_6_1_io_o_4_out[6] ,
    \cb_6_1_io_o_4_out[5] ,
    \cb_6_1_io_o_4_out[4] ,
    \cb_6_1_io_o_4_out[3] ,
    \cb_6_1_io_o_4_out[2] ,
    \cb_6_1_io_o_4_out[1] ,
    \cb_6_1_io_o_4_out[0] }),
    .io_o_5_out({\cb_6_1_io_o_5_out[7] ,
    \cb_6_1_io_o_5_out[6] ,
    \cb_6_1_io_o_5_out[5] ,
    \cb_6_1_io_o_5_out[4] ,
    \cb_6_1_io_o_5_out[3] ,
    \cb_6_1_io_o_5_out[2] ,
    \cb_6_1_io_o_5_out[1] ,
    \cb_6_1_io_o_5_out[0] }),
    .io_o_6_out({\cb_6_1_io_o_6_out[7] ,
    \cb_6_1_io_o_6_out[6] ,
    \cb_6_1_io_o_6_out[5] ,
    \cb_6_1_io_o_6_out[4] ,
    \cb_6_1_io_o_6_out[3] ,
    \cb_6_1_io_o_6_out[2] ,
    \cb_6_1_io_o_6_out[1] ,
    \cb_6_1_io_o_6_out[0] }),
    .io_o_7_out({\cb_6_1_io_o_7_out[7] ,
    \cb_6_1_io_o_7_out[6] ,
    \cb_6_1_io_o_7_out[5] ,
    \cb_6_1_io_o_7_out[4] ,
    \cb_6_1_io_o_7_out[3] ,
    \cb_6_1_io_o_7_out[2] ,
    \cb_6_1_io_o_7_out[1] ,
    \cb_6_1_io_o_7_out[0] }),
    .io_wo({\cb_6_0_io_eo[63] ,
    \cb_6_0_io_eo[62] ,
    \cb_6_0_io_eo[61] ,
    \cb_6_0_io_eo[60] ,
    \cb_6_0_io_eo[59] ,
    \cb_6_0_io_eo[58] ,
    \cb_6_0_io_eo[57] ,
    \cb_6_0_io_eo[56] ,
    \cb_6_0_io_eo[55] ,
    \cb_6_0_io_eo[54] ,
    \cb_6_0_io_eo[53] ,
    \cb_6_0_io_eo[52] ,
    \cb_6_0_io_eo[51] ,
    \cb_6_0_io_eo[50] ,
    \cb_6_0_io_eo[49] ,
    \cb_6_0_io_eo[48] ,
    \cb_6_0_io_eo[47] ,
    \cb_6_0_io_eo[46] ,
    \cb_6_0_io_eo[45] ,
    \cb_6_0_io_eo[44] ,
    \cb_6_0_io_eo[43] ,
    \cb_6_0_io_eo[42] ,
    \cb_6_0_io_eo[41] ,
    \cb_6_0_io_eo[40] ,
    \cb_6_0_io_eo[39] ,
    \cb_6_0_io_eo[38] ,
    \cb_6_0_io_eo[37] ,
    \cb_6_0_io_eo[36] ,
    \cb_6_0_io_eo[35] ,
    \cb_6_0_io_eo[34] ,
    \cb_6_0_io_eo[33] ,
    \cb_6_0_io_eo[32] ,
    \cb_6_0_io_eo[31] ,
    \cb_6_0_io_eo[30] ,
    \cb_6_0_io_eo[29] ,
    \cb_6_0_io_eo[28] ,
    \cb_6_0_io_eo[27] ,
    \cb_6_0_io_eo[26] ,
    \cb_6_0_io_eo[25] ,
    \cb_6_0_io_eo[24] ,
    \cb_6_0_io_eo[23] ,
    \cb_6_0_io_eo[22] ,
    \cb_6_0_io_eo[21] ,
    \cb_6_0_io_eo[20] ,
    \cb_6_0_io_eo[19] ,
    \cb_6_0_io_eo[18] ,
    \cb_6_0_io_eo[17] ,
    \cb_6_0_io_eo[16] ,
    \cb_6_0_io_eo[15] ,
    \cb_6_0_io_eo[14] ,
    \cb_6_0_io_eo[13] ,
    \cb_6_0_io_eo[12] ,
    \cb_6_0_io_eo[11] ,
    \cb_6_0_io_eo[10] ,
    \cb_6_0_io_eo[9] ,
    \cb_6_0_io_eo[8] ,
    \cb_6_0_io_eo[7] ,
    \cb_6_0_io_eo[6] ,
    \cb_6_0_io_eo[5] ,
    \cb_6_0_io_eo[4] ,
    \cb_6_0_io_eo[3] ,
    \cb_6_0_io_eo[2] ,
    \cb_6_0_io_eo[1] ,
    \cb_6_0_io_eo[0] }));
 cic_block cb_6_10 (.io_cs_i(cb_6_10_io_cs_i),
    .io_i_0_ci(cb_6_10_io_i_0_ci),
    .io_i_1_ci(cb_6_10_io_i_1_ci),
    .io_i_2_ci(cb_6_10_io_i_2_ci),
    .io_i_3_ci(cb_6_10_io_i_3_ci),
    .io_i_4_ci(cb_6_10_io_i_4_ci),
    .io_i_5_ci(cb_6_10_io_i_5_ci),
    .io_i_6_ci(cb_6_10_io_i_6_ci),
    .io_i_7_ci(cb_6_10_io_i_7_ci),
    .io_o_0_co(cb_6_10_io_o_0_co),
    .io_o_1_co(cb_6_10_io_o_1_co),
    .io_o_2_co(cb_6_10_io_o_2_co),
    .io_o_3_co(cb_6_10_io_o_3_co),
    .io_o_4_co(cb_6_10_io_o_4_co),
    .io_o_5_co(cb_6_10_io_o_5_co),
    .io_o_6_co(cb_6_10_io_o_6_co),
    .io_o_7_co(cb_6_10_io_o_7_co),
    .io_vci(cb_6_10_io_vci),
    .io_vco(cb_6_10_io_vco),
    .io_vi(cb_6_10_io_vi),
    .io_we_i(cb_6_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_6_0_io_adr_i[1] ,
    \cb_6_0_io_adr_i[0] }),
    .io_dat_i({\cb_6_0_io_dat_i[15] ,
    \cb_6_0_io_dat_i[14] ,
    \cb_6_0_io_dat_i[13] ,
    \cb_6_0_io_dat_i[12] ,
    \cb_6_0_io_dat_i[11] ,
    \cb_6_0_io_dat_i[10] ,
    \cb_6_0_io_dat_i[9] ,
    \cb_6_0_io_dat_i[8] ,
    \cb_6_0_io_dat_i[7] ,
    \cb_6_0_io_dat_i[6] ,
    \cb_6_0_io_dat_i[5] ,
    \cb_6_0_io_dat_i[4] ,
    \cb_6_0_io_dat_i[3] ,
    \cb_6_0_io_dat_i[2] ,
    \cb_6_0_io_dat_i[1] ,
    \cb_6_0_io_dat_i[0] }),
    .io_dat_o({\cb_6_10_io_dat_o[15] ,
    \cb_6_10_io_dat_o[14] ,
    \cb_6_10_io_dat_o[13] ,
    \cb_6_10_io_dat_o[12] ,
    \cb_6_10_io_dat_o[11] ,
    \cb_6_10_io_dat_o[10] ,
    \cb_6_10_io_dat_o[9] ,
    \cb_6_10_io_dat_o[8] ,
    \cb_6_10_io_dat_o[7] ,
    \cb_6_10_io_dat_o[6] ,
    \cb_6_10_io_dat_o[5] ,
    \cb_6_10_io_dat_o[4] ,
    \cb_6_10_io_dat_o[3] ,
    \cb_6_10_io_dat_o[2] ,
    \cb_6_10_io_dat_o[1] ,
    \cb_6_10_io_dat_o[0] }),
    .io_eo({\_T_142[31] ,
    \_T_142[30] ,
    \_T_142[29] ,
    \_T_142[28] ,
    \_T_142[27] ,
    \_T_142[26] ,
    \_T_142[25] ,
    \_T_142[24] ,
    \_T_142[23] ,
    \_T_142[22] ,
    \_T_142[21] ,
    \_T_142[20] ,
    \_T_142[19] ,
    \_T_142[18] ,
    \_T_142[17] ,
    \_T_142[16] ,
    \_T_142[15] ,
    \_T_142[14] ,
    \_T_142[13] ,
    \_T_142[12] ,
    \_T_142[11] ,
    \_T_142[10] ,
    \_T_142[9] ,
    \_T_142[8] ,
    \_T_142[7] ,
    \_T_142[6] ,
    \_T_142[5] ,
    \_T_142[4] ,
    \_T_142[3] ,
    \_T_142[2] ,
    \_T_142[1] ,
    \_T_142[0] ,
    \_T_139[31] ,
    \_T_139[30] ,
    \_T_139[29] ,
    \_T_139[28] ,
    \_T_139[27] ,
    \_T_139[26] ,
    \_T_139[25] ,
    \_T_139[24] ,
    \_T_139[23] ,
    \_T_139[22] ,
    \_T_139[21] ,
    \_T_139[20] ,
    \_T_139[19] ,
    \_T_139[18] ,
    \_T_139[17] ,
    \_T_139[16] ,
    \_T_139[15] ,
    \_T_139[14] ,
    \_T_139[13] ,
    \_T_139[12] ,
    \_T_139[11] ,
    \_T_139[10] ,
    \_T_139[9] ,
    \_T_139[8] ,
    \_T_139[7] ,
    \_T_139[6] ,
    \_T_139[5] ,
    \_T_139[4] ,
    \_T_139[3] ,
    \_T_139[2] ,
    \_T_139[1] ,
    \_T_139[0] }),
    .io_i_0_in1({\cb_6_10_io_i_0_in1[7] ,
    \cb_6_10_io_i_0_in1[6] ,
    \cb_6_10_io_i_0_in1[5] ,
    \cb_6_10_io_i_0_in1[4] ,
    \cb_6_10_io_i_0_in1[3] ,
    \cb_6_10_io_i_0_in1[2] ,
    \cb_6_10_io_i_0_in1[1] ,
    \cb_6_10_io_i_0_in1[0] }),
    .io_i_1_in1({\cb_6_10_io_i_1_in1[7] ,
    \cb_6_10_io_i_1_in1[6] ,
    \cb_6_10_io_i_1_in1[5] ,
    \cb_6_10_io_i_1_in1[4] ,
    \cb_6_10_io_i_1_in1[3] ,
    \cb_6_10_io_i_1_in1[2] ,
    \cb_6_10_io_i_1_in1[1] ,
    \cb_6_10_io_i_1_in1[0] }),
    .io_i_2_in1({\cb_6_10_io_i_2_in1[7] ,
    \cb_6_10_io_i_2_in1[6] ,
    \cb_6_10_io_i_2_in1[5] ,
    \cb_6_10_io_i_2_in1[4] ,
    \cb_6_10_io_i_2_in1[3] ,
    \cb_6_10_io_i_2_in1[2] ,
    \cb_6_10_io_i_2_in1[1] ,
    \cb_6_10_io_i_2_in1[0] }),
    .io_i_3_in1({\cb_6_10_io_i_3_in1[7] ,
    \cb_6_10_io_i_3_in1[6] ,
    \cb_6_10_io_i_3_in1[5] ,
    \cb_6_10_io_i_3_in1[4] ,
    \cb_6_10_io_i_3_in1[3] ,
    \cb_6_10_io_i_3_in1[2] ,
    \cb_6_10_io_i_3_in1[1] ,
    \cb_6_10_io_i_3_in1[0] }),
    .io_i_4_in1({\cb_6_10_io_i_4_in1[7] ,
    \cb_6_10_io_i_4_in1[6] ,
    \cb_6_10_io_i_4_in1[5] ,
    \cb_6_10_io_i_4_in1[4] ,
    \cb_6_10_io_i_4_in1[3] ,
    \cb_6_10_io_i_4_in1[2] ,
    \cb_6_10_io_i_4_in1[1] ,
    \cb_6_10_io_i_4_in1[0] }),
    .io_i_5_in1({\cb_6_10_io_i_5_in1[7] ,
    \cb_6_10_io_i_5_in1[6] ,
    \cb_6_10_io_i_5_in1[5] ,
    \cb_6_10_io_i_5_in1[4] ,
    \cb_6_10_io_i_5_in1[3] ,
    \cb_6_10_io_i_5_in1[2] ,
    \cb_6_10_io_i_5_in1[1] ,
    \cb_6_10_io_i_5_in1[0] }),
    .io_i_6_in1({\cb_6_10_io_i_6_in1[7] ,
    \cb_6_10_io_i_6_in1[6] ,
    \cb_6_10_io_i_6_in1[5] ,
    \cb_6_10_io_i_6_in1[4] ,
    \cb_6_10_io_i_6_in1[3] ,
    \cb_6_10_io_i_6_in1[2] ,
    \cb_6_10_io_i_6_in1[1] ,
    \cb_6_10_io_i_6_in1[0] }),
    .io_i_7_in1({\cb_6_10_io_i_7_in1[7] ,
    \cb_6_10_io_i_7_in1[6] ,
    \cb_6_10_io_i_7_in1[5] ,
    \cb_6_10_io_i_7_in1[4] ,
    \cb_6_10_io_i_7_in1[3] ,
    \cb_6_10_io_i_7_in1[2] ,
    \cb_6_10_io_i_7_in1[1] ,
    \cb_6_10_io_i_7_in1[0] }),
    .io_o_0_out({\_T_139[7] ,
    \_T_139[6] ,
    \_T_139[5] ,
    \_T_139[4] ,
    \_T_139[3] ,
    \_T_139[2] ,
    \_T_139[1] ,
    \_T_139[0] }),
    .io_o_1_out({\_T_139[15] ,
    \_T_139[14] ,
    \_T_139[13] ,
    \_T_139[12] ,
    \_T_139[11] ,
    \_T_139[10] ,
    \_T_139[9] ,
    \_T_139[8] }),
    .io_o_2_out({\_T_139[23] ,
    \_T_139[22] ,
    \_T_139[21] ,
    \_T_139[20] ,
    \_T_139[19] ,
    \_T_139[18] ,
    \_T_139[17] ,
    \_T_139[16] }),
    .io_o_3_out({\_T_139[31] ,
    \_T_139[30] ,
    \_T_139[29] ,
    \_T_139[28] ,
    \_T_139[27] ,
    \_T_139[26] ,
    \_T_139[25] ,
    \_T_139[24] }),
    .io_o_4_out({\_T_142[7] ,
    \_T_142[6] ,
    \_T_142[5] ,
    \_T_142[4] ,
    \_T_142[3] ,
    \_T_142[2] ,
    \_T_142[1] ,
    \_T_142[0] }),
    .io_o_5_out({\_T_142[15] ,
    \_T_142[14] ,
    \_T_142[13] ,
    \_T_142[12] ,
    \_T_142[11] ,
    \_T_142[10] ,
    \_T_142[9] ,
    \_T_142[8] }),
    .io_o_6_out({\_T_142[23] ,
    \_T_142[22] ,
    \_T_142[21] ,
    \_T_142[20] ,
    \_T_142[19] ,
    \_T_142[18] ,
    \_T_142[17] ,
    \_T_142[16] }),
    .io_o_7_out({\_T_142[31] ,
    \_T_142[30] ,
    \_T_142[29] ,
    \_T_142[28] ,
    \_T_142[27] ,
    \_T_142[26] ,
    \_T_142[25] ,
    \_T_142[24] }),
    .io_wo({\cb_6_10_io_wo[63] ,
    \cb_6_10_io_wo[62] ,
    \cb_6_10_io_wo[61] ,
    \cb_6_10_io_wo[60] ,
    \cb_6_10_io_wo[59] ,
    \cb_6_10_io_wo[58] ,
    \cb_6_10_io_wo[57] ,
    \cb_6_10_io_wo[56] ,
    \cb_6_10_io_wo[55] ,
    \cb_6_10_io_wo[54] ,
    \cb_6_10_io_wo[53] ,
    \cb_6_10_io_wo[52] ,
    \cb_6_10_io_wo[51] ,
    \cb_6_10_io_wo[50] ,
    \cb_6_10_io_wo[49] ,
    \cb_6_10_io_wo[48] ,
    \cb_6_10_io_wo[47] ,
    \cb_6_10_io_wo[46] ,
    \cb_6_10_io_wo[45] ,
    \cb_6_10_io_wo[44] ,
    \cb_6_10_io_wo[43] ,
    \cb_6_10_io_wo[42] ,
    \cb_6_10_io_wo[41] ,
    \cb_6_10_io_wo[40] ,
    \cb_6_10_io_wo[39] ,
    \cb_6_10_io_wo[38] ,
    \cb_6_10_io_wo[37] ,
    \cb_6_10_io_wo[36] ,
    \cb_6_10_io_wo[35] ,
    \cb_6_10_io_wo[34] ,
    \cb_6_10_io_wo[33] ,
    \cb_6_10_io_wo[32] ,
    \cb_6_10_io_wo[31] ,
    \cb_6_10_io_wo[30] ,
    \cb_6_10_io_wo[29] ,
    \cb_6_10_io_wo[28] ,
    \cb_6_10_io_wo[27] ,
    \cb_6_10_io_wo[26] ,
    \cb_6_10_io_wo[25] ,
    \cb_6_10_io_wo[24] ,
    \cb_6_10_io_wo[23] ,
    \cb_6_10_io_wo[22] ,
    \cb_6_10_io_wo[21] ,
    \cb_6_10_io_wo[20] ,
    \cb_6_10_io_wo[19] ,
    \cb_6_10_io_wo[18] ,
    \cb_6_10_io_wo[17] ,
    \cb_6_10_io_wo[16] ,
    \cb_6_10_io_wo[15] ,
    \cb_6_10_io_wo[14] ,
    \cb_6_10_io_wo[13] ,
    \cb_6_10_io_wo[12] ,
    \cb_6_10_io_wo[11] ,
    \cb_6_10_io_wo[10] ,
    \cb_6_10_io_wo[9] ,
    \cb_6_10_io_wo[8] ,
    \cb_6_10_io_wo[7] ,
    \cb_6_10_io_wo[6] ,
    \cb_6_10_io_wo[5] ,
    \cb_6_10_io_wo[4] ,
    \cb_6_10_io_wo[3] ,
    \cb_6_10_io_wo[2] ,
    \cb_6_10_io_wo[1] ,
    \cb_6_10_io_wo[0] }));
 cic_block cb_6_2 (.io_cs_i(cb_6_2_io_cs_i),
    .io_i_0_ci(cb_6_1_io_o_0_co),
    .io_i_1_ci(cb_6_1_io_o_1_co),
    .io_i_2_ci(cb_6_1_io_o_2_co),
    .io_i_3_ci(cb_6_1_io_o_3_co),
    .io_i_4_ci(cb_6_1_io_o_4_co),
    .io_i_5_ci(cb_6_1_io_o_5_co),
    .io_i_6_ci(cb_6_1_io_o_6_co),
    .io_i_7_ci(cb_6_1_io_o_7_co),
    .io_o_0_co(cb_6_2_io_o_0_co),
    .io_o_1_co(cb_6_2_io_o_1_co),
    .io_o_2_co(cb_6_2_io_o_2_co),
    .io_o_3_co(cb_6_2_io_o_3_co),
    .io_o_4_co(cb_6_2_io_o_4_co),
    .io_o_5_co(cb_6_2_io_o_5_co),
    .io_o_6_co(cb_6_2_io_o_6_co),
    .io_o_7_co(cb_6_2_io_o_7_co),
    .io_vci(cb_6_1_io_vco),
    .io_vco(cb_6_2_io_vco),
    .io_vi(cb_6_2_io_vi),
    .io_we_i(cb_6_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_6_0_io_adr_i[1] ,
    \cb_6_0_io_adr_i[0] }),
    .io_dat_i({\cb_6_0_io_dat_i[15] ,
    \cb_6_0_io_dat_i[14] ,
    \cb_6_0_io_dat_i[13] ,
    \cb_6_0_io_dat_i[12] ,
    \cb_6_0_io_dat_i[11] ,
    \cb_6_0_io_dat_i[10] ,
    \cb_6_0_io_dat_i[9] ,
    \cb_6_0_io_dat_i[8] ,
    \cb_6_0_io_dat_i[7] ,
    \cb_6_0_io_dat_i[6] ,
    \cb_6_0_io_dat_i[5] ,
    \cb_6_0_io_dat_i[4] ,
    \cb_6_0_io_dat_i[3] ,
    \cb_6_0_io_dat_i[2] ,
    \cb_6_0_io_dat_i[1] ,
    \cb_6_0_io_dat_i[0] }),
    .io_dat_o({\cb_6_2_io_dat_o[15] ,
    \cb_6_2_io_dat_o[14] ,
    \cb_6_2_io_dat_o[13] ,
    \cb_6_2_io_dat_o[12] ,
    \cb_6_2_io_dat_o[11] ,
    \cb_6_2_io_dat_o[10] ,
    \cb_6_2_io_dat_o[9] ,
    \cb_6_2_io_dat_o[8] ,
    \cb_6_2_io_dat_o[7] ,
    \cb_6_2_io_dat_o[6] ,
    \cb_6_2_io_dat_o[5] ,
    \cb_6_2_io_dat_o[4] ,
    \cb_6_2_io_dat_o[3] ,
    \cb_6_2_io_dat_o[2] ,
    \cb_6_2_io_dat_o[1] ,
    \cb_6_2_io_dat_o[0] }),
    .io_eo({\cb_6_2_io_eo[63] ,
    \cb_6_2_io_eo[62] ,
    \cb_6_2_io_eo[61] ,
    \cb_6_2_io_eo[60] ,
    \cb_6_2_io_eo[59] ,
    \cb_6_2_io_eo[58] ,
    \cb_6_2_io_eo[57] ,
    \cb_6_2_io_eo[56] ,
    \cb_6_2_io_eo[55] ,
    \cb_6_2_io_eo[54] ,
    \cb_6_2_io_eo[53] ,
    \cb_6_2_io_eo[52] ,
    \cb_6_2_io_eo[51] ,
    \cb_6_2_io_eo[50] ,
    \cb_6_2_io_eo[49] ,
    \cb_6_2_io_eo[48] ,
    \cb_6_2_io_eo[47] ,
    \cb_6_2_io_eo[46] ,
    \cb_6_2_io_eo[45] ,
    \cb_6_2_io_eo[44] ,
    \cb_6_2_io_eo[43] ,
    \cb_6_2_io_eo[42] ,
    \cb_6_2_io_eo[41] ,
    \cb_6_2_io_eo[40] ,
    \cb_6_2_io_eo[39] ,
    \cb_6_2_io_eo[38] ,
    \cb_6_2_io_eo[37] ,
    \cb_6_2_io_eo[36] ,
    \cb_6_2_io_eo[35] ,
    \cb_6_2_io_eo[34] ,
    \cb_6_2_io_eo[33] ,
    \cb_6_2_io_eo[32] ,
    \cb_6_2_io_eo[31] ,
    \cb_6_2_io_eo[30] ,
    \cb_6_2_io_eo[29] ,
    \cb_6_2_io_eo[28] ,
    \cb_6_2_io_eo[27] ,
    \cb_6_2_io_eo[26] ,
    \cb_6_2_io_eo[25] ,
    \cb_6_2_io_eo[24] ,
    \cb_6_2_io_eo[23] ,
    \cb_6_2_io_eo[22] ,
    \cb_6_2_io_eo[21] ,
    \cb_6_2_io_eo[20] ,
    \cb_6_2_io_eo[19] ,
    \cb_6_2_io_eo[18] ,
    \cb_6_2_io_eo[17] ,
    \cb_6_2_io_eo[16] ,
    \cb_6_2_io_eo[15] ,
    \cb_6_2_io_eo[14] ,
    \cb_6_2_io_eo[13] ,
    \cb_6_2_io_eo[12] ,
    \cb_6_2_io_eo[11] ,
    \cb_6_2_io_eo[10] ,
    \cb_6_2_io_eo[9] ,
    \cb_6_2_io_eo[8] ,
    \cb_6_2_io_eo[7] ,
    \cb_6_2_io_eo[6] ,
    \cb_6_2_io_eo[5] ,
    \cb_6_2_io_eo[4] ,
    \cb_6_2_io_eo[3] ,
    \cb_6_2_io_eo[2] ,
    \cb_6_2_io_eo[1] ,
    \cb_6_2_io_eo[0] }),
    .io_i_0_in1({\cb_6_1_io_o_0_out[7] ,
    \cb_6_1_io_o_0_out[6] ,
    \cb_6_1_io_o_0_out[5] ,
    \cb_6_1_io_o_0_out[4] ,
    \cb_6_1_io_o_0_out[3] ,
    \cb_6_1_io_o_0_out[2] ,
    \cb_6_1_io_o_0_out[1] ,
    \cb_6_1_io_o_0_out[0] }),
    .io_i_1_in1({\cb_6_1_io_o_1_out[7] ,
    \cb_6_1_io_o_1_out[6] ,
    \cb_6_1_io_o_1_out[5] ,
    \cb_6_1_io_o_1_out[4] ,
    \cb_6_1_io_o_1_out[3] ,
    \cb_6_1_io_o_1_out[2] ,
    \cb_6_1_io_o_1_out[1] ,
    \cb_6_1_io_o_1_out[0] }),
    .io_i_2_in1({\cb_6_1_io_o_2_out[7] ,
    \cb_6_1_io_o_2_out[6] ,
    \cb_6_1_io_o_2_out[5] ,
    \cb_6_1_io_o_2_out[4] ,
    \cb_6_1_io_o_2_out[3] ,
    \cb_6_1_io_o_2_out[2] ,
    \cb_6_1_io_o_2_out[1] ,
    \cb_6_1_io_o_2_out[0] }),
    .io_i_3_in1({\cb_6_1_io_o_3_out[7] ,
    \cb_6_1_io_o_3_out[6] ,
    \cb_6_1_io_o_3_out[5] ,
    \cb_6_1_io_o_3_out[4] ,
    \cb_6_1_io_o_3_out[3] ,
    \cb_6_1_io_o_3_out[2] ,
    \cb_6_1_io_o_3_out[1] ,
    \cb_6_1_io_o_3_out[0] }),
    .io_i_4_in1({\cb_6_1_io_o_4_out[7] ,
    \cb_6_1_io_o_4_out[6] ,
    \cb_6_1_io_o_4_out[5] ,
    \cb_6_1_io_o_4_out[4] ,
    \cb_6_1_io_o_4_out[3] ,
    \cb_6_1_io_o_4_out[2] ,
    \cb_6_1_io_o_4_out[1] ,
    \cb_6_1_io_o_4_out[0] }),
    .io_i_5_in1({\cb_6_1_io_o_5_out[7] ,
    \cb_6_1_io_o_5_out[6] ,
    \cb_6_1_io_o_5_out[5] ,
    \cb_6_1_io_o_5_out[4] ,
    \cb_6_1_io_o_5_out[3] ,
    \cb_6_1_io_o_5_out[2] ,
    \cb_6_1_io_o_5_out[1] ,
    \cb_6_1_io_o_5_out[0] }),
    .io_i_6_in1({\cb_6_1_io_o_6_out[7] ,
    \cb_6_1_io_o_6_out[6] ,
    \cb_6_1_io_o_6_out[5] ,
    \cb_6_1_io_o_6_out[4] ,
    \cb_6_1_io_o_6_out[3] ,
    \cb_6_1_io_o_6_out[2] ,
    \cb_6_1_io_o_6_out[1] ,
    \cb_6_1_io_o_6_out[0] }),
    .io_i_7_in1({\cb_6_1_io_o_7_out[7] ,
    \cb_6_1_io_o_7_out[6] ,
    \cb_6_1_io_o_7_out[5] ,
    \cb_6_1_io_o_7_out[4] ,
    \cb_6_1_io_o_7_out[3] ,
    \cb_6_1_io_o_7_out[2] ,
    \cb_6_1_io_o_7_out[1] ,
    \cb_6_1_io_o_7_out[0] }),
    .io_o_0_out({\cb_6_2_io_o_0_out[7] ,
    \cb_6_2_io_o_0_out[6] ,
    \cb_6_2_io_o_0_out[5] ,
    \cb_6_2_io_o_0_out[4] ,
    \cb_6_2_io_o_0_out[3] ,
    \cb_6_2_io_o_0_out[2] ,
    \cb_6_2_io_o_0_out[1] ,
    \cb_6_2_io_o_0_out[0] }),
    .io_o_1_out({\cb_6_2_io_o_1_out[7] ,
    \cb_6_2_io_o_1_out[6] ,
    \cb_6_2_io_o_1_out[5] ,
    \cb_6_2_io_o_1_out[4] ,
    \cb_6_2_io_o_1_out[3] ,
    \cb_6_2_io_o_1_out[2] ,
    \cb_6_2_io_o_1_out[1] ,
    \cb_6_2_io_o_1_out[0] }),
    .io_o_2_out({\cb_6_2_io_o_2_out[7] ,
    \cb_6_2_io_o_2_out[6] ,
    \cb_6_2_io_o_2_out[5] ,
    \cb_6_2_io_o_2_out[4] ,
    \cb_6_2_io_o_2_out[3] ,
    \cb_6_2_io_o_2_out[2] ,
    \cb_6_2_io_o_2_out[1] ,
    \cb_6_2_io_o_2_out[0] }),
    .io_o_3_out({\cb_6_2_io_o_3_out[7] ,
    \cb_6_2_io_o_3_out[6] ,
    \cb_6_2_io_o_3_out[5] ,
    \cb_6_2_io_o_3_out[4] ,
    \cb_6_2_io_o_3_out[3] ,
    \cb_6_2_io_o_3_out[2] ,
    \cb_6_2_io_o_3_out[1] ,
    \cb_6_2_io_o_3_out[0] }),
    .io_o_4_out({\cb_6_2_io_o_4_out[7] ,
    \cb_6_2_io_o_4_out[6] ,
    \cb_6_2_io_o_4_out[5] ,
    \cb_6_2_io_o_4_out[4] ,
    \cb_6_2_io_o_4_out[3] ,
    \cb_6_2_io_o_4_out[2] ,
    \cb_6_2_io_o_4_out[1] ,
    \cb_6_2_io_o_4_out[0] }),
    .io_o_5_out({\cb_6_2_io_o_5_out[7] ,
    \cb_6_2_io_o_5_out[6] ,
    \cb_6_2_io_o_5_out[5] ,
    \cb_6_2_io_o_5_out[4] ,
    \cb_6_2_io_o_5_out[3] ,
    \cb_6_2_io_o_5_out[2] ,
    \cb_6_2_io_o_5_out[1] ,
    \cb_6_2_io_o_5_out[0] }),
    .io_o_6_out({\cb_6_2_io_o_6_out[7] ,
    \cb_6_2_io_o_6_out[6] ,
    \cb_6_2_io_o_6_out[5] ,
    \cb_6_2_io_o_6_out[4] ,
    \cb_6_2_io_o_6_out[3] ,
    \cb_6_2_io_o_6_out[2] ,
    \cb_6_2_io_o_6_out[1] ,
    \cb_6_2_io_o_6_out[0] }),
    .io_o_7_out({\cb_6_2_io_o_7_out[7] ,
    \cb_6_2_io_o_7_out[6] ,
    \cb_6_2_io_o_7_out[5] ,
    \cb_6_2_io_o_7_out[4] ,
    \cb_6_2_io_o_7_out[3] ,
    \cb_6_2_io_o_7_out[2] ,
    \cb_6_2_io_o_7_out[1] ,
    \cb_6_2_io_o_7_out[0] }),
    .io_wo({\cb_6_1_io_eo[63] ,
    \cb_6_1_io_eo[62] ,
    \cb_6_1_io_eo[61] ,
    \cb_6_1_io_eo[60] ,
    \cb_6_1_io_eo[59] ,
    \cb_6_1_io_eo[58] ,
    \cb_6_1_io_eo[57] ,
    \cb_6_1_io_eo[56] ,
    \cb_6_1_io_eo[55] ,
    \cb_6_1_io_eo[54] ,
    \cb_6_1_io_eo[53] ,
    \cb_6_1_io_eo[52] ,
    \cb_6_1_io_eo[51] ,
    \cb_6_1_io_eo[50] ,
    \cb_6_1_io_eo[49] ,
    \cb_6_1_io_eo[48] ,
    \cb_6_1_io_eo[47] ,
    \cb_6_1_io_eo[46] ,
    \cb_6_1_io_eo[45] ,
    \cb_6_1_io_eo[44] ,
    \cb_6_1_io_eo[43] ,
    \cb_6_1_io_eo[42] ,
    \cb_6_1_io_eo[41] ,
    \cb_6_1_io_eo[40] ,
    \cb_6_1_io_eo[39] ,
    \cb_6_1_io_eo[38] ,
    \cb_6_1_io_eo[37] ,
    \cb_6_1_io_eo[36] ,
    \cb_6_1_io_eo[35] ,
    \cb_6_1_io_eo[34] ,
    \cb_6_1_io_eo[33] ,
    \cb_6_1_io_eo[32] ,
    \cb_6_1_io_eo[31] ,
    \cb_6_1_io_eo[30] ,
    \cb_6_1_io_eo[29] ,
    \cb_6_1_io_eo[28] ,
    \cb_6_1_io_eo[27] ,
    \cb_6_1_io_eo[26] ,
    \cb_6_1_io_eo[25] ,
    \cb_6_1_io_eo[24] ,
    \cb_6_1_io_eo[23] ,
    \cb_6_1_io_eo[22] ,
    \cb_6_1_io_eo[21] ,
    \cb_6_1_io_eo[20] ,
    \cb_6_1_io_eo[19] ,
    \cb_6_1_io_eo[18] ,
    \cb_6_1_io_eo[17] ,
    \cb_6_1_io_eo[16] ,
    \cb_6_1_io_eo[15] ,
    \cb_6_1_io_eo[14] ,
    \cb_6_1_io_eo[13] ,
    \cb_6_1_io_eo[12] ,
    \cb_6_1_io_eo[11] ,
    \cb_6_1_io_eo[10] ,
    \cb_6_1_io_eo[9] ,
    \cb_6_1_io_eo[8] ,
    \cb_6_1_io_eo[7] ,
    \cb_6_1_io_eo[6] ,
    \cb_6_1_io_eo[5] ,
    \cb_6_1_io_eo[4] ,
    \cb_6_1_io_eo[3] ,
    \cb_6_1_io_eo[2] ,
    \cb_6_1_io_eo[1] ,
    \cb_6_1_io_eo[0] }));
 cic_block cb_6_3 (.io_cs_i(cb_6_3_io_cs_i),
    .io_i_0_ci(cb_6_2_io_o_0_co),
    .io_i_1_ci(cb_6_2_io_o_1_co),
    .io_i_2_ci(cb_6_2_io_o_2_co),
    .io_i_3_ci(cb_6_2_io_o_3_co),
    .io_i_4_ci(cb_6_2_io_o_4_co),
    .io_i_5_ci(cb_6_2_io_o_5_co),
    .io_i_6_ci(cb_6_2_io_o_6_co),
    .io_i_7_ci(cb_6_2_io_o_7_co),
    .io_o_0_co(cb_6_3_io_o_0_co),
    .io_o_1_co(cb_6_3_io_o_1_co),
    .io_o_2_co(cb_6_3_io_o_2_co),
    .io_o_3_co(cb_6_3_io_o_3_co),
    .io_o_4_co(cb_6_3_io_o_4_co),
    .io_o_5_co(cb_6_3_io_o_5_co),
    .io_o_6_co(cb_6_3_io_o_6_co),
    .io_o_7_co(cb_6_3_io_o_7_co),
    .io_vci(cb_6_2_io_vco),
    .io_vco(cb_6_3_io_vco),
    .io_vi(cb_6_3_io_vi),
    .io_we_i(cb_6_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_6_0_io_adr_i[1] ,
    \cb_6_0_io_adr_i[0] }),
    .io_dat_i({\cb_6_0_io_dat_i[15] ,
    \cb_6_0_io_dat_i[14] ,
    \cb_6_0_io_dat_i[13] ,
    \cb_6_0_io_dat_i[12] ,
    \cb_6_0_io_dat_i[11] ,
    \cb_6_0_io_dat_i[10] ,
    \cb_6_0_io_dat_i[9] ,
    \cb_6_0_io_dat_i[8] ,
    \cb_6_0_io_dat_i[7] ,
    \cb_6_0_io_dat_i[6] ,
    \cb_6_0_io_dat_i[5] ,
    \cb_6_0_io_dat_i[4] ,
    \cb_6_0_io_dat_i[3] ,
    \cb_6_0_io_dat_i[2] ,
    \cb_6_0_io_dat_i[1] ,
    \cb_6_0_io_dat_i[0] }),
    .io_dat_o({\cb_6_3_io_dat_o[15] ,
    \cb_6_3_io_dat_o[14] ,
    \cb_6_3_io_dat_o[13] ,
    \cb_6_3_io_dat_o[12] ,
    \cb_6_3_io_dat_o[11] ,
    \cb_6_3_io_dat_o[10] ,
    \cb_6_3_io_dat_o[9] ,
    \cb_6_3_io_dat_o[8] ,
    \cb_6_3_io_dat_o[7] ,
    \cb_6_3_io_dat_o[6] ,
    \cb_6_3_io_dat_o[5] ,
    \cb_6_3_io_dat_o[4] ,
    \cb_6_3_io_dat_o[3] ,
    \cb_6_3_io_dat_o[2] ,
    \cb_6_3_io_dat_o[1] ,
    \cb_6_3_io_dat_o[0] }),
    .io_eo({\cb_6_3_io_eo[63] ,
    \cb_6_3_io_eo[62] ,
    \cb_6_3_io_eo[61] ,
    \cb_6_3_io_eo[60] ,
    \cb_6_3_io_eo[59] ,
    \cb_6_3_io_eo[58] ,
    \cb_6_3_io_eo[57] ,
    \cb_6_3_io_eo[56] ,
    \cb_6_3_io_eo[55] ,
    \cb_6_3_io_eo[54] ,
    \cb_6_3_io_eo[53] ,
    \cb_6_3_io_eo[52] ,
    \cb_6_3_io_eo[51] ,
    \cb_6_3_io_eo[50] ,
    \cb_6_3_io_eo[49] ,
    \cb_6_3_io_eo[48] ,
    \cb_6_3_io_eo[47] ,
    \cb_6_3_io_eo[46] ,
    \cb_6_3_io_eo[45] ,
    \cb_6_3_io_eo[44] ,
    \cb_6_3_io_eo[43] ,
    \cb_6_3_io_eo[42] ,
    \cb_6_3_io_eo[41] ,
    \cb_6_3_io_eo[40] ,
    \cb_6_3_io_eo[39] ,
    \cb_6_3_io_eo[38] ,
    \cb_6_3_io_eo[37] ,
    \cb_6_3_io_eo[36] ,
    \cb_6_3_io_eo[35] ,
    \cb_6_3_io_eo[34] ,
    \cb_6_3_io_eo[33] ,
    \cb_6_3_io_eo[32] ,
    \cb_6_3_io_eo[31] ,
    \cb_6_3_io_eo[30] ,
    \cb_6_3_io_eo[29] ,
    \cb_6_3_io_eo[28] ,
    \cb_6_3_io_eo[27] ,
    \cb_6_3_io_eo[26] ,
    \cb_6_3_io_eo[25] ,
    \cb_6_3_io_eo[24] ,
    \cb_6_3_io_eo[23] ,
    \cb_6_3_io_eo[22] ,
    \cb_6_3_io_eo[21] ,
    \cb_6_3_io_eo[20] ,
    \cb_6_3_io_eo[19] ,
    \cb_6_3_io_eo[18] ,
    \cb_6_3_io_eo[17] ,
    \cb_6_3_io_eo[16] ,
    \cb_6_3_io_eo[15] ,
    \cb_6_3_io_eo[14] ,
    \cb_6_3_io_eo[13] ,
    \cb_6_3_io_eo[12] ,
    \cb_6_3_io_eo[11] ,
    \cb_6_3_io_eo[10] ,
    \cb_6_3_io_eo[9] ,
    \cb_6_3_io_eo[8] ,
    \cb_6_3_io_eo[7] ,
    \cb_6_3_io_eo[6] ,
    \cb_6_3_io_eo[5] ,
    \cb_6_3_io_eo[4] ,
    \cb_6_3_io_eo[3] ,
    \cb_6_3_io_eo[2] ,
    \cb_6_3_io_eo[1] ,
    \cb_6_3_io_eo[0] }),
    .io_i_0_in1({\cb_6_2_io_o_0_out[7] ,
    \cb_6_2_io_o_0_out[6] ,
    \cb_6_2_io_o_0_out[5] ,
    \cb_6_2_io_o_0_out[4] ,
    \cb_6_2_io_o_0_out[3] ,
    \cb_6_2_io_o_0_out[2] ,
    \cb_6_2_io_o_0_out[1] ,
    \cb_6_2_io_o_0_out[0] }),
    .io_i_1_in1({\cb_6_2_io_o_1_out[7] ,
    \cb_6_2_io_o_1_out[6] ,
    \cb_6_2_io_o_1_out[5] ,
    \cb_6_2_io_o_1_out[4] ,
    \cb_6_2_io_o_1_out[3] ,
    \cb_6_2_io_o_1_out[2] ,
    \cb_6_2_io_o_1_out[1] ,
    \cb_6_2_io_o_1_out[0] }),
    .io_i_2_in1({\cb_6_2_io_o_2_out[7] ,
    \cb_6_2_io_o_2_out[6] ,
    \cb_6_2_io_o_2_out[5] ,
    \cb_6_2_io_o_2_out[4] ,
    \cb_6_2_io_o_2_out[3] ,
    \cb_6_2_io_o_2_out[2] ,
    \cb_6_2_io_o_2_out[1] ,
    \cb_6_2_io_o_2_out[0] }),
    .io_i_3_in1({\cb_6_2_io_o_3_out[7] ,
    \cb_6_2_io_o_3_out[6] ,
    \cb_6_2_io_o_3_out[5] ,
    \cb_6_2_io_o_3_out[4] ,
    \cb_6_2_io_o_3_out[3] ,
    \cb_6_2_io_o_3_out[2] ,
    \cb_6_2_io_o_3_out[1] ,
    \cb_6_2_io_o_3_out[0] }),
    .io_i_4_in1({\cb_6_2_io_o_4_out[7] ,
    \cb_6_2_io_o_4_out[6] ,
    \cb_6_2_io_o_4_out[5] ,
    \cb_6_2_io_o_4_out[4] ,
    \cb_6_2_io_o_4_out[3] ,
    \cb_6_2_io_o_4_out[2] ,
    \cb_6_2_io_o_4_out[1] ,
    \cb_6_2_io_o_4_out[0] }),
    .io_i_5_in1({\cb_6_2_io_o_5_out[7] ,
    \cb_6_2_io_o_5_out[6] ,
    \cb_6_2_io_o_5_out[5] ,
    \cb_6_2_io_o_5_out[4] ,
    \cb_6_2_io_o_5_out[3] ,
    \cb_6_2_io_o_5_out[2] ,
    \cb_6_2_io_o_5_out[1] ,
    \cb_6_2_io_o_5_out[0] }),
    .io_i_6_in1({\cb_6_2_io_o_6_out[7] ,
    \cb_6_2_io_o_6_out[6] ,
    \cb_6_2_io_o_6_out[5] ,
    \cb_6_2_io_o_6_out[4] ,
    \cb_6_2_io_o_6_out[3] ,
    \cb_6_2_io_o_6_out[2] ,
    \cb_6_2_io_o_6_out[1] ,
    \cb_6_2_io_o_6_out[0] }),
    .io_i_7_in1({\cb_6_2_io_o_7_out[7] ,
    \cb_6_2_io_o_7_out[6] ,
    \cb_6_2_io_o_7_out[5] ,
    \cb_6_2_io_o_7_out[4] ,
    \cb_6_2_io_o_7_out[3] ,
    \cb_6_2_io_o_7_out[2] ,
    \cb_6_2_io_o_7_out[1] ,
    \cb_6_2_io_o_7_out[0] }),
    .io_o_0_out({\cb_6_3_io_o_0_out[7] ,
    \cb_6_3_io_o_0_out[6] ,
    \cb_6_3_io_o_0_out[5] ,
    \cb_6_3_io_o_0_out[4] ,
    \cb_6_3_io_o_0_out[3] ,
    \cb_6_3_io_o_0_out[2] ,
    \cb_6_3_io_o_0_out[1] ,
    \cb_6_3_io_o_0_out[0] }),
    .io_o_1_out({\cb_6_3_io_o_1_out[7] ,
    \cb_6_3_io_o_1_out[6] ,
    \cb_6_3_io_o_1_out[5] ,
    \cb_6_3_io_o_1_out[4] ,
    \cb_6_3_io_o_1_out[3] ,
    \cb_6_3_io_o_1_out[2] ,
    \cb_6_3_io_o_1_out[1] ,
    \cb_6_3_io_o_1_out[0] }),
    .io_o_2_out({\cb_6_3_io_o_2_out[7] ,
    \cb_6_3_io_o_2_out[6] ,
    \cb_6_3_io_o_2_out[5] ,
    \cb_6_3_io_o_2_out[4] ,
    \cb_6_3_io_o_2_out[3] ,
    \cb_6_3_io_o_2_out[2] ,
    \cb_6_3_io_o_2_out[1] ,
    \cb_6_3_io_o_2_out[0] }),
    .io_o_3_out({\cb_6_3_io_o_3_out[7] ,
    \cb_6_3_io_o_3_out[6] ,
    \cb_6_3_io_o_3_out[5] ,
    \cb_6_3_io_o_3_out[4] ,
    \cb_6_3_io_o_3_out[3] ,
    \cb_6_3_io_o_3_out[2] ,
    \cb_6_3_io_o_3_out[1] ,
    \cb_6_3_io_o_3_out[0] }),
    .io_o_4_out({\cb_6_3_io_o_4_out[7] ,
    \cb_6_3_io_o_4_out[6] ,
    \cb_6_3_io_o_4_out[5] ,
    \cb_6_3_io_o_4_out[4] ,
    \cb_6_3_io_o_4_out[3] ,
    \cb_6_3_io_o_4_out[2] ,
    \cb_6_3_io_o_4_out[1] ,
    \cb_6_3_io_o_4_out[0] }),
    .io_o_5_out({\cb_6_3_io_o_5_out[7] ,
    \cb_6_3_io_o_5_out[6] ,
    \cb_6_3_io_o_5_out[5] ,
    \cb_6_3_io_o_5_out[4] ,
    \cb_6_3_io_o_5_out[3] ,
    \cb_6_3_io_o_5_out[2] ,
    \cb_6_3_io_o_5_out[1] ,
    \cb_6_3_io_o_5_out[0] }),
    .io_o_6_out({\cb_6_3_io_o_6_out[7] ,
    \cb_6_3_io_o_6_out[6] ,
    \cb_6_3_io_o_6_out[5] ,
    \cb_6_3_io_o_6_out[4] ,
    \cb_6_3_io_o_6_out[3] ,
    \cb_6_3_io_o_6_out[2] ,
    \cb_6_3_io_o_6_out[1] ,
    \cb_6_3_io_o_6_out[0] }),
    .io_o_7_out({\cb_6_3_io_o_7_out[7] ,
    \cb_6_3_io_o_7_out[6] ,
    \cb_6_3_io_o_7_out[5] ,
    \cb_6_3_io_o_7_out[4] ,
    \cb_6_3_io_o_7_out[3] ,
    \cb_6_3_io_o_7_out[2] ,
    \cb_6_3_io_o_7_out[1] ,
    \cb_6_3_io_o_7_out[0] }),
    .io_wo({\cb_6_2_io_eo[63] ,
    \cb_6_2_io_eo[62] ,
    \cb_6_2_io_eo[61] ,
    \cb_6_2_io_eo[60] ,
    \cb_6_2_io_eo[59] ,
    \cb_6_2_io_eo[58] ,
    \cb_6_2_io_eo[57] ,
    \cb_6_2_io_eo[56] ,
    \cb_6_2_io_eo[55] ,
    \cb_6_2_io_eo[54] ,
    \cb_6_2_io_eo[53] ,
    \cb_6_2_io_eo[52] ,
    \cb_6_2_io_eo[51] ,
    \cb_6_2_io_eo[50] ,
    \cb_6_2_io_eo[49] ,
    \cb_6_2_io_eo[48] ,
    \cb_6_2_io_eo[47] ,
    \cb_6_2_io_eo[46] ,
    \cb_6_2_io_eo[45] ,
    \cb_6_2_io_eo[44] ,
    \cb_6_2_io_eo[43] ,
    \cb_6_2_io_eo[42] ,
    \cb_6_2_io_eo[41] ,
    \cb_6_2_io_eo[40] ,
    \cb_6_2_io_eo[39] ,
    \cb_6_2_io_eo[38] ,
    \cb_6_2_io_eo[37] ,
    \cb_6_2_io_eo[36] ,
    \cb_6_2_io_eo[35] ,
    \cb_6_2_io_eo[34] ,
    \cb_6_2_io_eo[33] ,
    \cb_6_2_io_eo[32] ,
    \cb_6_2_io_eo[31] ,
    \cb_6_2_io_eo[30] ,
    \cb_6_2_io_eo[29] ,
    \cb_6_2_io_eo[28] ,
    \cb_6_2_io_eo[27] ,
    \cb_6_2_io_eo[26] ,
    \cb_6_2_io_eo[25] ,
    \cb_6_2_io_eo[24] ,
    \cb_6_2_io_eo[23] ,
    \cb_6_2_io_eo[22] ,
    \cb_6_2_io_eo[21] ,
    \cb_6_2_io_eo[20] ,
    \cb_6_2_io_eo[19] ,
    \cb_6_2_io_eo[18] ,
    \cb_6_2_io_eo[17] ,
    \cb_6_2_io_eo[16] ,
    \cb_6_2_io_eo[15] ,
    \cb_6_2_io_eo[14] ,
    \cb_6_2_io_eo[13] ,
    \cb_6_2_io_eo[12] ,
    \cb_6_2_io_eo[11] ,
    \cb_6_2_io_eo[10] ,
    \cb_6_2_io_eo[9] ,
    \cb_6_2_io_eo[8] ,
    \cb_6_2_io_eo[7] ,
    \cb_6_2_io_eo[6] ,
    \cb_6_2_io_eo[5] ,
    \cb_6_2_io_eo[4] ,
    \cb_6_2_io_eo[3] ,
    \cb_6_2_io_eo[2] ,
    \cb_6_2_io_eo[1] ,
    \cb_6_2_io_eo[0] }));
 cic_block cb_6_4 (.io_cs_i(cb_6_4_io_cs_i),
    .io_i_0_ci(cb_6_3_io_o_0_co),
    .io_i_1_ci(cb_6_3_io_o_1_co),
    .io_i_2_ci(cb_6_3_io_o_2_co),
    .io_i_3_ci(cb_6_3_io_o_3_co),
    .io_i_4_ci(cb_6_3_io_o_4_co),
    .io_i_5_ci(cb_6_3_io_o_5_co),
    .io_i_6_ci(cb_6_3_io_o_6_co),
    .io_i_7_ci(cb_6_3_io_o_7_co),
    .io_o_0_co(cb_6_4_io_o_0_co),
    .io_o_1_co(cb_6_4_io_o_1_co),
    .io_o_2_co(cb_6_4_io_o_2_co),
    .io_o_3_co(cb_6_4_io_o_3_co),
    .io_o_4_co(cb_6_4_io_o_4_co),
    .io_o_5_co(cb_6_4_io_o_5_co),
    .io_o_6_co(cb_6_4_io_o_6_co),
    .io_o_7_co(cb_6_4_io_o_7_co),
    .io_vci(cb_6_3_io_vco),
    .io_vco(cb_6_4_io_vco),
    .io_vi(cb_6_4_io_vi),
    .io_we_i(cb_6_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_6_0_io_adr_i[1] ,
    \cb_6_0_io_adr_i[0] }),
    .io_dat_i({\cb_6_0_io_dat_i[15] ,
    \cb_6_0_io_dat_i[14] ,
    \cb_6_0_io_dat_i[13] ,
    \cb_6_0_io_dat_i[12] ,
    \cb_6_0_io_dat_i[11] ,
    \cb_6_0_io_dat_i[10] ,
    \cb_6_0_io_dat_i[9] ,
    \cb_6_0_io_dat_i[8] ,
    \cb_6_0_io_dat_i[7] ,
    \cb_6_0_io_dat_i[6] ,
    \cb_6_0_io_dat_i[5] ,
    \cb_6_0_io_dat_i[4] ,
    \cb_6_0_io_dat_i[3] ,
    \cb_6_0_io_dat_i[2] ,
    \cb_6_0_io_dat_i[1] ,
    \cb_6_0_io_dat_i[0] }),
    .io_dat_o({\cb_6_4_io_dat_o[15] ,
    \cb_6_4_io_dat_o[14] ,
    \cb_6_4_io_dat_o[13] ,
    \cb_6_4_io_dat_o[12] ,
    \cb_6_4_io_dat_o[11] ,
    \cb_6_4_io_dat_o[10] ,
    \cb_6_4_io_dat_o[9] ,
    \cb_6_4_io_dat_o[8] ,
    \cb_6_4_io_dat_o[7] ,
    \cb_6_4_io_dat_o[6] ,
    \cb_6_4_io_dat_o[5] ,
    \cb_6_4_io_dat_o[4] ,
    \cb_6_4_io_dat_o[3] ,
    \cb_6_4_io_dat_o[2] ,
    \cb_6_4_io_dat_o[1] ,
    \cb_6_4_io_dat_o[0] }),
    .io_eo({\cb_6_4_io_eo[63] ,
    \cb_6_4_io_eo[62] ,
    \cb_6_4_io_eo[61] ,
    \cb_6_4_io_eo[60] ,
    \cb_6_4_io_eo[59] ,
    \cb_6_4_io_eo[58] ,
    \cb_6_4_io_eo[57] ,
    \cb_6_4_io_eo[56] ,
    \cb_6_4_io_eo[55] ,
    \cb_6_4_io_eo[54] ,
    \cb_6_4_io_eo[53] ,
    \cb_6_4_io_eo[52] ,
    \cb_6_4_io_eo[51] ,
    \cb_6_4_io_eo[50] ,
    \cb_6_4_io_eo[49] ,
    \cb_6_4_io_eo[48] ,
    \cb_6_4_io_eo[47] ,
    \cb_6_4_io_eo[46] ,
    \cb_6_4_io_eo[45] ,
    \cb_6_4_io_eo[44] ,
    \cb_6_4_io_eo[43] ,
    \cb_6_4_io_eo[42] ,
    \cb_6_4_io_eo[41] ,
    \cb_6_4_io_eo[40] ,
    \cb_6_4_io_eo[39] ,
    \cb_6_4_io_eo[38] ,
    \cb_6_4_io_eo[37] ,
    \cb_6_4_io_eo[36] ,
    \cb_6_4_io_eo[35] ,
    \cb_6_4_io_eo[34] ,
    \cb_6_4_io_eo[33] ,
    \cb_6_4_io_eo[32] ,
    \cb_6_4_io_eo[31] ,
    \cb_6_4_io_eo[30] ,
    \cb_6_4_io_eo[29] ,
    \cb_6_4_io_eo[28] ,
    \cb_6_4_io_eo[27] ,
    \cb_6_4_io_eo[26] ,
    \cb_6_4_io_eo[25] ,
    \cb_6_4_io_eo[24] ,
    \cb_6_4_io_eo[23] ,
    \cb_6_4_io_eo[22] ,
    \cb_6_4_io_eo[21] ,
    \cb_6_4_io_eo[20] ,
    \cb_6_4_io_eo[19] ,
    \cb_6_4_io_eo[18] ,
    \cb_6_4_io_eo[17] ,
    \cb_6_4_io_eo[16] ,
    \cb_6_4_io_eo[15] ,
    \cb_6_4_io_eo[14] ,
    \cb_6_4_io_eo[13] ,
    \cb_6_4_io_eo[12] ,
    \cb_6_4_io_eo[11] ,
    \cb_6_4_io_eo[10] ,
    \cb_6_4_io_eo[9] ,
    \cb_6_4_io_eo[8] ,
    \cb_6_4_io_eo[7] ,
    \cb_6_4_io_eo[6] ,
    \cb_6_4_io_eo[5] ,
    \cb_6_4_io_eo[4] ,
    \cb_6_4_io_eo[3] ,
    \cb_6_4_io_eo[2] ,
    \cb_6_4_io_eo[1] ,
    \cb_6_4_io_eo[0] }),
    .io_i_0_in1({\cb_6_3_io_o_0_out[7] ,
    \cb_6_3_io_o_0_out[6] ,
    \cb_6_3_io_o_0_out[5] ,
    \cb_6_3_io_o_0_out[4] ,
    \cb_6_3_io_o_0_out[3] ,
    \cb_6_3_io_o_0_out[2] ,
    \cb_6_3_io_o_0_out[1] ,
    \cb_6_3_io_o_0_out[0] }),
    .io_i_1_in1({\cb_6_3_io_o_1_out[7] ,
    \cb_6_3_io_o_1_out[6] ,
    \cb_6_3_io_o_1_out[5] ,
    \cb_6_3_io_o_1_out[4] ,
    \cb_6_3_io_o_1_out[3] ,
    \cb_6_3_io_o_1_out[2] ,
    \cb_6_3_io_o_1_out[1] ,
    \cb_6_3_io_o_1_out[0] }),
    .io_i_2_in1({\cb_6_3_io_o_2_out[7] ,
    \cb_6_3_io_o_2_out[6] ,
    \cb_6_3_io_o_2_out[5] ,
    \cb_6_3_io_o_2_out[4] ,
    \cb_6_3_io_o_2_out[3] ,
    \cb_6_3_io_o_2_out[2] ,
    \cb_6_3_io_o_2_out[1] ,
    \cb_6_3_io_o_2_out[0] }),
    .io_i_3_in1({\cb_6_3_io_o_3_out[7] ,
    \cb_6_3_io_o_3_out[6] ,
    \cb_6_3_io_o_3_out[5] ,
    \cb_6_3_io_o_3_out[4] ,
    \cb_6_3_io_o_3_out[3] ,
    \cb_6_3_io_o_3_out[2] ,
    \cb_6_3_io_o_3_out[1] ,
    \cb_6_3_io_o_3_out[0] }),
    .io_i_4_in1({\cb_6_3_io_o_4_out[7] ,
    \cb_6_3_io_o_4_out[6] ,
    \cb_6_3_io_o_4_out[5] ,
    \cb_6_3_io_o_4_out[4] ,
    \cb_6_3_io_o_4_out[3] ,
    \cb_6_3_io_o_4_out[2] ,
    \cb_6_3_io_o_4_out[1] ,
    \cb_6_3_io_o_4_out[0] }),
    .io_i_5_in1({\cb_6_3_io_o_5_out[7] ,
    \cb_6_3_io_o_5_out[6] ,
    \cb_6_3_io_o_5_out[5] ,
    \cb_6_3_io_o_5_out[4] ,
    \cb_6_3_io_o_5_out[3] ,
    \cb_6_3_io_o_5_out[2] ,
    \cb_6_3_io_o_5_out[1] ,
    \cb_6_3_io_o_5_out[0] }),
    .io_i_6_in1({\cb_6_3_io_o_6_out[7] ,
    \cb_6_3_io_o_6_out[6] ,
    \cb_6_3_io_o_6_out[5] ,
    \cb_6_3_io_o_6_out[4] ,
    \cb_6_3_io_o_6_out[3] ,
    \cb_6_3_io_o_6_out[2] ,
    \cb_6_3_io_o_6_out[1] ,
    \cb_6_3_io_o_6_out[0] }),
    .io_i_7_in1({\cb_6_3_io_o_7_out[7] ,
    \cb_6_3_io_o_7_out[6] ,
    \cb_6_3_io_o_7_out[5] ,
    \cb_6_3_io_o_7_out[4] ,
    \cb_6_3_io_o_7_out[3] ,
    \cb_6_3_io_o_7_out[2] ,
    \cb_6_3_io_o_7_out[1] ,
    \cb_6_3_io_o_7_out[0] }),
    .io_o_0_out({\cb_6_4_io_o_0_out[7] ,
    \cb_6_4_io_o_0_out[6] ,
    \cb_6_4_io_o_0_out[5] ,
    \cb_6_4_io_o_0_out[4] ,
    \cb_6_4_io_o_0_out[3] ,
    \cb_6_4_io_o_0_out[2] ,
    \cb_6_4_io_o_0_out[1] ,
    \cb_6_4_io_o_0_out[0] }),
    .io_o_1_out({\cb_6_4_io_o_1_out[7] ,
    \cb_6_4_io_o_1_out[6] ,
    \cb_6_4_io_o_1_out[5] ,
    \cb_6_4_io_o_1_out[4] ,
    \cb_6_4_io_o_1_out[3] ,
    \cb_6_4_io_o_1_out[2] ,
    \cb_6_4_io_o_1_out[1] ,
    \cb_6_4_io_o_1_out[0] }),
    .io_o_2_out({\cb_6_4_io_o_2_out[7] ,
    \cb_6_4_io_o_2_out[6] ,
    \cb_6_4_io_o_2_out[5] ,
    \cb_6_4_io_o_2_out[4] ,
    \cb_6_4_io_o_2_out[3] ,
    \cb_6_4_io_o_2_out[2] ,
    \cb_6_4_io_o_2_out[1] ,
    \cb_6_4_io_o_2_out[0] }),
    .io_o_3_out({\cb_6_4_io_o_3_out[7] ,
    \cb_6_4_io_o_3_out[6] ,
    \cb_6_4_io_o_3_out[5] ,
    \cb_6_4_io_o_3_out[4] ,
    \cb_6_4_io_o_3_out[3] ,
    \cb_6_4_io_o_3_out[2] ,
    \cb_6_4_io_o_3_out[1] ,
    \cb_6_4_io_o_3_out[0] }),
    .io_o_4_out({\cb_6_4_io_o_4_out[7] ,
    \cb_6_4_io_o_4_out[6] ,
    \cb_6_4_io_o_4_out[5] ,
    \cb_6_4_io_o_4_out[4] ,
    \cb_6_4_io_o_4_out[3] ,
    \cb_6_4_io_o_4_out[2] ,
    \cb_6_4_io_o_4_out[1] ,
    \cb_6_4_io_o_4_out[0] }),
    .io_o_5_out({\cb_6_4_io_o_5_out[7] ,
    \cb_6_4_io_o_5_out[6] ,
    \cb_6_4_io_o_5_out[5] ,
    \cb_6_4_io_o_5_out[4] ,
    \cb_6_4_io_o_5_out[3] ,
    \cb_6_4_io_o_5_out[2] ,
    \cb_6_4_io_o_5_out[1] ,
    \cb_6_4_io_o_5_out[0] }),
    .io_o_6_out({\cb_6_4_io_o_6_out[7] ,
    \cb_6_4_io_o_6_out[6] ,
    \cb_6_4_io_o_6_out[5] ,
    \cb_6_4_io_o_6_out[4] ,
    \cb_6_4_io_o_6_out[3] ,
    \cb_6_4_io_o_6_out[2] ,
    \cb_6_4_io_o_6_out[1] ,
    \cb_6_4_io_o_6_out[0] }),
    .io_o_7_out({\cb_6_4_io_o_7_out[7] ,
    \cb_6_4_io_o_7_out[6] ,
    \cb_6_4_io_o_7_out[5] ,
    \cb_6_4_io_o_7_out[4] ,
    \cb_6_4_io_o_7_out[3] ,
    \cb_6_4_io_o_7_out[2] ,
    \cb_6_4_io_o_7_out[1] ,
    \cb_6_4_io_o_7_out[0] }),
    .io_wo({\cb_6_3_io_eo[63] ,
    \cb_6_3_io_eo[62] ,
    \cb_6_3_io_eo[61] ,
    \cb_6_3_io_eo[60] ,
    \cb_6_3_io_eo[59] ,
    \cb_6_3_io_eo[58] ,
    \cb_6_3_io_eo[57] ,
    \cb_6_3_io_eo[56] ,
    \cb_6_3_io_eo[55] ,
    \cb_6_3_io_eo[54] ,
    \cb_6_3_io_eo[53] ,
    \cb_6_3_io_eo[52] ,
    \cb_6_3_io_eo[51] ,
    \cb_6_3_io_eo[50] ,
    \cb_6_3_io_eo[49] ,
    \cb_6_3_io_eo[48] ,
    \cb_6_3_io_eo[47] ,
    \cb_6_3_io_eo[46] ,
    \cb_6_3_io_eo[45] ,
    \cb_6_3_io_eo[44] ,
    \cb_6_3_io_eo[43] ,
    \cb_6_3_io_eo[42] ,
    \cb_6_3_io_eo[41] ,
    \cb_6_3_io_eo[40] ,
    \cb_6_3_io_eo[39] ,
    \cb_6_3_io_eo[38] ,
    \cb_6_3_io_eo[37] ,
    \cb_6_3_io_eo[36] ,
    \cb_6_3_io_eo[35] ,
    \cb_6_3_io_eo[34] ,
    \cb_6_3_io_eo[33] ,
    \cb_6_3_io_eo[32] ,
    \cb_6_3_io_eo[31] ,
    \cb_6_3_io_eo[30] ,
    \cb_6_3_io_eo[29] ,
    \cb_6_3_io_eo[28] ,
    \cb_6_3_io_eo[27] ,
    \cb_6_3_io_eo[26] ,
    \cb_6_3_io_eo[25] ,
    \cb_6_3_io_eo[24] ,
    \cb_6_3_io_eo[23] ,
    \cb_6_3_io_eo[22] ,
    \cb_6_3_io_eo[21] ,
    \cb_6_3_io_eo[20] ,
    \cb_6_3_io_eo[19] ,
    \cb_6_3_io_eo[18] ,
    \cb_6_3_io_eo[17] ,
    \cb_6_3_io_eo[16] ,
    \cb_6_3_io_eo[15] ,
    \cb_6_3_io_eo[14] ,
    \cb_6_3_io_eo[13] ,
    \cb_6_3_io_eo[12] ,
    \cb_6_3_io_eo[11] ,
    \cb_6_3_io_eo[10] ,
    \cb_6_3_io_eo[9] ,
    \cb_6_3_io_eo[8] ,
    \cb_6_3_io_eo[7] ,
    \cb_6_3_io_eo[6] ,
    \cb_6_3_io_eo[5] ,
    \cb_6_3_io_eo[4] ,
    \cb_6_3_io_eo[3] ,
    \cb_6_3_io_eo[2] ,
    \cb_6_3_io_eo[1] ,
    \cb_6_3_io_eo[0] }));
 cic_block cb_6_5 (.io_cs_i(cb_6_5_io_cs_i),
    .io_i_0_ci(cb_6_4_io_o_0_co),
    .io_i_1_ci(cb_6_4_io_o_1_co),
    .io_i_2_ci(cb_6_4_io_o_2_co),
    .io_i_3_ci(cb_6_4_io_o_3_co),
    .io_i_4_ci(cb_6_4_io_o_4_co),
    .io_i_5_ci(cb_6_4_io_o_5_co),
    .io_i_6_ci(cb_6_4_io_o_6_co),
    .io_i_7_ci(cb_6_4_io_o_7_co),
    .io_o_0_co(cb_6_5_io_o_0_co),
    .io_o_1_co(cb_6_5_io_o_1_co),
    .io_o_2_co(cb_6_5_io_o_2_co),
    .io_o_3_co(cb_6_5_io_o_3_co),
    .io_o_4_co(cb_6_5_io_o_4_co),
    .io_o_5_co(cb_6_5_io_o_5_co),
    .io_o_6_co(cb_6_5_io_o_6_co),
    .io_o_7_co(cb_6_5_io_o_7_co),
    .io_vci(cb_6_4_io_vco),
    .io_vco(cb_6_5_io_vco),
    .io_vi(cb_6_5_io_vi),
    .io_we_i(cb_6_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_6_0_io_adr_i[1] ,
    \cb_6_0_io_adr_i[0] }),
    .io_dat_i({\cb_6_0_io_dat_i[15] ,
    \cb_6_0_io_dat_i[14] ,
    \cb_6_0_io_dat_i[13] ,
    \cb_6_0_io_dat_i[12] ,
    \cb_6_0_io_dat_i[11] ,
    \cb_6_0_io_dat_i[10] ,
    \cb_6_0_io_dat_i[9] ,
    \cb_6_0_io_dat_i[8] ,
    \cb_6_0_io_dat_i[7] ,
    \cb_6_0_io_dat_i[6] ,
    \cb_6_0_io_dat_i[5] ,
    \cb_6_0_io_dat_i[4] ,
    \cb_6_0_io_dat_i[3] ,
    \cb_6_0_io_dat_i[2] ,
    \cb_6_0_io_dat_i[1] ,
    \cb_6_0_io_dat_i[0] }),
    .io_dat_o({\cb_6_5_io_dat_o[15] ,
    \cb_6_5_io_dat_o[14] ,
    \cb_6_5_io_dat_o[13] ,
    \cb_6_5_io_dat_o[12] ,
    \cb_6_5_io_dat_o[11] ,
    \cb_6_5_io_dat_o[10] ,
    \cb_6_5_io_dat_o[9] ,
    \cb_6_5_io_dat_o[8] ,
    \cb_6_5_io_dat_o[7] ,
    \cb_6_5_io_dat_o[6] ,
    \cb_6_5_io_dat_o[5] ,
    \cb_6_5_io_dat_o[4] ,
    \cb_6_5_io_dat_o[3] ,
    \cb_6_5_io_dat_o[2] ,
    \cb_6_5_io_dat_o[1] ,
    \cb_6_5_io_dat_o[0] }),
    .io_eo({\cb_6_5_io_eo[63] ,
    \cb_6_5_io_eo[62] ,
    \cb_6_5_io_eo[61] ,
    \cb_6_5_io_eo[60] ,
    \cb_6_5_io_eo[59] ,
    \cb_6_5_io_eo[58] ,
    \cb_6_5_io_eo[57] ,
    \cb_6_5_io_eo[56] ,
    \cb_6_5_io_eo[55] ,
    \cb_6_5_io_eo[54] ,
    \cb_6_5_io_eo[53] ,
    \cb_6_5_io_eo[52] ,
    \cb_6_5_io_eo[51] ,
    \cb_6_5_io_eo[50] ,
    \cb_6_5_io_eo[49] ,
    \cb_6_5_io_eo[48] ,
    \cb_6_5_io_eo[47] ,
    \cb_6_5_io_eo[46] ,
    \cb_6_5_io_eo[45] ,
    \cb_6_5_io_eo[44] ,
    \cb_6_5_io_eo[43] ,
    \cb_6_5_io_eo[42] ,
    \cb_6_5_io_eo[41] ,
    \cb_6_5_io_eo[40] ,
    \cb_6_5_io_eo[39] ,
    \cb_6_5_io_eo[38] ,
    \cb_6_5_io_eo[37] ,
    \cb_6_5_io_eo[36] ,
    \cb_6_5_io_eo[35] ,
    \cb_6_5_io_eo[34] ,
    \cb_6_5_io_eo[33] ,
    \cb_6_5_io_eo[32] ,
    \cb_6_5_io_eo[31] ,
    \cb_6_5_io_eo[30] ,
    \cb_6_5_io_eo[29] ,
    \cb_6_5_io_eo[28] ,
    \cb_6_5_io_eo[27] ,
    \cb_6_5_io_eo[26] ,
    \cb_6_5_io_eo[25] ,
    \cb_6_5_io_eo[24] ,
    \cb_6_5_io_eo[23] ,
    \cb_6_5_io_eo[22] ,
    \cb_6_5_io_eo[21] ,
    \cb_6_5_io_eo[20] ,
    \cb_6_5_io_eo[19] ,
    \cb_6_5_io_eo[18] ,
    \cb_6_5_io_eo[17] ,
    \cb_6_5_io_eo[16] ,
    \cb_6_5_io_eo[15] ,
    \cb_6_5_io_eo[14] ,
    \cb_6_5_io_eo[13] ,
    \cb_6_5_io_eo[12] ,
    \cb_6_5_io_eo[11] ,
    \cb_6_5_io_eo[10] ,
    \cb_6_5_io_eo[9] ,
    \cb_6_5_io_eo[8] ,
    \cb_6_5_io_eo[7] ,
    \cb_6_5_io_eo[6] ,
    \cb_6_5_io_eo[5] ,
    \cb_6_5_io_eo[4] ,
    \cb_6_5_io_eo[3] ,
    \cb_6_5_io_eo[2] ,
    \cb_6_5_io_eo[1] ,
    \cb_6_5_io_eo[0] }),
    .io_i_0_in1({\cb_6_4_io_o_0_out[7] ,
    \cb_6_4_io_o_0_out[6] ,
    \cb_6_4_io_o_0_out[5] ,
    \cb_6_4_io_o_0_out[4] ,
    \cb_6_4_io_o_0_out[3] ,
    \cb_6_4_io_o_0_out[2] ,
    \cb_6_4_io_o_0_out[1] ,
    \cb_6_4_io_o_0_out[0] }),
    .io_i_1_in1({\cb_6_4_io_o_1_out[7] ,
    \cb_6_4_io_o_1_out[6] ,
    \cb_6_4_io_o_1_out[5] ,
    \cb_6_4_io_o_1_out[4] ,
    \cb_6_4_io_o_1_out[3] ,
    \cb_6_4_io_o_1_out[2] ,
    \cb_6_4_io_o_1_out[1] ,
    \cb_6_4_io_o_1_out[0] }),
    .io_i_2_in1({\cb_6_4_io_o_2_out[7] ,
    \cb_6_4_io_o_2_out[6] ,
    \cb_6_4_io_o_2_out[5] ,
    \cb_6_4_io_o_2_out[4] ,
    \cb_6_4_io_o_2_out[3] ,
    \cb_6_4_io_o_2_out[2] ,
    \cb_6_4_io_o_2_out[1] ,
    \cb_6_4_io_o_2_out[0] }),
    .io_i_3_in1({\cb_6_4_io_o_3_out[7] ,
    \cb_6_4_io_o_3_out[6] ,
    \cb_6_4_io_o_3_out[5] ,
    \cb_6_4_io_o_3_out[4] ,
    \cb_6_4_io_o_3_out[3] ,
    \cb_6_4_io_o_3_out[2] ,
    \cb_6_4_io_o_3_out[1] ,
    \cb_6_4_io_o_3_out[0] }),
    .io_i_4_in1({\cb_6_4_io_o_4_out[7] ,
    \cb_6_4_io_o_4_out[6] ,
    \cb_6_4_io_o_4_out[5] ,
    \cb_6_4_io_o_4_out[4] ,
    \cb_6_4_io_o_4_out[3] ,
    \cb_6_4_io_o_4_out[2] ,
    \cb_6_4_io_o_4_out[1] ,
    \cb_6_4_io_o_4_out[0] }),
    .io_i_5_in1({\cb_6_4_io_o_5_out[7] ,
    \cb_6_4_io_o_5_out[6] ,
    \cb_6_4_io_o_5_out[5] ,
    \cb_6_4_io_o_5_out[4] ,
    \cb_6_4_io_o_5_out[3] ,
    \cb_6_4_io_o_5_out[2] ,
    \cb_6_4_io_o_5_out[1] ,
    \cb_6_4_io_o_5_out[0] }),
    .io_i_6_in1({\cb_6_4_io_o_6_out[7] ,
    \cb_6_4_io_o_6_out[6] ,
    \cb_6_4_io_o_6_out[5] ,
    \cb_6_4_io_o_6_out[4] ,
    \cb_6_4_io_o_6_out[3] ,
    \cb_6_4_io_o_6_out[2] ,
    \cb_6_4_io_o_6_out[1] ,
    \cb_6_4_io_o_6_out[0] }),
    .io_i_7_in1({\cb_6_4_io_o_7_out[7] ,
    \cb_6_4_io_o_7_out[6] ,
    \cb_6_4_io_o_7_out[5] ,
    \cb_6_4_io_o_7_out[4] ,
    \cb_6_4_io_o_7_out[3] ,
    \cb_6_4_io_o_7_out[2] ,
    \cb_6_4_io_o_7_out[1] ,
    \cb_6_4_io_o_7_out[0] }),
    .io_o_0_out({\cb_6_5_io_o_0_out[7] ,
    \cb_6_5_io_o_0_out[6] ,
    \cb_6_5_io_o_0_out[5] ,
    \cb_6_5_io_o_0_out[4] ,
    \cb_6_5_io_o_0_out[3] ,
    \cb_6_5_io_o_0_out[2] ,
    \cb_6_5_io_o_0_out[1] ,
    \cb_6_5_io_o_0_out[0] }),
    .io_o_1_out({\cb_6_5_io_o_1_out[7] ,
    \cb_6_5_io_o_1_out[6] ,
    \cb_6_5_io_o_1_out[5] ,
    \cb_6_5_io_o_1_out[4] ,
    \cb_6_5_io_o_1_out[3] ,
    \cb_6_5_io_o_1_out[2] ,
    \cb_6_5_io_o_1_out[1] ,
    \cb_6_5_io_o_1_out[0] }),
    .io_o_2_out({\cb_6_5_io_o_2_out[7] ,
    \cb_6_5_io_o_2_out[6] ,
    \cb_6_5_io_o_2_out[5] ,
    \cb_6_5_io_o_2_out[4] ,
    \cb_6_5_io_o_2_out[3] ,
    \cb_6_5_io_o_2_out[2] ,
    \cb_6_5_io_o_2_out[1] ,
    \cb_6_5_io_o_2_out[0] }),
    .io_o_3_out({\cb_6_5_io_o_3_out[7] ,
    \cb_6_5_io_o_3_out[6] ,
    \cb_6_5_io_o_3_out[5] ,
    \cb_6_5_io_o_3_out[4] ,
    \cb_6_5_io_o_3_out[3] ,
    \cb_6_5_io_o_3_out[2] ,
    \cb_6_5_io_o_3_out[1] ,
    \cb_6_5_io_o_3_out[0] }),
    .io_o_4_out({\cb_6_5_io_o_4_out[7] ,
    \cb_6_5_io_o_4_out[6] ,
    \cb_6_5_io_o_4_out[5] ,
    \cb_6_5_io_o_4_out[4] ,
    \cb_6_5_io_o_4_out[3] ,
    \cb_6_5_io_o_4_out[2] ,
    \cb_6_5_io_o_4_out[1] ,
    \cb_6_5_io_o_4_out[0] }),
    .io_o_5_out({\cb_6_5_io_o_5_out[7] ,
    \cb_6_5_io_o_5_out[6] ,
    \cb_6_5_io_o_5_out[5] ,
    \cb_6_5_io_o_5_out[4] ,
    \cb_6_5_io_o_5_out[3] ,
    \cb_6_5_io_o_5_out[2] ,
    \cb_6_5_io_o_5_out[1] ,
    \cb_6_5_io_o_5_out[0] }),
    .io_o_6_out({\cb_6_5_io_o_6_out[7] ,
    \cb_6_5_io_o_6_out[6] ,
    \cb_6_5_io_o_6_out[5] ,
    \cb_6_5_io_o_6_out[4] ,
    \cb_6_5_io_o_6_out[3] ,
    \cb_6_5_io_o_6_out[2] ,
    \cb_6_5_io_o_6_out[1] ,
    \cb_6_5_io_o_6_out[0] }),
    .io_o_7_out({\cb_6_5_io_o_7_out[7] ,
    \cb_6_5_io_o_7_out[6] ,
    \cb_6_5_io_o_7_out[5] ,
    \cb_6_5_io_o_7_out[4] ,
    \cb_6_5_io_o_7_out[3] ,
    \cb_6_5_io_o_7_out[2] ,
    \cb_6_5_io_o_7_out[1] ,
    \cb_6_5_io_o_7_out[0] }),
    .io_wo({\cb_6_4_io_eo[63] ,
    \cb_6_4_io_eo[62] ,
    \cb_6_4_io_eo[61] ,
    \cb_6_4_io_eo[60] ,
    \cb_6_4_io_eo[59] ,
    \cb_6_4_io_eo[58] ,
    \cb_6_4_io_eo[57] ,
    \cb_6_4_io_eo[56] ,
    \cb_6_4_io_eo[55] ,
    \cb_6_4_io_eo[54] ,
    \cb_6_4_io_eo[53] ,
    \cb_6_4_io_eo[52] ,
    \cb_6_4_io_eo[51] ,
    \cb_6_4_io_eo[50] ,
    \cb_6_4_io_eo[49] ,
    \cb_6_4_io_eo[48] ,
    \cb_6_4_io_eo[47] ,
    \cb_6_4_io_eo[46] ,
    \cb_6_4_io_eo[45] ,
    \cb_6_4_io_eo[44] ,
    \cb_6_4_io_eo[43] ,
    \cb_6_4_io_eo[42] ,
    \cb_6_4_io_eo[41] ,
    \cb_6_4_io_eo[40] ,
    \cb_6_4_io_eo[39] ,
    \cb_6_4_io_eo[38] ,
    \cb_6_4_io_eo[37] ,
    \cb_6_4_io_eo[36] ,
    \cb_6_4_io_eo[35] ,
    \cb_6_4_io_eo[34] ,
    \cb_6_4_io_eo[33] ,
    \cb_6_4_io_eo[32] ,
    \cb_6_4_io_eo[31] ,
    \cb_6_4_io_eo[30] ,
    \cb_6_4_io_eo[29] ,
    \cb_6_4_io_eo[28] ,
    \cb_6_4_io_eo[27] ,
    \cb_6_4_io_eo[26] ,
    \cb_6_4_io_eo[25] ,
    \cb_6_4_io_eo[24] ,
    \cb_6_4_io_eo[23] ,
    \cb_6_4_io_eo[22] ,
    \cb_6_4_io_eo[21] ,
    \cb_6_4_io_eo[20] ,
    \cb_6_4_io_eo[19] ,
    \cb_6_4_io_eo[18] ,
    \cb_6_4_io_eo[17] ,
    \cb_6_4_io_eo[16] ,
    \cb_6_4_io_eo[15] ,
    \cb_6_4_io_eo[14] ,
    \cb_6_4_io_eo[13] ,
    \cb_6_4_io_eo[12] ,
    \cb_6_4_io_eo[11] ,
    \cb_6_4_io_eo[10] ,
    \cb_6_4_io_eo[9] ,
    \cb_6_4_io_eo[8] ,
    \cb_6_4_io_eo[7] ,
    \cb_6_4_io_eo[6] ,
    \cb_6_4_io_eo[5] ,
    \cb_6_4_io_eo[4] ,
    \cb_6_4_io_eo[3] ,
    \cb_6_4_io_eo[2] ,
    \cb_6_4_io_eo[1] ,
    \cb_6_4_io_eo[0] }));
 cic_block cb_6_6 (.io_cs_i(cb_6_6_io_cs_i),
    .io_i_0_ci(cb_6_5_io_o_0_co),
    .io_i_1_ci(cb_6_5_io_o_1_co),
    .io_i_2_ci(cb_6_5_io_o_2_co),
    .io_i_3_ci(cb_6_5_io_o_3_co),
    .io_i_4_ci(cb_6_5_io_o_4_co),
    .io_i_5_ci(cb_6_5_io_o_5_co),
    .io_i_6_ci(cb_6_5_io_o_6_co),
    .io_i_7_ci(cb_6_5_io_o_7_co),
    .io_o_0_co(cb_6_6_io_o_0_co),
    .io_o_1_co(cb_6_6_io_o_1_co),
    .io_o_2_co(cb_6_6_io_o_2_co),
    .io_o_3_co(cb_6_6_io_o_3_co),
    .io_o_4_co(cb_6_6_io_o_4_co),
    .io_o_5_co(cb_6_6_io_o_5_co),
    .io_o_6_co(cb_6_6_io_o_6_co),
    .io_o_7_co(cb_6_6_io_o_7_co),
    .io_vci(cb_6_5_io_vco),
    .io_vco(cb_6_6_io_vco),
    .io_vi(cb_6_6_io_vi),
    .io_we_i(cb_6_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_6_0_io_adr_i[1] ,
    \cb_6_0_io_adr_i[0] }),
    .io_dat_i({\cb_6_0_io_dat_i[15] ,
    \cb_6_0_io_dat_i[14] ,
    \cb_6_0_io_dat_i[13] ,
    \cb_6_0_io_dat_i[12] ,
    \cb_6_0_io_dat_i[11] ,
    \cb_6_0_io_dat_i[10] ,
    \cb_6_0_io_dat_i[9] ,
    \cb_6_0_io_dat_i[8] ,
    \cb_6_0_io_dat_i[7] ,
    \cb_6_0_io_dat_i[6] ,
    \cb_6_0_io_dat_i[5] ,
    \cb_6_0_io_dat_i[4] ,
    \cb_6_0_io_dat_i[3] ,
    \cb_6_0_io_dat_i[2] ,
    \cb_6_0_io_dat_i[1] ,
    \cb_6_0_io_dat_i[0] }),
    .io_dat_o({\cb_6_6_io_dat_o[15] ,
    \cb_6_6_io_dat_o[14] ,
    \cb_6_6_io_dat_o[13] ,
    \cb_6_6_io_dat_o[12] ,
    \cb_6_6_io_dat_o[11] ,
    \cb_6_6_io_dat_o[10] ,
    \cb_6_6_io_dat_o[9] ,
    \cb_6_6_io_dat_o[8] ,
    \cb_6_6_io_dat_o[7] ,
    \cb_6_6_io_dat_o[6] ,
    \cb_6_6_io_dat_o[5] ,
    \cb_6_6_io_dat_o[4] ,
    \cb_6_6_io_dat_o[3] ,
    \cb_6_6_io_dat_o[2] ,
    \cb_6_6_io_dat_o[1] ,
    \cb_6_6_io_dat_o[0] }),
    .io_eo({\cb_6_6_io_eo[63] ,
    \cb_6_6_io_eo[62] ,
    \cb_6_6_io_eo[61] ,
    \cb_6_6_io_eo[60] ,
    \cb_6_6_io_eo[59] ,
    \cb_6_6_io_eo[58] ,
    \cb_6_6_io_eo[57] ,
    \cb_6_6_io_eo[56] ,
    \cb_6_6_io_eo[55] ,
    \cb_6_6_io_eo[54] ,
    \cb_6_6_io_eo[53] ,
    \cb_6_6_io_eo[52] ,
    \cb_6_6_io_eo[51] ,
    \cb_6_6_io_eo[50] ,
    \cb_6_6_io_eo[49] ,
    \cb_6_6_io_eo[48] ,
    \cb_6_6_io_eo[47] ,
    \cb_6_6_io_eo[46] ,
    \cb_6_6_io_eo[45] ,
    \cb_6_6_io_eo[44] ,
    \cb_6_6_io_eo[43] ,
    \cb_6_6_io_eo[42] ,
    \cb_6_6_io_eo[41] ,
    \cb_6_6_io_eo[40] ,
    \cb_6_6_io_eo[39] ,
    \cb_6_6_io_eo[38] ,
    \cb_6_6_io_eo[37] ,
    \cb_6_6_io_eo[36] ,
    \cb_6_6_io_eo[35] ,
    \cb_6_6_io_eo[34] ,
    \cb_6_6_io_eo[33] ,
    \cb_6_6_io_eo[32] ,
    \cb_6_6_io_eo[31] ,
    \cb_6_6_io_eo[30] ,
    \cb_6_6_io_eo[29] ,
    \cb_6_6_io_eo[28] ,
    \cb_6_6_io_eo[27] ,
    \cb_6_6_io_eo[26] ,
    \cb_6_6_io_eo[25] ,
    \cb_6_6_io_eo[24] ,
    \cb_6_6_io_eo[23] ,
    \cb_6_6_io_eo[22] ,
    \cb_6_6_io_eo[21] ,
    \cb_6_6_io_eo[20] ,
    \cb_6_6_io_eo[19] ,
    \cb_6_6_io_eo[18] ,
    \cb_6_6_io_eo[17] ,
    \cb_6_6_io_eo[16] ,
    \cb_6_6_io_eo[15] ,
    \cb_6_6_io_eo[14] ,
    \cb_6_6_io_eo[13] ,
    \cb_6_6_io_eo[12] ,
    \cb_6_6_io_eo[11] ,
    \cb_6_6_io_eo[10] ,
    \cb_6_6_io_eo[9] ,
    \cb_6_6_io_eo[8] ,
    \cb_6_6_io_eo[7] ,
    \cb_6_6_io_eo[6] ,
    \cb_6_6_io_eo[5] ,
    \cb_6_6_io_eo[4] ,
    \cb_6_6_io_eo[3] ,
    \cb_6_6_io_eo[2] ,
    \cb_6_6_io_eo[1] ,
    \cb_6_6_io_eo[0] }),
    .io_i_0_in1({\cb_6_5_io_o_0_out[7] ,
    \cb_6_5_io_o_0_out[6] ,
    \cb_6_5_io_o_0_out[5] ,
    \cb_6_5_io_o_0_out[4] ,
    \cb_6_5_io_o_0_out[3] ,
    \cb_6_5_io_o_0_out[2] ,
    \cb_6_5_io_o_0_out[1] ,
    \cb_6_5_io_o_0_out[0] }),
    .io_i_1_in1({\cb_6_5_io_o_1_out[7] ,
    \cb_6_5_io_o_1_out[6] ,
    \cb_6_5_io_o_1_out[5] ,
    \cb_6_5_io_o_1_out[4] ,
    \cb_6_5_io_o_1_out[3] ,
    \cb_6_5_io_o_1_out[2] ,
    \cb_6_5_io_o_1_out[1] ,
    \cb_6_5_io_o_1_out[0] }),
    .io_i_2_in1({\cb_6_5_io_o_2_out[7] ,
    \cb_6_5_io_o_2_out[6] ,
    \cb_6_5_io_o_2_out[5] ,
    \cb_6_5_io_o_2_out[4] ,
    \cb_6_5_io_o_2_out[3] ,
    \cb_6_5_io_o_2_out[2] ,
    \cb_6_5_io_o_2_out[1] ,
    \cb_6_5_io_o_2_out[0] }),
    .io_i_3_in1({\cb_6_5_io_o_3_out[7] ,
    \cb_6_5_io_o_3_out[6] ,
    \cb_6_5_io_o_3_out[5] ,
    \cb_6_5_io_o_3_out[4] ,
    \cb_6_5_io_o_3_out[3] ,
    \cb_6_5_io_o_3_out[2] ,
    \cb_6_5_io_o_3_out[1] ,
    \cb_6_5_io_o_3_out[0] }),
    .io_i_4_in1({\cb_6_5_io_o_4_out[7] ,
    \cb_6_5_io_o_4_out[6] ,
    \cb_6_5_io_o_4_out[5] ,
    \cb_6_5_io_o_4_out[4] ,
    \cb_6_5_io_o_4_out[3] ,
    \cb_6_5_io_o_4_out[2] ,
    \cb_6_5_io_o_4_out[1] ,
    \cb_6_5_io_o_4_out[0] }),
    .io_i_5_in1({\cb_6_5_io_o_5_out[7] ,
    \cb_6_5_io_o_5_out[6] ,
    \cb_6_5_io_o_5_out[5] ,
    \cb_6_5_io_o_5_out[4] ,
    \cb_6_5_io_o_5_out[3] ,
    \cb_6_5_io_o_5_out[2] ,
    \cb_6_5_io_o_5_out[1] ,
    \cb_6_5_io_o_5_out[0] }),
    .io_i_6_in1({\cb_6_5_io_o_6_out[7] ,
    \cb_6_5_io_o_6_out[6] ,
    \cb_6_5_io_o_6_out[5] ,
    \cb_6_5_io_o_6_out[4] ,
    \cb_6_5_io_o_6_out[3] ,
    \cb_6_5_io_o_6_out[2] ,
    \cb_6_5_io_o_6_out[1] ,
    \cb_6_5_io_o_6_out[0] }),
    .io_i_7_in1({\cb_6_5_io_o_7_out[7] ,
    \cb_6_5_io_o_7_out[6] ,
    \cb_6_5_io_o_7_out[5] ,
    \cb_6_5_io_o_7_out[4] ,
    \cb_6_5_io_o_7_out[3] ,
    \cb_6_5_io_o_7_out[2] ,
    \cb_6_5_io_o_7_out[1] ,
    \cb_6_5_io_o_7_out[0] }),
    .io_o_0_out({\cb_6_6_io_o_0_out[7] ,
    \cb_6_6_io_o_0_out[6] ,
    \cb_6_6_io_o_0_out[5] ,
    \cb_6_6_io_o_0_out[4] ,
    \cb_6_6_io_o_0_out[3] ,
    \cb_6_6_io_o_0_out[2] ,
    \cb_6_6_io_o_0_out[1] ,
    \cb_6_6_io_o_0_out[0] }),
    .io_o_1_out({\cb_6_6_io_o_1_out[7] ,
    \cb_6_6_io_o_1_out[6] ,
    \cb_6_6_io_o_1_out[5] ,
    \cb_6_6_io_o_1_out[4] ,
    \cb_6_6_io_o_1_out[3] ,
    \cb_6_6_io_o_1_out[2] ,
    \cb_6_6_io_o_1_out[1] ,
    \cb_6_6_io_o_1_out[0] }),
    .io_o_2_out({\cb_6_6_io_o_2_out[7] ,
    \cb_6_6_io_o_2_out[6] ,
    \cb_6_6_io_o_2_out[5] ,
    \cb_6_6_io_o_2_out[4] ,
    \cb_6_6_io_o_2_out[3] ,
    \cb_6_6_io_o_2_out[2] ,
    \cb_6_6_io_o_2_out[1] ,
    \cb_6_6_io_o_2_out[0] }),
    .io_o_3_out({\cb_6_6_io_o_3_out[7] ,
    \cb_6_6_io_o_3_out[6] ,
    \cb_6_6_io_o_3_out[5] ,
    \cb_6_6_io_o_3_out[4] ,
    \cb_6_6_io_o_3_out[3] ,
    \cb_6_6_io_o_3_out[2] ,
    \cb_6_6_io_o_3_out[1] ,
    \cb_6_6_io_o_3_out[0] }),
    .io_o_4_out({\cb_6_6_io_o_4_out[7] ,
    \cb_6_6_io_o_4_out[6] ,
    \cb_6_6_io_o_4_out[5] ,
    \cb_6_6_io_o_4_out[4] ,
    \cb_6_6_io_o_4_out[3] ,
    \cb_6_6_io_o_4_out[2] ,
    \cb_6_6_io_o_4_out[1] ,
    \cb_6_6_io_o_4_out[0] }),
    .io_o_5_out({\cb_6_6_io_o_5_out[7] ,
    \cb_6_6_io_o_5_out[6] ,
    \cb_6_6_io_o_5_out[5] ,
    \cb_6_6_io_o_5_out[4] ,
    \cb_6_6_io_o_5_out[3] ,
    \cb_6_6_io_o_5_out[2] ,
    \cb_6_6_io_o_5_out[1] ,
    \cb_6_6_io_o_5_out[0] }),
    .io_o_6_out({\cb_6_6_io_o_6_out[7] ,
    \cb_6_6_io_o_6_out[6] ,
    \cb_6_6_io_o_6_out[5] ,
    \cb_6_6_io_o_6_out[4] ,
    \cb_6_6_io_o_6_out[3] ,
    \cb_6_6_io_o_6_out[2] ,
    \cb_6_6_io_o_6_out[1] ,
    \cb_6_6_io_o_6_out[0] }),
    .io_o_7_out({\cb_6_6_io_o_7_out[7] ,
    \cb_6_6_io_o_7_out[6] ,
    \cb_6_6_io_o_7_out[5] ,
    \cb_6_6_io_o_7_out[4] ,
    \cb_6_6_io_o_7_out[3] ,
    \cb_6_6_io_o_7_out[2] ,
    \cb_6_6_io_o_7_out[1] ,
    \cb_6_6_io_o_7_out[0] }),
    .io_wo({\cb_6_5_io_eo[63] ,
    \cb_6_5_io_eo[62] ,
    \cb_6_5_io_eo[61] ,
    \cb_6_5_io_eo[60] ,
    \cb_6_5_io_eo[59] ,
    \cb_6_5_io_eo[58] ,
    \cb_6_5_io_eo[57] ,
    \cb_6_5_io_eo[56] ,
    \cb_6_5_io_eo[55] ,
    \cb_6_5_io_eo[54] ,
    \cb_6_5_io_eo[53] ,
    \cb_6_5_io_eo[52] ,
    \cb_6_5_io_eo[51] ,
    \cb_6_5_io_eo[50] ,
    \cb_6_5_io_eo[49] ,
    \cb_6_5_io_eo[48] ,
    \cb_6_5_io_eo[47] ,
    \cb_6_5_io_eo[46] ,
    \cb_6_5_io_eo[45] ,
    \cb_6_5_io_eo[44] ,
    \cb_6_5_io_eo[43] ,
    \cb_6_5_io_eo[42] ,
    \cb_6_5_io_eo[41] ,
    \cb_6_5_io_eo[40] ,
    \cb_6_5_io_eo[39] ,
    \cb_6_5_io_eo[38] ,
    \cb_6_5_io_eo[37] ,
    \cb_6_5_io_eo[36] ,
    \cb_6_5_io_eo[35] ,
    \cb_6_5_io_eo[34] ,
    \cb_6_5_io_eo[33] ,
    \cb_6_5_io_eo[32] ,
    \cb_6_5_io_eo[31] ,
    \cb_6_5_io_eo[30] ,
    \cb_6_5_io_eo[29] ,
    \cb_6_5_io_eo[28] ,
    \cb_6_5_io_eo[27] ,
    \cb_6_5_io_eo[26] ,
    \cb_6_5_io_eo[25] ,
    \cb_6_5_io_eo[24] ,
    \cb_6_5_io_eo[23] ,
    \cb_6_5_io_eo[22] ,
    \cb_6_5_io_eo[21] ,
    \cb_6_5_io_eo[20] ,
    \cb_6_5_io_eo[19] ,
    \cb_6_5_io_eo[18] ,
    \cb_6_5_io_eo[17] ,
    \cb_6_5_io_eo[16] ,
    \cb_6_5_io_eo[15] ,
    \cb_6_5_io_eo[14] ,
    \cb_6_5_io_eo[13] ,
    \cb_6_5_io_eo[12] ,
    \cb_6_5_io_eo[11] ,
    \cb_6_5_io_eo[10] ,
    \cb_6_5_io_eo[9] ,
    \cb_6_5_io_eo[8] ,
    \cb_6_5_io_eo[7] ,
    \cb_6_5_io_eo[6] ,
    \cb_6_5_io_eo[5] ,
    \cb_6_5_io_eo[4] ,
    \cb_6_5_io_eo[3] ,
    \cb_6_5_io_eo[2] ,
    \cb_6_5_io_eo[1] ,
    \cb_6_5_io_eo[0] }));
 cic_block cb_6_7 (.io_cs_i(cb_6_7_io_cs_i),
    .io_i_0_ci(cb_6_6_io_o_0_co),
    .io_i_1_ci(cb_6_6_io_o_1_co),
    .io_i_2_ci(cb_6_6_io_o_2_co),
    .io_i_3_ci(cb_6_6_io_o_3_co),
    .io_i_4_ci(cb_6_6_io_o_4_co),
    .io_i_5_ci(cb_6_6_io_o_5_co),
    .io_i_6_ci(cb_6_6_io_o_6_co),
    .io_i_7_ci(cb_6_6_io_o_7_co),
    .io_o_0_co(cb_6_7_io_o_0_co),
    .io_o_1_co(cb_6_7_io_o_1_co),
    .io_o_2_co(cb_6_7_io_o_2_co),
    .io_o_3_co(cb_6_7_io_o_3_co),
    .io_o_4_co(cb_6_7_io_o_4_co),
    .io_o_5_co(cb_6_7_io_o_5_co),
    .io_o_6_co(cb_6_7_io_o_6_co),
    .io_o_7_co(cb_6_7_io_o_7_co),
    .io_vci(cb_6_6_io_vco),
    .io_vco(cb_6_7_io_vco),
    .io_vi(cb_6_7_io_vi),
    .io_we_i(cb_6_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_6_0_io_adr_i[1] ,
    \cb_6_0_io_adr_i[0] }),
    .io_dat_i({\cb_6_0_io_dat_i[15] ,
    \cb_6_0_io_dat_i[14] ,
    \cb_6_0_io_dat_i[13] ,
    \cb_6_0_io_dat_i[12] ,
    \cb_6_0_io_dat_i[11] ,
    \cb_6_0_io_dat_i[10] ,
    \cb_6_0_io_dat_i[9] ,
    \cb_6_0_io_dat_i[8] ,
    \cb_6_0_io_dat_i[7] ,
    \cb_6_0_io_dat_i[6] ,
    \cb_6_0_io_dat_i[5] ,
    \cb_6_0_io_dat_i[4] ,
    \cb_6_0_io_dat_i[3] ,
    \cb_6_0_io_dat_i[2] ,
    \cb_6_0_io_dat_i[1] ,
    \cb_6_0_io_dat_i[0] }),
    .io_dat_o({\cb_6_7_io_dat_o[15] ,
    \cb_6_7_io_dat_o[14] ,
    \cb_6_7_io_dat_o[13] ,
    \cb_6_7_io_dat_o[12] ,
    \cb_6_7_io_dat_o[11] ,
    \cb_6_7_io_dat_o[10] ,
    \cb_6_7_io_dat_o[9] ,
    \cb_6_7_io_dat_o[8] ,
    \cb_6_7_io_dat_o[7] ,
    \cb_6_7_io_dat_o[6] ,
    \cb_6_7_io_dat_o[5] ,
    \cb_6_7_io_dat_o[4] ,
    \cb_6_7_io_dat_o[3] ,
    \cb_6_7_io_dat_o[2] ,
    \cb_6_7_io_dat_o[1] ,
    \cb_6_7_io_dat_o[0] }),
    .io_eo({\cb_6_7_io_eo[63] ,
    \cb_6_7_io_eo[62] ,
    \cb_6_7_io_eo[61] ,
    \cb_6_7_io_eo[60] ,
    \cb_6_7_io_eo[59] ,
    \cb_6_7_io_eo[58] ,
    \cb_6_7_io_eo[57] ,
    \cb_6_7_io_eo[56] ,
    \cb_6_7_io_eo[55] ,
    \cb_6_7_io_eo[54] ,
    \cb_6_7_io_eo[53] ,
    \cb_6_7_io_eo[52] ,
    \cb_6_7_io_eo[51] ,
    \cb_6_7_io_eo[50] ,
    \cb_6_7_io_eo[49] ,
    \cb_6_7_io_eo[48] ,
    \cb_6_7_io_eo[47] ,
    \cb_6_7_io_eo[46] ,
    \cb_6_7_io_eo[45] ,
    \cb_6_7_io_eo[44] ,
    \cb_6_7_io_eo[43] ,
    \cb_6_7_io_eo[42] ,
    \cb_6_7_io_eo[41] ,
    \cb_6_7_io_eo[40] ,
    \cb_6_7_io_eo[39] ,
    \cb_6_7_io_eo[38] ,
    \cb_6_7_io_eo[37] ,
    \cb_6_7_io_eo[36] ,
    \cb_6_7_io_eo[35] ,
    \cb_6_7_io_eo[34] ,
    \cb_6_7_io_eo[33] ,
    \cb_6_7_io_eo[32] ,
    \cb_6_7_io_eo[31] ,
    \cb_6_7_io_eo[30] ,
    \cb_6_7_io_eo[29] ,
    \cb_6_7_io_eo[28] ,
    \cb_6_7_io_eo[27] ,
    \cb_6_7_io_eo[26] ,
    \cb_6_7_io_eo[25] ,
    \cb_6_7_io_eo[24] ,
    \cb_6_7_io_eo[23] ,
    \cb_6_7_io_eo[22] ,
    \cb_6_7_io_eo[21] ,
    \cb_6_7_io_eo[20] ,
    \cb_6_7_io_eo[19] ,
    \cb_6_7_io_eo[18] ,
    \cb_6_7_io_eo[17] ,
    \cb_6_7_io_eo[16] ,
    \cb_6_7_io_eo[15] ,
    \cb_6_7_io_eo[14] ,
    \cb_6_7_io_eo[13] ,
    \cb_6_7_io_eo[12] ,
    \cb_6_7_io_eo[11] ,
    \cb_6_7_io_eo[10] ,
    \cb_6_7_io_eo[9] ,
    \cb_6_7_io_eo[8] ,
    \cb_6_7_io_eo[7] ,
    \cb_6_7_io_eo[6] ,
    \cb_6_7_io_eo[5] ,
    \cb_6_7_io_eo[4] ,
    \cb_6_7_io_eo[3] ,
    \cb_6_7_io_eo[2] ,
    \cb_6_7_io_eo[1] ,
    \cb_6_7_io_eo[0] }),
    .io_i_0_in1({\cb_6_6_io_o_0_out[7] ,
    \cb_6_6_io_o_0_out[6] ,
    \cb_6_6_io_o_0_out[5] ,
    \cb_6_6_io_o_0_out[4] ,
    \cb_6_6_io_o_0_out[3] ,
    \cb_6_6_io_o_0_out[2] ,
    \cb_6_6_io_o_0_out[1] ,
    \cb_6_6_io_o_0_out[0] }),
    .io_i_1_in1({\cb_6_6_io_o_1_out[7] ,
    \cb_6_6_io_o_1_out[6] ,
    \cb_6_6_io_o_1_out[5] ,
    \cb_6_6_io_o_1_out[4] ,
    \cb_6_6_io_o_1_out[3] ,
    \cb_6_6_io_o_1_out[2] ,
    \cb_6_6_io_o_1_out[1] ,
    \cb_6_6_io_o_1_out[0] }),
    .io_i_2_in1({\cb_6_6_io_o_2_out[7] ,
    \cb_6_6_io_o_2_out[6] ,
    \cb_6_6_io_o_2_out[5] ,
    \cb_6_6_io_o_2_out[4] ,
    \cb_6_6_io_o_2_out[3] ,
    \cb_6_6_io_o_2_out[2] ,
    \cb_6_6_io_o_2_out[1] ,
    \cb_6_6_io_o_2_out[0] }),
    .io_i_3_in1({\cb_6_6_io_o_3_out[7] ,
    \cb_6_6_io_o_3_out[6] ,
    \cb_6_6_io_o_3_out[5] ,
    \cb_6_6_io_o_3_out[4] ,
    \cb_6_6_io_o_3_out[3] ,
    \cb_6_6_io_o_3_out[2] ,
    \cb_6_6_io_o_3_out[1] ,
    \cb_6_6_io_o_3_out[0] }),
    .io_i_4_in1({\cb_6_6_io_o_4_out[7] ,
    \cb_6_6_io_o_4_out[6] ,
    \cb_6_6_io_o_4_out[5] ,
    \cb_6_6_io_o_4_out[4] ,
    \cb_6_6_io_o_4_out[3] ,
    \cb_6_6_io_o_4_out[2] ,
    \cb_6_6_io_o_4_out[1] ,
    \cb_6_6_io_o_4_out[0] }),
    .io_i_5_in1({\cb_6_6_io_o_5_out[7] ,
    \cb_6_6_io_o_5_out[6] ,
    \cb_6_6_io_o_5_out[5] ,
    \cb_6_6_io_o_5_out[4] ,
    \cb_6_6_io_o_5_out[3] ,
    \cb_6_6_io_o_5_out[2] ,
    \cb_6_6_io_o_5_out[1] ,
    \cb_6_6_io_o_5_out[0] }),
    .io_i_6_in1({\cb_6_6_io_o_6_out[7] ,
    \cb_6_6_io_o_6_out[6] ,
    \cb_6_6_io_o_6_out[5] ,
    \cb_6_6_io_o_6_out[4] ,
    \cb_6_6_io_o_6_out[3] ,
    \cb_6_6_io_o_6_out[2] ,
    \cb_6_6_io_o_6_out[1] ,
    \cb_6_6_io_o_6_out[0] }),
    .io_i_7_in1({\cb_6_6_io_o_7_out[7] ,
    \cb_6_6_io_o_7_out[6] ,
    \cb_6_6_io_o_7_out[5] ,
    \cb_6_6_io_o_7_out[4] ,
    \cb_6_6_io_o_7_out[3] ,
    \cb_6_6_io_o_7_out[2] ,
    \cb_6_6_io_o_7_out[1] ,
    \cb_6_6_io_o_7_out[0] }),
    .io_o_0_out({\cb_6_7_io_o_0_out[7] ,
    \cb_6_7_io_o_0_out[6] ,
    \cb_6_7_io_o_0_out[5] ,
    \cb_6_7_io_o_0_out[4] ,
    \cb_6_7_io_o_0_out[3] ,
    \cb_6_7_io_o_0_out[2] ,
    \cb_6_7_io_o_0_out[1] ,
    \cb_6_7_io_o_0_out[0] }),
    .io_o_1_out({\cb_6_7_io_o_1_out[7] ,
    \cb_6_7_io_o_1_out[6] ,
    \cb_6_7_io_o_1_out[5] ,
    \cb_6_7_io_o_1_out[4] ,
    \cb_6_7_io_o_1_out[3] ,
    \cb_6_7_io_o_1_out[2] ,
    \cb_6_7_io_o_1_out[1] ,
    \cb_6_7_io_o_1_out[0] }),
    .io_o_2_out({\cb_6_7_io_o_2_out[7] ,
    \cb_6_7_io_o_2_out[6] ,
    \cb_6_7_io_o_2_out[5] ,
    \cb_6_7_io_o_2_out[4] ,
    \cb_6_7_io_o_2_out[3] ,
    \cb_6_7_io_o_2_out[2] ,
    \cb_6_7_io_o_2_out[1] ,
    \cb_6_7_io_o_2_out[0] }),
    .io_o_3_out({\cb_6_7_io_o_3_out[7] ,
    \cb_6_7_io_o_3_out[6] ,
    \cb_6_7_io_o_3_out[5] ,
    \cb_6_7_io_o_3_out[4] ,
    \cb_6_7_io_o_3_out[3] ,
    \cb_6_7_io_o_3_out[2] ,
    \cb_6_7_io_o_3_out[1] ,
    \cb_6_7_io_o_3_out[0] }),
    .io_o_4_out({\cb_6_7_io_o_4_out[7] ,
    \cb_6_7_io_o_4_out[6] ,
    \cb_6_7_io_o_4_out[5] ,
    \cb_6_7_io_o_4_out[4] ,
    \cb_6_7_io_o_4_out[3] ,
    \cb_6_7_io_o_4_out[2] ,
    \cb_6_7_io_o_4_out[1] ,
    \cb_6_7_io_o_4_out[0] }),
    .io_o_5_out({\cb_6_7_io_o_5_out[7] ,
    \cb_6_7_io_o_5_out[6] ,
    \cb_6_7_io_o_5_out[5] ,
    \cb_6_7_io_o_5_out[4] ,
    \cb_6_7_io_o_5_out[3] ,
    \cb_6_7_io_o_5_out[2] ,
    \cb_6_7_io_o_5_out[1] ,
    \cb_6_7_io_o_5_out[0] }),
    .io_o_6_out({\cb_6_7_io_o_6_out[7] ,
    \cb_6_7_io_o_6_out[6] ,
    \cb_6_7_io_o_6_out[5] ,
    \cb_6_7_io_o_6_out[4] ,
    \cb_6_7_io_o_6_out[3] ,
    \cb_6_7_io_o_6_out[2] ,
    \cb_6_7_io_o_6_out[1] ,
    \cb_6_7_io_o_6_out[0] }),
    .io_o_7_out({\cb_6_7_io_o_7_out[7] ,
    \cb_6_7_io_o_7_out[6] ,
    \cb_6_7_io_o_7_out[5] ,
    \cb_6_7_io_o_7_out[4] ,
    \cb_6_7_io_o_7_out[3] ,
    \cb_6_7_io_o_7_out[2] ,
    \cb_6_7_io_o_7_out[1] ,
    \cb_6_7_io_o_7_out[0] }),
    .io_wo({\cb_6_6_io_eo[63] ,
    \cb_6_6_io_eo[62] ,
    \cb_6_6_io_eo[61] ,
    \cb_6_6_io_eo[60] ,
    \cb_6_6_io_eo[59] ,
    \cb_6_6_io_eo[58] ,
    \cb_6_6_io_eo[57] ,
    \cb_6_6_io_eo[56] ,
    \cb_6_6_io_eo[55] ,
    \cb_6_6_io_eo[54] ,
    \cb_6_6_io_eo[53] ,
    \cb_6_6_io_eo[52] ,
    \cb_6_6_io_eo[51] ,
    \cb_6_6_io_eo[50] ,
    \cb_6_6_io_eo[49] ,
    \cb_6_6_io_eo[48] ,
    \cb_6_6_io_eo[47] ,
    \cb_6_6_io_eo[46] ,
    \cb_6_6_io_eo[45] ,
    \cb_6_6_io_eo[44] ,
    \cb_6_6_io_eo[43] ,
    \cb_6_6_io_eo[42] ,
    \cb_6_6_io_eo[41] ,
    \cb_6_6_io_eo[40] ,
    \cb_6_6_io_eo[39] ,
    \cb_6_6_io_eo[38] ,
    \cb_6_6_io_eo[37] ,
    \cb_6_6_io_eo[36] ,
    \cb_6_6_io_eo[35] ,
    \cb_6_6_io_eo[34] ,
    \cb_6_6_io_eo[33] ,
    \cb_6_6_io_eo[32] ,
    \cb_6_6_io_eo[31] ,
    \cb_6_6_io_eo[30] ,
    \cb_6_6_io_eo[29] ,
    \cb_6_6_io_eo[28] ,
    \cb_6_6_io_eo[27] ,
    \cb_6_6_io_eo[26] ,
    \cb_6_6_io_eo[25] ,
    \cb_6_6_io_eo[24] ,
    \cb_6_6_io_eo[23] ,
    \cb_6_6_io_eo[22] ,
    \cb_6_6_io_eo[21] ,
    \cb_6_6_io_eo[20] ,
    \cb_6_6_io_eo[19] ,
    \cb_6_6_io_eo[18] ,
    \cb_6_6_io_eo[17] ,
    \cb_6_6_io_eo[16] ,
    \cb_6_6_io_eo[15] ,
    \cb_6_6_io_eo[14] ,
    \cb_6_6_io_eo[13] ,
    \cb_6_6_io_eo[12] ,
    \cb_6_6_io_eo[11] ,
    \cb_6_6_io_eo[10] ,
    \cb_6_6_io_eo[9] ,
    \cb_6_6_io_eo[8] ,
    \cb_6_6_io_eo[7] ,
    \cb_6_6_io_eo[6] ,
    \cb_6_6_io_eo[5] ,
    \cb_6_6_io_eo[4] ,
    \cb_6_6_io_eo[3] ,
    \cb_6_6_io_eo[2] ,
    \cb_6_6_io_eo[1] ,
    \cb_6_6_io_eo[0] }));
 cic_block cb_6_8 (.io_cs_i(cb_6_8_io_cs_i),
    .io_i_0_ci(cb_6_7_io_o_0_co),
    .io_i_1_ci(cb_6_7_io_o_1_co),
    .io_i_2_ci(cb_6_7_io_o_2_co),
    .io_i_3_ci(cb_6_7_io_o_3_co),
    .io_i_4_ci(cb_6_7_io_o_4_co),
    .io_i_5_ci(cb_6_7_io_o_5_co),
    .io_i_6_ci(cb_6_7_io_o_6_co),
    .io_i_7_ci(cb_6_7_io_o_7_co),
    .io_o_0_co(cb_6_8_io_o_0_co),
    .io_o_1_co(cb_6_8_io_o_1_co),
    .io_o_2_co(cb_6_8_io_o_2_co),
    .io_o_3_co(cb_6_8_io_o_3_co),
    .io_o_4_co(cb_6_8_io_o_4_co),
    .io_o_5_co(cb_6_8_io_o_5_co),
    .io_o_6_co(cb_6_8_io_o_6_co),
    .io_o_7_co(cb_6_8_io_o_7_co),
    .io_vci(cb_6_7_io_vco),
    .io_vco(cb_6_8_io_vco),
    .io_vi(cb_6_8_io_vi),
    .io_we_i(cb_6_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_6_0_io_adr_i[1] ,
    \cb_6_0_io_adr_i[0] }),
    .io_dat_i({\cb_6_0_io_dat_i[15] ,
    \cb_6_0_io_dat_i[14] ,
    \cb_6_0_io_dat_i[13] ,
    \cb_6_0_io_dat_i[12] ,
    \cb_6_0_io_dat_i[11] ,
    \cb_6_0_io_dat_i[10] ,
    \cb_6_0_io_dat_i[9] ,
    \cb_6_0_io_dat_i[8] ,
    \cb_6_0_io_dat_i[7] ,
    \cb_6_0_io_dat_i[6] ,
    \cb_6_0_io_dat_i[5] ,
    \cb_6_0_io_dat_i[4] ,
    \cb_6_0_io_dat_i[3] ,
    \cb_6_0_io_dat_i[2] ,
    \cb_6_0_io_dat_i[1] ,
    \cb_6_0_io_dat_i[0] }),
    .io_dat_o({\cb_6_8_io_dat_o[15] ,
    \cb_6_8_io_dat_o[14] ,
    \cb_6_8_io_dat_o[13] ,
    \cb_6_8_io_dat_o[12] ,
    \cb_6_8_io_dat_o[11] ,
    \cb_6_8_io_dat_o[10] ,
    \cb_6_8_io_dat_o[9] ,
    \cb_6_8_io_dat_o[8] ,
    \cb_6_8_io_dat_o[7] ,
    \cb_6_8_io_dat_o[6] ,
    \cb_6_8_io_dat_o[5] ,
    \cb_6_8_io_dat_o[4] ,
    \cb_6_8_io_dat_o[3] ,
    \cb_6_8_io_dat_o[2] ,
    \cb_6_8_io_dat_o[1] ,
    \cb_6_8_io_dat_o[0] }),
    .io_eo({\cb_6_8_io_eo[63] ,
    \cb_6_8_io_eo[62] ,
    \cb_6_8_io_eo[61] ,
    \cb_6_8_io_eo[60] ,
    \cb_6_8_io_eo[59] ,
    \cb_6_8_io_eo[58] ,
    \cb_6_8_io_eo[57] ,
    \cb_6_8_io_eo[56] ,
    \cb_6_8_io_eo[55] ,
    \cb_6_8_io_eo[54] ,
    \cb_6_8_io_eo[53] ,
    \cb_6_8_io_eo[52] ,
    \cb_6_8_io_eo[51] ,
    \cb_6_8_io_eo[50] ,
    \cb_6_8_io_eo[49] ,
    \cb_6_8_io_eo[48] ,
    \cb_6_8_io_eo[47] ,
    \cb_6_8_io_eo[46] ,
    \cb_6_8_io_eo[45] ,
    \cb_6_8_io_eo[44] ,
    \cb_6_8_io_eo[43] ,
    \cb_6_8_io_eo[42] ,
    \cb_6_8_io_eo[41] ,
    \cb_6_8_io_eo[40] ,
    \cb_6_8_io_eo[39] ,
    \cb_6_8_io_eo[38] ,
    \cb_6_8_io_eo[37] ,
    \cb_6_8_io_eo[36] ,
    \cb_6_8_io_eo[35] ,
    \cb_6_8_io_eo[34] ,
    \cb_6_8_io_eo[33] ,
    \cb_6_8_io_eo[32] ,
    \cb_6_8_io_eo[31] ,
    \cb_6_8_io_eo[30] ,
    \cb_6_8_io_eo[29] ,
    \cb_6_8_io_eo[28] ,
    \cb_6_8_io_eo[27] ,
    \cb_6_8_io_eo[26] ,
    \cb_6_8_io_eo[25] ,
    \cb_6_8_io_eo[24] ,
    \cb_6_8_io_eo[23] ,
    \cb_6_8_io_eo[22] ,
    \cb_6_8_io_eo[21] ,
    \cb_6_8_io_eo[20] ,
    \cb_6_8_io_eo[19] ,
    \cb_6_8_io_eo[18] ,
    \cb_6_8_io_eo[17] ,
    \cb_6_8_io_eo[16] ,
    \cb_6_8_io_eo[15] ,
    \cb_6_8_io_eo[14] ,
    \cb_6_8_io_eo[13] ,
    \cb_6_8_io_eo[12] ,
    \cb_6_8_io_eo[11] ,
    \cb_6_8_io_eo[10] ,
    \cb_6_8_io_eo[9] ,
    \cb_6_8_io_eo[8] ,
    \cb_6_8_io_eo[7] ,
    \cb_6_8_io_eo[6] ,
    \cb_6_8_io_eo[5] ,
    \cb_6_8_io_eo[4] ,
    \cb_6_8_io_eo[3] ,
    \cb_6_8_io_eo[2] ,
    \cb_6_8_io_eo[1] ,
    \cb_6_8_io_eo[0] }),
    .io_i_0_in1({\cb_6_7_io_o_0_out[7] ,
    \cb_6_7_io_o_0_out[6] ,
    \cb_6_7_io_o_0_out[5] ,
    \cb_6_7_io_o_0_out[4] ,
    \cb_6_7_io_o_0_out[3] ,
    \cb_6_7_io_o_0_out[2] ,
    \cb_6_7_io_o_0_out[1] ,
    \cb_6_7_io_o_0_out[0] }),
    .io_i_1_in1({\cb_6_7_io_o_1_out[7] ,
    \cb_6_7_io_o_1_out[6] ,
    \cb_6_7_io_o_1_out[5] ,
    \cb_6_7_io_o_1_out[4] ,
    \cb_6_7_io_o_1_out[3] ,
    \cb_6_7_io_o_1_out[2] ,
    \cb_6_7_io_o_1_out[1] ,
    \cb_6_7_io_o_1_out[0] }),
    .io_i_2_in1({\cb_6_7_io_o_2_out[7] ,
    \cb_6_7_io_o_2_out[6] ,
    \cb_6_7_io_o_2_out[5] ,
    \cb_6_7_io_o_2_out[4] ,
    \cb_6_7_io_o_2_out[3] ,
    \cb_6_7_io_o_2_out[2] ,
    \cb_6_7_io_o_2_out[1] ,
    \cb_6_7_io_o_2_out[0] }),
    .io_i_3_in1({\cb_6_7_io_o_3_out[7] ,
    \cb_6_7_io_o_3_out[6] ,
    \cb_6_7_io_o_3_out[5] ,
    \cb_6_7_io_o_3_out[4] ,
    \cb_6_7_io_o_3_out[3] ,
    \cb_6_7_io_o_3_out[2] ,
    \cb_6_7_io_o_3_out[1] ,
    \cb_6_7_io_o_3_out[0] }),
    .io_i_4_in1({\cb_6_7_io_o_4_out[7] ,
    \cb_6_7_io_o_4_out[6] ,
    \cb_6_7_io_o_4_out[5] ,
    \cb_6_7_io_o_4_out[4] ,
    \cb_6_7_io_o_4_out[3] ,
    \cb_6_7_io_o_4_out[2] ,
    \cb_6_7_io_o_4_out[1] ,
    \cb_6_7_io_o_4_out[0] }),
    .io_i_5_in1({\cb_6_7_io_o_5_out[7] ,
    \cb_6_7_io_o_5_out[6] ,
    \cb_6_7_io_o_5_out[5] ,
    \cb_6_7_io_o_5_out[4] ,
    \cb_6_7_io_o_5_out[3] ,
    \cb_6_7_io_o_5_out[2] ,
    \cb_6_7_io_o_5_out[1] ,
    \cb_6_7_io_o_5_out[0] }),
    .io_i_6_in1({\cb_6_7_io_o_6_out[7] ,
    \cb_6_7_io_o_6_out[6] ,
    \cb_6_7_io_o_6_out[5] ,
    \cb_6_7_io_o_6_out[4] ,
    \cb_6_7_io_o_6_out[3] ,
    \cb_6_7_io_o_6_out[2] ,
    \cb_6_7_io_o_6_out[1] ,
    \cb_6_7_io_o_6_out[0] }),
    .io_i_7_in1({\cb_6_7_io_o_7_out[7] ,
    \cb_6_7_io_o_7_out[6] ,
    \cb_6_7_io_o_7_out[5] ,
    \cb_6_7_io_o_7_out[4] ,
    \cb_6_7_io_o_7_out[3] ,
    \cb_6_7_io_o_7_out[2] ,
    \cb_6_7_io_o_7_out[1] ,
    \cb_6_7_io_o_7_out[0] }),
    .io_o_0_out({\cb_6_8_io_o_0_out[7] ,
    \cb_6_8_io_o_0_out[6] ,
    \cb_6_8_io_o_0_out[5] ,
    \cb_6_8_io_o_0_out[4] ,
    \cb_6_8_io_o_0_out[3] ,
    \cb_6_8_io_o_0_out[2] ,
    \cb_6_8_io_o_0_out[1] ,
    \cb_6_8_io_o_0_out[0] }),
    .io_o_1_out({\cb_6_8_io_o_1_out[7] ,
    \cb_6_8_io_o_1_out[6] ,
    \cb_6_8_io_o_1_out[5] ,
    \cb_6_8_io_o_1_out[4] ,
    \cb_6_8_io_o_1_out[3] ,
    \cb_6_8_io_o_1_out[2] ,
    \cb_6_8_io_o_1_out[1] ,
    \cb_6_8_io_o_1_out[0] }),
    .io_o_2_out({\cb_6_8_io_o_2_out[7] ,
    \cb_6_8_io_o_2_out[6] ,
    \cb_6_8_io_o_2_out[5] ,
    \cb_6_8_io_o_2_out[4] ,
    \cb_6_8_io_o_2_out[3] ,
    \cb_6_8_io_o_2_out[2] ,
    \cb_6_8_io_o_2_out[1] ,
    \cb_6_8_io_o_2_out[0] }),
    .io_o_3_out({\cb_6_8_io_o_3_out[7] ,
    \cb_6_8_io_o_3_out[6] ,
    \cb_6_8_io_o_3_out[5] ,
    \cb_6_8_io_o_3_out[4] ,
    \cb_6_8_io_o_3_out[3] ,
    \cb_6_8_io_o_3_out[2] ,
    \cb_6_8_io_o_3_out[1] ,
    \cb_6_8_io_o_3_out[0] }),
    .io_o_4_out({\cb_6_8_io_o_4_out[7] ,
    \cb_6_8_io_o_4_out[6] ,
    \cb_6_8_io_o_4_out[5] ,
    \cb_6_8_io_o_4_out[4] ,
    \cb_6_8_io_o_4_out[3] ,
    \cb_6_8_io_o_4_out[2] ,
    \cb_6_8_io_o_4_out[1] ,
    \cb_6_8_io_o_4_out[0] }),
    .io_o_5_out({\cb_6_8_io_o_5_out[7] ,
    \cb_6_8_io_o_5_out[6] ,
    \cb_6_8_io_o_5_out[5] ,
    \cb_6_8_io_o_5_out[4] ,
    \cb_6_8_io_o_5_out[3] ,
    \cb_6_8_io_o_5_out[2] ,
    \cb_6_8_io_o_5_out[1] ,
    \cb_6_8_io_o_5_out[0] }),
    .io_o_6_out({\cb_6_8_io_o_6_out[7] ,
    \cb_6_8_io_o_6_out[6] ,
    \cb_6_8_io_o_6_out[5] ,
    \cb_6_8_io_o_6_out[4] ,
    \cb_6_8_io_o_6_out[3] ,
    \cb_6_8_io_o_6_out[2] ,
    \cb_6_8_io_o_6_out[1] ,
    \cb_6_8_io_o_6_out[0] }),
    .io_o_7_out({\cb_6_8_io_o_7_out[7] ,
    \cb_6_8_io_o_7_out[6] ,
    \cb_6_8_io_o_7_out[5] ,
    \cb_6_8_io_o_7_out[4] ,
    \cb_6_8_io_o_7_out[3] ,
    \cb_6_8_io_o_7_out[2] ,
    \cb_6_8_io_o_7_out[1] ,
    \cb_6_8_io_o_7_out[0] }),
    .io_wo({\cb_6_7_io_eo[63] ,
    \cb_6_7_io_eo[62] ,
    \cb_6_7_io_eo[61] ,
    \cb_6_7_io_eo[60] ,
    \cb_6_7_io_eo[59] ,
    \cb_6_7_io_eo[58] ,
    \cb_6_7_io_eo[57] ,
    \cb_6_7_io_eo[56] ,
    \cb_6_7_io_eo[55] ,
    \cb_6_7_io_eo[54] ,
    \cb_6_7_io_eo[53] ,
    \cb_6_7_io_eo[52] ,
    \cb_6_7_io_eo[51] ,
    \cb_6_7_io_eo[50] ,
    \cb_6_7_io_eo[49] ,
    \cb_6_7_io_eo[48] ,
    \cb_6_7_io_eo[47] ,
    \cb_6_7_io_eo[46] ,
    \cb_6_7_io_eo[45] ,
    \cb_6_7_io_eo[44] ,
    \cb_6_7_io_eo[43] ,
    \cb_6_7_io_eo[42] ,
    \cb_6_7_io_eo[41] ,
    \cb_6_7_io_eo[40] ,
    \cb_6_7_io_eo[39] ,
    \cb_6_7_io_eo[38] ,
    \cb_6_7_io_eo[37] ,
    \cb_6_7_io_eo[36] ,
    \cb_6_7_io_eo[35] ,
    \cb_6_7_io_eo[34] ,
    \cb_6_7_io_eo[33] ,
    \cb_6_7_io_eo[32] ,
    \cb_6_7_io_eo[31] ,
    \cb_6_7_io_eo[30] ,
    \cb_6_7_io_eo[29] ,
    \cb_6_7_io_eo[28] ,
    \cb_6_7_io_eo[27] ,
    \cb_6_7_io_eo[26] ,
    \cb_6_7_io_eo[25] ,
    \cb_6_7_io_eo[24] ,
    \cb_6_7_io_eo[23] ,
    \cb_6_7_io_eo[22] ,
    \cb_6_7_io_eo[21] ,
    \cb_6_7_io_eo[20] ,
    \cb_6_7_io_eo[19] ,
    \cb_6_7_io_eo[18] ,
    \cb_6_7_io_eo[17] ,
    \cb_6_7_io_eo[16] ,
    \cb_6_7_io_eo[15] ,
    \cb_6_7_io_eo[14] ,
    \cb_6_7_io_eo[13] ,
    \cb_6_7_io_eo[12] ,
    \cb_6_7_io_eo[11] ,
    \cb_6_7_io_eo[10] ,
    \cb_6_7_io_eo[9] ,
    \cb_6_7_io_eo[8] ,
    \cb_6_7_io_eo[7] ,
    \cb_6_7_io_eo[6] ,
    \cb_6_7_io_eo[5] ,
    \cb_6_7_io_eo[4] ,
    \cb_6_7_io_eo[3] ,
    \cb_6_7_io_eo[2] ,
    \cb_6_7_io_eo[1] ,
    \cb_6_7_io_eo[0] }));
 cic_block cb_6_9 (.io_cs_i(cb_6_9_io_cs_i),
    .io_i_0_ci(cb_6_8_io_o_0_co),
    .io_i_1_ci(cb_6_8_io_o_1_co),
    .io_i_2_ci(cb_6_8_io_o_2_co),
    .io_i_3_ci(cb_6_8_io_o_3_co),
    .io_i_4_ci(cb_6_8_io_o_4_co),
    .io_i_5_ci(cb_6_8_io_o_5_co),
    .io_i_6_ci(cb_6_8_io_o_6_co),
    .io_i_7_ci(cb_6_8_io_o_7_co),
    .io_o_0_co(cb_6_10_io_i_0_ci),
    .io_o_1_co(cb_6_10_io_i_1_ci),
    .io_o_2_co(cb_6_10_io_i_2_ci),
    .io_o_3_co(cb_6_10_io_i_3_ci),
    .io_o_4_co(cb_6_10_io_i_4_ci),
    .io_o_5_co(cb_6_10_io_i_5_ci),
    .io_o_6_co(cb_6_10_io_i_6_ci),
    .io_o_7_co(cb_6_10_io_i_7_ci),
    .io_vci(cb_6_8_io_vco),
    .io_vco(cb_6_10_io_vci),
    .io_vi(cb_6_9_io_vi),
    .io_we_i(cb_6_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_6_0_io_adr_i[1] ,
    \cb_6_0_io_adr_i[0] }),
    .io_dat_i({\cb_6_0_io_dat_i[15] ,
    \cb_6_0_io_dat_i[14] ,
    \cb_6_0_io_dat_i[13] ,
    \cb_6_0_io_dat_i[12] ,
    \cb_6_0_io_dat_i[11] ,
    \cb_6_0_io_dat_i[10] ,
    \cb_6_0_io_dat_i[9] ,
    \cb_6_0_io_dat_i[8] ,
    \cb_6_0_io_dat_i[7] ,
    \cb_6_0_io_dat_i[6] ,
    \cb_6_0_io_dat_i[5] ,
    \cb_6_0_io_dat_i[4] ,
    \cb_6_0_io_dat_i[3] ,
    \cb_6_0_io_dat_i[2] ,
    \cb_6_0_io_dat_i[1] ,
    \cb_6_0_io_dat_i[0] }),
    .io_dat_o({\cb_6_9_io_dat_o[15] ,
    \cb_6_9_io_dat_o[14] ,
    \cb_6_9_io_dat_o[13] ,
    \cb_6_9_io_dat_o[12] ,
    \cb_6_9_io_dat_o[11] ,
    \cb_6_9_io_dat_o[10] ,
    \cb_6_9_io_dat_o[9] ,
    \cb_6_9_io_dat_o[8] ,
    \cb_6_9_io_dat_o[7] ,
    \cb_6_9_io_dat_o[6] ,
    \cb_6_9_io_dat_o[5] ,
    \cb_6_9_io_dat_o[4] ,
    \cb_6_9_io_dat_o[3] ,
    \cb_6_9_io_dat_o[2] ,
    \cb_6_9_io_dat_o[1] ,
    \cb_6_9_io_dat_o[0] }),
    .io_eo({\cb_6_10_io_wo[63] ,
    \cb_6_10_io_wo[62] ,
    \cb_6_10_io_wo[61] ,
    \cb_6_10_io_wo[60] ,
    \cb_6_10_io_wo[59] ,
    \cb_6_10_io_wo[58] ,
    \cb_6_10_io_wo[57] ,
    \cb_6_10_io_wo[56] ,
    \cb_6_10_io_wo[55] ,
    \cb_6_10_io_wo[54] ,
    \cb_6_10_io_wo[53] ,
    \cb_6_10_io_wo[52] ,
    \cb_6_10_io_wo[51] ,
    \cb_6_10_io_wo[50] ,
    \cb_6_10_io_wo[49] ,
    \cb_6_10_io_wo[48] ,
    \cb_6_10_io_wo[47] ,
    \cb_6_10_io_wo[46] ,
    \cb_6_10_io_wo[45] ,
    \cb_6_10_io_wo[44] ,
    \cb_6_10_io_wo[43] ,
    \cb_6_10_io_wo[42] ,
    \cb_6_10_io_wo[41] ,
    \cb_6_10_io_wo[40] ,
    \cb_6_10_io_wo[39] ,
    \cb_6_10_io_wo[38] ,
    \cb_6_10_io_wo[37] ,
    \cb_6_10_io_wo[36] ,
    \cb_6_10_io_wo[35] ,
    \cb_6_10_io_wo[34] ,
    \cb_6_10_io_wo[33] ,
    \cb_6_10_io_wo[32] ,
    \cb_6_10_io_wo[31] ,
    \cb_6_10_io_wo[30] ,
    \cb_6_10_io_wo[29] ,
    \cb_6_10_io_wo[28] ,
    \cb_6_10_io_wo[27] ,
    \cb_6_10_io_wo[26] ,
    \cb_6_10_io_wo[25] ,
    \cb_6_10_io_wo[24] ,
    \cb_6_10_io_wo[23] ,
    \cb_6_10_io_wo[22] ,
    \cb_6_10_io_wo[21] ,
    \cb_6_10_io_wo[20] ,
    \cb_6_10_io_wo[19] ,
    \cb_6_10_io_wo[18] ,
    \cb_6_10_io_wo[17] ,
    \cb_6_10_io_wo[16] ,
    \cb_6_10_io_wo[15] ,
    \cb_6_10_io_wo[14] ,
    \cb_6_10_io_wo[13] ,
    \cb_6_10_io_wo[12] ,
    \cb_6_10_io_wo[11] ,
    \cb_6_10_io_wo[10] ,
    \cb_6_10_io_wo[9] ,
    \cb_6_10_io_wo[8] ,
    \cb_6_10_io_wo[7] ,
    \cb_6_10_io_wo[6] ,
    \cb_6_10_io_wo[5] ,
    \cb_6_10_io_wo[4] ,
    \cb_6_10_io_wo[3] ,
    \cb_6_10_io_wo[2] ,
    \cb_6_10_io_wo[1] ,
    \cb_6_10_io_wo[0] }),
    .io_i_0_in1({\cb_6_8_io_o_0_out[7] ,
    \cb_6_8_io_o_0_out[6] ,
    \cb_6_8_io_o_0_out[5] ,
    \cb_6_8_io_o_0_out[4] ,
    \cb_6_8_io_o_0_out[3] ,
    \cb_6_8_io_o_0_out[2] ,
    \cb_6_8_io_o_0_out[1] ,
    \cb_6_8_io_o_0_out[0] }),
    .io_i_1_in1({\cb_6_8_io_o_1_out[7] ,
    \cb_6_8_io_o_1_out[6] ,
    \cb_6_8_io_o_1_out[5] ,
    \cb_6_8_io_o_1_out[4] ,
    \cb_6_8_io_o_1_out[3] ,
    \cb_6_8_io_o_1_out[2] ,
    \cb_6_8_io_o_1_out[1] ,
    \cb_6_8_io_o_1_out[0] }),
    .io_i_2_in1({\cb_6_8_io_o_2_out[7] ,
    \cb_6_8_io_o_2_out[6] ,
    \cb_6_8_io_o_2_out[5] ,
    \cb_6_8_io_o_2_out[4] ,
    \cb_6_8_io_o_2_out[3] ,
    \cb_6_8_io_o_2_out[2] ,
    \cb_6_8_io_o_2_out[1] ,
    \cb_6_8_io_o_2_out[0] }),
    .io_i_3_in1({\cb_6_8_io_o_3_out[7] ,
    \cb_6_8_io_o_3_out[6] ,
    \cb_6_8_io_o_3_out[5] ,
    \cb_6_8_io_o_3_out[4] ,
    \cb_6_8_io_o_3_out[3] ,
    \cb_6_8_io_o_3_out[2] ,
    \cb_6_8_io_o_3_out[1] ,
    \cb_6_8_io_o_3_out[0] }),
    .io_i_4_in1({\cb_6_8_io_o_4_out[7] ,
    \cb_6_8_io_o_4_out[6] ,
    \cb_6_8_io_o_4_out[5] ,
    \cb_6_8_io_o_4_out[4] ,
    \cb_6_8_io_o_4_out[3] ,
    \cb_6_8_io_o_4_out[2] ,
    \cb_6_8_io_o_4_out[1] ,
    \cb_6_8_io_o_4_out[0] }),
    .io_i_5_in1({\cb_6_8_io_o_5_out[7] ,
    \cb_6_8_io_o_5_out[6] ,
    \cb_6_8_io_o_5_out[5] ,
    \cb_6_8_io_o_5_out[4] ,
    \cb_6_8_io_o_5_out[3] ,
    \cb_6_8_io_o_5_out[2] ,
    \cb_6_8_io_o_5_out[1] ,
    \cb_6_8_io_o_5_out[0] }),
    .io_i_6_in1({\cb_6_8_io_o_6_out[7] ,
    \cb_6_8_io_o_6_out[6] ,
    \cb_6_8_io_o_6_out[5] ,
    \cb_6_8_io_o_6_out[4] ,
    \cb_6_8_io_o_6_out[3] ,
    \cb_6_8_io_o_6_out[2] ,
    \cb_6_8_io_o_6_out[1] ,
    \cb_6_8_io_o_6_out[0] }),
    .io_i_7_in1({\cb_6_8_io_o_7_out[7] ,
    \cb_6_8_io_o_7_out[6] ,
    \cb_6_8_io_o_7_out[5] ,
    \cb_6_8_io_o_7_out[4] ,
    \cb_6_8_io_o_7_out[3] ,
    \cb_6_8_io_o_7_out[2] ,
    \cb_6_8_io_o_7_out[1] ,
    \cb_6_8_io_o_7_out[0] }),
    .io_o_0_out({\cb_6_10_io_i_0_in1[7] ,
    \cb_6_10_io_i_0_in1[6] ,
    \cb_6_10_io_i_0_in1[5] ,
    \cb_6_10_io_i_0_in1[4] ,
    \cb_6_10_io_i_0_in1[3] ,
    \cb_6_10_io_i_0_in1[2] ,
    \cb_6_10_io_i_0_in1[1] ,
    \cb_6_10_io_i_0_in1[0] }),
    .io_o_1_out({\cb_6_10_io_i_1_in1[7] ,
    \cb_6_10_io_i_1_in1[6] ,
    \cb_6_10_io_i_1_in1[5] ,
    \cb_6_10_io_i_1_in1[4] ,
    \cb_6_10_io_i_1_in1[3] ,
    \cb_6_10_io_i_1_in1[2] ,
    \cb_6_10_io_i_1_in1[1] ,
    \cb_6_10_io_i_1_in1[0] }),
    .io_o_2_out({\cb_6_10_io_i_2_in1[7] ,
    \cb_6_10_io_i_2_in1[6] ,
    \cb_6_10_io_i_2_in1[5] ,
    \cb_6_10_io_i_2_in1[4] ,
    \cb_6_10_io_i_2_in1[3] ,
    \cb_6_10_io_i_2_in1[2] ,
    \cb_6_10_io_i_2_in1[1] ,
    \cb_6_10_io_i_2_in1[0] }),
    .io_o_3_out({\cb_6_10_io_i_3_in1[7] ,
    \cb_6_10_io_i_3_in1[6] ,
    \cb_6_10_io_i_3_in1[5] ,
    \cb_6_10_io_i_3_in1[4] ,
    \cb_6_10_io_i_3_in1[3] ,
    \cb_6_10_io_i_3_in1[2] ,
    \cb_6_10_io_i_3_in1[1] ,
    \cb_6_10_io_i_3_in1[0] }),
    .io_o_4_out({\cb_6_10_io_i_4_in1[7] ,
    \cb_6_10_io_i_4_in1[6] ,
    \cb_6_10_io_i_4_in1[5] ,
    \cb_6_10_io_i_4_in1[4] ,
    \cb_6_10_io_i_4_in1[3] ,
    \cb_6_10_io_i_4_in1[2] ,
    \cb_6_10_io_i_4_in1[1] ,
    \cb_6_10_io_i_4_in1[0] }),
    .io_o_5_out({\cb_6_10_io_i_5_in1[7] ,
    \cb_6_10_io_i_5_in1[6] ,
    \cb_6_10_io_i_5_in1[5] ,
    \cb_6_10_io_i_5_in1[4] ,
    \cb_6_10_io_i_5_in1[3] ,
    \cb_6_10_io_i_5_in1[2] ,
    \cb_6_10_io_i_5_in1[1] ,
    \cb_6_10_io_i_5_in1[0] }),
    .io_o_6_out({\cb_6_10_io_i_6_in1[7] ,
    \cb_6_10_io_i_6_in1[6] ,
    \cb_6_10_io_i_6_in1[5] ,
    \cb_6_10_io_i_6_in1[4] ,
    \cb_6_10_io_i_6_in1[3] ,
    \cb_6_10_io_i_6_in1[2] ,
    \cb_6_10_io_i_6_in1[1] ,
    \cb_6_10_io_i_6_in1[0] }),
    .io_o_7_out({\cb_6_10_io_i_7_in1[7] ,
    \cb_6_10_io_i_7_in1[6] ,
    \cb_6_10_io_i_7_in1[5] ,
    \cb_6_10_io_i_7_in1[4] ,
    \cb_6_10_io_i_7_in1[3] ,
    \cb_6_10_io_i_7_in1[2] ,
    \cb_6_10_io_i_7_in1[1] ,
    \cb_6_10_io_i_7_in1[0] }),
    .io_wo({\cb_6_8_io_eo[63] ,
    \cb_6_8_io_eo[62] ,
    \cb_6_8_io_eo[61] ,
    \cb_6_8_io_eo[60] ,
    \cb_6_8_io_eo[59] ,
    \cb_6_8_io_eo[58] ,
    \cb_6_8_io_eo[57] ,
    \cb_6_8_io_eo[56] ,
    \cb_6_8_io_eo[55] ,
    \cb_6_8_io_eo[54] ,
    \cb_6_8_io_eo[53] ,
    \cb_6_8_io_eo[52] ,
    \cb_6_8_io_eo[51] ,
    \cb_6_8_io_eo[50] ,
    \cb_6_8_io_eo[49] ,
    \cb_6_8_io_eo[48] ,
    \cb_6_8_io_eo[47] ,
    \cb_6_8_io_eo[46] ,
    \cb_6_8_io_eo[45] ,
    \cb_6_8_io_eo[44] ,
    \cb_6_8_io_eo[43] ,
    \cb_6_8_io_eo[42] ,
    \cb_6_8_io_eo[41] ,
    \cb_6_8_io_eo[40] ,
    \cb_6_8_io_eo[39] ,
    \cb_6_8_io_eo[38] ,
    \cb_6_8_io_eo[37] ,
    \cb_6_8_io_eo[36] ,
    \cb_6_8_io_eo[35] ,
    \cb_6_8_io_eo[34] ,
    \cb_6_8_io_eo[33] ,
    \cb_6_8_io_eo[32] ,
    \cb_6_8_io_eo[31] ,
    \cb_6_8_io_eo[30] ,
    \cb_6_8_io_eo[29] ,
    \cb_6_8_io_eo[28] ,
    \cb_6_8_io_eo[27] ,
    \cb_6_8_io_eo[26] ,
    \cb_6_8_io_eo[25] ,
    \cb_6_8_io_eo[24] ,
    \cb_6_8_io_eo[23] ,
    \cb_6_8_io_eo[22] ,
    \cb_6_8_io_eo[21] ,
    \cb_6_8_io_eo[20] ,
    \cb_6_8_io_eo[19] ,
    \cb_6_8_io_eo[18] ,
    \cb_6_8_io_eo[17] ,
    \cb_6_8_io_eo[16] ,
    \cb_6_8_io_eo[15] ,
    \cb_6_8_io_eo[14] ,
    \cb_6_8_io_eo[13] ,
    \cb_6_8_io_eo[12] ,
    \cb_6_8_io_eo[11] ,
    \cb_6_8_io_eo[10] ,
    \cb_6_8_io_eo[9] ,
    \cb_6_8_io_eo[8] ,
    \cb_6_8_io_eo[7] ,
    \cb_6_8_io_eo[6] ,
    \cb_6_8_io_eo[5] ,
    \cb_6_8_io_eo[4] ,
    \cb_6_8_io_eo[3] ,
    \cb_6_8_io_eo[2] ,
    \cb_6_8_io_eo[1] ,
    \cb_6_8_io_eo[0] }));
 cic_block cb_7_0 (.io_cs_i(cb_7_0_io_cs_i),
    .io_i_0_ci(cb_7_0_io_i_0_ci),
    .io_o_0_co(cb_7_0_io_o_0_co),
    .io_o_1_co(cb_7_0_io_o_1_co),
    .io_o_2_co(cb_7_0_io_o_2_co),
    .io_o_3_co(cb_7_0_io_o_3_co),
    .io_o_4_co(cb_7_0_io_o_4_co),
    .io_o_5_co(cb_7_0_io_o_5_co),
    .io_o_6_co(cb_7_0_io_o_6_co),
    .io_o_7_co(cb_7_0_io_o_7_co),
    .io_vco(cb_7_0_io_vco),
    .io_vi(cb_7_0_io_vi),
    .io_we_i(cb_7_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_7_0_io_adr_i[1] ,
    \cb_7_0_io_adr_i[0] }),
    .io_dat_i({\cb_7_0_io_dat_i[15] ,
    \cb_7_0_io_dat_i[14] ,
    \cb_7_0_io_dat_i[13] ,
    \cb_7_0_io_dat_i[12] ,
    \cb_7_0_io_dat_i[11] ,
    \cb_7_0_io_dat_i[10] ,
    \cb_7_0_io_dat_i[9] ,
    \cb_7_0_io_dat_i[8] ,
    \cb_7_0_io_dat_i[7] ,
    \cb_7_0_io_dat_i[6] ,
    \cb_7_0_io_dat_i[5] ,
    \cb_7_0_io_dat_i[4] ,
    \cb_7_0_io_dat_i[3] ,
    \cb_7_0_io_dat_i[2] ,
    \cb_7_0_io_dat_i[1] ,
    \cb_7_0_io_dat_i[0] }),
    .io_dat_o({\cb_7_0_io_dat_o[15] ,
    \cb_7_0_io_dat_o[14] ,
    \cb_7_0_io_dat_o[13] ,
    \cb_7_0_io_dat_o[12] ,
    \cb_7_0_io_dat_o[11] ,
    \cb_7_0_io_dat_o[10] ,
    \cb_7_0_io_dat_o[9] ,
    \cb_7_0_io_dat_o[8] ,
    \cb_7_0_io_dat_o[7] ,
    \cb_7_0_io_dat_o[6] ,
    \cb_7_0_io_dat_o[5] ,
    \cb_7_0_io_dat_o[4] ,
    \cb_7_0_io_dat_o[3] ,
    \cb_7_0_io_dat_o[2] ,
    \cb_7_0_io_dat_o[1] ,
    \cb_7_0_io_dat_o[0] }),
    .io_eo({\cb_7_0_io_eo[63] ,
    \cb_7_0_io_eo[62] ,
    \cb_7_0_io_eo[61] ,
    \cb_7_0_io_eo[60] ,
    \cb_7_0_io_eo[59] ,
    \cb_7_0_io_eo[58] ,
    \cb_7_0_io_eo[57] ,
    \cb_7_0_io_eo[56] ,
    \cb_7_0_io_eo[55] ,
    \cb_7_0_io_eo[54] ,
    \cb_7_0_io_eo[53] ,
    \cb_7_0_io_eo[52] ,
    \cb_7_0_io_eo[51] ,
    \cb_7_0_io_eo[50] ,
    \cb_7_0_io_eo[49] ,
    \cb_7_0_io_eo[48] ,
    \cb_7_0_io_eo[47] ,
    \cb_7_0_io_eo[46] ,
    \cb_7_0_io_eo[45] ,
    \cb_7_0_io_eo[44] ,
    \cb_7_0_io_eo[43] ,
    \cb_7_0_io_eo[42] ,
    \cb_7_0_io_eo[41] ,
    \cb_7_0_io_eo[40] ,
    \cb_7_0_io_eo[39] ,
    \cb_7_0_io_eo[38] ,
    \cb_7_0_io_eo[37] ,
    \cb_7_0_io_eo[36] ,
    \cb_7_0_io_eo[35] ,
    \cb_7_0_io_eo[34] ,
    \cb_7_0_io_eo[33] ,
    \cb_7_0_io_eo[32] ,
    \cb_7_0_io_eo[31] ,
    \cb_7_0_io_eo[30] ,
    \cb_7_0_io_eo[29] ,
    \cb_7_0_io_eo[28] ,
    \cb_7_0_io_eo[27] ,
    \cb_7_0_io_eo[26] ,
    \cb_7_0_io_eo[25] ,
    \cb_7_0_io_eo[24] ,
    \cb_7_0_io_eo[23] ,
    \cb_7_0_io_eo[22] ,
    \cb_7_0_io_eo[21] ,
    \cb_7_0_io_eo[20] ,
    \cb_7_0_io_eo[19] ,
    \cb_7_0_io_eo[18] ,
    \cb_7_0_io_eo[17] ,
    \cb_7_0_io_eo[16] ,
    \cb_7_0_io_eo[15] ,
    \cb_7_0_io_eo[14] ,
    \cb_7_0_io_eo[13] ,
    \cb_7_0_io_eo[12] ,
    \cb_7_0_io_eo[11] ,
    \cb_7_0_io_eo[10] ,
    \cb_7_0_io_eo[9] ,
    \cb_7_0_io_eo[8] ,
    \cb_7_0_io_eo[7] ,
    \cb_7_0_io_eo[6] ,
    \cb_7_0_io_eo[5] ,
    \cb_7_0_io_eo[4] ,
    \cb_7_0_io_eo[3] ,
    \cb_7_0_io_eo[2] ,
    \cb_7_0_io_eo[1] ,
    \cb_7_0_io_eo[0] }),
    .io_i_0_in1({_NC449,
    _NC450,
    _NC451,
    _NC452,
    _NC453,
    _NC454,
    _NC455,
    _NC456}),
    .io_i_1_in1({_NC457,
    _NC458,
    _NC459,
    _NC460,
    _NC461,
    _NC462,
    _NC463,
    _NC464}),
    .io_i_2_in1({_NC465,
    _NC466,
    _NC467,
    _NC468,
    _NC469,
    _NC470,
    _NC471,
    _NC472}),
    .io_i_3_in1({_NC473,
    _NC474,
    _NC475,
    _NC476,
    _NC477,
    _NC478,
    _NC479,
    _NC480}),
    .io_i_4_in1({_NC481,
    _NC482,
    _NC483,
    _NC484,
    _NC485,
    _NC486,
    _NC487,
    _NC488}),
    .io_i_5_in1({_NC489,
    _NC490,
    _NC491,
    _NC492,
    _NC493,
    _NC494,
    _NC495,
    _NC496}),
    .io_i_6_in1({_NC497,
    _NC498,
    _NC499,
    _NC500,
    _NC501,
    _NC502,
    _NC503,
    _NC504}),
    .io_i_7_in1({_NC505,
    _NC506,
    _NC507,
    _NC508,
    _NC509,
    _NC510,
    _NC511,
    _NC512}),
    .io_o_0_out({\cb_7_0_io_o_0_out[7] ,
    \cb_7_0_io_o_0_out[6] ,
    \cb_7_0_io_o_0_out[5] ,
    \cb_7_0_io_o_0_out[4] ,
    \cb_7_0_io_o_0_out[3] ,
    \cb_7_0_io_o_0_out[2] ,
    \cb_7_0_io_o_0_out[1] ,
    \cb_7_0_io_o_0_out[0] }),
    .io_o_1_out({\cb_7_0_io_o_1_out[7] ,
    \cb_7_0_io_o_1_out[6] ,
    \cb_7_0_io_o_1_out[5] ,
    \cb_7_0_io_o_1_out[4] ,
    \cb_7_0_io_o_1_out[3] ,
    \cb_7_0_io_o_1_out[2] ,
    \cb_7_0_io_o_1_out[1] ,
    \cb_7_0_io_o_1_out[0] }),
    .io_o_2_out({\cb_7_0_io_o_2_out[7] ,
    \cb_7_0_io_o_2_out[6] ,
    \cb_7_0_io_o_2_out[5] ,
    \cb_7_0_io_o_2_out[4] ,
    \cb_7_0_io_o_2_out[3] ,
    \cb_7_0_io_o_2_out[2] ,
    \cb_7_0_io_o_2_out[1] ,
    \cb_7_0_io_o_2_out[0] }),
    .io_o_3_out({\cb_7_0_io_o_3_out[7] ,
    \cb_7_0_io_o_3_out[6] ,
    \cb_7_0_io_o_3_out[5] ,
    \cb_7_0_io_o_3_out[4] ,
    \cb_7_0_io_o_3_out[3] ,
    \cb_7_0_io_o_3_out[2] ,
    \cb_7_0_io_o_3_out[1] ,
    \cb_7_0_io_o_3_out[0] }),
    .io_o_4_out({\cb_7_0_io_o_4_out[7] ,
    \cb_7_0_io_o_4_out[6] ,
    \cb_7_0_io_o_4_out[5] ,
    \cb_7_0_io_o_4_out[4] ,
    \cb_7_0_io_o_4_out[3] ,
    \cb_7_0_io_o_4_out[2] ,
    \cb_7_0_io_o_4_out[1] ,
    \cb_7_0_io_o_4_out[0] }),
    .io_o_5_out({\cb_7_0_io_o_5_out[7] ,
    \cb_7_0_io_o_5_out[6] ,
    \cb_7_0_io_o_5_out[5] ,
    \cb_7_0_io_o_5_out[4] ,
    \cb_7_0_io_o_5_out[3] ,
    \cb_7_0_io_o_5_out[2] ,
    \cb_7_0_io_o_5_out[1] ,
    \cb_7_0_io_o_5_out[0] }),
    .io_o_6_out({\cb_7_0_io_o_6_out[7] ,
    \cb_7_0_io_o_6_out[6] ,
    \cb_7_0_io_o_6_out[5] ,
    \cb_7_0_io_o_6_out[4] ,
    \cb_7_0_io_o_6_out[3] ,
    \cb_7_0_io_o_6_out[2] ,
    \cb_7_0_io_o_6_out[1] ,
    \cb_7_0_io_o_6_out[0] }),
    .io_o_7_out({\cb_7_0_io_o_7_out[7] ,
    \cb_7_0_io_o_7_out[6] ,
    \cb_7_0_io_o_7_out[5] ,
    \cb_7_0_io_o_7_out[4] ,
    \cb_7_0_io_o_7_out[3] ,
    \cb_7_0_io_o_7_out[2] ,
    \cb_7_0_io_o_7_out[1] ,
    \cb_7_0_io_o_7_out[0] }),
    .io_wo({\cb_7_0_io_wo[63] ,
    \cb_7_0_io_wo[62] ,
    \cb_7_0_io_wo[61] ,
    \cb_7_0_io_wo[60] ,
    \cb_7_0_io_wo[59] ,
    \cb_7_0_io_wo[58] ,
    \cb_7_0_io_wo[57] ,
    \cb_7_0_io_wo[56] ,
    \cb_7_0_io_wo[55] ,
    \cb_7_0_io_wo[54] ,
    \cb_7_0_io_wo[53] ,
    \cb_7_0_io_wo[52] ,
    \cb_7_0_io_wo[51] ,
    \cb_7_0_io_wo[50] ,
    \cb_7_0_io_wo[49] ,
    \cb_7_0_io_wo[48] ,
    \cb_7_0_io_wo[47] ,
    \cb_7_0_io_wo[46] ,
    \cb_7_0_io_wo[45] ,
    \cb_7_0_io_wo[44] ,
    \cb_7_0_io_wo[43] ,
    \cb_7_0_io_wo[42] ,
    \cb_7_0_io_wo[41] ,
    \cb_7_0_io_wo[40] ,
    \cb_7_0_io_wo[39] ,
    \cb_7_0_io_wo[38] ,
    \cb_7_0_io_wo[37] ,
    \cb_7_0_io_wo[36] ,
    \cb_7_0_io_wo[35] ,
    \cb_7_0_io_wo[34] ,
    \cb_7_0_io_wo[33] ,
    \cb_7_0_io_wo[32] ,
    \cb_7_0_io_wo[31] ,
    \cb_7_0_io_wo[30] ,
    \cb_7_0_io_wo[29] ,
    \cb_7_0_io_wo[28] ,
    \cb_7_0_io_wo[27] ,
    \cb_7_0_io_wo[26] ,
    \cb_7_0_io_wo[25] ,
    \cb_7_0_io_wo[24] ,
    \cb_7_0_io_wo[23] ,
    \cb_7_0_io_wo[22] ,
    \cb_7_0_io_wo[21] ,
    \cb_7_0_io_wo[20] ,
    \cb_7_0_io_wo[19] ,
    \cb_7_0_io_wo[18] ,
    \cb_7_0_io_wo[17] ,
    \cb_7_0_io_wo[16] ,
    \cb_7_0_io_wo[15] ,
    \cb_7_0_io_wo[14] ,
    \cb_7_0_io_wo[13] ,
    \cb_7_0_io_wo[12] ,
    \cb_7_0_io_wo[11] ,
    \cb_7_0_io_wo[10] ,
    \cb_7_0_io_wo[9] ,
    \cb_7_0_io_wo[8] ,
    \cb_7_0_io_wo[7] ,
    \cb_7_0_io_wo[6] ,
    \cb_7_0_io_wo[5] ,
    \cb_7_0_io_wo[4] ,
    \cb_7_0_io_wo[3] ,
    \cb_7_0_io_wo[2] ,
    \cb_7_0_io_wo[1] ,
    \cb_7_0_io_wo[0] }));
 cic_block cb_7_1 (.io_cs_i(cb_7_1_io_cs_i),
    .io_i_0_ci(cb_7_0_io_o_0_co),
    .io_i_1_ci(cb_7_0_io_o_1_co),
    .io_i_2_ci(cb_7_0_io_o_2_co),
    .io_i_3_ci(cb_7_0_io_o_3_co),
    .io_i_4_ci(cb_7_0_io_o_4_co),
    .io_i_5_ci(cb_7_0_io_o_5_co),
    .io_i_6_ci(cb_7_0_io_o_6_co),
    .io_i_7_ci(cb_7_0_io_o_7_co),
    .io_o_0_co(cb_7_1_io_o_0_co),
    .io_o_1_co(cb_7_1_io_o_1_co),
    .io_o_2_co(cb_7_1_io_o_2_co),
    .io_o_3_co(cb_7_1_io_o_3_co),
    .io_o_4_co(cb_7_1_io_o_4_co),
    .io_o_5_co(cb_7_1_io_o_5_co),
    .io_o_6_co(cb_7_1_io_o_6_co),
    .io_o_7_co(cb_7_1_io_o_7_co),
    .io_vci(cb_7_0_io_vco),
    .io_vco(cb_7_1_io_vco),
    .io_vi(cb_7_1_io_vi),
    .io_we_i(cb_7_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_7_0_io_adr_i[1] ,
    \cb_7_0_io_adr_i[0] }),
    .io_dat_i({\cb_7_0_io_dat_i[15] ,
    \cb_7_0_io_dat_i[14] ,
    \cb_7_0_io_dat_i[13] ,
    \cb_7_0_io_dat_i[12] ,
    \cb_7_0_io_dat_i[11] ,
    \cb_7_0_io_dat_i[10] ,
    \cb_7_0_io_dat_i[9] ,
    \cb_7_0_io_dat_i[8] ,
    \cb_7_0_io_dat_i[7] ,
    \cb_7_0_io_dat_i[6] ,
    \cb_7_0_io_dat_i[5] ,
    \cb_7_0_io_dat_i[4] ,
    \cb_7_0_io_dat_i[3] ,
    \cb_7_0_io_dat_i[2] ,
    \cb_7_0_io_dat_i[1] ,
    \cb_7_0_io_dat_i[0] }),
    .io_dat_o({\cb_7_1_io_dat_o[15] ,
    \cb_7_1_io_dat_o[14] ,
    \cb_7_1_io_dat_o[13] ,
    \cb_7_1_io_dat_o[12] ,
    \cb_7_1_io_dat_o[11] ,
    \cb_7_1_io_dat_o[10] ,
    \cb_7_1_io_dat_o[9] ,
    \cb_7_1_io_dat_o[8] ,
    \cb_7_1_io_dat_o[7] ,
    \cb_7_1_io_dat_o[6] ,
    \cb_7_1_io_dat_o[5] ,
    \cb_7_1_io_dat_o[4] ,
    \cb_7_1_io_dat_o[3] ,
    \cb_7_1_io_dat_o[2] ,
    \cb_7_1_io_dat_o[1] ,
    \cb_7_1_io_dat_o[0] }),
    .io_eo({\cb_7_1_io_eo[63] ,
    \cb_7_1_io_eo[62] ,
    \cb_7_1_io_eo[61] ,
    \cb_7_1_io_eo[60] ,
    \cb_7_1_io_eo[59] ,
    \cb_7_1_io_eo[58] ,
    \cb_7_1_io_eo[57] ,
    \cb_7_1_io_eo[56] ,
    \cb_7_1_io_eo[55] ,
    \cb_7_1_io_eo[54] ,
    \cb_7_1_io_eo[53] ,
    \cb_7_1_io_eo[52] ,
    \cb_7_1_io_eo[51] ,
    \cb_7_1_io_eo[50] ,
    \cb_7_1_io_eo[49] ,
    \cb_7_1_io_eo[48] ,
    \cb_7_1_io_eo[47] ,
    \cb_7_1_io_eo[46] ,
    \cb_7_1_io_eo[45] ,
    \cb_7_1_io_eo[44] ,
    \cb_7_1_io_eo[43] ,
    \cb_7_1_io_eo[42] ,
    \cb_7_1_io_eo[41] ,
    \cb_7_1_io_eo[40] ,
    \cb_7_1_io_eo[39] ,
    \cb_7_1_io_eo[38] ,
    \cb_7_1_io_eo[37] ,
    \cb_7_1_io_eo[36] ,
    \cb_7_1_io_eo[35] ,
    \cb_7_1_io_eo[34] ,
    \cb_7_1_io_eo[33] ,
    \cb_7_1_io_eo[32] ,
    \cb_7_1_io_eo[31] ,
    \cb_7_1_io_eo[30] ,
    \cb_7_1_io_eo[29] ,
    \cb_7_1_io_eo[28] ,
    \cb_7_1_io_eo[27] ,
    \cb_7_1_io_eo[26] ,
    \cb_7_1_io_eo[25] ,
    \cb_7_1_io_eo[24] ,
    \cb_7_1_io_eo[23] ,
    \cb_7_1_io_eo[22] ,
    \cb_7_1_io_eo[21] ,
    \cb_7_1_io_eo[20] ,
    \cb_7_1_io_eo[19] ,
    \cb_7_1_io_eo[18] ,
    \cb_7_1_io_eo[17] ,
    \cb_7_1_io_eo[16] ,
    \cb_7_1_io_eo[15] ,
    \cb_7_1_io_eo[14] ,
    \cb_7_1_io_eo[13] ,
    \cb_7_1_io_eo[12] ,
    \cb_7_1_io_eo[11] ,
    \cb_7_1_io_eo[10] ,
    \cb_7_1_io_eo[9] ,
    \cb_7_1_io_eo[8] ,
    \cb_7_1_io_eo[7] ,
    \cb_7_1_io_eo[6] ,
    \cb_7_1_io_eo[5] ,
    \cb_7_1_io_eo[4] ,
    \cb_7_1_io_eo[3] ,
    \cb_7_1_io_eo[2] ,
    \cb_7_1_io_eo[1] ,
    \cb_7_1_io_eo[0] }),
    .io_i_0_in1({\cb_7_0_io_o_0_out[7] ,
    \cb_7_0_io_o_0_out[6] ,
    \cb_7_0_io_o_0_out[5] ,
    \cb_7_0_io_o_0_out[4] ,
    \cb_7_0_io_o_0_out[3] ,
    \cb_7_0_io_o_0_out[2] ,
    \cb_7_0_io_o_0_out[1] ,
    \cb_7_0_io_o_0_out[0] }),
    .io_i_1_in1({\cb_7_0_io_o_1_out[7] ,
    \cb_7_0_io_o_1_out[6] ,
    \cb_7_0_io_o_1_out[5] ,
    \cb_7_0_io_o_1_out[4] ,
    \cb_7_0_io_o_1_out[3] ,
    \cb_7_0_io_o_1_out[2] ,
    \cb_7_0_io_o_1_out[1] ,
    \cb_7_0_io_o_1_out[0] }),
    .io_i_2_in1({\cb_7_0_io_o_2_out[7] ,
    \cb_7_0_io_o_2_out[6] ,
    \cb_7_0_io_o_2_out[5] ,
    \cb_7_0_io_o_2_out[4] ,
    \cb_7_0_io_o_2_out[3] ,
    \cb_7_0_io_o_2_out[2] ,
    \cb_7_0_io_o_2_out[1] ,
    \cb_7_0_io_o_2_out[0] }),
    .io_i_3_in1({\cb_7_0_io_o_3_out[7] ,
    \cb_7_0_io_o_3_out[6] ,
    \cb_7_0_io_o_3_out[5] ,
    \cb_7_0_io_o_3_out[4] ,
    \cb_7_0_io_o_3_out[3] ,
    \cb_7_0_io_o_3_out[2] ,
    \cb_7_0_io_o_3_out[1] ,
    \cb_7_0_io_o_3_out[0] }),
    .io_i_4_in1({\cb_7_0_io_o_4_out[7] ,
    \cb_7_0_io_o_4_out[6] ,
    \cb_7_0_io_o_4_out[5] ,
    \cb_7_0_io_o_4_out[4] ,
    \cb_7_0_io_o_4_out[3] ,
    \cb_7_0_io_o_4_out[2] ,
    \cb_7_0_io_o_4_out[1] ,
    \cb_7_0_io_o_4_out[0] }),
    .io_i_5_in1({\cb_7_0_io_o_5_out[7] ,
    \cb_7_0_io_o_5_out[6] ,
    \cb_7_0_io_o_5_out[5] ,
    \cb_7_0_io_o_5_out[4] ,
    \cb_7_0_io_o_5_out[3] ,
    \cb_7_0_io_o_5_out[2] ,
    \cb_7_0_io_o_5_out[1] ,
    \cb_7_0_io_o_5_out[0] }),
    .io_i_6_in1({\cb_7_0_io_o_6_out[7] ,
    \cb_7_0_io_o_6_out[6] ,
    \cb_7_0_io_o_6_out[5] ,
    \cb_7_0_io_o_6_out[4] ,
    \cb_7_0_io_o_6_out[3] ,
    \cb_7_0_io_o_6_out[2] ,
    \cb_7_0_io_o_6_out[1] ,
    \cb_7_0_io_o_6_out[0] }),
    .io_i_7_in1({\cb_7_0_io_o_7_out[7] ,
    \cb_7_0_io_o_7_out[6] ,
    \cb_7_0_io_o_7_out[5] ,
    \cb_7_0_io_o_7_out[4] ,
    \cb_7_0_io_o_7_out[3] ,
    \cb_7_0_io_o_7_out[2] ,
    \cb_7_0_io_o_7_out[1] ,
    \cb_7_0_io_o_7_out[0] }),
    .io_o_0_out({\cb_7_1_io_o_0_out[7] ,
    \cb_7_1_io_o_0_out[6] ,
    \cb_7_1_io_o_0_out[5] ,
    \cb_7_1_io_o_0_out[4] ,
    \cb_7_1_io_o_0_out[3] ,
    \cb_7_1_io_o_0_out[2] ,
    \cb_7_1_io_o_0_out[1] ,
    \cb_7_1_io_o_0_out[0] }),
    .io_o_1_out({\cb_7_1_io_o_1_out[7] ,
    \cb_7_1_io_o_1_out[6] ,
    \cb_7_1_io_o_1_out[5] ,
    \cb_7_1_io_o_1_out[4] ,
    \cb_7_1_io_o_1_out[3] ,
    \cb_7_1_io_o_1_out[2] ,
    \cb_7_1_io_o_1_out[1] ,
    \cb_7_1_io_o_1_out[0] }),
    .io_o_2_out({\cb_7_1_io_o_2_out[7] ,
    \cb_7_1_io_o_2_out[6] ,
    \cb_7_1_io_o_2_out[5] ,
    \cb_7_1_io_o_2_out[4] ,
    \cb_7_1_io_o_2_out[3] ,
    \cb_7_1_io_o_2_out[2] ,
    \cb_7_1_io_o_2_out[1] ,
    \cb_7_1_io_o_2_out[0] }),
    .io_o_3_out({\cb_7_1_io_o_3_out[7] ,
    \cb_7_1_io_o_3_out[6] ,
    \cb_7_1_io_o_3_out[5] ,
    \cb_7_1_io_o_3_out[4] ,
    \cb_7_1_io_o_3_out[3] ,
    \cb_7_1_io_o_3_out[2] ,
    \cb_7_1_io_o_3_out[1] ,
    \cb_7_1_io_o_3_out[0] }),
    .io_o_4_out({\cb_7_1_io_o_4_out[7] ,
    \cb_7_1_io_o_4_out[6] ,
    \cb_7_1_io_o_4_out[5] ,
    \cb_7_1_io_o_4_out[4] ,
    \cb_7_1_io_o_4_out[3] ,
    \cb_7_1_io_o_4_out[2] ,
    \cb_7_1_io_o_4_out[1] ,
    \cb_7_1_io_o_4_out[0] }),
    .io_o_5_out({\cb_7_1_io_o_5_out[7] ,
    \cb_7_1_io_o_5_out[6] ,
    \cb_7_1_io_o_5_out[5] ,
    \cb_7_1_io_o_5_out[4] ,
    \cb_7_1_io_o_5_out[3] ,
    \cb_7_1_io_o_5_out[2] ,
    \cb_7_1_io_o_5_out[1] ,
    \cb_7_1_io_o_5_out[0] }),
    .io_o_6_out({\cb_7_1_io_o_6_out[7] ,
    \cb_7_1_io_o_6_out[6] ,
    \cb_7_1_io_o_6_out[5] ,
    \cb_7_1_io_o_6_out[4] ,
    \cb_7_1_io_o_6_out[3] ,
    \cb_7_1_io_o_6_out[2] ,
    \cb_7_1_io_o_6_out[1] ,
    \cb_7_1_io_o_6_out[0] }),
    .io_o_7_out({\cb_7_1_io_o_7_out[7] ,
    \cb_7_1_io_o_7_out[6] ,
    \cb_7_1_io_o_7_out[5] ,
    \cb_7_1_io_o_7_out[4] ,
    \cb_7_1_io_o_7_out[3] ,
    \cb_7_1_io_o_7_out[2] ,
    \cb_7_1_io_o_7_out[1] ,
    \cb_7_1_io_o_7_out[0] }),
    .io_wo({\cb_7_0_io_eo[63] ,
    \cb_7_0_io_eo[62] ,
    \cb_7_0_io_eo[61] ,
    \cb_7_0_io_eo[60] ,
    \cb_7_0_io_eo[59] ,
    \cb_7_0_io_eo[58] ,
    \cb_7_0_io_eo[57] ,
    \cb_7_0_io_eo[56] ,
    \cb_7_0_io_eo[55] ,
    \cb_7_0_io_eo[54] ,
    \cb_7_0_io_eo[53] ,
    \cb_7_0_io_eo[52] ,
    \cb_7_0_io_eo[51] ,
    \cb_7_0_io_eo[50] ,
    \cb_7_0_io_eo[49] ,
    \cb_7_0_io_eo[48] ,
    \cb_7_0_io_eo[47] ,
    \cb_7_0_io_eo[46] ,
    \cb_7_0_io_eo[45] ,
    \cb_7_0_io_eo[44] ,
    \cb_7_0_io_eo[43] ,
    \cb_7_0_io_eo[42] ,
    \cb_7_0_io_eo[41] ,
    \cb_7_0_io_eo[40] ,
    \cb_7_0_io_eo[39] ,
    \cb_7_0_io_eo[38] ,
    \cb_7_0_io_eo[37] ,
    \cb_7_0_io_eo[36] ,
    \cb_7_0_io_eo[35] ,
    \cb_7_0_io_eo[34] ,
    \cb_7_0_io_eo[33] ,
    \cb_7_0_io_eo[32] ,
    \cb_7_0_io_eo[31] ,
    \cb_7_0_io_eo[30] ,
    \cb_7_0_io_eo[29] ,
    \cb_7_0_io_eo[28] ,
    \cb_7_0_io_eo[27] ,
    \cb_7_0_io_eo[26] ,
    \cb_7_0_io_eo[25] ,
    \cb_7_0_io_eo[24] ,
    \cb_7_0_io_eo[23] ,
    \cb_7_0_io_eo[22] ,
    \cb_7_0_io_eo[21] ,
    \cb_7_0_io_eo[20] ,
    \cb_7_0_io_eo[19] ,
    \cb_7_0_io_eo[18] ,
    \cb_7_0_io_eo[17] ,
    \cb_7_0_io_eo[16] ,
    \cb_7_0_io_eo[15] ,
    \cb_7_0_io_eo[14] ,
    \cb_7_0_io_eo[13] ,
    \cb_7_0_io_eo[12] ,
    \cb_7_0_io_eo[11] ,
    \cb_7_0_io_eo[10] ,
    \cb_7_0_io_eo[9] ,
    \cb_7_0_io_eo[8] ,
    \cb_7_0_io_eo[7] ,
    \cb_7_0_io_eo[6] ,
    \cb_7_0_io_eo[5] ,
    \cb_7_0_io_eo[4] ,
    \cb_7_0_io_eo[3] ,
    \cb_7_0_io_eo[2] ,
    \cb_7_0_io_eo[1] ,
    \cb_7_0_io_eo[0] }));
 cic_block cb_7_10 (.io_cs_i(cb_7_10_io_cs_i),
    .io_i_0_ci(cb_7_10_io_i_0_ci),
    .io_i_1_ci(cb_7_10_io_i_1_ci),
    .io_i_2_ci(cb_7_10_io_i_2_ci),
    .io_i_3_ci(cb_7_10_io_i_3_ci),
    .io_i_4_ci(cb_7_10_io_i_4_ci),
    .io_i_5_ci(cb_7_10_io_i_5_ci),
    .io_i_6_ci(cb_7_10_io_i_6_ci),
    .io_i_7_ci(cb_7_10_io_i_7_ci),
    .io_o_0_co(cb_7_10_io_o_0_co),
    .io_o_1_co(cb_7_10_io_o_1_co),
    .io_o_2_co(cb_7_10_io_o_2_co),
    .io_o_3_co(cb_7_10_io_o_3_co),
    .io_o_4_co(cb_7_10_io_o_4_co),
    .io_o_5_co(cb_7_10_io_o_5_co),
    .io_o_6_co(cb_7_10_io_o_6_co),
    .io_o_7_co(cb_7_10_io_o_7_co),
    .io_vci(cb_7_10_io_vci),
    .io_vco(cb_7_10_io_vco),
    .io_vi(cb_7_10_io_vi),
    .io_we_i(cb_7_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_7_0_io_adr_i[1] ,
    \cb_7_0_io_adr_i[0] }),
    .io_dat_i({\cb_7_0_io_dat_i[15] ,
    \cb_7_0_io_dat_i[14] ,
    \cb_7_0_io_dat_i[13] ,
    \cb_7_0_io_dat_i[12] ,
    \cb_7_0_io_dat_i[11] ,
    \cb_7_0_io_dat_i[10] ,
    \cb_7_0_io_dat_i[9] ,
    \cb_7_0_io_dat_i[8] ,
    \cb_7_0_io_dat_i[7] ,
    \cb_7_0_io_dat_i[6] ,
    \cb_7_0_io_dat_i[5] ,
    \cb_7_0_io_dat_i[4] ,
    \cb_7_0_io_dat_i[3] ,
    \cb_7_0_io_dat_i[2] ,
    \cb_7_0_io_dat_i[1] ,
    \cb_7_0_io_dat_i[0] }),
    .io_dat_o({\cb_7_10_io_dat_o[15] ,
    \cb_7_10_io_dat_o[14] ,
    \cb_7_10_io_dat_o[13] ,
    \cb_7_10_io_dat_o[12] ,
    \cb_7_10_io_dat_o[11] ,
    \cb_7_10_io_dat_o[10] ,
    \cb_7_10_io_dat_o[9] ,
    \cb_7_10_io_dat_o[8] ,
    \cb_7_10_io_dat_o[7] ,
    \cb_7_10_io_dat_o[6] ,
    \cb_7_10_io_dat_o[5] ,
    \cb_7_10_io_dat_o[4] ,
    \cb_7_10_io_dat_o[3] ,
    \cb_7_10_io_dat_o[2] ,
    \cb_7_10_io_dat_o[1] ,
    \cb_7_10_io_dat_o[0] }),
    .io_eo({\_T_161[31] ,
    \_T_161[30] ,
    \_T_161[29] ,
    \_T_161[28] ,
    \_T_161[27] ,
    \_T_161[26] ,
    \_T_161[25] ,
    \_T_161[24] ,
    \_T_161[23] ,
    \_T_161[22] ,
    \_T_161[21] ,
    \_T_161[20] ,
    \_T_161[19] ,
    \_T_161[18] ,
    \_T_161[17] ,
    \_T_161[16] ,
    \_T_161[15] ,
    \_T_161[14] ,
    \_T_161[13] ,
    \_T_161[12] ,
    \_T_161[11] ,
    \_T_161[10] ,
    \_T_161[9] ,
    \_T_161[8] ,
    \_T_161[7] ,
    \_T_161[6] ,
    \_T_161[5] ,
    \_T_161[4] ,
    \_T_161[3] ,
    \_T_161[2] ,
    \_T_161[1] ,
    \_T_161[0] ,
    \_T_158[31] ,
    \_T_158[30] ,
    \_T_158[29] ,
    \_T_158[28] ,
    \_T_158[27] ,
    \_T_158[26] ,
    \_T_158[25] ,
    \_T_158[24] ,
    \_T_158[23] ,
    \_T_158[22] ,
    \_T_158[21] ,
    \_T_158[20] ,
    \_T_158[19] ,
    \_T_158[18] ,
    \_T_158[17] ,
    \_T_158[16] ,
    \_T_158[15] ,
    \_T_158[14] ,
    \_T_158[13] ,
    \_T_158[12] ,
    \_T_158[11] ,
    \_T_158[10] ,
    \_T_158[9] ,
    \_T_158[8] ,
    \_T_158[7] ,
    \_T_158[6] ,
    \_T_158[5] ,
    \_T_158[4] ,
    \_T_158[3] ,
    \_T_158[2] ,
    \_T_158[1] ,
    \_T_158[0] }),
    .io_i_0_in1({\cb_7_10_io_i_0_in1[7] ,
    \cb_7_10_io_i_0_in1[6] ,
    \cb_7_10_io_i_0_in1[5] ,
    \cb_7_10_io_i_0_in1[4] ,
    \cb_7_10_io_i_0_in1[3] ,
    \cb_7_10_io_i_0_in1[2] ,
    \cb_7_10_io_i_0_in1[1] ,
    \cb_7_10_io_i_0_in1[0] }),
    .io_i_1_in1({\cb_7_10_io_i_1_in1[7] ,
    \cb_7_10_io_i_1_in1[6] ,
    \cb_7_10_io_i_1_in1[5] ,
    \cb_7_10_io_i_1_in1[4] ,
    \cb_7_10_io_i_1_in1[3] ,
    \cb_7_10_io_i_1_in1[2] ,
    \cb_7_10_io_i_1_in1[1] ,
    \cb_7_10_io_i_1_in1[0] }),
    .io_i_2_in1({\cb_7_10_io_i_2_in1[7] ,
    \cb_7_10_io_i_2_in1[6] ,
    \cb_7_10_io_i_2_in1[5] ,
    \cb_7_10_io_i_2_in1[4] ,
    \cb_7_10_io_i_2_in1[3] ,
    \cb_7_10_io_i_2_in1[2] ,
    \cb_7_10_io_i_2_in1[1] ,
    \cb_7_10_io_i_2_in1[0] }),
    .io_i_3_in1({\cb_7_10_io_i_3_in1[7] ,
    \cb_7_10_io_i_3_in1[6] ,
    \cb_7_10_io_i_3_in1[5] ,
    \cb_7_10_io_i_3_in1[4] ,
    \cb_7_10_io_i_3_in1[3] ,
    \cb_7_10_io_i_3_in1[2] ,
    \cb_7_10_io_i_3_in1[1] ,
    \cb_7_10_io_i_3_in1[0] }),
    .io_i_4_in1({\cb_7_10_io_i_4_in1[7] ,
    \cb_7_10_io_i_4_in1[6] ,
    \cb_7_10_io_i_4_in1[5] ,
    \cb_7_10_io_i_4_in1[4] ,
    \cb_7_10_io_i_4_in1[3] ,
    \cb_7_10_io_i_4_in1[2] ,
    \cb_7_10_io_i_4_in1[1] ,
    \cb_7_10_io_i_4_in1[0] }),
    .io_i_5_in1({\cb_7_10_io_i_5_in1[7] ,
    \cb_7_10_io_i_5_in1[6] ,
    \cb_7_10_io_i_5_in1[5] ,
    \cb_7_10_io_i_5_in1[4] ,
    \cb_7_10_io_i_5_in1[3] ,
    \cb_7_10_io_i_5_in1[2] ,
    \cb_7_10_io_i_5_in1[1] ,
    \cb_7_10_io_i_5_in1[0] }),
    .io_i_6_in1({\cb_7_10_io_i_6_in1[7] ,
    \cb_7_10_io_i_6_in1[6] ,
    \cb_7_10_io_i_6_in1[5] ,
    \cb_7_10_io_i_6_in1[4] ,
    \cb_7_10_io_i_6_in1[3] ,
    \cb_7_10_io_i_6_in1[2] ,
    \cb_7_10_io_i_6_in1[1] ,
    \cb_7_10_io_i_6_in1[0] }),
    .io_i_7_in1({\cb_7_10_io_i_7_in1[7] ,
    \cb_7_10_io_i_7_in1[6] ,
    \cb_7_10_io_i_7_in1[5] ,
    \cb_7_10_io_i_7_in1[4] ,
    \cb_7_10_io_i_7_in1[3] ,
    \cb_7_10_io_i_7_in1[2] ,
    \cb_7_10_io_i_7_in1[1] ,
    \cb_7_10_io_i_7_in1[0] }),
    .io_o_0_out({\_T_158[7] ,
    \_T_158[6] ,
    \_T_158[5] ,
    \_T_158[4] ,
    \_T_158[3] ,
    \_T_158[2] ,
    \_T_158[1] ,
    \_T_158[0] }),
    .io_o_1_out({\_T_158[15] ,
    \_T_158[14] ,
    \_T_158[13] ,
    \_T_158[12] ,
    \_T_158[11] ,
    \_T_158[10] ,
    \_T_158[9] ,
    \_T_158[8] }),
    .io_o_2_out({\_T_158[23] ,
    \_T_158[22] ,
    \_T_158[21] ,
    \_T_158[20] ,
    \_T_158[19] ,
    \_T_158[18] ,
    \_T_158[17] ,
    \_T_158[16] }),
    .io_o_3_out({\_T_158[31] ,
    \_T_158[30] ,
    \_T_158[29] ,
    \_T_158[28] ,
    \_T_158[27] ,
    \_T_158[26] ,
    \_T_158[25] ,
    \_T_158[24] }),
    .io_o_4_out({\_T_161[7] ,
    \_T_161[6] ,
    \_T_161[5] ,
    \_T_161[4] ,
    \_T_161[3] ,
    \_T_161[2] ,
    \_T_161[1] ,
    \_T_161[0] }),
    .io_o_5_out({\_T_161[15] ,
    \_T_161[14] ,
    \_T_161[13] ,
    \_T_161[12] ,
    \_T_161[11] ,
    \_T_161[10] ,
    \_T_161[9] ,
    \_T_161[8] }),
    .io_o_6_out({\_T_161[23] ,
    \_T_161[22] ,
    \_T_161[21] ,
    \_T_161[20] ,
    \_T_161[19] ,
    \_T_161[18] ,
    \_T_161[17] ,
    \_T_161[16] }),
    .io_o_7_out({\_T_161[31] ,
    \_T_161[30] ,
    \_T_161[29] ,
    \_T_161[28] ,
    \_T_161[27] ,
    \_T_161[26] ,
    \_T_161[25] ,
    \_T_161[24] }),
    .io_wo({\cb_7_10_io_wo[63] ,
    \cb_7_10_io_wo[62] ,
    \cb_7_10_io_wo[61] ,
    \cb_7_10_io_wo[60] ,
    \cb_7_10_io_wo[59] ,
    \cb_7_10_io_wo[58] ,
    \cb_7_10_io_wo[57] ,
    \cb_7_10_io_wo[56] ,
    \cb_7_10_io_wo[55] ,
    \cb_7_10_io_wo[54] ,
    \cb_7_10_io_wo[53] ,
    \cb_7_10_io_wo[52] ,
    \cb_7_10_io_wo[51] ,
    \cb_7_10_io_wo[50] ,
    \cb_7_10_io_wo[49] ,
    \cb_7_10_io_wo[48] ,
    \cb_7_10_io_wo[47] ,
    \cb_7_10_io_wo[46] ,
    \cb_7_10_io_wo[45] ,
    \cb_7_10_io_wo[44] ,
    \cb_7_10_io_wo[43] ,
    \cb_7_10_io_wo[42] ,
    \cb_7_10_io_wo[41] ,
    \cb_7_10_io_wo[40] ,
    \cb_7_10_io_wo[39] ,
    \cb_7_10_io_wo[38] ,
    \cb_7_10_io_wo[37] ,
    \cb_7_10_io_wo[36] ,
    \cb_7_10_io_wo[35] ,
    \cb_7_10_io_wo[34] ,
    \cb_7_10_io_wo[33] ,
    \cb_7_10_io_wo[32] ,
    \cb_7_10_io_wo[31] ,
    \cb_7_10_io_wo[30] ,
    \cb_7_10_io_wo[29] ,
    \cb_7_10_io_wo[28] ,
    \cb_7_10_io_wo[27] ,
    \cb_7_10_io_wo[26] ,
    \cb_7_10_io_wo[25] ,
    \cb_7_10_io_wo[24] ,
    \cb_7_10_io_wo[23] ,
    \cb_7_10_io_wo[22] ,
    \cb_7_10_io_wo[21] ,
    \cb_7_10_io_wo[20] ,
    \cb_7_10_io_wo[19] ,
    \cb_7_10_io_wo[18] ,
    \cb_7_10_io_wo[17] ,
    \cb_7_10_io_wo[16] ,
    \cb_7_10_io_wo[15] ,
    \cb_7_10_io_wo[14] ,
    \cb_7_10_io_wo[13] ,
    \cb_7_10_io_wo[12] ,
    \cb_7_10_io_wo[11] ,
    \cb_7_10_io_wo[10] ,
    \cb_7_10_io_wo[9] ,
    \cb_7_10_io_wo[8] ,
    \cb_7_10_io_wo[7] ,
    \cb_7_10_io_wo[6] ,
    \cb_7_10_io_wo[5] ,
    \cb_7_10_io_wo[4] ,
    \cb_7_10_io_wo[3] ,
    \cb_7_10_io_wo[2] ,
    \cb_7_10_io_wo[1] ,
    \cb_7_10_io_wo[0] }));
 cic_block cb_7_2 (.io_cs_i(cb_7_2_io_cs_i),
    .io_i_0_ci(cb_7_1_io_o_0_co),
    .io_i_1_ci(cb_7_1_io_o_1_co),
    .io_i_2_ci(cb_7_1_io_o_2_co),
    .io_i_3_ci(cb_7_1_io_o_3_co),
    .io_i_4_ci(cb_7_1_io_o_4_co),
    .io_i_5_ci(cb_7_1_io_o_5_co),
    .io_i_6_ci(cb_7_1_io_o_6_co),
    .io_i_7_ci(cb_7_1_io_o_7_co),
    .io_o_0_co(cb_7_2_io_o_0_co),
    .io_o_1_co(cb_7_2_io_o_1_co),
    .io_o_2_co(cb_7_2_io_o_2_co),
    .io_o_3_co(cb_7_2_io_o_3_co),
    .io_o_4_co(cb_7_2_io_o_4_co),
    .io_o_5_co(cb_7_2_io_o_5_co),
    .io_o_6_co(cb_7_2_io_o_6_co),
    .io_o_7_co(cb_7_2_io_o_7_co),
    .io_vci(cb_7_1_io_vco),
    .io_vco(cb_7_2_io_vco),
    .io_vi(cb_7_2_io_vi),
    .io_we_i(cb_7_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_7_0_io_adr_i[1] ,
    \cb_7_0_io_adr_i[0] }),
    .io_dat_i({\cb_7_0_io_dat_i[15] ,
    \cb_7_0_io_dat_i[14] ,
    \cb_7_0_io_dat_i[13] ,
    \cb_7_0_io_dat_i[12] ,
    \cb_7_0_io_dat_i[11] ,
    \cb_7_0_io_dat_i[10] ,
    \cb_7_0_io_dat_i[9] ,
    \cb_7_0_io_dat_i[8] ,
    \cb_7_0_io_dat_i[7] ,
    \cb_7_0_io_dat_i[6] ,
    \cb_7_0_io_dat_i[5] ,
    \cb_7_0_io_dat_i[4] ,
    \cb_7_0_io_dat_i[3] ,
    \cb_7_0_io_dat_i[2] ,
    \cb_7_0_io_dat_i[1] ,
    \cb_7_0_io_dat_i[0] }),
    .io_dat_o({\cb_7_2_io_dat_o[15] ,
    \cb_7_2_io_dat_o[14] ,
    \cb_7_2_io_dat_o[13] ,
    \cb_7_2_io_dat_o[12] ,
    \cb_7_2_io_dat_o[11] ,
    \cb_7_2_io_dat_o[10] ,
    \cb_7_2_io_dat_o[9] ,
    \cb_7_2_io_dat_o[8] ,
    \cb_7_2_io_dat_o[7] ,
    \cb_7_2_io_dat_o[6] ,
    \cb_7_2_io_dat_o[5] ,
    \cb_7_2_io_dat_o[4] ,
    \cb_7_2_io_dat_o[3] ,
    \cb_7_2_io_dat_o[2] ,
    \cb_7_2_io_dat_o[1] ,
    \cb_7_2_io_dat_o[0] }),
    .io_eo({\cb_7_2_io_eo[63] ,
    \cb_7_2_io_eo[62] ,
    \cb_7_2_io_eo[61] ,
    \cb_7_2_io_eo[60] ,
    \cb_7_2_io_eo[59] ,
    \cb_7_2_io_eo[58] ,
    \cb_7_2_io_eo[57] ,
    \cb_7_2_io_eo[56] ,
    \cb_7_2_io_eo[55] ,
    \cb_7_2_io_eo[54] ,
    \cb_7_2_io_eo[53] ,
    \cb_7_2_io_eo[52] ,
    \cb_7_2_io_eo[51] ,
    \cb_7_2_io_eo[50] ,
    \cb_7_2_io_eo[49] ,
    \cb_7_2_io_eo[48] ,
    \cb_7_2_io_eo[47] ,
    \cb_7_2_io_eo[46] ,
    \cb_7_2_io_eo[45] ,
    \cb_7_2_io_eo[44] ,
    \cb_7_2_io_eo[43] ,
    \cb_7_2_io_eo[42] ,
    \cb_7_2_io_eo[41] ,
    \cb_7_2_io_eo[40] ,
    \cb_7_2_io_eo[39] ,
    \cb_7_2_io_eo[38] ,
    \cb_7_2_io_eo[37] ,
    \cb_7_2_io_eo[36] ,
    \cb_7_2_io_eo[35] ,
    \cb_7_2_io_eo[34] ,
    \cb_7_2_io_eo[33] ,
    \cb_7_2_io_eo[32] ,
    \cb_7_2_io_eo[31] ,
    \cb_7_2_io_eo[30] ,
    \cb_7_2_io_eo[29] ,
    \cb_7_2_io_eo[28] ,
    \cb_7_2_io_eo[27] ,
    \cb_7_2_io_eo[26] ,
    \cb_7_2_io_eo[25] ,
    \cb_7_2_io_eo[24] ,
    \cb_7_2_io_eo[23] ,
    \cb_7_2_io_eo[22] ,
    \cb_7_2_io_eo[21] ,
    \cb_7_2_io_eo[20] ,
    \cb_7_2_io_eo[19] ,
    \cb_7_2_io_eo[18] ,
    \cb_7_2_io_eo[17] ,
    \cb_7_2_io_eo[16] ,
    \cb_7_2_io_eo[15] ,
    \cb_7_2_io_eo[14] ,
    \cb_7_2_io_eo[13] ,
    \cb_7_2_io_eo[12] ,
    \cb_7_2_io_eo[11] ,
    \cb_7_2_io_eo[10] ,
    \cb_7_2_io_eo[9] ,
    \cb_7_2_io_eo[8] ,
    \cb_7_2_io_eo[7] ,
    \cb_7_2_io_eo[6] ,
    \cb_7_2_io_eo[5] ,
    \cb_7_2_io_eo[4] ,
    \cb_7_2_io_eo[3] ,
    \cb_7_2_io_eo[2] ,
    \cb_7_2_io_eo[1] ,
    \cb_7_2_io_eo[0] }),
    .io_i_0_in1({\cb_7_1_io_o_0_out[7] ,
    \cb_7_1_io_o_0_out[6] ,
    \cb_7_1_io_o_0_out[5] ,
    \cb_7_1_io_o_0_out[4] ,
    \cb_7_1_io_o_0_out[3] ,
    \cb_7_1_io_o_0_out[2] ,
    \cb_7_1_io_o_0_out[1] ,
    \cb_7_1_io_o_0_out[0] }),
    .io_i_1_in1({\cb_7_1_io_o_1_out[7] ,
    \cb_7_1_io_o_1_out[6] ,
    \cb_7_1_io_o_1_out[5] ,
    \cb_7_1_io_o_1_out[4] ,
    \cb_7_1_io_o_1_out[3] ,
    \cb_7_1_io_o_1_out[2] ,
    \cb_7_1_io_o_1_out[1] ,
    \cb_7_1_io_o_1_out[0] }),
    .io_i_2_in1({\cb_7_1_io_o_2_out[7] ,
    \cb_7_1_io_o_2_out[6] ,
    \cb_7_1_io_o_2_out[5] ,
    \cb_7_1_io_o_2_out[4] ,
    \cb_7_1_io_o_2_out[3] ,
    \cb_7_1_io_o_2_out[2] ,
    \cb_7_1_io_o_2_out[1] ,
    \cb_7_1_io_o_2_out[0] }),
    .io_i_3_in1({\cb_7_1_io_o_3_out[7] ,
    \cb_7_1_io_o_3_out[6] ,
    \cb_7_1_io_o_3_out[5] ,
    \cb_7_1_io_o_3_out[4] ,
    \cb_7_1_io_o_3_out[3] ,
    \cb_7_1_io_o_3_out[2] ,
    \cb_7_1_io_o_3_out[1] ,
    \cb_7_1_io_o_3_out[0] }),
    .io_i_4_in1({\cb_7_1_io_o_4_out[7] ,
    \cb_7_1_io_o_4_out[6] ,
    \cb_7_1_io_o_4_out[5] ,
    \cb_7_1_io_o_4_out[4] ,
    \cb_7_1_io_o_4_out[3] ,
    \cb_7_1_io_o_4_out[2] ,
    \cb_7_1_io_o_4_out[1] ,
    \cb_7_1_io_o_4_out[0] }),
    .io_i_5_in1({\cb_7_1_io_o_5_out[7] ,
    \cb_7_1_io_o_5_out[6] ,
    \cb_7_1_io_o_5_out[5] ,
    \cb_7_1_io_o_5_out[4] ,
    \cb_7_1_io_o_5_out[3] ,
    \cb_7_1_io_o_5_out[2] ,
    \cb_7_1_io_o_5_out[1] ,
    \cb_7_1_io_o_5_out[0] }),
    .io_i_6_in1({\cb_7_1_io_o_6_out[7] ,
    \cb_7_1_io_o_6_out[6] ,
    \cb_7_1_io_o_6_out[5] ,
    \cb_7_1_io_o_6_out[4] ,
    \cb_7_1_io_o_6_out[3] ,
    \cb_7_1_io_o_6_out[2] ,
    \cb_7_1_io_o_6_out[1] ,
    \cb_7_1_io_o_6_out[0] }),
    .io_i_7_in1({\cb_7_1_io_o_7_out[7] ,
    \cb_7_1_io_o_7_out[6] ,
    \cb_7_1_io_o_7_out[5] ,
    \cb_7_1_io_o_7_out[4] ,
    \cb_7_1_io_o_7_out[3] ,
    \cb_7_1_io_o_7_out[2] ,
    \cb_7_1_io_o_7_out[1] ,
    \cb_7_1_io_o_7_out[0] }),
    .io_o_0_out({\cb_7_2_io_o_0_out[7] ,
    \cb_7_2_io_o_0_out[6] ,
    \cb_7_2_io_o_0_out[5] ,
    \cb_7_2_io_o_0_out[4] ,
    \cb_7_2_io_o_0_out[3] ,
    \cb_7_2_io_o_0_out[2] ,
    \cb_7_2_io_o_0_out[1] ,
    \cb_7_2_io_o_0_out[0] }),
    .io_o_1_out({\cb_7_2_io_o_1_out[7] ,
    \cb_7_2_io_o_1_out[6] ,
    \cb_7_2_io_o_1_out[5] ,
    \cb_7_2_io_o_1_out[4] ,
    \cb_7_2_io_o_1_out[3] ,
    \cb_7_2_io_o_1_out[2] ,
    \cb_7_2_io_o_1_out[1] ,
    \cb_7_2_io_o_1_out[0] }),
    .io_o_2_out({\cb_7_2_io_o_2_out[7] ,
    \cb_7_2_io_o_2_out[6] ,
    \cb_7_2_io_o_2_out[5] ,
    \cb_7_2_io_o_2_out[4] ,
    \cb_7_2_io_o_2_out[3] ,
    \cb_7_2_io_o_2_out[2] ,
    \cb_7_2_io_o_2_out[1] ,
    \cb_7_2_io_o_2_out[0] }),
    .io_o_3_out({\cb_7_2_io_o_3_out[7] ,
    \cb_7_2_io_o_3_out[6] ,
    \cb_7_2_io_o_3_out[5] ,
    \cb_7_2_io_o_3_out[4] ,
    \cb_7_2_io_o_3_out[3] ,
    \cb_7_2_io_o_3_out[2] ,
    \cb_7_2_io_o_3_out[1] ,
    \cb_7_2_io_o_3_out[0] }),
    .io_o_4_out({\cb_7_2_io_o_4_out[7] ,
    \cb_7_2_io_o_4_out[6] ,
    \cb_7_2_io_o_4_out[5] ,
    \cb_7_2_io_o_4_out[4] ,
    \cb_7_2_io_o_4_out[3] ,
    \cb_7_2_io_o_4_out[2] ,
    \cb_7_2_io_o_4_out[1] ,
    \cb_7_2_io_o_4_out[0] }),
    .io_o_5_out({\cb_7_2_io_o_5_out[7] ,
    \cb_7_2_io_o_5_out[6] ,
    \cb_7_2_io_o_5_out[5] ,
    \cb_7_2_io_o_5_out[4] ,
    \cb_7_2_io_o_5_out[3] ,
    \cb_7_2_io_o_5_out[2] ,
    \cb_7_2_io_o_5_out[1] ,
    \cb_7_2_io_o_5_out[0] }),
    .io_o_6_out({\cb_7_2_io_o_6_out[7] ,
    \cb_7_2_io_o_6_out[6] ,
    \cb_7_2_io_o_6_out[5] ,
    \cb_7_2_io_o_6_out[4] ,
    \cb_7_2_io_o_6_out[3] ,
    \cb_7_2_io_o_6_out[2] ,
    \cb_7_2_io_o_6_out[1] ,
    \cb_7_2_io_o_6_out[0] }),
    .io_o_7_out({\cb_7_2_io_o_7_out[7] ,
    \cb_7_2_io_o_7_out[6] ,
    \cb_7_2_io_o_7_out[5] ,
    \cb_7_2_io_o_7_out[4] ,
    \cb_7_2_io_o_7_out[3] ,
    \cb_7_2_io_o_7_out[2] ,
    \cb_7_2_io_o_7_out[1] ,
    \cb_7_2_io_o_7_out[0] }),
    .io_wo({\cb_7_1_io_eo[63] ,
    \cb_7_1_io_eo[62] ,
    \cb_7_1_io_eo[61] ,
    \cb_7_1_io_eo[60] ,
    \cb_7_1_io_eo[59] ,
    \cb_7_1_io_eo[58] ,
    \cb_7_1_io_eo[57] ,
    \cb_7_1_io_eo[56] ,
    \cb_7_1_io_eo[55] ,
    \cb_7_1_io_eo[54] ,
    \cb_7_1_io_eo[53] ,
    \cb_7_1_io_eo[52] ,
    \cb_7_1_io_eo[51] ,
    \cb_7_1_io_eo[50] ,
    \cb_7_1_io_eo[49] ,
    \cb_7_1_io_eo[48] ,
    \cb_7_1_io_eo[47] ,
    \cb_7_1_io_eo[46] ,
    \cb_7_1_io_eo[45] ,
    \cb_7_1_io_eo[44] ,
    \cb_7_1_io_eo[43] ,
    \cb_7_1_io_eo[42] ,
    \cb_7_1_io_eo[41] ,
    \cb_7_1_io_eo[40] ,
    \cb_7_1_io_eo[39] ,
    \cb_7_1_io_eo[38] ,
    \cb_7_1_io_eo[37] ,
    \cb_7_1_io_eo[36] ,
    \cb_7_1_io_eo[35] ,
    \cb_7_1_io_eo[34] ,
    \cb_7_1_io_eo[33] ,
    \cb_7_1_io_eo[32] ,
    \cb_7_1_io_eo[31] ,
    \cb_7_1_io_eo[30] ,
    \cb_7_1_io_eo[29] ,
    \cb_7_1_io_eo[28] ,
    \cb_7_1_io_eo[27] ,
    \cb_7_1_io_eo[26] ,
    \cb_7_1_io_eo[25] ,
    \cb_7_1_io_eo[24] ,
    \cb_7_1_io_eo[23] ,
    \cb_7_1_io_eo[22] ,
    \cb_7_1_io_eo[21] ,
    \cb_7_1_io_eo[20] ,
    \cb_7_1_io_eo[19] ,
    \cb_7_1_io_eo[18] ,
    \cb_7_1_io_eo[17] ,
    \cb_7_1_io_eo[16] ,
    \cb_7_1_io_eo[15] ,
    \cb_7_1_io_eo[14] ,
    \cb_7_1_io_eo[13] ,
    \cb_7_1_io_eo[12] ,
    \cb_7_1_io_eo[11] ,
    \cb_7_1_io_eo[10] ,
    \cb_7_1_io_eo[9] ,
    \cb_7_1_io_eo[8] ,
    \cb_7_1_io_eo[7] ,
    \cb_7_1_io_eo[6] ,
    \cb_7_1_io_eo[5] ,
    \cb_7_1_io_eo[4] ,
    \cb_7_1_io_eo[3] ,
    \cb_7_1_io_eo[2] ,
    \cb_7_1_io_eo[1] ,
    \cb_7_1_io_eo[0] }));
 cic_block cb_7_3 (.io_cs_i(cb_7_3_io_cs_i),
    .io_i_0_ci(cb_7_2_io_o_0_co),
    .io_i_1_ci(cb_7_2_io_o_1_co),
    .io_i_2_ci(cb_7_2_io_o_2_co),
    .io_i_3_ci(cb_7_2_io_o_3_co),
    .io_i_4_ci(cb_7_2_io_o_4_co),
    .io_i_5_ci(cb_7_2_io_o_5_co),
    .io_i_6_ci(cb_7_2_io_o_6_co),
    .io_i_7_ci(cb_7_2_io_o_7_co),
    .io_o_0_co(cb_7_3_io_o_0_co),
    .io_o_1_co(cb_7_3_io_o_1_co),
    .io_o_2_co(cb_7_3_io_o_2_co),
    .io_o_3_co(cb_7_3_io_o_3_co),
    .io_o_4_co(cb_7_3_io_o_4_co),
    .io_o_5_co(cb_7_3_io_o_5_co),
    .io_o_6_co(cb_7_3_io_o_6_co),
    .io_o_7_co(cb_7_3_io_o_7_co),
    .io_vci(cb_7_2_io_vco),
    .io_vco(cb_7_3_io_vco),
    .io_vi(cb_7_3_io_vi),
    .io_we_i(cb_7_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_7_0_io_adr_i[1] ,
    \cb_7_0_io_adr_i[0] }),
    .io_dat_i({\cb_7_0_io_dat_i[15] ,
    \cb_7_0_io_dat_i[14] ,
    \cb_7_0_io_dat_i[13] ,
    \cb_7_0_io_dat_i[12] ,
    \cb_7_0_io_dat_i[11] ,
    \cb_7_0_io_dat_i[10] ,
    \cb_7_0_io_dat_i[9] ,
    \cb_7_0_io_dat_i[8] ,
    \cb_7_0_io_dat_i[7] ,
    \cb_7_0_io_dat_i[6] ,
    \cb_7_0_io_dat_i[5] ,
    \cb_7_0_io_dat_i[4] ,
    \cb_7_0_io_dat_i[3] ,
    \cb_7_0_io_dat_i[2] ,
    \cb_7_0_io_dat_i[1] ,
    \cb_7_0_io_dat_i[0] }),
    .io_dat_o({\cb_7_3_io_dat_o[15] ,
    \cb_7_3_io_dat_o[14] ,
    \cb_7_3_io_dat_o[13] ,
    \cb_7_3_io_dat_o[12] ,
    \cb_7_3_io_dat_o[11] ,
    \cb_7_3_io_dat_o[10] ,
    \cb_7_3_io_dat_o[9] ,
    \cb_7_3_io_dat_o[8] ,
    \cb_7_3_io_dat_o[7] ,
    \cb_7_3_io_dat_o[6] ,
    \cb_7_3_io_dat_o[5] ,
    \cb_7_3_io_dat_o[4] ,
    \cb_7_3_io_dat_o[3] ,
    \cb_7_3_io_dat_o[2] ,
    \cb_7_3_io_dat_o[1] ,
    \cb_7_3_io_dat_o[0] }),
    .io_eo({\cb_7_3_io_eo[63] ,
    \cb_7_3_io_eo[62] ,
    \cb_7_3_io_eo[61] ,
    \cb_7_3_io_eo[60] ,
    \cb_7_3_io_eo[59] ,
    \cb_7_3_io_eo[58] ,
    \cb_7_3_io_eo[57] ,
    \cb_7_3_io_eo[56] ,
    \cb_7_3_io_eo[55] ,
    \cb_7_3_io_eo[54] ,
    \cb_7_3_io_eo[53] ,
    \cb_7_3_io_eo[52] ,
    \cb_7_3_io_eo[51] ,
    \cb_7_3_io_eo[50] ,
    \cb_7_3_io_eo[49] ,
    \cb_7_3_io_eo[48] ,
    \cb_7_3_io_eo[47] ,
    \cb_7_3_io_eo[46] ,
    \cb_7_3_io_eo[45] ,
    \cb_7_3_io_eo[44] ,
    \cb_7_3_io_eo[43] ,
    \cb_7_3_io_eo[42] ,
    \cb_7_3_io_eo[41] ,
    \cb_7_3_io_eo[40] ,
    \cb_7_3_io_eo[39] ,
    \cb_7_3_io_eo[38] ,
    \cb_7_3_io_eo[37] ,
    \cb_7_3_io_eo[36] ,
    \cb_7_3_io_eo[35] ,
    \cb_7_3_io_eo[34] ,
    \cb_7_3_io_eo[33] ,
    \cb_7_3_io_eo[32] ,
    \cb_7_3_io_eo[31] ,
    \cb_7_3_io_eo[30] ,
    \cb_7_3_io_eo[29] ,
    \cb_7_3_io_eo[28] ,
    \cb_7_3_io_eo[27] ,
    \cb_7_3_io_eo[26] ,
    \cb_7_3_io_eo[25] ,
    \cb_7_3_io_eo[24] ,
    \cb_7_3_io_eo[23] ,
    \cb_7_3_io_eo[22] ,
    \cb_7_3_io_eo[21] ,
    \cb_7_3_io_eo[20] ,
    \cb_7_3_io_eo[19] ,
    \cb_7_3_io_eo[18] ,
    \cb_7_3_io_eo[17] ,
    \cb_7_3_io_eo[16] ,
    \cb_7_3_io_eo[15] ,
    \cb_7_3_io_eo[14] ,
    \cb_7_3_io_eo[13] ,
    \cb_7_3_io_eo[12] ,
    \cb_7_3_io_eo[11] ,
    \cb_7_3_io_eo[10] ,
    \cb_7_3_io_eo[9] ,
    \cb_7_3_io_eo[8] ,
    \cb_7_3_io_eo[7] ,
    \cb_7_3_io_eo[6] ,
    \cb_7_3_io_eo[5] ,
    \cb_7_3_io_eo[4] ,
    \cb_7_3_io_eo[3] ,
    \cb_7_3_io_eo[2] ,
    \cb_7_3_io_eo[1] ,
    \cb_7_3_io_eo[0] }),
    .io_i_0_in1({\cb_7_2_io_o_0_out[7] ,
    \cb_7_2_io_o_0_out[6] ,
    \cb_7_2_io_o_0_out[5] ,
    \cb_7_2_io_o_0_out[4] ,
    \cb_7_2_io_o_0_out[3] ,
    \cb_7_2_io_o_0_out[2] ,
    \cb_7_2_io_o_0_out[1] ,
    \cb_7_2_io_o_0_out[0] }),
    .io_i_1_in1({\cb_7_2_io_o_1_out[7] ,
    \cb_7_2_io_o_1_out[6] ,
    \cb_7_2_io_o_1_out[5] ,
    \cb_7_2_io_o_1_out[4] ,
    \cb_7_2_io_o_1_out[3] ,
    \cb_7_2_io_o_1_out[2] ,
    \cb_7_2_io_o_1_out[1] ,
    \cb_7_2_io_o_1_out[0] }),
    .io_i_2_in1({\cb_7_2_io_o_2_out[7] ,
    \cb_7_2_io_o_2_out[6] ,
    \cb_7_2_io_o_2_out[5] ,
    \cb_7_2_io_o_2_out[4] ,
    \cb_7_2_io_o_2_out[3] ,
    \cb_7_2_io_o_2_out[2] ,
    \cb_7_2_io_o_2_out[1] ,
    \cb_7_2_io_o_2_out[0] }),
    .io_i_3_in1({\cb_7_2_io_o_3_out[7] ,
    \cb_7_2_io_o_3_out[6] ,
    \cb_7_2_io_o_3_out[5] ,
    \cb_7_2_io_o_3_out[4] ,
    \cb_7_2_io_o_3_out[3] ,
    \cb_7_2_io_o_3_out[2] ,
    \cb_7_2_io_o_3_out[1] ,
    \cb_7_2_io_o_3_out[0] }),
    .io_i_4_in1({\cb_7_2_io_o_4_out[7] ,
    \cb_7_2_io_o_4_out[6] ,
    \cb_7_2_io_o_4_out[5] ,
    \cb_7_2_io_o_4_out[4] ,
    \cb_7_2_io_o_4_out[3] ,
    \cb_7_2_io_o_4_out[2] ,
    \cb_7_2_io_o_4_out[1] ,
    \cb_7_2_io_o_4_out[0] }),
    .io_i_5_in1({\cb_7_2_io_o_5_out[7] ,
    \cb_7_2_io_o_5_out[6] ,
    \cb_7_2_io_o_5_out[5] ,
    \cb_7_2_io_o_5_out[4] ,
    \cb_7_2_io_o_5_out[3] ,
    \cb_7_2_io_o_5_out[2] ,
    \cb_7_2_io_o_5_out[1] ,
    \cb_7_2_io_o_5_out[0] }),
    .io_i_6_in1({\cb_7_2_io_o_6_out[7] ,
    \cb_7_2_io_o_6_out[6] ,
    \cb_7_2_io_o_6_out[5] ,
    \cb_7_2_io_o_6_out[4] ,
    \cb_7_2_io_o_6_out[3] ,
    \cb_7_2_io_o_6_out[2] ,
    \cb_7_2_io_o_6_out[1] ,
    \cb_7_2_io_o_6_out[0] }),
    .io_i_7_in1({\cb_7_2_io_o_7_out[7] ,
    \cb_7_2_io_o_7_out[6] ,
    \cb_7_2_io_o_7_out[5] ,
    \cb_7_2_io_o_7_out[4] ,
    \cb_7_2_io_o_7_out[3] ,
    \cb_7_2_io_o_7_out[2] ,
    \cb_7_2_io_o_7_out[1] ,
    \cb_7_2_io_o_7_out[0] }),
    .io_o_0_out({\cb_7_3_io_o_0_out[7] ,
    \cb_7_3_io_o_0_out[6] ,
    \cb_7_3_io_o_0_out[5] ,
    \cb_7_3_io_o_0_out[4] ,
    \cb_7_3_io_o_0_out[3] ,
    \cb_7_3_io_o_0_out[2] ,
    \cb_7_3_io_o_0_out[1] ,
    \cb_7_3_io_o_0_out[0] }),
    .io_o_1_out({\cb_7_3_io_o_1_out[7] ,
    \cb_7_3_io_o_1_out[6] ,
    \cb_7_3_io_o_1_out[5] ,
    \cb_7_3_io_o_1_out[4] ,
    \cb_7_3_io_o_1_out[3] ,
    \cb_7_3_io_o_1_out[2] ,
    \cb_7_3_io_o_1_out[1] ,
    \cb_7_3_io_o_1_out[0] }),
    .io_o_2_out({\cb_7_3_io_o_2_out[7] ,
    \cb_7_3_io_o_2_out[6] ,
    \cb_7_3_io_o_2_out[5] ,
    \cb_7_3_io_o_2_out[4] ,
    \cb_7_3_io_o_2_out[3] ,
    \cb_7_3_io_o_2_out[2] ,
    \cb_7_3_io_o_2_out[1] ,
    \cb_7_3_io_o_2_out[0] }),
    .io_o_3_out({\cb_7_3_io_o_3_out[7] ,
    \cb_7_3_io_o_3_out[6] ,
    \cb_7_3_io_o_3_out[5] ,
    \cb_7_3_io_o_3_out[4] ,
    \cb_7_3_io_o_3_out[3] ,
    \cb_7_3_io_o_3_out[2] ,
    \cb_7_3_io_o_3_out[1] ,
    \cb_7_3_io_o_3_out[0] }),
    .io_o_4_out({\cb_7_3_io_o_4_out[7] ,
    \cb_7_3_io_o_4_out[6] ,
    \cb_7_3_io_o_4_out[5] ,
    \cb_7_3_io_o_4_out[4] ,
    \cb_7_3_io_o_4_out[3] ,
    \cb_7_3_io_o_4_out[2] ,
    \cb_7_3_io_o_4_out[1] ,
    \cb_7_3_io_o_4_out[0] }),
    .io_o_5_out({\cb_7_3_io_o_5_out[7] ,
    \cb_7_3_io_o_5_out[6] ,
    \cb_7_3_io_o_5_out[5] ,
    \cb_7_3_io_o_5_out[4] ,
    \cb_7_3_io_o_5_out[3] ,
    \cb_7_3_io_o_5_out[2] ,
    \cb_7_3_io_o_5_out[1] ,
    \cb_7_3_io_o_5_out[0] }),
    .io_o_6_out({\cb_7_3_io_o_6_out[7] ,
    \cb_7_3_io_o_6_out[6] ,
    \cb_7_3_io_o_6_out[5] ,
    \cb_7_3_io_o_6_out[4] ,
    \cb_7_3_io_o_6_out[3] ,
    \cb_7_3_io_o_6_out[2] ,
    \cb_7_3_io_o_6_out[1] ,
    \cb_7_3_io_o_6_out[0] }),
    .io_o_7_out({\cb_7_3_io_o_7_out[7] ,
    \cb_7_3_io_o_7_out[6] ,
    \cb_7_3_io_o_7_out[5] ,
    \cb_7_3_io_o_7_out[4] ,
    \cb_7_3_io_o_7_out[3] ,
    \cb_7_3_io_o_7_out[2] ,
    \cb_7_3_io_o_7_out[1] ,
    \cb_7_3_io_o_7_out[0] }),
    .io_wo({\cb_7_2_io_eo[63] ,
    \cb_7_2_io_eo[62] ,
    \cb_7_2_io_eo[61] ,
    \cb_7_2_io_eo[60] ,
    \cb_7_2_io_eo[59] ,
    \cb_7_2_io_eo[58] ,
    \cb_7_2_io_eo[57] ,
    \cb_7_2_io_eo[56] ,
    \cb_7_2_io_eo[55] ,
    \cb_7_2_io_eo[54] ,
    \cb_7_2_io_eo[53] ,
    \cb_7_2_io_eo[52] ,
    \cb_7_2_io_eo[51] ,
    \cb_7_2_io_eo[50] ,
    \cb_7_2_io_eo[49] ,
    \cb_7_2_io_eo[48] ,
    \cb_7_2_io_eo[47] ,
    \cb_7_2_io_eo[46] ,
    \cb_7_2_io_eo[45] ,
    \cb_7_2_io_eo[44] ,
    \cb_7_2_io_eo[43] ,
    \cb_7_2_io_eo[42] ,
    \cb_7_2_io_eo[41] ,
    \cb_7_2_io_eo[40] ,
    \cb_7_2_io_eo[39] ,
    \cb_7_2_io_eo[38] ,
    \cb_7_2_io_eo[37] ,
    \cb_7_2_io_eo[36] ,
    \cb_7_2_io_eo[35] ,
    \cb_7_2_io_eo[34] ,
    \cb_7_2_io_eo[33] ,
    \cb_7_2_io_eo[32] ,
    \cb_7_2_io_eo[31] ,
    \cb_7_2_io_eo[30] ,
    \cb_7_2_io_eo[29] ,
    \cb_7_2_io_eo[28] ,
    \cb_7_2_io_eo[27] ,
    \cb_7_2_io_eo[26] ,
    \cb_7_2_io_eo[25] ,
    \cb_7_2_io_eo[24] ,
    \cb_7_2_io_eo[23] ,
    \cb_7_2_io_eo[22] ,
    \cb_7_2_io_eo[21] ,
    \cb_7_2_io_eo[20] ,
    \cb_7_2_io_eo[19] ,
    \cb_7_2_io_eo[18] ,
    \cb_7_2_io_eo[17] ,
    \cb_7_2_io_eo[16] ,
    \cb_7_2_io_eo[15] ,
    \cb_7_2_io_eo[14] ,
    \cb_7_2_io_eo[13] ,
    \cb_7_2_io_eo[12] ,
    \cb_7_2_io_eo[11] ,
    \cb_7_2_io_eo[10] ,
    \cb_7_2_io_eo[9] ,
    \cb_7_2_io_eo[8] ,
    \cb_7_2_io_eo[7] ,
    \cb_7_2_io_eo[6] ,
    \cb_7_2_io_eo[5] ,
    \cb_7_2_io_eo[4] ,
    \cb_7_2_io_eo[3] ,
    \cb_7_2_io_eo[2] ,
    \cb_7_2_io_eo[1] ,
    \cb_7_2_io_eo[0] }));
 cic_block cb_7_4 (.io_cs_i(cb_7_4_io_cs_i),
    .io_i_0_ci(cb_7_3_io_o_0_co),
    .io_i_1_ci(cb_7_3_io_o_1_co),
    .io_i_2_ci(cb_7_3_io_o_2_co),
    .io_i_3_ci(cb_7_3_io_o_3_co),
    .io_i_4_ci(cb_7_3_io_o_4_co),
    .io_i_5_ci(cb_7_3_io_o_5_co),
    .io_i_6_ci(cb_7_3_io_o_6_co),
    .io_i_7_ci(cb_7_3_io_o_7_co),
    .io_o_0_co(cb_7_4_io_o_0_co),
    .io_o_1_co(cb_7_4_io_o_1_co),
    .io_o_2_co(cb_7_4_io_o_2_co),
    .io_o_3_co(cb_7_4_io_o_3_co),
    .io_o_4_co(cb_7_4_io_o_4_co),
    .io_o_5_co(cb_7_4_io_o_5_co),
    .io_o_6_co(cb_7_4_io_o_6_co),
    .io_o_7_co(cb_7_4_io_o_7_co),
    .io_vci(cb_7_3_io_vco),
    .io_vco(cb_7_4_io_vco),
    .io_vi(cb_7_4_io_vi),
    .io_we_i(cb_7_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_7_0_io_adr_i[1] ,
    \cb_7_0_io_adr_i[0] }),
    .io_dat_i({\cb_7_0_io_dat_i[15] ,
    \cb_7_0_io_dat_i[14] ,
    \cb_7_0_io_dat_i[13] ,
    \cb_7_0_io_dat_i[12] ,
    \cb_7_0_io_dat_i[11] ,
    \cb_7_0_io_dat_i[10] ,
    \cb_7_0_io_dat_i[9] ,
    \cb_7_0_io_dat_i[8] ,
    \cb_7_0_io_dat_i[7] ,
    \cb_7_0_io_dat_i[6] ,
    \cb_7_0_io_dat_i[5] ,
    \cb_7_0_io_dat_i[4] ,
    \cb_7_0_io_dat_i[3] ,
    \cb_7_0_io_dat_i[2] ,
    \cb_7_0_io_dat_i[1] ,
    \cb_7_0_io_dat_i[0] }),
    .io_dat_o({\cb_7_4_io_dat_o[15] ,
    \cb_7_4_io_dat_o[14] ,
    \cb_7_4_io_dat_o[13] ,
    \cb_7_4_io_dat_o[12] ,
    \cb_7_4_io_dat_o[11] ,
    \cb_7_4_io_dat_o[10] ,
    \cb_7_4_io_dat_o[9] ,
    \cb_7_4_io_dat_o[8] ,
    \cb_7_4_io_dat_o[7] ,
    \cb_7_4_io_dat_o[6] ,
    \cb_7_4_io_dat_o[5] ,
    \cb_7_4_io_dat_o[4] ,
    \cb_7_4_io_dat_o[3] ,
    \cb_7_4_io_dat_o[2] ,
    \cb_7_4_io_dat_o[1] ,
    \cb_7_4_io_dat_o[0] }),
    .io_eo({\cb_7_4_io_eo[63] ,
    \cb_7_4_io_eo[62] ,
    \cb_7_4_io_eo[61] ,
    \cb_7_4_io_eo[60] ,
    \cb_7_4_io_eo[59] ,
    \cb_7_4_io_eo[58] ,
    \cb_7_4_io_eo[57] ,
    \cb_7_4_io_eo[56] ,
    \cb_7_4_io_eo[55] ,
    \cb_7_4_io_eo[54] ,
    \cb_7_4_io_eo[53] ,
    \cb_7_4_io_eo[52] ,
    \cb_7_4_io_eo[51] ,
    \cb_7_4_io_eo[50] ,
    \cb_7_4_io_eo[49] ,
    \cb_7_4_io_eo[48] ,
    \cb_7_4_io_eo[47] ,
    \cb_7_4_io_eo[46] ,
    \cb_7_4_io_eo[45] ,
    \cb_7_4_io_eo[44] ,
    \cb_7_4_io_eo[43] ,
    \cb_7_4_io_eo[42] ,
    \cb_7_4_io_eo[41] ,
    \cb_7_4_io_eo[40] ,
    \cb_7_4_io_eo[39] ,
    \cb_7_4_io_eo[38] ,
    \cb_7_4_io_eo[37] ,
    \cb_7_4_io_eo[36] ,
    \cb_7_4_io_eo[35] ,
    \cb_7_4_io_eo[34] ,
    \cb_7_4_io_eo[33] ,
    \cb_7_4_io_eo[32] ,
    \cb_7_4_io_eo[31] ,
    \cb_7_4_io_eo[30] ,
    \cb_7_4_io_eo[29] ,
    \cb_7_4_io_eo[28] ,
    \cb_7_4_io_eo[27] ,
    \cb_7_4_io_eo[26] ,
    \cb_7_4_io_eo[25] ,
    \cb_7_4_io_eo[24] ,
    \cb_7_4_io_eo[23] ,
    \cb_7_4_io_eo[22] ,
    \cb_7_4_io_eo[21] ,
    \cb_7_4_io_eo[20] ,
    \cb_7_4_io_eo[19] ,
    \cb_7_4_io_eo[18] ,
    \cb_7_4_io_eo[17] ,
    \cb_7_4_io_eo[16] ,
    \cb_7_4_io_eo[15] ,
    \cb_7_4_io_eo[14] ,
    \cb_7_4_io_eo[13] ,
    \cb_7_4_io_eo[12] ,
    \cb_7_4_io_eo[11] ,
    \cb_7_4_io_eo[10] ,
    \cb_7_4_io_eo[9] ,
    \cb_7_4_io_eo[8] ,
    \cb_7_4_io_eo[7] ,
    \cb_7_4_io_eo[6] ,
    \cb_7_4_io_eo[5] ,
    \cb_7_4_io_eo[4] ,
    \cb_7_4_io_eo[3] ,
    \cb_7_4_io_eo[2] ,
    \cb_7_4_io_eo[1] ,
    \cb_7_4_io_eo[0] }),
    .io_i_0_in1({\cb_7_3_io_o_0_out[7] ,
    \cb_7_3_io_o_0_out[6] ,
    \cb_7_3_io_o_0_out[5] ,
    \cb_7_3_io_o_0_out[4] ,
    \cb_7_3_io_o_0_out[3] ,
    \cb_7_3_io_o_0_out[2] ,
    \cb_7_3_io_o_0_out[1] ,
    \cb_7_3_io_o_0_out[0] }),
    .io_i_1_in1({\cb_7_3_io_o_1_out[7] ,
    \cb_7_3_io_o_1_out[6] ,
    \cb_7_3_io_o_1_out[5] ,
    \cb_7_3_io_o_1_out[4] ,
    \cb_7_3_io_o_1_out[3] ,
    \cb_7_3_io_o_1_out[2] ,
    \cb_7_3_io_o_1_out[1] ,
    \cb_7_3_io_o_1_out[0] }),
    .io_i_2_in1({\cb_7_3_io_o_2_out[7] ,
    \cb_7_3_io_o_2_out[6] ,
    \cb_7_3_io_o_2_out[5] ,
    \cb_7_3_io_o_2_out[4] ,
    \cb_7_3_io_o_2_out[3] ,
    \cb_7_3_io_o_2_out[2] ,
    \cb_7_3_io_o_2_out[1] ,
    \cb_7_3_io_o_2_out[0] }),
    .io_i_3_in1({\cb_7_3_io_o_3_out[7] ,
    \cb_7_3_io_o_3_out[6] ,
    \cb_7_3_io_o_3_out[5] ,
    \cb_7_3_io_o_3_out[4] ,
    \cb_7_3_io_o_3_out[3] ,
    \cb_7_3_io_o_3_out[2] ,
    \cb_7_3_io_o_3_out[1] ,
    \cb_7_3_io_o_3_out[0] }),
    .io_i_4_in1({\cb_7_3_io_o_4_out[7] ,
    \cb_7_3_io_o_4_out[6] ,
    \cb_7_3_io_o_4_out[5] ,
    \cb_7_3_io_o_4_out[4] ,
    \cb_7_3_io_o_4_out[3] ,
    \cb_7_3_io_o_4_out[2] ,
    \cb_7_3_io_o_4_out[1] ,
    \cb_7_3_io_o_4_out[0] }),
    .io_i_5_in1({\cb_7_3_io_o_5_out[7] ,
    \cb_7_3_io_o_5_out[6] ,
    \cb_7_3_io_o_5_out[5] ,
    \cb_7_3_io_o_5_out[4] ,
    \cb_7_3_io_o_5_out[3] ,
    \cb_7_3_io_o_5_out[2] ,
    \cb_7_3_io_o_5_out[1] ,
    \cb_7_3_io_o_5_out[0] }),
    .io_i_6_in1({\cb_7_3_io_o_6_out[7] ,
    \cb_7_3_io_o_6_out[6] ,
    \cb_7_3_io_o_6_out[5] ,
    \cb_7_3_io_o_6_out[4] ,
    \cb_7_3_io_o_6_out[3] ,
    \cb_7_3_io_o_6_out[2] ,
    \cb_7_3_io_o_6_out[1] ,
    \cb_7_3_io_o_6_out[0] }),
    .io_i_7_in1({\cb_7_3_io_o_7_out[7] ,
    \cb_7_3_io_o_7_out[6] ,
    \cb_7_3_io_o_7_out[5] ,
    \cb_7_3_io_o_7_out[4] ,
    \cb_7_3_io_o_7_out[3] ,
    \cb_7_3_io_o_7_out[2] ,
    \cb_7_3_io_o_7_out[1] ,
    \cb_7_3_io_o_7_out[0] }),
    .io_o_0_out({\cb_7_4_io_o_0_out[7] ,
    \cb_7_4_io_o_0_out[6] ,
    \cb_7_4_io_o_0_out[5] ,
    \cb_7_4_io_o_0_out[4] ,
    \cb_7_4_io_o_0_out[3] ,
    \cb_7_4_io_o_0_out[2] ,
    \cb_7_4_io_o_0_out[1] ,
    \cb_7_4_io_o_0_out[0] }),
    .io_o_1_out({\cb_7_4_io_o_1_out[7] ,
    \cb_7_4_io_o_1_out[6] ,
    \cb_7_4_io_o_1_out[5] ,
    \cb_7_4_io_o_1_out[4] ,
    \cb_7_4_io_o_1_out[3] ,
    \cb_7_4_io_o_1_out[2] ,
    \cb_7_4_io_o_1_out[1] ,
    \cb_7_4_io_o_1_out[0] }),
    .io_o_2_out({\cb_7_4_io_o_2_out[7] ,
    \cb_7_4_io_o_2_out[6] ,
    \cb_7_4_io_o_2_out[5] ,
    \cb_7_4_io_o_2_out[4] ,
    \cb_7_4_io_o_2_out[3] ,
    \cb_7_4_io_o_2_out[2] ,
    \cb_7_4_io_o_2_out[1] ,
    \cb_7_4_io_o_2_out[0] }),
    .io_o_3_out({\cb_7_4_io_o_3_out[7] ,
    \cb_7_4_io_o_3_out[6] ,
    \cb_7_4_io_o_3_out[5] ,
    \cb_7_4_io_o_3_out[4] ,
    \cb_7_4_io_o_3_out[3] ,
    \cb_7_4_io_o_3_out[2] ,
    \cb_7_4_io_o_3_out[1] ,
    \cb_7_4_io_o_3_out[0] }),
    .io_o_4_out({\cb_7_4_io_o_4_out[7] ,
    \cb_7_4_io_o_4_out[6] ,
    \cb_7_4_io_o_4_out[5] ,
    \cb_7_4_io_o_4_out[4] ,
    \cb_7_4_io_o_4_out[3] ,
    \cb_7_4_io_o_4_out[2] ,
    \cb_7_4_io_o_4_out[1] ,
    \cb_7_4_io_o_4_out[0] }),
    .io_o_5_out({\cb_7_4_io_o_5_out[7] ,
    \cb_7_4_io_o_5_out[6] ,
    \cb_7_4_io_o_5_out[5] ,
    \cb_7_4_io_o_5_out[4] ,
    \cb_7_4_io_o_5_out[3] ,
    \cb_7_4_io_o_5_out[2] ,
    \cb_7_4_io_o_5_out[1] ,
    \cb_7_4_io_o_5_out[0] }),
    .io_o_6_out({\cb_7_4_io_o_6_out[7] ,
    \cb_7_4_io_o_6_out[6] ,
    \cb_7_4_io_o_6_out[5] ,
    \cb_7_4_io_o_6_out[4] ,
    \cb_7_4_io_o_6_out[3] ,
    \cb_7_4_io_o_6_out[2] ,
    \cb_7_4_io_o_6_out[1] ,
    \cb_7_4_io_o_6_out[0] }),
    .io_o_7_out({\cb_7_4_io_o_7_out[7] ,
    \cb_7_4_io_o_7_out[6] ,
    \cb_7_4_io_o_7_out[5] ,
    \cb_7_4_io_o_7_out[4] ,
    \cb_7_4_io_o_7_out[3] ,
    \cb_7_4_io_o_7_out[2] ,
    \cb_7_4_io_o_7_out[1] ,
    \cb_7_4_io_o_7_out[0] }),
    .io_wo({\cb_7_3_io_eo[63] ,
    \cb_7_3_io_eo[62] ,
    \cb_7_3_io_eo[61] ,
    \cb_7_3_io_eo[60] ,
    \cb_7_3_io_eo[59] ,
    \cb_7_3_io_eo[58] ,
    \cb_7_3_io_eo[57] ,
    \cb_7_3_io_eo[56] ,
    \cb_7_3_io_eo[55] ,
    \cb_7_3_io_eo[54] ,
    \cb_7_3_io_eo[53] ,
    \cb_7_3_io_eo[52] ,
    \cb_7_3_io_eo[51] ,
    \cb_7_3_io_eo[50] ,
    \cb_7_3_io_eo[49] ,
    \cb_7_3_io_eo[48] ,
    \cb_7_3_io_eo[47] ,
    \cb_7_3_io_eo[46] ,
    \cb_7_3_io_eo[45] ,
    \cb_7_3_io_eo[44] ,
    \cb_7_3_io_eo[43] ,
    \cb_7_3_io_eo[42] ,
    \cb_7_3_io_eo[41] ,
    \cb_7_3_io_eo[40] ,
    \cb_7_3_io_eo[39] ,
    \cb_7_3_io_eo[38] ,
    \cb_7_3_io_eo[37] ,
    \cb_7_3_io_eo[36] ,
    \cb_7_3_io_eo[35] ,
    \cb_7_3_io_eo[34] ,
    \cb_7_3_io_eo[33] ,
    \cb_7_3_io_eo[32] ,
    \cb_7_3_io_eo[31] ,
    \cb_7_3_io_eo[30] ,
    \cb_7_3_io_eo[29] ,
    \cb_7_3_io_eo[28] ,
    \cb_7_3_io_eo[27] ,
    \cb_7_3_io_eo[26] ,
    \cb_7_3_io_eo[25] ,
    \cb_7_3_io_eo[24] ,
    \cb_7_3_io_eo[23] ,
    \cb_7_3_io_eo[22] ,
    \cb_7_3_io_eo[21] ,
    \cb_7_3_io_eo[20] ,
    \cb_7_3_io_eo[19] ,
    \cb_7_3_io_eo[18] ,
    \cb_7_3_io_eo[17] ,
    \cb_7_3_io_eo[16] ,
    \cb_7_3_io_eo[15] ,
    \cb_7_3_io_eo[14] ,
    \cb_7_3_io_eo[13] ,
    \cb_7_3_io_eo[12] ,
    \cb_7_3_io_eo[11] ,
    \cb_7_3_io_eo[10] ,
    \cb_7_3_io_eo[9] ,
    \cb_7_3_io_eo[8] ,
    \cb_7_3_io_eo[7] ,
    \cb_7_3_io_eo[6] ,
    \cb_7_3_io_eo[5] ,
    \cb_7_3_io_eo[4] ,
    \cb_7_3_io_eo[3] ,
    \cb_7_3_io_eo[2] ,
    \cb_7_3_io_eo[1] ,
    \cb_7_3_io_eo[0] }));
 cic_block cb_7_5 (.io_cs_i(cb_7_5_io_cs_i),
    .io_i_0_ci(cb_7_4_io_o_0_co),
    .io_i_1_ci(cb_7_4_io_o_1_co),
    .io_i_2_ci(cb_7_4_io_o_2_co),
    .io_i_3_ci(cb_7_4_io_o_3_co),
    .io_i_4_ci(cb_7_4_io_o_4_co),
    .io_i_5_ci(cb_7_4_io_o_5_co),
    .io_i_6_ci(cb_7_4_io_o_6_co),
    .io_i_7_ci(cb_7_4_io_o_7_co),
    .io_o_0_co(cb_7_5_io_o_0_co),
    .io_o_1_co(cb_7_5_io_o_1_co),
    .io_o_2_co(cb_7_5_io_o_2_co),
    .io_o_3_co(cb_7_5_io_o_3_co),
    .io_o_4_co(cb_7_5_io_o_4_co),
    .io_o_5_co(cb_7_5_io_o_5_co),
    .io_o_6_co(cb_7_5_io_o_6_co),
    .io_o_7_co(cb_7_5_io_o_7_co),
    .io_vci(cb_7_4_io_vco),
    .io_vco(cb_7_5_io_vco),
    .io_vi(cb_7_5_io_vi),
    .io_we_i(cb_7_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_7_0_io_adr_i[1] ,
    \cb_7_0_io_adr_i[0] }),
    .io_dat_i({\cb_7_0_io_dat_i[15] ,
    \cb_7_0_io_dat_i[14] ,
    \cb_7_0_io_dat_i[13] ,
    \cb_7_0_io_dat_i[12] ,
    \cb_7_0_io_dat_i[11] ,
    \cb_7_0_io_dat_i[10] ,
    \cb_7_0_io_dat_i[9] ,
    \cb_7_0_io_dat_i[8] ,
    \cb_7_0_io_dat_i[7] ,
    \cb_7_0_io_dat_i[6] ,
    \cb_7_0_io_dat_i[5] ,
    \cb_7_0_io_dat_i[4] ,
    \cb_7_0_io_dat_i[3] ,
    \cb_7_0_io_dat_i[2] ,
    \cb_7_0_io_dat_i[1] ,
    \cb_7_0_io_dat_i[0] }),
    .io_dat_o({\cb_7_5_io_dat_o[15] ,
    \cb_7_5_io_dat_o[14] ,
    \cb_7_5_io_dat_o[13] ,
    \cb_7_5_io_dat_o[12] ,
    \cb_7_5_io_dat_o[11] ,
    \cb_7_5_io_dat_o[10] ,
    \cb_7_5_io_dat_o[9] ,
    \cb_7_5_io_dat_o[8] ,
    \cb_7_5_io_dat_o[7] ,
    \cb_7_5_io_dat_o[6] ,
    \cb_7_5_io_dat_o[5] ,
    \cb_7_5_io_dat_o[4] ,
    \cb_7_5_io_dat_o[3] ,
    \cb_7_5_io_dat_o[2] ,
    \cb_7_5_io_dat_o[1] ,
    \cb_7_5_io_dat_o[0] }),
    .io_eo({\cb_7_5_io_eo[63] ,
    \cb_7_5_io_eo[62] ,
    \cb_7_5_io_eo[61] ,
    \cb_7_5_io_eo[60] ,
    \cb_7_5_io_eo[59] ,
    \cb_7_5_io_eo[58] ,
    \cb_7_5_io_eo[57] ,
    \cb_7_5_io_eo[56] ,
    \cb_7_5_io_eo[55] ,
    \cb_7_5_io_eo[54] ,
    \cb_7_5_io_eo[53] ,
    \cb_7_5_io_eo[52] ,
    \cb_7_5_io_eo[51] ,
    \cb_7_5_io_eo[50] ,
    \cb_7_5_io_eo[49] ,
    \cb_7_5_io_eo[48] ,
    \cb_7_5_io_eo[47] ,
    \cb_7_5_io_eo[46] ,
    \cb_7_5_io_eo[45] ,
    \cb_7_5_io_eo[44] ,
    \cb_7_5_io_eo[43] ,
    \cb_7_5_io_eo[42] ,
    \cb_7_5_io_eo[41] ,
    \cb_7_5_io_eo[40] ,
    \cb_7_5_io_eo[39] ,
    \cb_7_5_io_eo[38] ,
    \cb_7_5_io_eo[37] ,
    \cb_7_5_io_eo[36] ,
    \cb_7_5_io_eo[35] ,
    \cb_7_5_io_eo[34] ,
    \cb_7_5_io_eo[33] ,
    \cb_7_5_io_eo[32] ,
    \cb_7_5_io_eo[31] ,
    \cb_7_5_io_eo[30] ,
    \cb_7_5_io_eo[29] ,
    \cb_7_5_io_eo[28] ,
    \cb_7_5_io_eo[27] ,
    \cb_7_5_io_eo[26] ,
    \cb_7_5_io_eo[25] ,
    \cb_7_5_io_eo[24] ,
    \cb_7_5_io_eo[23] ,
    \cb_7_5_io_eo[22] ,
    \cb_7_5_io_eo[21] ,
    \cb_7_5_io_eo[20] ,
    \cb_7_5_io_eo[19] ,
    \cb_7_5_io_eo[18] ,
    \cb_7_5_io_eo[17] ,
    \cb_7_5_io_eo[16] ,
    \cb_7_5_io_eo[15] ,
    \cb_7_5_io_eo[14] ,
    \cb_7_5_io_eo[13] ,
    \cb_7_5_io_eo[12] ,
    \cb_7_5_io_eo[11] ,
    \cb_7_5_io_eo[10] ,
    \cb_7_5_io_eo[9] ,
    \cb_7_5_io_eo[8] ,
    \cb_7_5_io_eo[7] ,
    \cb_7_5_io_eo[6] ,
    \cb_7_5_io_eo[5] ,
    \cb_7_5_io_eo[4] ,
    \cb_7_5_io_eo[3] ,
    \cb_7_5_io_eo[2] ,
    \cb_7_5_io_eo[1] ,
    \cb_7_5_io_eo[0] }),
    .io_i_0_in1({\cb_7_4_io_o_0_out[7] ,
    \cb_7_4_io_o_0_out[6] ,
    \cb_7_4_io_o_0_out[5] ,
    \cb_7_4_io_o_0_out[4] ,
    \cb_7_4_io_o_0_out[3] ,
    \cb_7_4_io_o_0_out[2] ,
    \cb_7_4_io_o_0_out[1] ,
    \cb_7_4_io_o_0_out[0] }),
    .io_i_1_in1({\cb_7_4_io_o_1_out[7] ,
    \cb_7_4_io_o_1_out[6] ,
    \cb_7_4_io_o_1_out[5] ,
    \cb_7_4_io_o_1_out[4] ,
    \cb_7_4_io_o_1_out[3] ,
    \cb_7_4_io_o_1_out[2] ,
    \cb_7_4_io_o_1_out[1] ,
    \cb_7_4_io_o_1_out[0] }),
    .io_i_2_in1({\cb_7_4_io_o_2_out[7] ,
    \cb_7_4_io_o_2_out[6] ,
    \cb_7_4_io_o_2_out[5] ,
    \cb_7_4_io_o_2_out[4] ,
    \cb_7_4_io_o_2_out[3] ,
    \cb_7_4_io_o_2_out[2] ,
    \cb_7_4_io_o_2_out[1] ,
    \cb_7_4_io_o_2_out[0] }),
    .io_i_3_in1({\cb_7_4_io_o_3_out[7] ,
    \cb_7_4_io_o_3_out[6] ,
    \cb_7_4_io_o_3_out[5] ,
    \cb_7_4_io_o_3_out[4] ,
    \cb_7_4_io_o_3_out[3] ,
    \cb_7_4_io_o_3_out[2] ,
    \cb_7_4_io_o_3_out[1] ,
    \cb_7_4_io_o_3_out[0] }),
    .io_i_4_in1({\cb_7_4_io_o_4_out[7] ,
    \cb_7_4_io_o_4_out[6] ,
    \cb_7_4_io_o_4_out[5] ,
    \cb_7_4_io_o_4_out[4] ,
    \cb_7_4_io_o_4_out[3] ,
    \cb_7_4_io_o_4_out[2] ,
    \cb_7_4_io_o_4_out[1] ,
    \cb_7_4_io_o_4_out[0] }),
    .io_i_5_in1({\cb_7_4_io_o_5_out[7] ,
    \cb_7_4_io_o_5_out[6] ,
    \cb_7_4_io_o_5_out[5] ,
    \cb_7_4_io_o_5_out[4] ,
    \cb_7_4_io_o_5_out[3] ,
    \cb_7_4_io_o_5_out[2] ,
    \cb_7_4_io_o_5_out[1] ,
    \cb_7_4_io_o_5_out[0] }),
    .io_i_6_in1({\cb_7_4_io_o_6_out[7] ,
    \cb_7_4_io_o_6_out[6] ,
    \cb_7_4_io_o_6_out[5] ,
    \cb_7_4_io_o_6_out[4] ,
    \cb_7_4_io_o_6_out[3] ,
    \cb_7_4_io_o_6_out[2] ,
    \cb_7_4_io_o_6_out[1] ,
    \cb_7_4_io_o_6_out[0] }),
    .io_i_7_in1({\cb_7_4_io_o_7_out[7] ,
    \cb_7_4_io_o_7_out[6] ,
    \cb_7_4_io_o_7_out[5] ,
    \cb_7_4_io_o_7_out[4] ,
    \cb_7_4_io_o_7_out[3] ,
    \cb_7_4_io_o_7_out[2] ,
    \cb_7_4_io_o_7_out[1] ,
    \cb_7_4_io_o_7_out[0] }),
    .io_o_0_out({\cb_7_5_io_o_0_out[7] ,
    \cb_7_5_io_o_0_out[6] ,
    \cb_7_5_io_o_0_out[5] ,
    \cb_7_5_io_o_0_out[4] ,
    \cb_7_5_io_o_0_out[3] ,
    \cb_7_5_io_o_0_out[2] ,
    \cb_7_5_io_o_0_out[1] ,
    \cb_7_5_io_o_0_out[0] }),
    .io_o_1_out({\cb_7_5_io_o_1_out[7] ,
    \cb_7_5_io_o_1_out[6] ,
    \cb_7_5_io_o_1_out[5] ,
    \cb_7_5_io_o_1_out[4] ,
    \cb_7_5_io_o_1_out[3] ,
    \cb_7_5_io_o_1_out[2] ,
    \cb_7_5_io_o_1_out[1] ,
    \cb_7_5_io_o_1_out[0] }),
    .io_o_2_out({\cb_7_5_io_o_2_out[7] ,
    \cb_7_5_io_o_2_out[6] ,
    \cb_7_5_io_o_2_out[5] ,
    \cb_7_5_io_o_2_out[4] ,
    \cb_7_5_io_o_2_out[3] ,
    \cb_7_5_io_o_2_out[2] ,
    \cb_7_5_io_o_2_out[1] ,
    \cb_7_5_io_o_2_out[0] }),
    .io_o_3_out({\cb_7_5_io_o_3_out[7] ,
    \cb_7_5_io_o_3_out[6] ,
    \cb_7_5_io_o_3_out[5] ,
    \cb_7_5_io_o_3_out[4] ,
    \cb_7_5_io_o_3_out[3] ,
    \cb_7_5_io_o_3_out[2] ,
    \cb_7_5_io_o_3_out[1] ,
    \cb_7_5_io_o_3_out[0] }),
    .io_o_4_out({\cb_7_5_io_o_4_out[7] ,
    \cb_7_5_io_o_4_out[6] ,
    \cb_7_5_io_o_4_out[5] ,
    \cb_7_5_io_o_4_out[4] ,
    \cb_7_5_io_o_4_out[3] ,
    \cb_7_5_io_o_4_out[2] ,
    \cb_7_5_io_o_4_out[1] ,
    \cb_7_5_io_o_4_out[0] }),
    .io_o_5_out({\cb_7_5_io_o_5_out[7] ,
    \cb_7_5_io_o_5_out[6] ,
    \cb_7_5_io_o_5_out[5] ,
    \cb_7_5_io_o_5_out[4] ,
    \cb_7_5_io_o_5_out[3] ,
    \cb_7_5_io_o_5_out[2] ,
    \cb_7_5_io_o_5_out[1] ,
    \cb_7_5_io_o_5_out[0] }),
    .io_o_6_out({\cb_7_5_io_o_6_out[7] ,
    \cb_7_5_io_o_6_out[6] ,
    \cb_7_5_io_o_6_out[5] ,
    \cb_7_5_io_o_6_out[4] ,
    \cb_7_5_io_o_6_out[3] ,
    \cb_7_5_io_o_6_out[2] ,
    \cb_7_5_io_o_6_out[1] ,
    \cb_7_5_io_o_6_out[0] }),
    .io_o_7_out({\cb_7_5_io_o_7_out[7] ,
    \cb_7_5_io_o_7_out[6] ,
    \cb_7_5_io_o_7_out[5] ,
    \cb_7_5_io_o_7_out[4] ,
    \cb_7_5_io_o_7_out[3] ,
    \cb_7_5_io_o_7_out[2] ,
    \cb_7_5_io_o_7_out[1] ,
    \cb_7_5_io_o_7_out[0] }),
    .io_wo({\cb_7_4_io_eo[63] ,
    \cb_7_4_io_eo[62] ,
    \cb_7_4_io_eo[61] ,
    \cb_7_4_io_eo[60] ,
    \cb_7_4_io_eo[59] ,
    \cb_7_4_io_eo[58] ,
    \cb_7_4_io_eo[57] ,
    \cb_7_4_io_eo[56] ,
    \cb_7_4_io_eo[55] ,
    \cb_7_4_io_eo[54] ,
    \cb_7_4_io_eo[53] ,
    \cb_7_4_io_eo[52] ,
    \cb_7_4_io_eo[51] ,
    \cb_7_4_io_eo[50] ,
    \cb_7_4_io_eo[49] ,
    \cb_7_4_io_eo[48] ,
    \cb_7_4_io_eo[47] ,
    \cb_7_4_io_eo[46] ,
    \cb_7_4_io_eo[45] ,
    \cb_7_4_io_eo[44] ,
    \cb_7_4_io_eo[43] ,
    \cb_7_4_io_eo[42] ,
    \cb_7_4_io_eo[41] ,
    \cb_7_4_io_eo[40] ,
    \cb_7_4_io_eo[39] ,
    \cb_7_4_io_eo[38] ,
    \cb_7_4_io_eo[37] ,
    \cb_7_4_io_eo[36] ,
    \cb_7_4_io_eo[35] ,
    \cb_7_4_io_eo[34] ,
    \cb_7_4_io_eo[33] ,
    \cb_7_4_io_eo[32] ,
    \cb_7_4_io_eo[31] ,
    \cb_7_4_io_eo[30] ,
    \cb_7_4_io_eo[29] ,
    \cb_7_4_io_eo[28] ,
    \cb_7_4_io_eo[27] ,
    \cb_7_4_io_eo[26] ,
    \cb_7_4_io_eo[25] ,
    \cb_7_4_io_eo[24] ,
    \cb_7_4_io_eo[23] ,
    \cb_7_4_io_eo[22] ,
    \cb_7_4_io_eo[21] ,
    \cb_7_4_io_eo[20] ,
    \cb_7_4_io_eo[19] ,
    \cb_7_4_io_eo[18] ,
    \cb_7_4_io_eo[17] ,
    \cb_7_4_io_eo[16] ,
    \cb_7_4_io_eo[15] ,
    \cb_7_4_io_eo[14] ,
    \cb_7_4_io_eo[13] ,
    \cb_7_4_io_eo[12] ,
    \cb_7_4_io_eo[11] ,
    \cb_7_4_io_eo[10] ,
    \cb_7_4_io_eo[9] ,
    \cb_7_4_io_eo[8] ,
    \cb_7_4_io_eo[7] ,
    \cb_7_4_io_eo[6] ,
    \cb_7_4_io_eo[5] ,
    \cb_7_4_io_eo[4] ,
    \cb_7_4_io_eo[3] ,
    \cb_7_4_io_eo[2] ,
    \cb_7_4_io_eo[1] ,
    \cb_7_4_io_eo[0] }));
 cic_block cb_7_6 (.io_cs_i(cb_7_6_io_cs_i),
    .io_i_0_ci(cb_7_5_io_o_0_co),
    .io_i_1_ci(cb_7_5_io_o_1_co),
    .io_i_2_ci(cb_7_5_io_o_2_co),
    .io_i_3_ci(cb_7_5_io_o_3_co),
    .io_i_4_ci(cb_7_5_io_o_4_co),
    .io_i_5_ci(cb_7_5_io_o_5_co),
    .io_i_6_ci(cb_7_5_io_o_6_co),
    .io_i_7_ci(cb_7_5_io_o_7_co),
    .io_o_0_co(cb_7_6_io_o_0_co),
    .io_o_1_co(cb_7_6_io_o_1_co),
    .io_o_2_co(cb_7_6_io_o_2_co),
    .io_o_3_co(cb_7_6_io_o_3_co),
    .io_o_4_co(cb_7_6_io_o_4_co),
    .io_o_5_co(cb_7_6_io_o_5_co),
    .io_o_6_co(cb_7_6_io_o_6_co),
    .io_o_7_co(cb_7_6_io_o_7_co),
    .io_vci(cb_7_5_io_vco),
    .io_vco(cb_7_6_io_vco),
    .io_vi(cb_7_6_io_vi),
    .io_we_i(cb_7_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_7_0_io_adr_i[1] ,
    \cb_7_0_io_adr_i[0] }),
    .io_dat_i({\cb_7_0_io_dat_i[15] ,
    \cb_7_0_io_dat_i[14] ,
    \cb_7_0_io_dat_i[13] ,
    \cb_7_0_io_dat_i[12] ,
    \cb_7_0_io_dat_i[11] ,
    \cb_7_0_io_dat_i[10] ,
    \cb_7_0_io_dat_i[9] ,
    \cb_7_0_io_dat_i[8] ,
    \cb_7_0_io_dat_i[7] ,
    \cb_7_0_io_dat_i[6] ,
    \cb_7_0_io_dat_i[5] ,
    \cb_7_0_io_dat_i[4] ,
    \cb_7_0_io_dat_i[3] ,
    \cb_7_0_io_dat_i[2] ,
    \cb_7_0_io_dat_i[1] ,
    \cb_7_0_io_dat_i[0] }),
    .io_dat_o({\cb_7_6_io_dat_o[15] ,
    \cb_7_6_io_dat_o[14] ,
    \cb_7_6_io_dat_o[13] ,
    \cb_7_6_io_dat_o[12] ,
    \cb_7_6_io_dat_o[11] ,
    \cb_7_6_io_dat_o[10] ,
    \cb_7_6_io_dat_o[9] ,
    \cb_7_6_io_dat_o[8] ,
    \cb_7_6_io_dat_o[7] ,
    \cb_7_6_io_dat_o[6] ,
    \cb_7_6_io_dat_o[5] ,
    \cb_7_6_io_dat_o[4] ,
    \cb_7_6_io_dat_o[3] ,
    \cb_7_6_io_dat_o[2] ,
    \cb_7_6_io_dat_o[1] ,
    \cb_7_6_io_dat_o[0] }),
    .io_eo({\cb_7_6_io_eo[63] ,
    \cb_7_6_io_eo[62] ,
    \cb_7_6_io_eo[61] ,
    \cb_7_6_io_eo[60] ,
    \cb_7_6_io_eo[59] ,
    \cb_7_6_io_eo[58] ,
    \cb_7_6_io_eo[57] ,
    \cb_7_6_io_eo[56] ,
    \cb_7_6_io_eo[55] ,
    \cb_7_6_io_eo[54] ,
    \cb_7_6_io_eo[53] ,
    \cb_7_6_io_eo[52] ,
    \cb_7_6_io_eo[51] ,
    \cb_7_6_io_eo[50] ,
    \cb_7_6_io_eo[49] ,
    \cb_7_6_io_eo[48] ,
    \cb_7_6_io_eo[47] ,
    \cb_7_6_io_eo[46] ,
    \cb_7_6_io_eo[45] ,
    \cb_7_6_io_eo[44] ,
    \cb_7_6_io_eo[43] ,
    \cb_7_6_io_eo[42] ,
    \cb_7_6_io_eo[41] ,
    \cb_7_6_io_eo[40] ,
    \cb_7_6_io_eo[39] ,
    \cb_7_6_io_eo[38] ,
    \cb_7_6_io_eo[37] ,
    \cb_7_6_io_eo[36] ,
    \cb_7_6_io_eo[35] ,
    \cb_7_6_io_eo[34] ,
    \cb_7_6_io_eo[33] ,
    \cb_7_6_io_eo[32] ,
    \cb_7_6_io_eo[31] ,
    \cb_7_6_io_eo[30] ,
    \cb_7_6_io_eo[29] ,
    \cb_7_6_io_eo[28] ,
    \cb_7_6_io_eo[27] ,
    \cb_7_6_io_eo[26] ,
    \cb_7_6_io_eo[25] ,
    \cb_7_6_io_eo[24] ,
    \cb_7_6_io_eo[23] ,
    \cb_7_6_io_eo[22] ,
    \cb_7_6_io_eo[21] ,
    \cb_7_6_io_eo[20] ,
    \cb_7_6_io_eo[19] ,
    \cb_7_6_io_eo[18] ,
    \cb_7_6_io_eo[17] ,
    \cb_7_6_io_eo[16] ,
    \cb_7_6_io_eo[15] ,
    \cb_7_6_io_eo[14] ,
    \cb_7_6_io_eo[13] ,
    \cb_7_6_io_eo[12] ,
    \cb_7_6_io_eo[11] ,
    \cb_7_6_io_eo[10] ,
    \cb_7_6_io_eo[9] ,
    \cb_7_6_io_eo[8] ,
    \cb_7_6_io_eo[7] ,
    \cb_7_6_io_eo[6] ,
    \cb_7_6_io_eo[5] ,
    \cb_7_6_io_eo[4] ,
    \cb_7_6_io_eo[3] ,
    \cb_7_6_io_eo[2] ,
    \cb_7_6_io_eo[1] ,
    \cb_7_6_io_eo[0] }),
    .io_i_0_in1({\cb_7_5_io_o_0_out[7] ,
    \cb_7_5_io_o_0_out[6] ,
    \cb_7_5_io_o_0_out[5] ,
    \cb_7_5_io_o_0_out[4] ,
    \cb_7_5_io_o_0_out[3] ,
    \cb_7_5_io_o_0_out[2] ,
    \cb_7_5_io_o_0_out[1] ,
    \cb_7_5_io_o_0_out[0] }),
    .io_i_1_in1({\cb_7_5_io_o_1_out[7] ,
    \cb_7_5_io_o_1_out[6] ,
    \cb_7_5_io_o_1_out[5] ,
    \cb_7_5_io_o_1_out[4] ,
    \cb_7_5_io_o_1_out[3] ,
    \cb_7_5_io_o_1_out[2] ,
    \cb_7_5_io_o_1_out[1] ,
    \cb_7_5_io_o_1_out[0] }),
    .io_i_2_in1({\cb_7_5_io_o_2_out[7] ,
    \cb_7_5_io_o_2_out[6] ,
    \cb_7_5_io_o_2_out[5] ,
    \cb_7_5_io_o_2_out[4] ,
    \cb_7_5_io_o_2_out[3] ,
    \cb_7_5_io_o_2_out[2] ,
    \cb_7_5_io_o_2_out[1] ,
    \cb_7_5_io_o_2_out[0] }),
    .io_i_3_in1({\cb_7_5_io_o_3_out[7] ,
    \cb_7_5_io_o_3_out[6] ,
    \cb_7_5_io_o_3_out[5] ,
    \cb_7_5_io_o_3_out[4] ,
    \cb_7_5_io_o_3_out[3] ,
    \cb_7_5_io_o_3_out[2] ,
    \cb_7_5_io_o_3_out[1] ,
    \cb_7_5_io_o_3_out[0] }),
    .io_i_4_in1({\cb_7_5_io_o_4_out[7] ,
    \cb_7_5_io_o_4_out[6] ,
    \cb_7_5_io_o_4_out[5] ,
    \cb_7_5_io_o_4_out[4] ,
    \cb_7_5_io_o_4_out[3] ,
    \cb_7_5_io_o_4_out[2] ,
    \cb_7_5_io_o_4_out[1] ,
    \cb_7_5_io_o_4_out[0] }),
    .io_i_5_in1({\cb_7_5_io_o_5_out[7] ,
    \cb_7_5_io_o_5_out[6] ,
    \cb_7_5_io_o_5_out[5] ,
    \cb_7_5_io_o_5_out[4] ,
    \cb_7_5_io_o_5_out[3] ,
    \cb_7_5_io_o_5_out[2] ,
    \cb_7_5_io_o_5_out[1] ,
    \cb_7_5_io_o_5_out[0] }),
    .io_i_6_in1({\cb_7_5_io_o_6_out[7] ,
    \cb_7_5_io_o_6_out[6] ,
    \cb_7_5_io_o_6_out[5] ,
    \cb_7_5_io_o_6_out[4] ,
    \cb_7_5_io_o_6_out[3] ,
    \cb_7_5_io_o_6_out[2] ,
    \cb_7_5_io_o_6_out[1] ,
    \cb_7_5_io_o_6_out[0] }),
    .io_i_7_in1({\cb_7_5_io_o_7_out[7] ,
    \cb_7_5_io_o_7_out[6] ,
    \cb_7_5_io_o_7_out[5] ,
    \cb_7_5_io_o_7_out[4] ,
    \cb_7_5_io_o_7_out[3] ,
    \cb_7_5_io_o_7_out[2] ,
    \cb_7_5_io_o_7_out[1] ,
    \cb_7_5_io_o_7_out[0] }),
    .io_o_0_out({\cb_7_6_io_o_0_out[7] ,
    \cb_7_6_io_o_0_out[6] ,
    \cb_7_6_io_o_0_out[5] ,
    \cb_7_6_io_o_0_out[4] ,
    \cb_7_6_io_o_0_out[3] ,
    \cb_7_6_io_o_0_out[2] ,
    \cb_7_6_io_o_0_out[1] ,
    \cb_7_6_io_o_0_out[0] }),
    .io_o_1_out({\cb_7_6_io_o_1_out[7] ,
    \cb_7_6_io_o_1_out[6] ,
    \cb_7_6_io_o_1_out[5] ,
    \cb_7_6_io_o_1_out[4] ,
    \cb_7_6_io_o_1_out[3] ,
    \cb_7_6_io_o_1_out[2] ,
    \cb_7_6_io_o_1_out[1] ,
    \cb_7_6_io_o_1_out[0] }),
    .io_o_2_out({\cb_7_6_io_o_2_out[7] ,
    \cb_7_6_io_o_2_out[6] ,
    \cb_7_6_io_o_2_out[5] ,
    \cb_7_6_io_o_2_out[4] ,
    \cb_7_6_io_o_2_out[3] ,
    \cb_7_6_io_o_2_out[2] ,
    \cb_7_6_io_o_2_out[1] ,
    \cb_7_6_io_o_2_out[0] }),
    .io_o_3_out({\cb_7_6_io_o_3_out[7] ,
    \cb_7_6_io_o_3_out[6] ,
    \cb_7_6_io_o_3_out[5] ,
    \cb_7_6_io_o_3_out[4] ,
    \cb_7_6_io_o_3_out[3] ,
    \cb_7_6_io_o_3_out[2] ,
    \cb_7_6_io_o_3_out[1] ,
    \cb_7_6_io_o_3_out[0] }),
    .io_o_4_out({\cb_7_6_io_o_4_out[7] ,
    \cb_7_6_io_o_4_out[6] ,
    \cb_7_6_io_o_4_out[5] ,
    \cb_7_6_io_o_4_out[4] ,
    \cb_7_6_io_o_4_out[3] ,
    \cb_7_6_io_o_4_out[2] ,
    \cb_7_6_io_o_4_out[1] ,
    \cb_7_6_io_o_4_out[0] }),
    .io_o_5_out({\cb_7_6_io_o_5_out[7] ,
    \cb_7_6_io_o_5_out[6] ,
    \cb_7_6_io_o_5_out[5] ,
    \cb_7_6_io_o_5_out[4] ,
    \cb_7_6_io_o_5_out[3] ,
    \cb_7_6_io_o_5_out[2] ,
    \cb_7_6_io_o_5_out[1] ,
    \cb_7_6_io_o_5_out[0] }),
    .io_o_6_out({\cb_7_6_io_o_6_out[7] ,
    \cb_7_6_io_o_6_out[6] ,
    \cb_7_6_io_o_6_out[5] ,
    \cb_7_6_io_o_6_out[4] ,
    \cb_7_6_io_o_6_out[3] ,
    \cb_7_6_io_o_6_out[2] ,
    \cb_7_6_io_o_6_out[1] ,
    \cb_7_6_io_o_6_out[0] }),
    .io_o_7_out({\cb_7_6_io_o_7_out[7] ,
    \cb_7_6_io_o_7_out[6] ,
    \cb_7_6_io_o_7_out[5] ,
    \cb_7_6_io_o_7_out[4] ,
    \cb_7_6_io_o_7_out[3] ,
    \cb_7_6_io_o_7_out[2] ,
    \cb_7_6_io_o_7_out[1] ,
    \cb_7_6_io_o_7_out[0] }),
    .io_wo({\cb_7_5_io_eo[63] ,
    \cb_7_5_io_eo[62] ,
    \cb_7_5_io_eo[61] ,
    \cb_7_5_io_eo[60] ,
    \cb_7_5_io_eo[59] ,
    \cb_7_5_io_eo[58] ,
    \cb_7_5_io_eo[57] ,
    \cb_7_5_io_eo[56] ,
    \cb_7_5_io_eo[55] ,
    \cb_7_5_io_eo[54] ,
    \cb_7_5_io_eo[53] ,
    \cb_7_5_io_eo[52] ,
    \cb_7_5_io_eo[51] ,
    \cb_7_5_io_eo[50] ,
    \cb_7_5_io_eo[49] ,
    \cb_7_5_io_eo[48] ,
    \cb_7_5_io_eo[47] ,
    \cb_7_5_io_eo[46] ,
    \cb_7_5_io_eo[45] ,
    \cb_7_5_io_eo[44] ,
    \cb_7_5_io_eo[43] ,
    \cb_7_5_io_eo[42] ,
    \cb_7_5_io_eo[41] ,
    \cb_7_5_io_eo[40] ,
    \cb_7_5_io_eo[39] ,
    \cb_7_5_io_eo[38] ,
    \cb_7_5_io_eo[37] ,
    \cb_7_5_io_eo[36] ,
    \cb_7_5_io_eo[35] ,
    \cb_7_5_io_eo[34] ,
    \cb_7_5_io_eo[33] ,
    \cb_7_5_io_eo[32] ,
    \cb_7_5_io_eo[31] ,
    \cb_7_5_io_eo[30] ,
    \cb_7_5_io_eo[29] ,
    \cb_7_5_io_eo[28] ,
    \cb_7_5_io_eo[27] ,
    \cb_7_5_io_eo[26] ,
    \cb_7_5_io_eo[25] ,
    \cb_7_5_io_eo[24] ,
    \cb_7_5_io_eo[23] ,
    \cb_7_5_io_eo[22] ,
    \cb_7_5_io_eo[21] ,
    \cb_7_5_io_eo[20] ,
    \cb_7_5_io_eo[19] ,
    \cb_7_5_io_eo[18] ,
    \cb_7_5_io_eo[17] ,
    \cb_7_5_io_eo[16] ,
    \cb_7_5_io_eo[15] ,
    \cb_7_5_io_eo[14] ,
    \cb_7_5_io_eo[13] ,
    \cb_7_5_io_eo[12] ,
    \cb_7_5_io_eo[11] ,
    \cb_7_5_io_eo[10] ,
    \cb_7_5_io_eo[9] ,
    \cb_7_5_io_eo[8] ,
    \cb_7_5_io_eo[7] ,
    \cb_7_5_io_eo[6] ,
    \cb_7_5_io_eo[5] ,
    \cb_7_5_io_eo[4] ,
    \cb_7_5_io_eo[3] ,
    \cb_7_5_io_eo[2] ,
    \cb_7_5_io_eo[1] ,
    \cb_7_5_io_eo[0] }));
 cic_block cb_7_7 (.io_cs_i(cb_7_7_io_cs_i),
    .io_i_0_ci(cb_7_6_io_o_0_co),
    .io_i_1_ci(cb_7_6_io_o_1_co),
    .io_i_2_ci(cb_7_6_io_o_2_co),
    .io_i_3_ci(cb_7_6_io_o_3_co),
    .io_i_4_ci(cb_7_6_io_o_4_co),
    .io_i_5_ci(cb_7_6_io_o_5_co),
    .io_i_6_ci(cb_7_6_io_o_6_co),
    .io_i_7_ci(cb_7_6_io_o_7_co),
    .io_o_0_co(cb_7_7_io_o_0_co),
    .io_o_1_co(cb_7_7_io_o_1_co),
    .io_o_2_co(cb_7_7_io_o_2_co),
    .io_o_3_co(cb_7_7_io_o_3_co),
    .io_o_4_co(cb_7_7_io_o_4_co),
    .io_o_5_co(cb_7_7_io_o_5_co),
    .io_o_6_co(cb_7_7_io_o_6_co),
    .io_o_7_co(cb_7_7_io_o_7_co),
    .io_vci(cb_7_6_io_vco),
    .io_vco(cb_7_7_io_vco),
    .io_vi(cb_7_7_io_vi),
    .io_we_i(cb_7_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_7_0_io_adr_i[1] ,
    \cb_7_0_io_adr_i[0] }),
    .io_dat_i({\cb_7_0_io_dat_i[15] ,
    \cb_7_0_io_dat_i[14] ,
    \cb_7_0_io_dat_i[13] ,
    \cb_7_0_io_dat_i[12] ,
    \cb_7_0_io_dat_i[11] ,
    \cb_7_0_io_dat_i[10] ,
    \cb_7_0_io_dat_i[9] ,
    \cb_7_0_io_dat_i[8] ,
    \cb_7_0_io_dat_i[7] ,
    \cb_7_0_io_dat_i[6] ,
    \cb_7_0_io_dat_i[5] ,
    \cb_7_0_io_dat_i[4] ,
    \cb_7_0_io_dat_i[3] ,
    \cb_7_0_io_dat_i[2] ,
    \cb_7_0_io_dat_i[1] ,
    \cb_7_0_io_dat_i[0] }),
    .io_dat_o({\cb_7_7_io_dat_o[15] ,
    \cb_7_7_io_dat_o[14] ,
    \cb_7_7_io_dat_o[13] ,
    \cb_7_7_io_dat_o[12] ,
    \cb_7_7_io_dat_o[11] ,
    \cb_7_7_io_dat_o[10] ,
    \cb_7_7_io_dat_o[9] ,
    \cb_7_7_io_dat_o[8] ,
    \cb_7_7_io_dat_o[7] ,
    \cb_7_7_io_dat_o[6] ,
    \cb_7_7_io_dat_o[5] ,
    \cb_7_7_io_dat_o[4] ,
    \cb_7_7_io_dat_o[3] ,
    \cb_7_7_io_dat_o[2] ,
    \cb_7_7_io_dat_o[1] ,
    \cb_7_7_io_dat_o[0] }),
    .io_eo({\cb_7_7_io_eo[63] ,
    \cb_7_7_io_eo[62] ,
    \cb_7_7_io_eo[61] ,
    \cb_7_7_io_eo[60] ,
    \cb_7_7_io_eo[59] ,
    \cb_7_7_io_eo[58] ,
    \cb_7_7_io_eo[57] ,
    \cb_7_7_io_eo[56] ,
    \cb_7_7_io_eo[55] ,
    \cb_7_7_io_eo[54] ,
    \cb_7_7_io_eo[53] ,
    \cb_7_7_io_eo[52] ,
    \cb_7_7_io_eo[51] ,
    \cb_7_7_io_eo[50] ,
    \cb_7_7_io_eo[49] ,
    \cb_7_7_io_eo[48] ,
    \cb_7_7_io_eo[47] ,
    \cb_7_7_io_eo[46] ,
    \cb_7_7_io_eo[45] ,
    \cb_7_7_io_eo[44] ,
    \cb_7_7_io_eo[43] ,
    \cb_7_7_io_eo[42] ,
    \cb_7_7_io_eo[41] ,
    \cb_7_7_io_eo[40] ,
    \cb_7_7_io_eo[39] ,
    \cb_7_7_io_eo[38] ,
    \cb_7_7_io_eo[37] ,
    \cb_7_7_io_eo[36] ,
    \cb_7_7_io_eo[35] ,
    \cb_7_7_io_eo[34] ,
    \cb_7_7_io_eo[33] ,
    \cb_7_7_io_eo[32] ,
    \cb_7_7_io_eo[31] ,
    \cb_7_7_io_eo[30] ,
    \cb_7_7_io_eo[29] ,
    \cb_7_7_io_eo[28] ,
    \cb_7_7_io_eo[27] ,
    \cb_7_7_io_eo[26] ,
    \cb_7_7_io_eo[25] ,
    \cb_7_7_io_eo[24] ,
    \cb_7_7_io_eo[23] ,
    \cb_7_7_io_eo[22] ,
    \cb_7_7_io_eo[21] ,
    \cb_7_7_io_eo[20] ,
    \cb_7_7_io_eo[19] ,
    \cb_7_7_io_eo[18] ,
    \cb_7_7_io_eo[17] ,
    \cb_7_7_io_eo[16] ,
    \cb_7_7_io_eo[15] ,
    \cb_7_7_io_eo[14] ,
    \cb_7_7_io_eo[13] ,
    \cb_7_7_io_eo[12] ,
    \cb_7_7_io_eo[11] ,
    \cb_7_7_io_eo[10] ,
    \cb_7_7_io_eo[9] ,
    \cb_7_7_io_eo[8] ,
    \cb_7_7_io_eo[7] ,
    \cb_7_7_io_eo[6] ,
    \cb_7_7_io_eo[5] ,
    \cb_7_7_io_eo[4] ,
    \cb_7_7_io_eo[3] ,
    \cb_7_7_io_eo[2] ,
    \cb_7_7_io_eo[1] ,
    \cb_7_7_io_eo[0] }),
    .io_i_0_in1({\cb_7_6_io_o_0_out[7] ,
    \cb_7_6_io_o_0_out[6] ,
    \cb_7_6_io_o_0_out[5] ,
    \cb_7_6_io_o_0_out[4] ,
    \cb_7_6_io_o_0_out[3] ,
    \cb_7_6_io_o_0_out[2] ,
    \cb_7_6_io_o_0_out[1] ,
    \cb_7_6_io_o_0_out[0] }),
    .io_i_1_in1({\cb_7_6_io_o_1_out[7] ,
    \cb_7_6_io_o_1_out[6] ,
    \cb_7_6_io_o_1_out[5] ,
    \cb_7_6_io_o_1_out[4] ,
    \cb_7_6_io_o_1_out[3] ,
    \cb_7_6_io_o_1_out[2] ,
    \cb_7_6_io_o_1_out[1] ,
    \cb_7_6_io_o_1_out[0] }),
    .io_i_2_in1({\cb_7_6_io_o_2_out[7] ,
    \cb_7_6_io_o_2_out[6] ,
    \cb_7_6_io_o_2_out[5] ,
    \cb_7_6_io_o_2_out[4] ,
    \cb_7_6_io_o_2_out[3] ,
    \cb_7_6_io_o_2_out[2] ,
    \cb_7_6_io_o_2_out[1] ,
    \cb_7_6_io_o_2_out[0] }),
    .io_i_3_in1({\cb_7_6_io_o_3_out[7] ,
    \cb_7_6_io_o_3_out[6] ,
    \cb_7_6_io_o_3_out[5] ,
    \cb_7_6_io_o_3_out[4] ,
    \cb_7_6_io_o_3_out[3] ,
    \cb_7_6_io_o_3_out[2] ,
    \cb_7_6_io_o_3_out[1] ,
    \cb_7_6_io_o_3_out[0] }),
    .io_i_4_in1({\cb_7_6_io_o_4_out[7] ,
    \cb_7_6_io_o_4_out[6] ,
    \cb_7_6_io_o_4_out[5] ,
    \cb_7_6_io_o_4_out[4] ,
    \cb_7_6_io_o_4_out[3] ,
    \cb_7_6_io_o_4_out[2] ,
    \cb_7_6_io_o_4_out[1] ,
    \cb_7_6_io_o_4_out[0] }),
    .io_i_5_in1({\cb_7_6_io_o_5_out[7] ,
    \cb_7_6_io_o_5_out[6] ,
    \cb_7_6_io_o_5_out[5] ,
    \cb_7_6_io_o_5_out[4] ,
    \cb_7_6_io_o_5_out[3] ,
    \cb_7_6_io_o_5_out[2] ,
    \cb_7_6_io_o_5_out[1] ,
    \cb_7_6_io_o_5_out[0] }),
    .io_i_6_in1({\cb_7_6_io_o_6_out[7] ,
    \cb_7_6_io_o_6_out[6] ,
    \cb_7_6_io_o_6_out[5] ,
    \cb_7_6_io_o_6_out[4] ,
    \cb_7_6_io_o_6_out[3] ,
    \cb_7_6_io_o_6_out[2] ,
    \cb_7_6_io_o_6_out[1] ,
    \cb_7_6_io_o_6_out[0] }),
    .io_i_7_in1({\cb_7_6_io_o_7_out[7] ,
    \cb_7_6_io_o_7_out[6] ,
    \cb_7_6_io_o_7_out[5] ,
    \cb_7_6_io_o_7_out[4] ,
    \cb_7_6_io_o_7_out[3] ,
    \cb_7_6_io_o_7_out[2] ,
    \cb_7_6_io_o_7_out[1] ,
    \cb_7_6_io_o_7_out[0] }),
    .io_o_0_out({\cb_7_7_io_o_0_out[7] ,
    \cb_7_7_io_o_0_out[6] ,
    \cb_7_7_io_o_0_out[5] ,
    \cb_7_7_io_o_0_out[4] ,
    \cb_7_7_io_o_0_out[3] ,
    \cb_7_7_io_o_0_out[2] ,
    \cb_7_7_io_o_0_out[1] ,
    \cb_7_7_io_o_0_out[0] }),
    .io_o_1_out({\cb_7_7_io_o_1_out[7] ,
    \cb_7_7_io_o_1_out[6] ,
    \cb_7_7_io_o_1_out[5] ,
    \cb_7_7_io_o_1_out[4] ,
    \cb_7_7_io_o_1_out[3] ,
    \cb_7_7_io_o_1_out[2] ,
    \cb_7_7_io_o_1_out[1] ,
    \cb_7_7_io_o_1_out[0] }),
    .io_o_2_out({\cb_7_7_io_o_2_out[7] ,
    \cb_7_7_io_o_2_out[6] ,
    \cb_7_7_io_o_2_out[5] ,
    \cb_7_7_io_o_2_out[4] ,
    \cb_7_7_io_o_2_out[3] ,
    \cb_7_7_io_o_2_out[2] ,
    \cb_7_7_io_o_2_out[1] ,
    \cb_7_7_io_o_2_out[0] }),
    .io_o_3_out({\cb_7_7_io_o_3_out[7] ,
    \cb_7_7_io_o_3_out[6] ,
    \cb_7_7_io_o_3_out[5] ,
    \cb_7_7_io_o_3_out[4] ,
    \cb_7_7_io_o_3_out[3] ,
    \cb_7_7_io_o_3_out[2] ,
    \cb_7_7_io_o_3_out[1] ,
    \cb_7_7_io_o_3_out[0] }),
    .io_o_4_out({\cb_7_7_io_o_4_out[7] ,
    \cb_7_7_io_o_4_out[6] ,
    \cb_7_7_io_o_4_out[5] ,
    \cb_7_7_io_o_4_out[4] ,
    \cb_7_7_io_o_4_out[3] ,
    \cb_7_7_io_o_4_out[2] ,
    \cb_7_7_io_o_4_out[1] ,
    \cb_7_7_io_o_4_out[0] }),
    .io_o_5_out({\cb_7_7_io_o_5_out[7] ,
    \cb_7_7_io_o_5_out[6] ,
    \cb_7_7_io_o_5_out[5] ,
    \cb_7_7_io_o_5_out[4] ,
    \cb_7_7_io_o_5_out[3] ,
    \cb_7_7_io_o_5_out[2] ,
    \cb_7_7_io_o_5_out[1] ,
    \cb_7_7_io_o_5_out[0] }),
    .io_o_6_out({\cb_7_7_io_o_6_out[7] ,
    \cb_7_7_io_o_6_out[6] ,
    \cb_7_7_io_o_6_out[5] ,
    \cb_7_7_io_o_6_out[4] ,
    \cb_7_7_io_o_6_out[3] ,
    \cb_7_7_io_o_6_out[2] ,
    \cb_7_7_io_o_6_out[1] ,
    \cb_7_7_io_o_6_out[0] }),
    .io_o_7_out({\cb_7_7_io_o_7_out[7] ,
    \cb_7_7_io_o_7_out[6] ,
    \cb_7_7_io_o_7_out[5] ,
    \cb_7_7_io_o_7_out[4] ,
    \cb_7_7_io_o_7_out[3] ,
    \cb_7_7_io_o_7_out[2] ,
    \cb_7_7_io_o_7_out[1] ,
    \cb_7_7_io_o_7_out[0] }),
    .io_wo({\cb_7_6_io_eo[63] ,
    \cb_7_6_io_eo[62] ,
    \cb_7_6_io_eo[61] ,
    \cb_7_6_io_eo[60] ,
    \cb_7_6_io_eo[59] ,
    \cb_7_6_io_eo[58] ,
    \cb_7_6_io_eo[57] ,
    \cb_7_6_io_eo[56] ,
    \cb_7_6_io_eo[55] ,
    \cb_7_6_io_eo[54] ,
    \cb_7_6_io_eo[53] ,
    \cb_7_6_io_eo[52] ,
    \cb_7_6_io_eo[51] ,
    \cb_7_6_io_eo[50] ,
    \cb_7_6_io_eo[49] ,
    \cb_7_6_io_eo[48] ,
    \cb_7_6_io_eo[47] ,
    \cb_7_6_io_eo[46] ,
    \cb_7_6_io_eo[45] ,
    \cb_7_6_io_eo[44] ,
    \cb_7_6_io_eo[43] ,
    \cb_7_6_io_eo[42] ,
    \cb_7_6_io_eo[41] ,
    \cb_7_6_io_eo[40] ,
    \cb_7_6_io_eo[39] ,
    \cb_7_6_io_eo[38] ,
    \cb_7_6_io_eo[37] ,
    \cb_7_6_io_eo[36] ,
    \cb_7_6_io_eo[35] ,
    \cb_7_6_io_eo[34] ,
    \cb_7_6_io_eo[33] ,
    \cb_7_6_io_eo[32] ,
    \cb_7_6_io_eo[31] ,
    \cb_7_6_io_eo[30] ,
    \cb_7_6_io_eo[29] ,
    \cb_7_6_io_eo[28] ,
    \cb_7_6_io_eo[27] ,
    \cb_7_6_io_eo[26] ,
    \cb_7_6_io_eo[25] ,
    \cb_7_6_io_eo[24] ,
    \cb_7_6_io_eo[23] ,
    \cb_7_6_io_eo[22] ,
    \cb_7_6_io_eo[21] ,
    \cb_7_6_io_eo[20] ,
    \cb_7_6_io_eo[19] ,
    \cb_7_6_io_eo[18] ,
    \cb_7_6_io_eo[17] ,
    \cb_7_6_io_eo[16] ,
    \cb_7_6_io_eo[15] ,
    \cb_7_6_io_eo[14] ,
    \cb_7_6_io_eo[13] ,
    \cb_7_6_io_eo[12] ,
    \cb_7_6_io_eo[11] ,
    \cb_7_6_io_eo[10] ,
    \cb_7_6_io_eo[9] ,
    \cb_7_6_io_eo[8] ,
    \cb_7_6_io_eo[7] ,
    \cb_7_6_io_eo[6] ,
    \cb_7_6_io_eo[5] ,
    \cb_7_6_io_eo[4] ,
    \cb_7_6_io_eo[3] ,
    \cb_7_6_io_eo[2] ,
    \cb_7_6_io_eo[1] ,
    \cb_7_6_io_eo[0] }));
 cic_block cb_7_8 (.io_cs_i(cb_7_8_io_cs_i),
    .io_i_0_ci(cb_7_7_io_o_0_co),
    .io_i_1_ci(cb_7_7_io_o_1_co),
    .io_i_2_ci(cb_7_7_io_o_2_co),
    .io_i_3_ci(cb_7_7_io_o_3_co),
    .io_i_4_ci(cb_7_7_io_o_4_co),
    .io_i_5_ci(cb_7_7_io_o_5_co),
    .io_i_6_ci(cb_7_7_io_o_6_co),
    .io_i_7_ci(cb_7_7_io_o_7_co),
    .io_o_0_co(cb_7_8_io_o_0_co),
    .io_o_1_co(cb_7_8_io_o_1_co),
    .io_o_2_co(cb_7_8_io_o_2_co),
    .io_o_3_co(cb_7_8_io_o_3_co),
    .io_o_4_co(cb_7_8_io_o_4_co),
    .io_o_5_co(cb_7_8_io_o_5_co),
    .io_o_6_co(cb_7_8_io_o_6_co),
    .io_o_7_co(cb_7_8_io_o_7_co),
    .io_vci(cb_7_7_io_vco),
    .io_vco(cb_7_8_io_vco),
    .io_vi(cb_7_8_io_vi),
    .io_we_i(cb_7_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_7_0_io_adr_i[1] ,
    \cb_7_0_io_adr_i[0] }),
    .io_dat_i({\cb_7_0_io_dat_i[15] ,
    \cb_7_0_io_dat_i[14] ,
    \cb_7_0_io_dat_i[13] ,
    \cb_7_0_io_dat_i[12] ,
    \cb_7_0_io_dat_i[11] ,
    \cb_7_0_io_dat_i[10] ,
    \cb_7_0_io_dat_i[9] ,
    \cb_7_0_io_dat_i[8] ,
    \cb_7_0_io_dat_i[7] ,
    \cb_7_0_io_dat_i[6] ,
    \cb_7_0_io_dat_i[5] ,
    \cb_7_0_io_dat_i[4] ,
    \cb_7_0_io_dat_i[3] ,
    \cb_7_0_io_dat_i[2] ,
    \cb_7_0_io_dat_i[1] ,
    \cb_7_0_io_dat_i[0] }),
    .io_dat_o({\cb_7_8_io_dat_o[15] ,
    \cb_7_8_io_dat_o[14] ,
    \cb_7_8_io_dat_o[13] ,
    \cb_7_8_io_dat_o[12] ,
    \cb_7_8_io_dat_o[11] ,
    \cb_7_8_io_dat_o[10] ,
    \cb_7_8_io_dat_o[9] ,
    \cb_7_8_io_dat_o[8] ,
    \cb_7_8_io_dat_o[7] ,
    \cb_7_8_io_dat_o[6] ,
    \cb_7_8_io_dat_o[5] ,
    \cb_7_8_io_dat_o[4] ,
    \cb_7_8_io_dat_o[3] ,
    \cb_7_8_io_dat_o[2] ,
    \cb_7_8_io_dat_o[1] ,
    \cb_7_8_io_dat_o[0] }),
    .io_eo({\cb_7_8_io_eo[63] ,
    \cb_7_8_io_eo[62] ,
    \cb_7_8_io_eo[61] ,
    \cb_7_8_io_eo[60] ,
    \cb_7_8_io_eo[59] ,
    \cb_7_8_io_eo[58] ,
    \cb_7_8_io_eo[57] ,
    \cb_7_8_io_eo[56] ,
    \cb_7_8_io_eo[55] ,
    \cb_7_8_io_eo[54] ,
    \cb_7_8_io_eo[53] ,
    \cb_7_8_io_eo[52] ,
    \cb_7_8_io_eo[51] ,
    \cb_7_8_io_eo[50] ,
    \cb_7_8_io_eo[49] ,
    \cb_7_8_io_eo[48] ,
    \cb_7_8_io_eo[47] ,
    \cb_7_8_io_eo[46] ,
    \cb_7_8_io_eo[45] ,
    \cb_7_8_io_eo[44] ,
    \cb_7_8_io_eo[43] ,
    \cb_7_8_io_eo[42] ,
    \cb_7_8_io_eo[41] ,
    \cb_7_8_io_eo[40] ,
    \cb_7_8_io_eo[39] ,
    \cb_7_8_io_eo[38] ,
    \cb_7_8_io_eo[37] ,
    \cb_7_8_io_eo[36] ,
    \cb_7_8_io_eo[35] ,
    \cb_7_8_io_eo[34] ,
    \cb_7_8_io_eo[33] ,
    \cb_7_8_io_eo[32] ,
    \cb_7_8_io_eo[31] ,
    \cb_7_8_io_eo[30] ,
    \cb_7_8_io_eo[29] ,
    \cb_7_8_io_eo[28] ,
    \cb_7_8_io_eo[27] ,
    \cb_7_8_io_eo[26] ,
    \cb_7_8_io_eo[25] ,
    \cb_7_8_io_eo[24] ,
    \cb_7_8_io_eo[23] ,
    \cb_7_8_io_eo[22] ,
    \cb_7_8_io_eo[21] ,
    \cb_7_8_io_eo[20] ,
    \cb_7_8_io_eo[19] ,
    \cb_7_8_io_eo[18] ,
    \cb_7_8_io_eo[17] ,
    \cb_7_8_io_eo[16] ,
    \cb_7_8_io_eo[15] ,
    \cb_7_8_io_eo[14] ,
    \cb_7_8_io_eo[13] ,
    \cb_7_8_io_eo[12] ,
    \cb_7_8_io_eo[11] ,
    \cb_7_8_io_eo[10] ,
    \cb_7_8_io_eo[9] ,
    \cb_7_8_io_eo[8] ,
    \cb_7_8_io_eo[7] ,
    \cb_7_8_io_eo[6] ,
    \cb_7_8_io_eo[5] ,
    \cb_7_8_io_eo[4] ,
    \cb_7_8_io_eo[3] ,
    \cb_7_8_io_eo[2] ,
    \cb_7_8_io_eo[1] ,
    \cb_7_8_io_eo[0] }),
    .io_i_0_in1({\cb_7_7_io_o_0_out[7] ,
    \cb_7_7_io_o_0_out[6] ,
    \cb_7_7_io_o_0_out[5] ,
    \cb_7_7_io_o_0_out[4] ,
    \cb_7_7_io_o_0_out[3] ,
    \cb_7_7_io_o_0_out[2] ,
    \cb_7_7_io_o_0_out[1] ,
    \cb_7_7_io_o_0_out[0] }),
    .io_i_1_in1({\cb_7_7_io_o_1_out[7] ,
    \cb_7_7_io_o_1_out[6] ,
    \cb_7_7_io_o_1_out[5] ,
    \cb_7_7_io_o_1_out[4] ,
    \cb_7_7_io_o_1_out[3] ,
    \cb_7_7_io_o_1_out[2] ,
    \cb_7_7_io_o_1_out[1] ,
    \cb_7_7_io_o_1_out[0] }),
    .io_i_2_in1({\cb_7_7_io_o_2_out[7] ,
    \cb_7_7_io_o_2_out[6] ,
    \cb_7_7_io_o_2_out[5] ,
    \cb_7_7_io_o_2_out[4] ,
    \cb_7_7_io_o_2_out[3] ,
    \cb_7_7_io_o_2_out[2] ,
    \cb_7_7_io_o_2_out[1] ,
    \cb_7_7_io_o_2_out[0] }),
    .io_i_3_in1({\cb_7_7_io_o_3_out[7] ,
    \cb_7_7_io_o_3_out[6] ,
    \cb_7_7_io_o_3_out[5] ,
    \cb_7_7_io_o_3_out[4] ,
    \cb_7_7_io_o_3_out[3] ,
    \cb_7_7_io_o_3_out[2] ,
    \cb_7_7_io_o_3_out[1] ,
    \cb_7_7_io_o_3_out[0] }),
    .io_i_4_in1({\cb_7_7_io_o_4_out[7] ,
    \cb_7_7_io_o_4_out[6] ,
    \cb_7_7_io_o_4_out[5] ,
    \cb_7_7_io_o_4_out[4] ,
    \cb_7_7_io_o_4_out[3] ,
    \cb_7_7_io_o_4_out[2] ,
    \cb_7_7_io_o_4_out[1] ,
    \cb_7_7_io_o_4_out[0] }),
    .io_i_5_in1({\cb_7_7_io_o_5_out[7] ,
    \cb_7_7_io_o_5_out[6] ,
    \cb_7_7_io_o_5_out[5] ,
    \cb_7_7_io_o_5_out[4] ,
    \cb_7_7_io_o_5_out[3] ,
    \cb_7_7_io_o_5_out[2] ,
    \cb_7_7_io_o_5_out[1] ,
    \cb_7_7_io_o_5_out[0] }),
    .io_i_6_in1({\cb_7_7_io_o_6_out[7] ,
    \cb_7_7_io_o_6_out[6] ,
    \cb_7_7_io_o_6_out[5] ,
    \cb_7_7_io_o_6_out[4] ,
    \cb_7_7_io_o_6_out[3] ,
    \cb_7_7_io_o_6_out[2] ,
    \cb_7_7_io_o_6_out[1] ,
    \cb_7_7_io_o_6_out[0] }),
    .io_i_7_in1({\cb_7_7_io_o_7_out[7] ,
    \cb_7_7_io_o_7_out[6] ,
    \cb_7_7_io_o_7_out[5] ,
    \cb_7_7_io_o_7_out[4] ,
    \cb_7_7_io_o_7_out[3] ,
    \cb_7_7_io_o_7_out[2] ,
    \cb_7_7_io_o_7_out[1] ,
    \cb_7_7_io_o_7_out[0] }),
    .io_o_0_out({\cb_7_8_io_o_0_out[7] ,
    \cb_7_8_io_o_0_out[6] ,
    \cb_7_8_io_o_0_out[5] ,
    \cb_7_8_io_o_0_out[4] ,
    \cb_7_8_io_o_0_out[3] ,
    \cb_7_8_io_o_0_out[2] ,
    \cb_7_8_io_o_0_out[1] ,
    \cb_7_8_io_o_0_out[0] }),
    .io_o_1_out({\cb_7_8_io_o_1_out[7] ,
    \cb_7_8_io_o_1_out[6] ,
    \cb_7_8_io_o_1_out[5] ,
    \cb_7_8_io_o_1_out[4] ,
    \cb_7_8_io_o_1_out[3] ,
    \cb_7_8_io_o_1_out[2] ,
    \cb_7_8_io_o_1_out[1] ,
    \cb_7_8_io_o_1_out[0] }),
    .io_o_2_out({\cb_7_8_io_o_2_out[7] ,
    \cb_7_8_io_o_2_out[6] ,
    \cb_7_8_io_o_2_out[5] ,
    \cb_7_8_io_o_2_out[4] ,
    \cb_7_8_io_o_2_out[3] ,
    \cb_7_8_io_o_2_out[2] ,
    \cb_7_8_io_o_2_out[1] ,
    \cb_7_8_io_o_2_out[0] }),
    .io_o_3_out({\cb_7_8_io_o_3_out[7] ,
    \cb_7_8_io_o_3_out[6] ,
    \cb_7_8_io_o_3_out[5] ,
    \cb_7_8_io_o_3_out[4] ,
    \cb_7_8_io_o_3_out[3] ,
    \cb_7_8_io_o_3_out[2] ,
    \cb_7_8_io_o_3_out[1] ,
    \cb_7_8_io_o_3_out[0] }),
    .io_o_4_out({\cb_7_8_io_o_4_out[7] ,
    \cb_7_8_io_o_4_out[6] ,
    \cb_7_8_io_o_4_out[5] ,
    \cb_7_8_io_o_4_out[4] ,
    \cb_7_8_io_o_4_out[3] ,
    \cb_7_8_io_o_4_out[2] ,
    \cb_7_8_io_o_4_out[1] ,
    \cb_7_8_io_o_4_out[0] }),
    .io_o_5_out({\cb_7_8_io_o_5_out[7] ,
    \cb_7_8_io_o_5_out[6] ,
    \cb_7_8_io_o_5_out[5] ,
    \cb_7_8_io_o_5_out[4] ,
    \cb_7_8_io_o_5_out[3] ,
    \cb_7_8_io_o_5_out[2] ,
    \cb_7_8_io_o_5_out[1] ,
    \cb_7_8_io_o_5_out[0] }),
    .io_o_6_out({\cb_7_8_io_o_6_out[7] ,
    \cb_7_8_io_o_6_out[6] ,
    \cb_7_8_io_o_6_out[5] ,
    \cb_7_8_io_o_6_out[4] ,
    \cb_7_8_io_o_6_out[3] ,
    \cb_7_8_io_o_6_out[2] ,
    \cb_7_8_io_o_6_out[1] ,
    \cb_7_8_io_o_6_out[0] }),
    .io_o_7_out({\cb_7_8_io_o_7_out[7] ,
    \cb_7_8_io_o_7_out[6] ,
    \cb_7_8_io_o_7_out[5] ,
    \cb_7_8_io_o_7_out[4] ,
    \cb_7_8_io_o_7_out[3] ,
    \cb_7_8_io_o_7_out[2] ,
    \cb_7_8_io_o_7_out[1] ,
    \cb_7_8_io_o_7_out[0] }),
    .io_wo({\cb_7_7_io_eo[63] ,
    \cb_7_7_io_eo[62] ,
    \cb_7_7_io_eo[61] ,
    \cb_7_7_io_eo[60] ,
    \cb_7_7_io_eo[59] ,
    \cb_7_7_io_eo[58] ,
    \cb_7_7_io_eo[57] ,
    \cb_7_7_io_eo[56] ,
    \cb_7_7_io_eo[55] ,
    \cb_7_7_io_eo[54] ,
    \cb_7_7_io_eo[53] ,
    \cb_7_7_io_eo[52] ,
    \cb_7_7_io_eo[51] ,
    \cb_7_7_io_eo[50] ,
    \cb_7_7_io_eo[49] ,
    \cb_7_7_io_eo[48] ,
    \cb_7_7_io_eo[47] ,
    \cb_7_7_io_eo[46] ,
    \cb_7_7_io_eo[45] ,
    \cb_7_7_io_eo[44] ,
    \cb_7_7_io_eo[43] ,
    \cb_7_7_io_eo[42] ,
    \cb_7_7_io_eo[41] ,
    \cb_7_7_io_eo[40] ,
    \cb_7_7_io_eo[39] ,
    \cb_7_7_io_eo[38] ,
    \cb_7_7_io_eo[37] ,
    \cb_7_7_io_eo[36] ,
    \cb_7_7_io_eo[35] ,
    \cb_7_7_io_eo[34] ,
    \cb_7_7_io_eo[33] ,
    \cb_7_7_io_eo[32] ,
    \cb_7_7_io_eo[31] ,
    \cb_7_7_io_eo[30] ,
    \cb_7_7_io_eo[29] ,
    \cb_7_7_io_eo[28] ,
    \cb_7_7_io_eo[27] ,
    \cb_7_7_io_eo[26] ,
    \cb_7_7_io_eo[25] ,
    \cb_7_7_io_eo[24] ,
    \cb_7_7_io_eo[23] ,
    \cb_7_7_io_eo[22] ,
    \cb_7_7_io_eo[21] ,
    \cb_7_7_io_eo[20] ,
    \cb_7_7_io_eo[19] ,
    \cb_7_7_io_eo[18] ,
    \cb_7_7_io_eo[17] ,
    \cb_7_7_io_eo[16] ,
    \cb_7_7_io_eo[15] ,
    \cb_7_7_io_eo[14] ,
    \cb_7_7_io_eo[13] ,
    \cb_7_7_io_eo[12] ,
    \cb_7_7_io_eo[11] ,
    \cb_7_7_io_eo[10] ,
    \cb_7_7_io_eo[9] ,
    \cb_7_7_io_eo[8] ,
    \cb_7_7_io_eo[7] ,
    \cb_7_7_io_eo[6] ,
    \cb_7_7_io_eo[5] ,
    \cb_7_7_io_eo[4] ,
    \cb_7_7_io_eo[3] ,
    \cb_7_7_io_eo[2] ,
    \cb_7_7_io_eo[1] ,
    \cb_7_7_io_eo[0] }));
 cic_block cb_7_9 (.io_cs_i(cb_7_9_io_cs_i),
    .io_i_0_ci(cb_7_8_io_o_0_co),
    .io_i_1_ci(cb_7_8_io_o_1_co),
    .io_i_2_ci(cb_7_8_io_o_2_co),
    .io_i_3_ci(cb_7_8_io_o_3_co),
    .io_i_4_ci(cb_7_8_io_o_4_co),
    .io_i_5_ci(cb_7_8_io_o_5_co),
    .io_i_6_ci(cb_7_8_io_o_6_co),
    .io_i_7_ci(cb_7_8_io_o_7_co),
    .io_o_0_co(cb_7_10_io_i_0_ci),
    .io_o_1_co(cb_7_10_io_i_1_ci),
    .io_o_2_co(cb_7_10_io_i_2_ci),
    .io_o_3_co(cb_7_10_io_i_3_ci),
    .io_o_4_co(cb_7_10_io_i_4_ci),
    .io_o_5_co(cb_7_10_io_i_5_ci),
    .io_o_6_co(cb_7_10_io_i_6_ci),
    .io_o_7_co(cb_7_10_io_i_7_ci),
    .io_vci(cb_7_8_io_vco),
    .io_vco(cb_7_10_io_vci),
    .io_vi(cb_7_9_io_vi),
    .io_we_i(cb_7_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\cb_7_0_io_adr_i[1] ,
    \cb_7_0_io_adr_i[0] }),
    .io_dat_i({\cb_7_0_io_dat_i[15] ,
    \cb_7_0_io_dat_i[14] ,
    \cb_7_0_io_dat_i[13] ,
    \cb_7_0_io_dat_i[12] ,
    \cb_7_0_io_dat_i[11] ,
    \cb_7_0_io_dat_i[10] ,
    \cb_7_0_io_dat_i[9] ,
    \cb_7_0_io_dat_i[8] ,
    \cb_7_0_io_dat_i[7] ,
    \cb_7_0_io_dat_i[6] ,
    \cb_7_0_io_dat_i[5] ,
    \cb_7_0_io_dat_i[4] ,
    \cb_7_0_io_dat_i[3] ,
    \cb_7_0_io_dat_i[2] ,
    \cb_7_0_io_dat_i[1] ,
    \cb_7_0_io_dat_i[0] }),
    .io_dat_o({\cb_7_9_io_dat_o[15] ,
    \cb_7_9_io_dat_o[14] ,
    \cb_7_9_io_dat_o[13] ,
    \cb_7_9_io_dat_o[12] ,
    \cb_7_9_io_dat_o[11] ,
    \cb_7_9_io_dat_o[10] ,
    \cb_7_9_io_dat_o[9] ,
    \cb_7_9_io_dat_o[8] ,
    \cb_7_9_io_dat_o[7] ,
    \cb_7_9_io_dat_o[6] ,
    \cb_7_9_io_dat_o[5] ,
    \cb_7_9_io_dat_o[4] ,
    \cb_7_9_io_dat_o[3] ,
    \cb_7_9_io_dat_o[2] ,
    \cb_7_9_io_dat_o[1] ,
    \cb_7_9_io_dat_o[0] }),
    .io_eo({\cb_7_10_io_wo[63] ,
    \cb_7_10_io_wo[62] ,
    \cb_7_10_io_wo[61] ,
    \cb_7_10_io_wo[60] ,
    \cb_7_10_io_wo[59] ,
    \cb_7_10_io_wo[58] ,
    \cb_7_10_io_wo[57] ,
    \cb_7_10_io_wo[56] ,
    \cb_7_10_io_wo[55] ,
    \cb_7_10_io_wo[54] ,
    \cb_7_10_io_wo[53] ,
    \cb_7_10_io_wo[52] ,
    \cb_7_10_io_wo[51] ,
    \cb_7_10_io_wo[50] ,
    \cb_7_10_io_wo[49] ,
    \cb_7_10_io_wo[48] ,
    \cb_7_10_io_wo[47] ,
    \cb_7_10_io_wo[46] ,
    \cb_7_10_io_wo[45] ,
    \cb_7_10_io_wo[44] ,
    \cb_7_10_io_wo[43] ,
    \cb_7_10_io_wo[42] ,
    \cb_7_10_io_wo[41] ,
    \cb_7_10_io_wo[40] ,
    \cb_7_10_io_wo[39] ,
    \cb_7_10_io_wo[38] ,
    \cb_7_10_io_wo[37] ,
    \cb_7_10_io_wo[36] ,
    \cb_7_10_io_wo[35] ,
    \cb_7_10_io_wo[34] ,
    \cb_7_10_io_wo[33] ,
    \cb_7_10_io_wo[32] ,
    \cb_7_10_io_wo[31] ,
    \cb_7_10_io_wo[30] ,
    \cb_7_10_io_wo[29] ,
    \cb_7_10_io_wo[28] ,
    \cb_7_10_io_wo[27] ,
    \cb_7_10_io_wo[26] ,
    \cb_7_10_io_wo[25] ,
    \cb_7_10_io_wo[24] ,
    \cb_7_10_io_wo[23] ,
    \cb_7_10_io_wo[22] ,
    \cb_7_10_io_wo[21] ,
    \cb_7_10_io_wo[20] ,
    \cb_7_10_io_wo[19] ,
    \cb_7_10_io_wo[18] ,
    \cb_7_10_io_wo[17] ,
    \cb_7_10_io_wo[16] ,
    \cb_7_10_io_wo[15] ,
    \cb_7_10_io_wo[14] ,
    \cb_7_10_io_wo[13] ,
    \cb_7_10_io_wo[12] ,
    \cb_7_10_io_wo[11] ,
    \cb_7_10_io_wo[10] ,
    \cb_7_10_io_wo[9] ,
    \cb_7_10_io_wo[8] ,
    \cb_7_10_io_wo[7] ,
    \cb_7_10_io_wo[6] ,
    \cb_7_10_io_wo[5] ,
    \cb_7_10_io_wo[4] ,
    \cb_7_10_io_wo[3] ,
    \cb_7_10_io_wo[2] ,
    \cb_7_10_io_wo[1] ,
    \cb_7_10_io_wo[0] }),
    .io_i_0_in1({\cb_7_8_io_o_0_out[7] ,
    \cb_7_8_io_o_0_out[6] ,
    \cb_7_8_io_o_0_out[5] ,
    \cb_7_8_io_o_0_out[4] ,
    \cb_7_8_io_o_0_out[3] ,
    \cb_7_8_io_o_0_out[2] ,
    \cb_7_8_io_o_0_out[1] ,
    \cb_7_8_io_o_0_out[0] }),
    .io_i_1_in1({\cb_7_8_io_o_1_out[7] ,
    \cb_7_8_io_o_1_out[6] ,
    \cb_7_8_io_o_1_out[5] ,
    \cb_7_8_io_o_1_out[4] ,
    \cb_7_8_io_o_1_out[3] ,
    \cb_7_8_io_o_1_out[2] ,
    \cb_7_8_io_o_1_out[1] ,
    \cb_7_8_io_o_1_out[0] }),
    .io_i_2_in1({\cb_7_8_io_o_2_out[7] ,
    \cb_7_8_io_o_2_out[6] ,
    \cb_7_8_io_o_2_out[5] ,
    \cb_7_8_io_o_2_out[4] ,
    \cb_7_8_io_o_2_out[3] ,
    \cb_7_8_io_o_2_out[2] ,
    \cb_7_8_io_o_2_out[1] ,
    \cb_7_8_io_o_2_out[0] }),
    .io_i_3_in1({\cb_7_8_io_o_3_out[7] ,
    \cb_7_8_io_o_3_out[6] ,
    \cb_7_8_io_o_3_out[5] ,
    \cb_7_8_io_o_3_out[4] ,
    \cb_7_8_io_o_3_out[3] ,
    \cb_7_8_io_o_3_out[2] ,
    \cb_7_8_io_o_3_out[1] ,
    \cb_7_8_io_o_3_out[0] }),
    .io_i_4_in1({\cb_7_8_io_o_4_out[7] ,
    \cb_7_8_io_o_4_out[6] ,
    \cb_7_8_io_o_4_out[5] ,
    \cb_7_8_io_o_4_out[4] ,
    \cb_7_8_io_o_4_out[3] ,
    \cb_7_8_io_o_4_out[2] ,
    \cb_7_8_io_o_4_out[1] ,
    \cb_7_8_io_o_4_out[0] }),
    .io_i_5_in1({\cb_7_8_io_o_5_out[7] ,
    \cb_7_8_io_o_5_out[6] ,
    \cb_7_8_io_o_5_out[5] ,
    \cb_7_8_io_o_5_out[4] ,
    \cb_7_8_io_o_5_out[3] ,
    \cb_7_8_io_o_5_out[2] ,
    \cb_7_8_io_o_5_out[1] ,
    \cb_7_8_io_o_5_out[0] }),
    .io_i_6_in1({\cb_7_8_io_o_6_out[7] ,
    \cb_7_8_io_o_6_out[6] ,
    \cb_7_8_io_o_6_out[5] ,
    \cb_7_8_io_o_6_out[4] ,
    \cb_7_8_io_o_6_out[3] ,
    \cb_7_8_io_o_6_out[2] ,
    \cb_7_8_io_o_6_out[1] ,
    \cb_7_8_io_o_6_out[0] }),
    .io_i_7_in1({\cb_7_8_io_o_7_out[7] ,
    \cb_7_8_io_o_7_out[6] ,
    \cb_7_8_io_o_7_out[5] ,
    \cb_7_8_io_o_7_out[4] ,
    \cb_7_8_io_o_7_out[3] ,
    \cb_7_8_io_o_7_out[2] ,
    \cb_7_8_io_o_7_out[1] ,
    \cb_7_8_io_o_7_out[0] }),
    .io_o_0_out({\cb_7_10_io_i_0_in1[7] ,
    \cb_7_10_io_i_0_in1[6] ,
    \cb_7_10_io_i_0_in1[5] ,
    \cb_7_10_io_i_0_in1[4] ,
    \cb_7_10_io_i_0_in1[3] ,
    \cb_7_10_io_i_0_in1[2] ,
    \cb_7_10_io_i_0_in1[1] ,
    \cb_7_10_io_i_0_in1[0] }),
    .io_o_1_out({\cb_7_10_io_i_1_in1[7] ,
    \cb_7_10_io_i_1_in1[6] ,
    \cb_7_10_io_i_1_in1[5] ,
    \cb_7_10_io_i_1_in1[4] ,
    \cb_7_10_io_i_1_in1[3] ,
    \cb_7_10_io_i_1_in1[2] ,
    \cb_7_10_io_i_1_in1[1] ,
    \cb_7_10_io_i_1_in1[0] }),
    .io_o_2_out({\cb_7_10_io_i_2_in1[7] ,
    \cb_7_10_io_i_2_in1[6] ,
    \cb_7_10_io_i_2_in1[5] ,
    \cb_7_10_io_i_2_in1[4] ,
    \cb_7_10_io_i_2_in1[3] ,
    \cb_7_10_io_i_2_in1[2] ,
    \cb_7_10_io_i_2_in1[1] ,
    \cb_7_10_io_i_2_in1[0] }),
    .io_o_3_out({\cb_7_10_io_i_3_in1[7] ,
    \cb_7_10_io_i_3_in1[6] ,
    \cb_7_10_io_i_3_in1[5] ,
    \cb_7_10_io_i_3_in1[4] ,
    \cb_7_10_io_i_3_in1[3] ,
    \cb_7_10_io_i_3_in1[2] ,
    \cb_7_10_io_i_3_in1[1] ,
    \cb_7_10_io_i_3_in1[0] }),
    .io_o_4_out({\cb_7_10_io_i_4_in1[7] ,
    \cb_7_10_io_i_4_in1[6] ,
    \cb_7_10_io_i_4_in1[5] ,
    \cb_7_10_io_i_4_in1[4] ,
    \cb_7_10_io_i_4_in1[3] ,
    \cb_7_10_io_i_4_in1[2] ,
    \cb_7_10_io_i_4_in1[1] ,
    \cb_7_10_io_i_4_in1[0] }),
    .io_o_5_out({\cb_7_10_io_i_5_in1[7] ,
    \cb_7_10_io_i_5_in1[6] ,
    \cb_7_10_io_i_5_in1[5] ,
    \cb_7_10_io_i_5_in1[4] ,
    \cb_7_10_io_i_5_in1[3] ,
    \cb_7_10_io_i_5_in1[2] ,
    \cb_7_10_io_i_5_in1[1] ,
    \cb_7_10_io_i_5_in1[0] }),
    .io_o_6_out({\cb_7_10_io_i_6_in1[7] ,
    \cb_7_10_io_i_6_in1[6] ,
    \cb_7_10_io_i_6_in1[5] ,
    \cb_7_10_io_i_6_in1[4] ,
    \cb_7_10_io_i_6_in1[3] ,
    \cb_7_10_io_i_6_in1[2] ,
    \cb_7_10_io_i_6_in1[1] ,
    \cb_7_10_io_i_6_in1[0] }),
    .io_o_7_out({\cb_7_10_io_i_7_in1[7] ,
    \cb_7_10_io_i_7_in1[6] ,
    \cb_7_10_io_i_7_in1[5] ,
    \cb_7_10_io_i_7_in1[4] ,
    \cb_7_10_io_i_7_in1[3] ,
    \cb_7_10_io_i_7_in1[2] ,
    \cb_7_10_io_i_7_in1[1] ,
    \cb_7_10_io_i_7_in1[0] }),
    .io_wo({\cb_7_8_io_eo[63] ,
    \cb_7_8_io_eo[62] ,
    \cb_7_8_io_eo[61] ,
    \cb_7_8_io_eo[60] ,
    \cb_7_8_io_eo[59] ,
    \cb_7_8_io_eo[58] ,
    \cb_7_8_io_eo[57] ,
    \cb_7_8_io_eo[56] ,
    \cb_7_8_io_eo[55] ,
    \cb_7_8_io_eo[54] ,
    \cb_7_8_io_eo[53] ,
    \cb_7_8_io_eo[52] ,
    \cb_7_8_io_eo[51] ,
    \cb_7_8_io_eo[50] ,
    \cb_7_8_io_eo[49] ,
    \cb_7_8_io_eo[48] ,
    \cb_7_8_io_eo[47] ,
    \cb_7_8_io_eo[46] ,
    \cb_7_8_io_eo[45] ,
    \cb_7_8_io_eo[44] ,
    \cb_7_8_io_eo[43] ,
    \cb_7_8_io_eo[42] ,
    \cb_7_8_io_eo[41] ,
    \cb_7_8_io_eo[40] ,
    \cb_7_8_io_eo[39] ,
    \cb_7_8_io_eo[38] ,
    \cb_7_8_io_eo[37] ,
    \cb_7_8_io_eo[36] ,
    \cb_7_8_io_eo[35] ,
    \cb_7_8_io_eo[34] ,
    \cb_7_8_io_eo[33] ,
    \cb_7_8_io_eo[32] ,
    \cb_7_8_io_eo[31] ,
    \cb_7_8_io_eo[30] ,
    \cb_7_8_io_eo[29] ,
    \cb_7_8_io_eo[28] ,
    \cb_7_8_io_eo[27] ,
    \cb_7_8_io_eo[26] ,
    \cb_7_8_io_eo[25] ,
    \cb_7_8_io_eo[24] ,
    \cb_7_8_io_eo[23] ,
    \cb_7_8_io_eo[22] ,
    \cb_7_8_io_eo[21] ,
    \cb_7_8_io_eo[20] ,
    \cb_7_8_io_eo[19] ,
    \cb_7_8_io_eo[18] ,
    \cb_7_8_io_eo[17] ,
    \cb_7_8_io_eo[16] ,
    \cb_7_8_io_eo[15] ,
    \cb_7_8_io_eo[14] ,
    \cb_7_8_io_eo[13] ,
    \cb_7_8_io_eo[12] ,
    \cb_7_8_io_eo[11] ,
    \cb_7_8_io_eo[10] ,
    \cb_7_8_io_eo[9] ,
    \cb_7_8_io_eo[8] ,
    \cb_7_8_io_eo[7] ,
    \cb_7_8_io_eo[6] ,
    \cb_7_8_io_eo[5] ,
    \cb_7_8_io_eo[4] ,
    \cb_7_8_io_eo[3] ,
    \cb_7_8_io_eo[2] ,
    \cb_7_8_io_eo[1] ,
    \cb_7_8_io_eo[0] }));
 cic_con ccon_0 (.io_ack_o(\_T_167[4] ),
    .io_b_cs_i_0(cb_0_0_io_cs_i),
    .io_b_cs_i_1(cb_0_1_io_cs_i),
    .io_b_cs_i_10(cb_0_10_io_cs_i),
    .io_b_cs_i_2(cb_0_2_io_cs_i),
    .io_b_cs_i_3(cb_0_3_io_cs_i),
    .io_b_cs_i_4(cb_0_4_io_cs_i),
    .io_b_cs_i_5(cb_0_5_io_cs_i),
    .io_b_cs_i_6(cb_0_6_io_cs_i),
    .io_b_cs_i_7(cb_0_7_io_cs_i),
    .io_b_cs_i_8(cb_0_8_io_cs_i),
    .io_b_cs_i_9(cb_0_9_io_cs_i),
    .io_b_we_i(cb_0_0_io_we_i),
    .io_cs_i(ccon_0_io_cs_i),
    .io_dsi_o(cb_0_0_io_i_0_ci),
    .io_irq(\_T_178[4] ),
    .io_we_i(ccon_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\ccon_0_io_adr_i[11] ,
    \ccon_0_io_adr_i[10] ,
    \ccon_0_io_adr_i[9] ,
    \ccon_0_io_adr_i[8] ,
    \ccon_0_io_adr_i[7] ,
    \ccon_0_io_adr_i[6] ,
    \ccon_0_io_adr_i[5] ,
    \ccon_0_io_adr_i[4] ,
    \ccon_0_io_adr_i[3] ,
    \ccon_0_io_adr_i[2] ,
    \ccon_0_io_adr_i[1] ,
    \ccon_0_io_adr_i[0] }),
    .io_b_adr_i({\cb_0_0_io_adr_i[1] ,
    \cb_0_0_io_adr_i[0] }),
    .io_b_dat_i({\cb_0_0_io_dat_i[15] ,
    \cb_0_0_io_dat_i[14] ,
    \cb_0_0_io_dat_i[13] ,
    \cb_0_0_io_dat_i[12] ,
    \cb_0_0_io_dat_i[11] ,
    \cb_0_0_io_dat_i[10] ,
    \cb_0_0_io_dat_i[9] ,
    \cb_0_0_io_dat_i[8] ,
    \cb_0_0_io_dat_i[7] ,
    \cb_0_0_io_dat_i[6] ,
    \cb_0_0_io_dat_i[5] ,
    \cb_0_0_io_dat_i[4] ,
    \cb_0_0_io_dat_i[3] ,
    \cb_0_0_io_dat_i[2] ,
    \cb_0_0_io_dat_i[1] ,
    \cb_0_0_io_dat_i[0] }),
    .io_b_dat_o_0({\cb_0_0_io_dat_o[15] ,
    \cb_0_0_io_dat_o[14] ,
    \cb_0_0_io_dat_o[13] ,
    \cb_0_0_io_dat_o[12] ,
    \cb_0_0_io_dat_o[11] ,
    \cb_0_0_io_dat_o[10] ,
    \cb_0_0_io_dat_o[9] ,
    \cb_0_0_io_dat_o[8] ,
    \cb_0_0_io_dat_o[7] ,
    \cb_0_0_io_dat_o[6] ,
    \cb_0_0_io_dat_o[5] ,
    \cb_0_0_io_dat_o[4] ,
    \cb_0_0_io_dat_o[3] ,
    \cb_0_0_io_dat_o[2] ,
    \cb_0_0_io_dat_o[1] ,
    \cb_0_0_io_dat_o[0] }),
    .io_b_dat_o_1({\cb_0_1_io_dat_o[15] ,
    \cb_0_1_io_dat_o[14] ,
    \cb_0_1_io_dat_o[13] ,
    \cb_0_1_io_dat_o[12] ,
    \cb_0_1_io_dat_o[11] ,
    \cb_0_1_io_dat_o[10] ,
    \cb_0_1_io_dat_o[9] ,
    \cb_0_1_io_dat_o[8] ,
    \cb_0_1_io_dat_o[7] ,
    \cb_0_1_io_dat_o[6] ,
    \cb_0_1_io_dat_o[5] ,
    \cb_0_1_io_dat_o[4] ,
    \cb_0_1_io_dat_o[3] ,
    \cb_0_1_io_dat_o[2] ,
    \cb_0_1_io_dat_o[1] ,
    \cb_0_1_io_dat_o[0] }),
    .io_b_dat_o_10({\cb_0_10_io_dat_o[15] ,
    \cb_0_10_io_dat_o[14] ,
    \cb_0_10_io_dat_o[13] ,
    \cb_0_10_io_dat_o[12] ,
    \cb_0_10_io_dat_o[11] ,
    \cb_0_10_io_dat_o[10] ,
    \cb_0_10_io_dat_o[9] ,
    \cb_0_10_io_dat_o[8] ,
    \cb_0_10_io_dat_o[7] ,
    \cb_0_10_io_dat_o[6] ,
    \cb_0_10_io_dat_o[5] ,
    \cb_0_10_io_dat_o[4] ,
    \cb_0_10_io_dat_o[3] ,
    \cb_0_10_io_dat_o[2] ,
    \cb_0_10_io_dat_o[1] ,
    \cb_0_10_io_dat_o[0] }),
    .io_b_dat_o_2({\cb_0_2_io_dat_o[15] ,
    \cb_0_2_io_dat_o[14] ,
    \cb_0_2_io_dat_o[13] ,
    \cb_0_2_io_dat_o[12] ,
    \cb_0_2_io_dat_o[11] ,
    \cb_0_2_io_dat_o[10] ,
    \cb_0_2_io_dat_o[9] ,
    \cb_0_2_io_dat_o[8] ,
    \cb_0_2_io_dat_o[7] ,
    \cb_0_2_io_dat_o[6] ,
    \cb_0_2_io_dat_o[5] ,
    \cb_0_2_io_dat_o[4] ,
    \cb_0_2_io_dat_o[3] ,
    \cb_0_2_io_dat_o[2] ,
    \cb_0_2_io_dat_o[1] ,
    \cb_0_2_io_dat_o[0] }),
    .io_b_dat_o_3({\cb_0_3_io_dat_o[15] ,
    \cb_0_3_io_dat_o[14] ,
    \cb_0_3_io_dat_o[13] ,
    \cb_0_3_io_dat_o[12] ,
    \cb_0_3_io_dat_o[11] ,
    \cb_0_3_io_dat_o[10] ,
    \cb_0_3_io_dat_o[9] ,
    \cb_0_3_io_dat_o[8] ,
    \cb_0_3_io_dat_o[7] ,
    \cb_0_3_io_dat_o[6] ,
    \cb_0_3_io_dat_o[5] ,
    \cb_0_3_io_dat_o[4] ,
    \cb_0_3_io_dat_o[3] ,
    \cb_0_3_io_dat_o[2] ,
    \cb_0_3_io_dat_o[1] ,
    \cb_0_3_io_dat_o[0] }),
    .io_b_dat_o_4({\cb_0_4_io_dat_o[15] ,
    \cb_0_4_io_dat_o[14] ,
    \cb_0_4_io_dat_o[13] ,
    \cb_0_4_io_dat_o[12] ,
    \cb_0_4_io_dat_o[11] ,
    \cb_0_4_io_dat_o[10] ,
    \cb_0_4_io_dat_o[9] ,
    \cb_0_4_io_dat_o[8] ,
    \cb_0_4_io_dat_o[7] ,
    \cb_0_4_io_dat_o[6] ,
    \cb_0_4_io_dat_o[5] ,
    \cb_0_4_io_dat_o[4] ,
    \cb_0_4_io_dat_o[3] ,
    \cb_0_4_io_dat_o[2] ,
    \cb_0_4_io_dat_o[1] ,
    \cb_0_4_io_dat_o[0] }),
    .io_b_dat_o_5({\cb_0_5_io_dat_o[15] ,
    \cb_0_5_io_dat_o[14] ,
    \cb_0_5_io_dat_o[13] ,
    \cb_0_5_io_dat_o[12] ,
    \cb_0_5_io_dat_o[11] ,
    \cb_0_5_io_dat_o[10] ,
    \cb_0_5_io_dat_o[9] ,
    \cb_0_5_io_dat_o[8] ,
    \cb_0_5_io_dat_o[7] ,
    \cb_0_5_io_dat_o[6] ,
    \cb_0_5_io_dat_o[5] ,
    \cb_0_5_io_dat_o[4] ,
    \cb_0_5_io_dat_o[3] ,
    \cb_0_5_io_dat_o[2] ,
    \cb_0_5_io_dat_o[1] ,
    \cb_0_5_io_dat_o[0] }),
    .io_b_dat_o_6({\cb_0_6_io_dat_o[15] ,
    \cb_0_6_io_dat_o[14] ,
    \cb_0_6_io_dat_o[13] ,
    \cb_0_6_io_dat_o[12] ,
    \cb_0_6_io_dat_o[11] ,
    \cb_0_6_io_dat_o[10] ,
    \cb_0_6_io_dat_o[9] ,
    \cb_0_6_io_dat_o[8] ,
    \cb_0_6_io_dat_o[7] ,
    \cb_0_6_io_dat_o[6] ,
    \cb_0_6_io_dat_o[5] ,
    \cb_0_6_io_dat_o[4] ,
    \cb_0_6_io_dat_o[3] ,
    \cb_0_6_io_dat_o[2] ,
    \cb_0_6_io_dat_o[1] ,
    \cb_0_6_io_dat_o[0] }),
    .io_b_dat_o_7({\cb_0_7_io_dat_o[15] ,
    \cb_0_7_io_dat_o[14] ,
    \cb_0_7_io_dat_o[13] ,
    \cb_0_7_io_dat_o[12] ,
    \cb_0_7_io_dat_o[11] ,
    \cb_0_7_io_dat_o[10] ,
    \cb_0_7_io_dat_o[9] ,
    \cb_0_7_io_dat_o[8] ,
    \cb_0_7_io_dat_o[7] ,
    \cb_0_7_io_dat_o[6] ,
    \cb_0_7_io_dat_o[5] ,
    \cb_0_7_io_dat_o[4] ,
    \cb_0_7_io_dat_o[3] ,
    \cb_0_7_io_dat_o[2] ,
    \cb_0_7_io_dat_o[1] ,
    \cb_0_7_io_dat_o[0] }),
    .io_b_dat_o_8({\cb_0_8_io_dat_o[15] ,
    \cb_0_8_io_dat_o[14] ,
    \cb_0_8_io_dat_o[13] ,
    \cb_0_8_io_dat_o[12] ,
    \cb_0_8_io_dat_o[11] ,
    \cb_0_8_io_dat_o[10] ,
    \cb_0_8_io_dat_o[9] ,
    \cb_0_8_io_dat_o[8] ,
    \cb_0_8_io_dat_o[7] ,
    \cb_0_8_io_dat_o[6] ,
    \cb_0_8_io_dat_o[5] ,
    \cb_0_8_io_dat_o[4] ,
    \cb_0_8_io_dat_o[3] ,
    \cb_0_8_io_dat_o[2] ,
    \cb_0_8_io_dat_o[1] ,
    \cb_0_8_io_dat_o[0] }),
    .io_b_dat_o_9({\cb_0_9_io_dat_o[15] ,
    \cb_0_9_io_dat_o[14] ,
    \cb_0_9_io_dat_o[13] ,
    \cb_0_9_io_dat_o[12] ,
    \cb_0_9_io_dat_o[11] ,
    \cb_0_9_io_dat_o[10] ,
    \cb_0_9_io_dat_o[9] ,
    \cb_0_9_io_dat_o[8] ,
    \cb_0_9_io_dat_o[7] ,
    \cb_0_9_io_dat_o[6] ,
    \cb_0_9_io_dat_o[5] ,
    \cb_0_9_io_dat_o[4] ,
    \cb_0_9_io_dat_o[3] ,
    \cb_0_9_io_dat_o[2] ,
    \cb_0_9_io_dat_o[1] ,
    \cb_0_9_io_dat_o[0] }),
    .io_dat_i({\ccon_0_io_dat_i[31] ,
    \ccon_0_io_dat_i[30] ,
    \ccon_0_io_dat_i[29] ,
    \ccon_0_io_dat_i[28] ,
    \ccon_0_io_dat_i[27] ,
    \ccon_0_io_dat_i[26] ,
    \ccon_0_io_dat_i[25] ,
    \ccon_0_io_dat_i[24] ,
    \ccon_0_io_dat_i[23] ,
    \ccon_0_io_dat_i[22] ,
    \ccon_0_io_dat_i[21] ,
    \ccon_0_io_dat_i[20] ,
    \ccon_0_io_dat_i[19] ,
    \ccon_0_io_dat_i[18] ,
    \ccon_0_io_dat_i[17] ,
    \ccon_0_io_dat_i[16] ,
    \ccon_0_io_dat_i[15] ,
    \ccon_0_io_dat_i[14] ,
    \ccon_0_io_dat_i[13] ,
    \ccon_0_io_dat_i[12] ,
    \ccon_0_io_dat_i[11] ,
    \ccon_0_io_dat_i[10] ,
    \ccon_0_io_dat_i[9] ,
    \ccon_0_io_dat_i[8] ,
    \ccon_0_io_dat_i[7] ,
    \ccon_0_io_dat_i[6] ,
    \ccon_0_io_dat_i[5] ,
    \ccon_0_io_dat_i[4] ,
    \ccon_0_io_dat_i[3] ,
    \ccon_0_io_dat_i[2] ,
    \ccon_0_io_dat_i[1] ,
    \ccon_0_io_dat_i[0] }),
    .io_dat_o({\ccon_0_io_dat_o[31] ,
    \ccon_0_io_dat_o[30] ,
    \ccon_0_io_dat_o[29] ,
    \ccon_0_io_dat_o[28] ,
    \ccon_0_io_dat_o[27] ,
    \ccon_0_io_dat_o[26] ,
    \ccon_0_io_dat_o[25] ,
    \ccon_0_io_dat_o[24] ,
    \ccon_0_io_dat_o[23] ,
    \ccon_0_io_dat_o[22] ,
    \ccon_0_io_dat_o[21] ,
    \ccon_0_io_dat_o[20] ,
    \ccon_0_io_dat_o[19] ,
    \ccon_0_io_dat_o[18] ,
    \ccon_0_io_dat_o[17] ,
    \ccon_0_io_dat_o[16] ,
    \ccon_0_io_dat_o[15] ,
    \ccon_0_io_dat_o[14] ,
    \ccon_0_io_dat_o[13] ,
    \ccon_0_io_dat_o[12] ,
    \ccon_0_io_dat_o[11] ,
    \ccon_0_io_dat_o[10] ,
    \ccon_0_io_dat_o[9] ,
    \ccon_0_io_dat_o[8] ,
    \ccon_0_io_dat_o[7] ,
    \ccon_0_io_dat_o[6] ,
    \ccon_0_io_dat_o[5] ,
    \ccon_0_io_dat_o[4] ,
    \ccon_0_io_dat_o[3] ,
    \ccon_0_io_dat_o[2] ,
    \ccon_0_io_dat_o[1] ,
    \ccon_0_io_dat_o[0] }),
    .io_dataLastBlock({\cb_0_0_io_wo[63] ,
    \cb_0_0_io_wo[62] ,
    \cb_0_0_io_wo[61] ,
    \cb_0_0_io_wo[60] ,
    \cb_0_0_io_wo[59] ,
    \cb_0_0_io_wo[58] ,
    \cb_0_0_io_wo[57] ,
    \cb_0_0_io_wo[56] ,
    \cb_0_0_io_wo[55] ,
    \cb_0_0_io_wo[54] ,
    \cb_0_0_io_wo[53] ,
    \cb_0_0_io_wo[52] ,
    \cb_0_0_io_wo[51] ,
    \cb_0_0_io_wo[50] ,
    \cb_0_0_io_wo[49] ,
    \cb_0_0_io_wo[48] ,
    \cb_0_0_io_wo[47] ,
    \cb_0_0_io_wo[46] ,
    \cb_0_0_io_wo[45] ,
    \cb_0_0_io_wo[44] ,
    \cb_0_0_io_wo[43] ,
    \cb_0_0_io_wo[42] ,
    \cb_0_0_io_wo[41] ,
    \cb_0_0_io_wo[40] ,
    \cb_0_0_io_wo[39] ,
    \cb_0_0_io_wo[38] ,
    \cb_0_0_io_wo[37] ,
    \cb_0_0_io_wo[36] ,
    \cb_0_0_io_wo[35] ,
    \cb_0_0_io_wo[34] ,
    \cb_0_0_io_wo[33] ,
    \cb_0_0_io_wo[32] ,
    \cb_0_0_io_wo[31] ,
    \cb_0_0_io_wo[30] ,
    \cb_0_0_io_wo[29] ,
    \cb_0_0_io_wo[28] ,
    \cb_0_0_io_wo[27] ,
    \cb_0_0_io_wo[26] ,
    \cb_0_0_io_wo[25] ,
    \cb_0_0_io_wo[24] ,
    \cb_0_0_io_wo[23] ,
    \cb_0_0_io_wo[22] ,
    \cb_0_0_io_wo[21] ,
    \cb_0_0_io_wo[20] ,
    \cb_0_0_io_wo[19] ,
    \cb_0_0_io_wo[18] ,
    \cb_0_0_io_wo[17] ,
    \cb_0_0_io_wo[16] ,
    \cb_0_0_io_wo[15] ,
    \cb_0_0_io_wo[14] ,
    \cb_0_0_io_wo[13] ,
    \cb_0_0_io_wo[12] ,
    \cb_0_0_io_wo[11] ,
    \cb_0_0_io_wo[10] ,
    \cb_0_0_io_wo[9] ,
    \cb_0_0_io_wo[8] ,
    \cb_0_0_io_wo[7] ,
    \cb_0_0_io_wo[6] ,
    \cb_0_0_io_wo[5] ,
    \cb_0_0_io_wo[4] ,
    \cb_0_0_io_wo[3] ,
    \cb_0_0_io_wo[2] ,
    \cb_0_0_io_wo[1] ,
    \cb_0_0_io_wo[0] }),
    .io_dsi_in({\ccon_0_io_dsi_in[7] ,
    \ccon_0_io_dsi_in[6] ,
    \ccon_0_io_dsi_in[5] ,
    \ccon_0_io_dsi_in[4] ,
    \ccon_0_io_dsi_in[3] ,
    \ccon_0_io_dsi_in[2] ,
    \ccon_0_io_dsi_in[1] ,
    \ccon_0_io_dsi_in[0] }),
    .io_vout({cb_0_10_io_vi,
    cb_0_9_io_vi,
    cb_0_8_io_vi,
    cb_0_7_io_vi,
    cb_0_6_io_vi,
    cb_0_5_io_vi,
    cb_0_4_io_vi,
    cb_0_3_io_vi,
    cb_0_2_io_vi,
    cb_0_1_io_vi,
    cb_0_0_io_vi}));
 cic_con ccon_1 (.io_ack_o(\_T_167[5] ),
    .io_b_cs_i_0(cb_1_0_io_cs_i),
    .io_b_cs_i_1(cb_1_1_io_cs_i),
    .io_b_cs_i_10(cb_1_10_io_cs_i),
    .io_b_cs_i_2(cb_1_2_io_cs_i),
    .io_b_cs_i_3(cb_1_3_io_cs_i),
    .io_b_cs_i_4(cb_1_4_io_cs_i),
    .io_b_cs_i_5(cb_1_5_io_cs_i),
    .io_b_cs_i_6(cb_1_6_io_cs_i),
    .io_b_cs_i_7(cb_1_7_io_cs_i),
    .io_b_cs_i_8(cb_1_8_io_cs_i),
    .io_b_cs_i_9(cb_1_9_io_cs_i),
    .io_b_we_i(cb_1_0_io_we_i),
    .io_cs_i(ccon_1_io_cs_i),
    .io_dsi_o(cb_1_0_io_i_0_ci),
    .io_irq(\_T_178[5] ),
    .io_we_i(ccon_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\ccon_0_io_adr_i[11] ,
    \ccon_0_io_adr_i[10] ,
    \ccon_0_io_adr_i[9] ,
    \ccon_0_io_adr_i[8] ,
    \ccon_0_io_adr_i[7] ,
    \ccon_0_io_adr_i[6] ,
    \ccon_0_io_adr_i[5] ,
    \ccon_0_io_adr_i[4] ,
    \ccon_0_io_adr_i[3] ,
    \ccon_0_io_adr_i[2] ,
    \ccon_0_io_adr_i[1] ,
    \ccon_0_io_adr_i[0] }),
    .io_b_adr_i({\cb_1_0_io_adr_i[1] ,
    \cb_1_0_io_adr_i[0] }),
    .io_b_dat_i({\cb_1_0_io_dat_i[15] ,
    \cb_1_0_io_dat_i[14] ,
    \cb_1_0_io_dat_i[13] ,
    \cb_1_0_io_dat_i[12] ,
    \cb_1_0_io_dat_i[11] ,
    \cb_1_0_io_dat_i[10] ,
    \cb_1_0_io_dat_i[9] ,
    \cb_1_0_io_dat_i[8] ,
    \cb_1_0_io_dat_i[7] ,
    \cb_1_0_io_dat_i[6] ,
    \cb_1_0_io_dat_i[5] ,
    \cb_1_0_io_dat_i[4] ,
    \cb_1_0_io_dat_i[3] ,
    \cb_1_0_io_dat_i[2] ,
    \cb_1_0_io_dat_i[1] ,
    \cb_1_0_io_dat_i[0] }),
    .io_b_dat_o_0({\cb_1_0_io_dat_o[15] ,
    \cb_1_0_io_dat_o[14] ,
    \cb_1_0_io_dat_o[13] ,
    \cb_1_0_io_dat_o[12] ,
    \cb_1_0_io_dat_o[11] ,
    \cb_1_0_io_dat_o[10] ,
    \cb_1_0_io_dat_o[9] ,
    \cb_1_0_io_dat_o[8] ,
    \cb_1_0_io_dat_o[7] ,
    \cb_1_0_io_dat_o[6] ,
    \cb_1_0_io_dat_o[5] ,
    \cb_1_0_io_dat_o[4] ,
    \cb_1_0_io_dat_o[3] ,
    \cb_1_0_io_dat_o[2] ,
    \cb_1_0_io_dat_o[1] ,
    \cb_1_0_io_dat_o[0] }),
    .io_b_dat_o_1({\cb_1_1_io_dat_o[15] ,
    \cb_1_1_io_dat_o[14] ,
    \cb_1_1_io_dat_o[13] ,
    \cb_1_1_io_dat_o[12] ,
    \cb_1_1_io_dat_o[11] ,
    \cb_1_1_io_dat_o[10] ,
    \cb_1_1_io_dat_o[9] ,
    \cb_1_1_io_dat_o[8] ,
    \cb_1_1_io_dat_o[7] ,
    \cb_1_1_io_dat_o[6] ,
    \cb_1_1_io_dat_o[5] ,
    \cb_1_1_io_dat_o[4] ,
    \cb_1_1_io_dat_o[3] ,
    \cb_1_1_io_dat_o[2] ,
    \cb_1_1_io_dat_o[1] ,
    \cb_1_1_io_dat_o[0] }),
    .io_b_dat_o_10({\cb_1_10_io_dat_o[15] ,
    \cb_1_10_io_dat_o[14] ,
    \cb_1_10_io_dat_o[13] ,
    \cb_1_10_io_dat_o[12] ,
    \cb_1_10_io_dat_o[11] ,
    \cb_1_10_io_dat_o[10] ,
    \cb_1_10_io_dat_o[9] ,
    \cb_1_10_io_dat_o[8] ,
    \cb_1_10_io_dat_o[7] ,
    \cb_1_10_io_dat_o[6] ,
    \cb_1_10_io_dat_o[5] ,
    \cb_1_10_io_dat_o[4] ,
    \cb_1_10_io_dat_o[3] ,
    \cb_1_10_io_dat_o[2] ,
    \cb_1_10_io_dat_o[1] ,
    \cb_1_10_io_dat_o[0] }),
    .io_b_dat_o_2({\cb_1_2_io_dat_o[15] ,
    \cb_1_2_io_dat_o[14] ,
    \cb_1_2_io_dat_o[13] ,
    \cb_1_2_io_dat_o[12] ,
    \cb_1_2_io_dat_o[11] ,
    \cb_1_2_io_dat_o[10] ,
    \cb_1_2_io_dat_o[9] ,
    \cb_1_2_io_dat_o[8] ,
    \cb_1_2_io_dat_o[7] ,
    \cb_1_2_io_dat_o[6] ,
    \cb_1_2_io_dat_o[5] ,
    \cb_1_2_io_dat_o[4] ,
    \cb_1_2_io_dat_o[3] ,
    \cb_1_2_io_dat_o[2] ,
    \cb_1_2_io_dat_o[1] ,
    \cb_1_2_io_dat_o[0] }),
    .io_b_dat_o_3({\cb_1_3_io_dat_o[15] ,
    \cb_1_3_io_dat_o[14] ,
    \cb_1_3_io_dat_o[13] ,
    \cb_1_3_io_dat_o[12] ,
    \cb_1_3_io_dat_o[11] ,
    \cb_1_3_io_dat_o[10] ,
    \cb_1_3_io_dat_o[9] ,
    \cb_1_3_io_dat_o[8] ,
    \cb_1_3_io_dat_o[7] ,
    \cb_1_3_io_dat_o[6] ,
    \cb_1_3_io_dat_o[5] ,
    \cb_1_3_io_dat_o[4] ,
    \cb_1_3_io_dat_o[3] ,
    \cb_1_3_io_dat_o[2] ,
    \cb_1_3_io_dat_o[1] ,
    \cb_1_3_io_dat_o[0] }),
    .io_b_dat_o_4({\cb_1_4_io_dat_o[15] ,
    \cb_1_4_io_dat_o[14] ,
    \cb_1_4_io_dat_o[13] ,
    \cb_1_4_io_dat_o[12] ,
    \cb_1_4_io_dat_o[11] ,
    \cb_1_4_io_dat_o[10] ,
    \cb_1_4_io_dat_o[9] ,
    \cb_1_4_io_dat_o[8] ,
    \cb_1_4_io_dat_o[7] ,
    \cb_1_4_io_dat_o[6] ,
    \cb_1_4_io_dat_o[5] ,
    \cb_1_4_io_dat_o[4] ,
    \cb_1_4_io_dat_o[3] ,
    \cb_1_4_io_dat_o[2] ,
    \cb_1_4_io_dat_o[1] ,
    \cb_1_4_io_dat_o[0] }),
    .io_b_dat_o_5({\cb_1_5_io_dat_o[15] ,
    \cb_1_5_io_dat_o[14] ,
    \cb_1_5_io_dat_o[13] ,
    \cb_1_5_io_dat_o[12] ,
    \cb_1_5_io_dat_o[11] ,
    \cb_1_5_io_dat_o[10] ,
    \cb_1_5_io_dat_o[9] ,
    \cb_1_5_io_dat_o[8] ,
    \cb_1_5_io_dat_o[7] ,
    \cb_1_5_io_dat_o[6] ,
    \cb_1_5_io_dat_o[5] ,
    \cb_1_5_io_dat_o[4] ,
    \cb_1_5_io_dat_o[3] ,
    \cb_1_5_io_dat_o[2] ,
    \cb_1_5_io_dat_o[1] ,
    \cb_1_5_io_dat_o[0] }),
    .io_b_dat_o_6({\cb_1_6_io_dat_o[15] ,
    \cb_1_6_io_dat_o[14] ,
    \cb_1_6_io_dat_o[13] ,
    \cb_1_6_io_dat_o[12] ,
    \cb_1_6_io_dat_o[11] ,
    \cb_1_6_io_dat_o[10] ,
    \cb_1_6_io_dat_o[9] ,
    \cb_1_6_io_dat_o[8] ,
    \cb_1_6_io_dat_o[7] ,
    \cb_1_6_io_dat_o[6] ,
    \cb_1_6_io_dat_o[5] ,
    \cb_1_6_io_dat_o[4] ,
    \cb_1_6_io_dat_o[3] ,
    \cb_1_6_io_dat_o[2] ,
    \cb_1_6_io_dat_o[1] ,
    \cb_1_6_io_dat_o[0] }),
    .io_b_dat_o_7({\cb_1_7_io_dat_o[15] ,
    \cb_1_7_io_dat_o[14] ,
    \cb_1_7_io_dat_o[13] ,
    \cb_1_7_io_dat_o[12] ,
    \cb_1_7_io_dat_o[11] ,
    \cb_1_7_io_dat_o[10] ,
    \cb_1_7_io_dat_o[9] ,
    \cb_1_7_io_dat_o[8] ,
    \cb_1_7_io_dat_o[7] ,
    \cb_1_7_io_dat_o[6] ,
    \cb_1_7_io_dat_o[5] ,
    \cb_1_7_io_dat_o[4] ,
    \cb_1_7_io_dat_o[3] ,
    \cb_1_7_io_dat_o[2] ,
    \cb_1_7_io_dat_o[1] ,
    \cb_1_7_io_dat_o[0] }),
    .io_b_dat_o_8({\cb_1_8_io_dat_o[15] ,
    \cb_1_8_io_dat_o[14] ,
    \cb_1_8_io_dat_o[13] ,
    \cb_1_8_io_dat_o[12] ,
    \cb_1_8_io_dat_o[11] ,
    \cb_1_8_io_dat_o[10] ,
    \cb_1_8_io_dat_o[9] ,
    \cb_1_8_io_dat_o[8] ,
    \cb_1_8_io_dat_o[7] ,
    \cb_1_8_io_dat_o[6] ,
    \cb_1_8_io_dat_o[5] ,
    \cb_1_8_io_dat_o[4] ,
    \cb_1_8_io_dat_o[3] ,
    \cb_1_8_io_dat_o[2] ,
    \cb_1_8_io_dat_o[1] ,
    \cb_1_8_io_dat_o[0] }),
    .io_b_dat_o_9({\cb_1_9_io_dat_o[15] ,
    \cb_1_9_io_dat_o[14] ,
    \cb_1_9_io_dat_o[13] ,
    \cb_1_9_io_dat_o[12] ,
    \cb_1_9_io_dat_o[11] ,
    \cb_1_9_io_dat_o[10] ,
    \cb_1_9_io_dat_o[9] ,
    \cb_1_9_io_dat_o[8] ,
    \cb_1_9_io_dat_o[7] ,
    \cb_1_9_io_dat_o[6] ,
    \cb_1_9_io_dat_o[5] ,
    \cb_1_9_io_dat_o[4] ,
    \cb_1_9_io_dat_o[3] ,
    \cb_1_9_io_dat_o[2] ,
    \cb_1_9_io_dat_o[1] ,
    \cb_1_9_io_dat_o[0] }),
    .io_dat_i({\ccon_0_io_dat_i[31] ,
    \ccon_0_io_dat_i[30] ,
    \ccon_0_io_dat_i[29] ,
    \ccon_0_io_dat_i[28] ,
    \ccon_0_io_dat_i[27] ,
    \ccon_0_io_dat_i[26] ,
    \ccon_0_io_dat_i[25] ,
    \ccon_0_io_dat_i[24] ,
    \ccon_0_io_dat_i[23] ,
    \ccon_0_io_dat_i[22] ,
    \ccon_0_io_dat_i[21] ,
    \ccon_0_io_dat_i[20] ,
    \ccon_0_io_dat_i[19] ,
    \ccon_0_io_dat_i[18] ,
    \ccon_0_io_dat_i[17] ,
    \ccon_0_io_dat_i[16] ,
    \ccon_0_io_dat_i[15] ,
    \ccon_0_io_dat_i[14] ,
    \ccon_0_io_dat_i[13] ,
    \ccon_0_io_dat_i[12] ,
    \ccon_0_io_dat_i[11] ,
    \ccon_0_io_dat_i[10] ,
    \ccon_0_io_dat_i[9] ,
    \ccon_0_io_dat_i[8] ,
    \ccon_0_io_dat_i[7] ,
    \ccon_0_io_dat_i[6] ,
    \ccon_0_io_dat_i[5] ,
    \ccon_0_io_dat_i[4] ,
    \ccon_0_io_dat_i[3] ,
    \ccon_0_io_dat_i[2] ,
    \ccon_0_io_dat_i[1] ,
    \ccon_0_io_dat_i[0] }),
    .io_dat_o({\ccon_1_io_dat_o[31] ,
    \ccon_1_io_dat_o[30] ,
    \ccon_1_io_dat_o[29] ,
    \ccon_1_io_dat_o[28] ,
    \ccon_1_io_dat_o[27] ,
    \ccon_1_io_dat_o[26] ,
    \ccon_1_io_dat_o[25] ,
    \ccon_1_io_dat_o[24] ,
    \ccon_1_io_dat_o[23] ,
    \ccon_1_io_dat_o[22] ,
    \ccon_1_io_dat_o[21] ,
    \ccon_1_io_dat_o[20] ,
    \ccon_1_io_dat_o[19] ,
    \ccon_1_io_dat_o[18] ,
    \ccon_1_io_dat_o[17] ,
    \ccon_1_io_dat_o[16] ,
    \ccon_1_io_dat_o[15] ,
    \ccon_1_io_dat_o[14] ,
    \ccon_1_io_dat_o[13] ,
    \ccon_1_io_dat_o[12] ,
    \ccon_1_io_dat_o[11] ,
    \ccon_1_io_dat_o[10] ,
    \ccon_1_io_dat_o[9] ,
    \ccon_1_io_dat_o[8] ,
    \ccon_1_io_dat_o[7] ,
    \ccon_1_io_dat_o[6] ,
    \ccon_1_io_dat_o[5] ,
    \ccon_1_io_dat_o[4] ,
    \ccon_1_io_dat_o[3] ,
    \ccon_1_io_dat_o[2] ,
    \ccon_1_io_dat_o[1] ,
    \ccon_1_io_dat_o[0] }),
    .io_dataLastBlock({\cb_1_0_io_wo[63] ,
    \cb_1_0_io_wo[62] ,
    \cb_1_0_io_wo[61] ,
    \cb_1_0_io_wo[60] ,
    \cb_1_0_io_wo[59] ,
    \cb_1_0_io_wo[58] ,
    \cb_1_0_io_wo[57] ,
    \cb_1_0_io_wo[56] ,
    \cb_1_0_io_wo[55] ,
    \cb_1_0_io_wo[54] ,
    \cb_1_0_io_wo[53] ,
    \cb_1_0_io_wo[52] ,
    \cb_1_0_io_wo[51] ,
    \cb_1_0_io_wo[50] ,
    \cb_1_0_io_wo[49] ,
    \cb_1_0_io_wo[48] ,
    \cb_1_0_io_wo[47] ,
    \cb_1_0_io_wo[46] ,
    \cb_1_0_io_wo[45] ,
    \cb_1_0_io_wo[44] ,
    \cb_1_0_io_wo[43] ,
    \cb_1_0_io_wo[42] ,
    \cb_1_0_io_wo[41] ,
    \cb_1_0_io_wo[40] ,
    \cb_1_0_io_wo[39] ,
    \cb_1_0_io_wo[38] ,
    \cb_1_0_io_wo[37] ,
    \cb_1_0_io_wo[36] ,
    \cb_1_0_io_wo[35] ,
    \cb_1_0_io_wo[34] ,
    \cb_1_0_io_wo[33] ,
    \cb_1_0_io_wo[32] ,
    \cb_1_0_io_wo[31] ,
    \cb_1_0_io_wo[30] ,
    \cb_1_0_io_wo[29] ,
    \cb_1_0_io_wo[28] ,
    \cb_1_0_io_wo[27] ,
    \cb_1_0_io_wo[26] ,
    \cb_1_0_io_wo[25] ,
    \cb_1_0_io_wo[24] ,
    \cb_1_0_io_wo[23] ,
    \cb_1_0_io_wo[22] ,
    \cb_1_0_io_wo[21] ,
    \cb_1_0_io_wo[20] ,
    \cb_1_0_io_wo[19] ,
    \cb_1_0_io_wo[18] ,
    \cb_1_0_io_wo[17] ,
    \cb_1_0_io_wo[16] ,
    \cb_1_0_io_wo[15] ,
    \cb_1_0_io_wo[14] ,
    \cb_1_0_io_wo[13] ,
    \cb_1_0_io_wo[12] ,
    \cb_1_0_io_wo[11] ,
    \cb_1_0_io_wo[10] ,
    \cb_1_0_io_wo[9] ,
    \cb_1_0_io_wo[8] ,
    \cb_1_0_io_wo[7] ,
    \cb_1_0_io_wo[6] ,
    \cb_1_0_io_wo[5] ,
    \cb_1_0_io_wo[4] ,
    \cb_1_0_io_wo[3] ,
    \cb_1_0_io_wo[2] ,
    \cb_1_0_io_wo[1] ,
    \cb_1_0_io_wo[0] }),
    .io_dsi_in({\ccon_0_io_dsi_in[7] ,
    \ccon_0_io_dsi_in[6] ,
    \ccon_0_io_dsi_in[5] ,
    \ccon_0_io_dsi_in[4] ,
    \ccon_0_io_dsi_in[3] ,
    \ccon_0_io_dsi_in[2] ,
    \ccon_0_io_dsi_in[1] ,
    \ccon_0_io_dsi_in[0] }),
    .io_vout({cb_1_10_io_vi,
    cb_1_9_io_vi,
    cb_1_8_io_vi,
    cb_1_7_io_vi,
    cb_1_6_io_vi,
    cb_1_5_io_vi,
    cb_1_4_io_vi,
    cb_1_3_io_vi,
    cb_1_2_io_vi,
    cb_1_1_io_vi,
    cb_1_0_io_vi}));
 cic_con ccon_2 (.io_ack_o(\_T_172[0] ),
    .io_b_cs_i_0(cb_2_0_io_cs_i),
    .io_b_cs_i_1(cb_2_1_io_cs_i),
    .io_b_cs_i_10(cb_2_10_io_cs_i),
    .io_b_cs_i_2(cb_2_2_io_cs_i),
    .io_b_cs_i_3(cb_2_3_io_cs_i),
    .io_b_cs_i_4(cb_2_4_io_cs_i),
    .io_b_cs_i_5(cb_2_5_io_cs_i),
    .io_b_cs_i_6(cb_2_6_io_cs_i),
    .io_b_cs_i_7(cb_2_7_io_cs_i),
    .io_b_cs_i_8(cb_2_8_io_cs_i),
    .io_b_cs_i_9(cb_2_9_io_cs_i),
    .io_b_we_i(cb_2_0_io_we_i),
    .io_cs_i(ccon_2_io_cs_i),
    .io_dsi_o(cb_2_0_io_i_0_ci),
    .io_irq(\_T_183[0] ),
    .io_we_i(ccon_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\ccon_0_io_adr_i[11] ,
    \ccon_0_io_adr_i[10] ,
    \ccon_0_io_adr_i[9] ,
    \ccon_0_io_adr_i[8] ,
    \ccon_0_io_adr_i[7] ,
    \ccon_0_io_adr_i[6] ,
    \ccon_0_io_adr_i[5] ,
    \ccon_0_io_adr_i[4] ,
    \ccon_0_io_adr_i[3] ,
    \ccon_0_io_adr_i[2] ,
    \ccon_0_io_adr_i[1] ,
    \ccon_0_io_adr_i[0] }),
    .io_b_adr_i({\cb_2_0_io_adr_i[1] ,
    \cb_2_0_io_adr_i[0] }),
    .io_b_dat_i({\cb_2_0_io_dat_i[15] ,
    \cb_2_0_io_dat_i[14] ,
    \cb_2_0_io_dat_i[13] ,
    \cb_2_0_io_dat_i[12] ,
    \cb_2_0_io_dat_i[11] ,
    \cb_2_0_io_dat_i[10] ,
    \cb_2_0_io_dat_i[9] ,
    \cb_2_0_io_dat_i[8] ,
    \cb_2_0_io_dat_i[7] ,
    \cb_2_0_io_dat_i[6] ,
    \cb_2_0_io_dat_i[5] ,
    \cb_2_0_io_dat_i[4] ,
    \cb_2_0_io_dat_i[3] ,
    \cb_2_0_io_dat_i[2] ,
    \cb_2_0_io_dat_i[1] ,
    \cb_2_0_io_dat_i[0] }),
    .io_b_dat_o_0({\cb_2_0_io_dat_o[15] ,
    \cb_2_0_io_dat_o[14] ,
    \cb_2_0_io_dat_o[13] ,
    \cb_2_0_io_dat_o[12] ,
    \cb_2_0_io_dat_o[11] ,
    \cb_2_0_io_dat_o[10] ,
    \cb_2_0_io_dat_o[9] ,
    \cb_2_0_io_dat_o[8] ,
    \cb_2_0_io_dat_o[7] ,
    \cb_2_0_io_dat_o[6] ,
    \cb_2_0_io_dat_o[5] ,
    \cb_2_0_io_dat_o[4] ,
    \cb_2_0_io_dat_o[3] ,
    \cb_2_0_io_dat_o[2] ,
    \cb_2_0_io_dat_o[1] ,
    \cb_2_0_io_dat_o[0] }),
    .io_b_dat_o_1({\cb_2_1_io_dat_o[15] ,
    \cb_2_1_io_dat_o[14] ,
    \cb_2_1_io_dat_o[13] ,
    \cb_2_1_io_dat_o[12] ,
    \cb_2_1_io_dat_o[11] ,
    \cb_2_1_io_dat_o[10] ,
    \cb_2_1_io_dat_o[9] ,
    \cb_2_1_io_dat_o[8] ,
    \cb_2_1_io_dat_o[7] ,
    \cb_2_1_io_dat_o[6] ,
    \cb_2_1_io_dat_o[5] ,
    \cb_2_1_io_dat_o[4] ,
    \cb_2_1_io_dat_o[3] ,
    \cb_2_1_io_dat_o[2] ,
    \cb_2_1_io_dat_o[1] ,
    \cb_2_1_io_dat_o[0] }),
    .io_b_dat_o_10({\cb_2_10_io_dat_o[15] ,
    \cb_2_10_io_dat_o[14] ,
    \cb_2_10_io_dat_o[13] ,
    \cb_2_10_io_dat_o[12] ,
    \cb_2_10_io_dat_o[11] ,
    \cb_2_10_io_dat_o[10] ,
    \cb_2_10_io_dat_o[9] ,
    \cb_2_10_io_dat_o[8] ,
    \cb_2_10_io_dat_o[7] ,
    \cb_2_10_io_dat_o[6] ,
    \cb_2_10_io_dat_o[5] ,
    \cb_2_10_io_dat_o[4] ,
    \cb_2_10_io_dat_o[3] ,
    \cb_2_10_io_dat_o[2] ,
    \cb_2_10_io_dat_o[1] ,
    \cb_2_10_io_dat_o[0] }),
    .io_b_dat_o_2({\cb_2_2_io_dat_o[15] ,
    \cb_2_2_io_dat_o[14] ,
    \cb_2_2_io_dat_o[13] ,
    \cb_2_2_io_dat_o[12] ,
    \cb_2_2_io_dat_o[11] ,
    \cb_2_2_io_dat_o[10] ,
    \cb_2_2_io_dat_o[9] ,
    \cb_2_2_io_dat_o[8] ,
    \cb_2_2_io_dat_o[7] ,
    \cb_2_2_io_dat_o[6] ,
    \cb_2_2_io_dat_o[5] ,
    \cb_2_2_io_dat_o[4] ,
    \cb_2_2_io_dat_o[3] ,
    \cb_2_2_io_dat_o[2] ,
    \cb_2_2_io_dat_o[1] ,
    \cb_2_2_io_dat_o[0] }),
    .io_b_dat_o_3({\cb_2_3_io_dat_o[15] ,
    \cb_2_3_io_dat_o[14] ,
    \cb_2_3_io_dat_o[13] ,
    \cb_2_3_io_dat_o[12] ,
    \cb_2_3_io_dat_o[11] ,
    \cb_2_3_io_dat_o[10] ,
    \cb_2_3_io_dat_o[9] ,
    \cb_2_3_io_dat_o[8] ,
    \cb_2_3_io_dat_o[7] ,
    \cb_2_3_io_dat_o[6] ,
    \cb_2_3_io_dat_o[5] ,
    \cb_2_3_io_dat_o[4] ,
    \cb_2_3_io_dat_o[3] ,
    \cb_2_3_io_dat_o[2] ,
    \cb_2_3_io_dat_o[1] ,
    \cb_2_3_io_dat_o[0] }),
    .io_b_dat_o_4({\cb_2_4_io_dat_o[15] ,
    \cb_2_4_io_dat_o[14] ,
    \cb_2_4_io_dat_o[13] ,
    \cb_2_4_io_dat_o[12] ,
    \cb_2_4_io_dat_o[11] ,
    \cb_2_4_io_dat_o[10] ,
    \cb_2_4_io_dat_o[9] ,
    \cb_2_4_io_dat_o[8] ,
    \cb_2_4_io_dat_o[7] ,
    \cb_2_4_io_dat_o[6] ,
    \cb_2_4_io_dat_o[5] ,
    \cb_2_4_io_dat_o[4] ,
    \cb_2_4_io_dat_o[3] ,
    \cb_2_4_io_dat_o[2] ,
    \cb_2_4_io_dat_o[1] ,
    \cb_2_4_io_dat_o[0] }),
    .io_b_dat_o_5({\cb_2_5_io_dat_o[15] ,
    \cb_2_5_io_dat_o[14] ,
    \cb_2_5_io_dat_o[13] ,
    \cb_2_5_io_dat_o[12] ,
    \cb_2_5_io_dat_o[11] ,
    \cb_2_5_io_dat_o[10] ,
    \cb_2_5_io_dat_o[9] ,
    \cb_2_5_io_dat_o[8] ,
    \cb_2_5_io_dat_o[7] ,
    \cb_2_5_io_dat_o[6] ,
    \cb_2_5_io_dat_o[5] ,
    \cb_2_5_io_dat_o[4] ,
    \cb_2_5_io_dat_o[3] ,
    \cb_2_5_io_dat_o[2] ,
    \cb_2_5_io_dat_o[1] ,
    \cb_2_5_io_dat_o[0] }),
    .io_b_dat_o_6({\cb_2_6_io_dat_o[15] ,
    \cb_2_6_io_dat_o[14] ,
    \cb_2_6_io_dat_o[13] ,
    \cb_2_6_io_dat_o[12] ,
    \cb_2_6_io_dat_o[11] ,
    \cb_2_6_io_dat_o[10] ,
    \cb_2_6_io_dat_o[9] ,
    \cb_2_6_io_dat_o[8] ,
    \cb_2_6_io_dat_o[7] ,
    \cb_2_6_io_dat_o[6] ,
    \cb_2_6_io_dat_o[5] ,
    \cb_2_6_io_dat_o[4] ,
    \cb_2_6_io_dat_o[3] ,
    \cb_2_6_io_dat_o[2] ,
    \cb_2_6_io_dat_o[1] ,
    \cb_2_6_io_dat_o[0] }),
    .io_b_dat_o_7({\cb_2_7_io_dat_o[15] ,
    \cb_2_7_io_dat_o[14] ,
    \cb_2_7_io_dat_o[13] ,
    \cb_2_7_io_dat_o[12] ,
    \cb_2_7_io_dat_o[11] ,
    \cb_2_7_io_dat_o[10] ,
    \cb_2_7_io_dat_o[9] ,
    \cb_2_7_io_dat_o[8] ,
    \cb_2_7_io_dat_o[7] ,
    \cb_2_7_io_dat_o[6] ,
    \cb_2_7_io_dat_o[5] ,
    \cb_2_7_io_dat_o[4] ,
    \cb_2_7_io_dat_o[3] ,
    \cb_2_7_io_dat_o[2] ,
    \cb_2_7_io_dat_o[1] ,
    \cb_2_7_io_dat_o[0] }),
    .io_b_dat_o_8({\cb_2_8_io_dat_o[15] ,
    \cb_2_8_io_dat_o[14] ,
    \cb_2_8_io_dat_o[13] ,
    \cb_2_8_io_dat_o[12] ,
    \cb_2_8_io_dat_o[11] ,
    \cb_2_8_io_dat_o[10] ,
    \cb_2_8_io_dat_o[9] ,
    \cb_2_8_io_dat_o[8] ,
    \cb_2_8_io_dat_o[7] ,
    \cb_2_8_io_dat_o[6] ,
    \cb_2_8_io_dat_o[5] ,
    \cb_2_8_io_dat_o[4] ,
    \cb_2_8_io_dat_o[3] ,
    \cb_2_8_io_dat_o[2] ,
    \cb_2_8_io_dat_o[1] ,
    \cb_2_8_io_dat_o[0] }),
    .io_b_dat_o_9({\cb_2_9_io_dat_o[15] ,
    \cb_2_9_io_dat_o[14] ,
    \cb_2_9_io_dat_o[13] ,
    \cb_2_9_io_dat_o[12] ,
    \cb_2_9_io_dat_o[11] ,
    \cb_2_9_io_dat_o[10] ,
    \cb_2_9_io_dat_o[9] ,
    \cb_2_9_io_dat_o[8] ,
    \cb_2_9_io_dat_o[7] ,
    \cb_2_9_io_dat_o[6] ,
    \cb_2_9_io_dat_o[5] ,
    \cb_2_9_io_dat_o[4] ,
    \cb_2_9_io_dat_o[3] ,
    \cb_2_9_io_dat_o[2] ,
    \cb_2_9_io_dat_o[1] ,
    \cb_2_9_io_dat_o[0] }),
    .io_dat_i({\ccon_0_io_dat_i[31] ,
    \ccon_0_io_dat_i[30] ,
    \ccon_0_io_dat_i[29] ,
    \ccon_0_io_dat_i[28] ,
    \ccon_0_io_dat_i[27] ,
    \ccon_0_io_dat_i[26] ,
    \ccon_0_io_dat_i[25] ,
    \ccon_0_io_dat_i[24] ,
    \ccon_0_io_dat_i[23] ,
    \ccon_0_io_dat_i[22] ,
    \ccon_0_io_dat_i[21] ,
    \ccon_0_io_dat_i[20] ,
    \ccon_0_io_dat_i[19] ,
    \ccon_0_io_dat_i[18] ,
    \ccon_0_io_dat_i[17] ,
    \ccon_0_io_dat_i[16] ,
    \ccon_0_io_dat_i[15] ,
    \ccon_0_io_dat_i[14] ,
    \ccon_0_io_dat_i[13] ,
    \ccon_0_io_dat_i[12] ,
    \ccon_0_io_dat_i[11] ,
    \ccon_0_io_dat_i[10] ,
    \ccon_0_io_dat_i[9] ,
    \ccon_0_io_dat_i[8] ,
    \ccon_0_io_dat_i[7] ,
    \ccon_0_io_dat_i[6] ,
    \ccon_0_io_dat_i[5] ,
    \ccon_0_io_dat_i[4] ,
    \ccon_0_io_dat_i[3] ,
    \ccon_0_io_dat_i[2] ,
    \ccon_0_io_dat_i[1] ,
    \ccon_0_io_dat_i[0] }),
    .io_dat_o({\ccon_2_io_dat_o[31] ,
    \ccon_2_io_dat_o[30] ,
    \ccon_2_io_dat_o[29] ,
    \ccon_2_io_dat_o[28] ,
    \ccon_2_io_dat_o[27] ,
    \ccon_2_io_dat_o[26] ,
    \ccon_2_io_dat_o[25] ,
    \ccon_2_io_dat_o[24] ,
    \ccon_2_io_dat_o[23] ,
    \ccon_2_io_dat_o[22] ,
    \ccon_2_io_dat_o[21] ,
    \ccon_2_io_dat_o[20] ,
    \ccon_2_io_dat_o[19] ,
    \ccon_2_io_dat_o[18] ,
    \ccon_2_io_dat_o[17] ,
    \ccon_2_io_dat_o[16] ,
    \ccon_2_io_dat_o[15] ,
    \ccon_2_io_dat_o[14] ,
    \ccon_2_io_dat_o[13] ,
    \ccon_2_io_dat_o[12] ,
    \ccon_2_io_dat_o[11] ,
    \ccon_2_io_dat_o[10] ,
    \ccon_2_io_dat_o[9] ,
    \ccon_2_io_dat_o[8] ,
    \ccon_2_io_dat_o[7] ,
    \ccon_2_io_dat_o[6] ,
    \ccon_2_io_dat_o[5] ,
    \ccon_2_io_dat_o[4] ,
    \ccon_2_io_dat_o[3] ,
    \ccon_2_io_dat_o[2] ,
    \ccon_2_io_dat_o[1] ,
    \ccon_2_io_dat_o[0] }),
    .io_dataLastBlock({\cb_2_0_io_wo[63] ,
    \cb_2_0_io_wo[62] ,
    \cb_2_0_io_wo[61] ,
    \cb_2_0_io_wo[60] ,
    \cb_2_0_io_wo[59] ,
    \cb_2_0_io_wo[58] ,
    \cb_2_0_io_wo[57] ,
    \cb_2_0_io_wo[56] ,
    \cb_2_0_io_wo[55] ,
    \cb_2_0_io_wo[54] ,
    \cb_2_0_io_wo[53] ,
    \cb_2_0_io_wo[52] ,
    \cb_2_0_io_wo[51] ,
    \cb_2_0_io_wo[50] ,
    \cb_2_0_io_wo[49] ,
    \cb_2_0_io_wo[48] ,
    \cb_2_0_io_wo[47] ,
    \cb_2_0_io_wo[46] ,
    \cb_2_0_io_wo[45] ,
    \cb_2_0_io_wo[44] ,
    \cb_2_0_io_wo[43] ,
    \cb_2_0_io_wo[42] ,
    \cb_2_0_io_wo[41] ,
    \cb_2_0_io_wo[40] ,
    \cb_2_0_io_wo[39] ,
    \cb_2_0_io_wo[38] ,
    \cb_2_0_io_wo[37] ,
    \cb_2_0_io_wo[36] ,
    \cb_2_0_io_wo[35] ,
    \cb_2_0_io_wo[34] ,
    \cb_2_0_io_wo[33] ,
    \cb_2_0_io_wo[32] ,
    \cb_2_0_io_wo[31] ,
    \cb_2_0_io_wo[30] ,
    \cb_2_0_io_wo[29] ,
    \cb_2_0_io_wo[28] ,
    \cb_2_0_io_wo[27] ,
    \cb_2_0_io_wo[26] ,
    \cb_2_0_io_wo[25] ,
    \cb_2_0_io_wo[24] ,
    \cb_2_0_io_wo[23] ,
    \cb_2_0_io_wo[22] ,
    \cb_2_0_io_wo[21] ,
    \cb_2_0_io_wo[20] ,
    \cb_2_0_io_wo[19] ,
    \cb_2_0_io_wo[18] ,
    \cb_2_0_io_wo[17] ,
    \cb_2_0_io_wo[16] ,
    \cb_2_0_io_wo[15] ,
    \cb_2_0_io_wo[14] ,
    \cb_2_0_io_wo[13] ,
    \cb_2_0_io_wo[12] ,
    \cb_2_0_io_wo[11] ,
    \cb_2_0_io_wo[10] ,
    \cb_2_0_io_wo[9] ,
    \cb_2_0_io_wo[8] ,
    \cb_2_0_io_wo[7] ,
    \cb_2_0_io_wo[6] ,
    \cb_2_0_io_wo[5] ,
    \cb_2_0_io_wo[4] ,
    \cb_2_0_io_wo[3] ,
    \cb_2_0_io_wo[2] ,
    \cb_2_0_io_wo[1] ,
    \cb_2_0_io_wo[0] }),
    .io_dsi_in({\ccon_0_io_dsi_in[7] ,
    \ccon_0_io_dsi_in[6] ,
    \ccon_0_io_dsi_in[5] ,
    \ccon_0_io_dsi_in[4] ,
    \ccon_0_io_dsi_in[3] ,
    \ccon_0_io_dsi_in[2] ,
    \ccon_0_io_dsi_in[1] ,
    \ccon_0_io_dsi_in[0] }),
    .io_vout({cb_2_10_io_vi,
    cb_2_9_io_vi,
    cb_2_8_io_vi,
    cb_2_7_io_vi,
    cb_2_6_io_vi,
    cb_2_5_io_vi,
    cb_2_4_io_vi,
    cb_2_3_io_vi,
    cb_2_2_io_vi,
    cb_2_1_io_vi,
    cb_2_0_io_vi}));
 cic_con ccon_3 (.io_ack_o(\_T_172[1] ),
    .io_b_cs_i_0(cb_3_0_io_cs_i),
    .io_b_cs_i_1(cb_3_1_io_cs_i),
    .io_b_cs_i_10(cb_3_10_io_cs_i),
    .io_b_cs_i_2(cb_3_2_io_cs_i),
    .io_b_cs_i_3(cb_3_3_io_cs_i),
    .io_b_cs_i_4(cb_3_4_io_cs_i),
    .io_b_cs_i_5(cb_3_5_io_cs_i),
    .io_b_cs_i_6(cb_3_6_io_cs_i),
    .io_b_cs_i_7(cb_3_7_io_cs_i),
    .io_b_cs_i_8(cb_3_8_io_cs_i),
    .io_b_cs_i_9(cb_3_9_io_cs_i),
    .io_b_we_i(cb_3_0_io_we_i),
    .io_cs_i(ccon_3_io_cs_i),
    .io_dsi_o(cb_3_0_io_i_0_ci),
    .io_irq(\_T_183[1] ),
    .io_we_i(ccon_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\ccon_0_io_adr_i[11] ,
    \ccon_0_io_adr_i[10] ,
    \ccon_0_io_adr_i[9] ,
    \ccon_0_io_adr_i[8] ,
    \ccon_0_io_adr_i[7] ,
    \ccon_0_io_adr_i[6] ,
    \ccon_0_io_adr_i[5] ,
    \ccon_0_io_adr_i[4] ,
    \ccon_0_io_adr_i[3] ,
    \ccon_0_io_adr_i[2] ,
    \ccon_0_io_adr_i[1] ,
    \ccon_0_io_adr_i[0] }),
    .io_b_adr_i({\cb_3_0_io_adr_i[1] ,
    \cb_3_0_io_adr_i[0] }),
    .io_b_dat_i({\cb_3_0_io_dat_i[15] ,
    \cb_3_0_io_dat_i[14] ,
    \cb_3_0_io_dat_i[13] ,
    \cb_3_0_io_dat_i[12] ,
    \cb_3_0_io_dat_i[11] ,
    \cb_3_0_io_dat_i[10] ,
    \cb_3_0_io_dat_i[9] ,
    \cb_3_0_io_dat_i[8] ,
    \cb_3_0_io_dat_i[7] ,
    \cb_3_0_io_dat_i[6] ,
    \cb_3_0_io_dat_i[5] ,
    \cb_3_0_io_dat_i[4] ,
    \cb_3_0_io_dat_i[3] ,
    \cb_3_0_io_dat_i[2] ,
    \cb_3_0_io_dat_i[1] ,
    \cb_3_0_io_dat_i[0] }),
    .io_b_dat_o_0({\cb_3_0_io_dat_o[15] ,
    \cb_3_0_io_dat_o[14] ,
    \cb_3_0_io_dat_o[13] ,
    \cb_3_0_io_dat_o[12] ,
    \cb_3_0_io_dat_o[11] ,
    \cb_3_0_io_dat_o[10] ,
    \cb_3_0_io_dat_o[9] ,
    \cb_3_0_io_dat_o[8] ,
    \cb_3_0_io_dat_o[7] ,
    \cb_3_0_io_dat_o[6] ,
    \cb_3_0_io_dat_o[5] ,
    \cb_3_0_io_dat_o[4] ,
    \cb_3_0_io_dat_o[3] ,
    \cb_3_0_io_dat_o[2] ,
    \cb_3_0_io_dat_o[1] ,
    \cb_3_0_io_dat_o[0] }),
    .io_b_dat_o_1({\cb_3_1_io_dat_o[15] ,
    \cb_3_1_io_dat_o[14] ,
    \cb_3_1_io_dat_o[13] ,
    \cb_3_1_io_dat_o[12] ,
    \cb_3_1_io_dat_o[11] ,
    \cb_3_1_io_dat_o[10] ,
    \cb_3_1_io_dat_o[9] ,
    \cb_3_1_io_dat_o[8] ,
    \cb_3_1_io_dat_o[7] ,
    \cb_3_1_io_dat_o[6] ,
    \cb_3_1_io_dat_o[5] ,
    \cb_3_1_io_dat_o[4] ,
    \cb_3_1_io_dat_o[3] ,
    \cb_3_1_io_dat_o[2] ,
    \cb_3_1_io_dat_o[1] ,
    \cb_3_1_io_dat_o[0] }),
    .io_b_dat_o_10({\cb_3_10_io_dat_o[15] ,
    \cb_3_10_io_dat_o[14] ,
    \cb_3_10_io_dat_o[13] ,
    \cb_3_10_io_dat_o[12] ,
    \cb_3_10_io_dat_o[11] ,
    \cb_3_10_io_dat_o[10] ,
    \cb_3_10_io_dat_o[9] ,
    \cb_3_10_io_dat_o[8] ,
    \cb_3_10_io_dat_o[7] ,
    \cb_3_10_io_dat_o[6] ,
    \cb_3_10_io_dat_o[5] ,
    \cb_3_10_io_dat_o[4] ,
    \cb_3_10_io_dat_o[3] ,
    \cb_3_10_io_dat_o[2] ,
    \cb_3_10_io_dat_o[1] ,
    \cb_3_10_io_dat_o[0] }),
    .io_b_dat_o_2({\cb_3_2_io_dat_o[15] ,
    \cb_3_2_io_dat_o[14] ,
    \cb_3_2_io_dat_o[13] ,
    \cb_3_2_io_dat_o[12] ,
    \cb_3_2_io_dat_o[11] ,
    \cb_3_2_io_dat_o[10] ,
    \cb_3_2_io_dat_o[9] ,
    \cb_3_2_io_dat_o[8] ,
    \cb_3_2_io_dat_o[7] ,
    \cb_3_2_io_dat_o[6] ,
    \cb_3_2_io_dat_o[5] ,
    \cb_3_2_io_dat_o[4] ,
    \cb_3_2_io_dat_o[3] ,
    \cb_3_2_io_dat_o[2] ,
    \cb_3_2_io_dat_o[1] ,
    \cb_3_2_io_dat_o[0] }),
    .io_b_dat_o_3({\cb_3_3_io_dat_o[15] ,
    \cb_3_3_io_dat_o[14] ,
    \cb_3_3_io_dat_o[13] ,
    \cb_3_3_io_dat_o[12] ,
    \cb_3_3_io_dat_o[11] ,
    \cb_3_3_io_dat_o[10] ,
    \cb_3_3_io_dat_o[9] ,
    \cb_3_3_io_dat_o[8] ,
    \cb_3_3_io_dat_o[7] ,
    \cb_3_3_io_dat_o[6] ,
    \cb_3_3_io_dat_o[5] ,
    \cb_3_3_io_dat_o[4] ,
    \cb_3_3_io_dat_o[3] ,
    \cb_3_3_io_dat_o[2] ,
    \cb_3_3_io_dat_o[1] ,
    \cb_3_3_io_dat_o[0] }),
    .io_b_dat_o_4({\cb_3_4_io_dat_o[15] ,
    \cb_3_4_io_dat_o[14] ,
    \cb_3_4_io_dat_o[13] ,
    \cb_3_4_io_dat_o[12] ,
    \cb_3_4_io_dat_o[11] ,
    \cb_3_4_io_dat_o[10] ,
    \cb_3_4_io_dat_o[9] ,
    \cb_3_4_io_dat_o[8] ,
    \cb_3_4_io_dat_o[7] ,
    \cb_3_4_io_dat_o[6] ,
    \cb_3_4_io_dat_o[5] ,
    \cb_3_4_io_dat_o[4] ,
    \cb_3_4_io_dat_o[3] ,
    \cb_3_4_io_dat_o[2] ,
    \cb_3_4_io_dat_o[1] ,
    \cb_3_4_io_dat_o[0] }),
    .io_b_dat_o_5({\cb_3_5_io_dat_o[15] ,
    \cb_3_5_io_dat_o[14] ,
    \cb_3_5_io_dat_o[13] ,
    \cb_3_5_io_dat_o[12] ,
    \cb_3_5_io_dat_o[11] ,
    \cb_3_5_io_dat_o[10] ,
    \cb_3_5_io_dat_o[9] ,
    \cb_3_5_io_dat_o[8] ,
    \cb_3_5_io_dat_o[7] ,
    \cb_3_5_io_dat_o[6] ,
    \cb_3_5_io_dat_o[5] ,
    \cb_3_5_io_dat_o[4] ,
    \cb_3_5_io_dat_o[3] ,
    \cb_3_5_io_dat_o[2] ,
    \cb_3_5_io_dat_o[1] ,
    \cb_3_5_io_dat_o[0] }),
    .io_b_dat_o_6({\cb_3_6_io_dat_o[15] ,
    \cb_3_6_io_dat_o[14] ,
    \cb_3_6_io_dat_o[13] ,
    \cb_3_6_io_dat_o[12] ,
    \cb_3_6_io_dat_o[11] ,
    \cb_3_6_io_dat_o[10] ,
    \cb_3_6_io_dat_o[9] ,
    \cb_3_6_io_dat_o[8] ,
    \cb_3_6_io_dat_o[7] ,
    \cb_3_6_io_dat_o[6] ,
    \cb_3_6_io_dat_o[5] ,
    \cb_3_6_io_dat_o[4] ,
    \cb_3_6_io_dat_o[3] ,
    \cb_3_6_io_dat_o[2] ,
    \cb_3_6_io_dat_o[1] ,
    \cb_3_6_io_dat_o[0] }),
    .io_b_dat_o_7({\cb_3_7_io_dat_o[15] ,
    \cb_3_7_io_dat_o[14] ,
    \cb_3_7_io_dat_o[13] ,
    \cb_3_7_io_dat_o[12] ,
    \cb_3_7_io_dat_o[11] ,
    \cb_3_7_io_dat_o[10] ,
    \cb_3_7_io_dat_o[9] ,
    \cb_3_7_io_dat_o[8] ,
    \cb_3_7_io_dat_o[7] ,
    \cb_3_7_io_dat_o[6] ,
    \cb_3_7_io_dat_o[5] ,
    \cb_3_7_io_dat_o[4] ,
    \cb_3_7_io_dat_o[3] ,
    \cb_3_7_io_dat_o[2] ,
    \cb_3_7_io_dat_o[1] ,
    \cb_3_7_io_dat_o[0] }),
    .io_b_dat_o_8({\cb_3_8_io_dat_o[15] ,
    \cb_3_8_io_dat_o[14] ,
    \cb_3_8_io_dat_o[13] ,
    \cb_3_8_io_dat_o[12] ,
    \cb_3_8_io_dat_o[11] ,
    \cb_3_8_io_dat_o[10] ,
    \cb_3_8_io_dat_o[9] ,
    \cb_3_8_io_dat_o[8] ,
    \cb_3_8_io_dat_o[7] ,
    \cb_3_8_io_dat_o[6] ,
    \cb_3_8_io_dat_o[5] ,
    \cb_3_8_io_dat_o[4] ,
    \cb_3_8_io_dat_o[3] ,
    \cb_3_8_io_dat_o[2] ,
    \cb_3_8_io_dat_o[1] ,
    \cb_3_8_io_dat_o[0] }),
    .io_b_dat_o_9({\cb_3_9_io_dat_o[15] ,
    \cb_3_9_io_dat_o[14] ,
    \cb_3_9_io_dat_o[13] ,
    \cb_3_9_io_dat_o[12] ,
    \cb_3_9_io_dat_o[11] ,
    \cb_3_9_io_dat_o[10] ,
    \cb_3_9_io_dat_o[9] ,
    \cb_3_9_io_dat_o[8] ,
    \cb_3_9_io_dat_o[7] ,
    \cb_3_9_io_dat_o[6] ,
    \cb_3_9_io_dat_o[5] ,
    \cb_3_9_io_dat_o[4] ,
    \cb_3_9_io_dat_o[3] ,
    \cb_3_9_io_dat_o[2] ,
    \cb_3_9_io_dat_o[1] ,
    \cb_3_9_io_dat_o[0] }),
    .io_dat_i({\ccon_0_io_dat_i[31] ,
    \ccon_0_io_dat_i[30] ,
    \ccon_0_io_dat_i[29] ,
    \ccon_0_io_dat_i[28] ,
    \ccon_0_io_dat_i[27] ,
    \ccon_0_io_dat_i[26] ,
    \ccon_0_io_dat_i[25] ,
    \ccon_0_io_dat_i[24] ,
    \ccon_0_io_dat_i[23] ,
    \ccon_0_io_dat_i[22] ,
    \ccon_0_io_dat_i[21] ,
    \ccon_0_io_dat_i[20] ,
    \ccon_0_io_dat_i[19] ,
    \ccon_0_io_dat_i[18] ,
    \ccon_0_io_dat_i[17] ,
    \ccon_0_io_dat_i[16] ,
    \ccon_0_io_dat_i[15] ,
    \ccon_0_io_dat_i[14] ,
    \ccon_0_io_dat_i[13] ,
    \ccon_0_io_dat_i[12] ,
    \ccon_0_io_dat_i[11] ,
    \ccon_0_io_dat_i[10] ,
    \ccon_0_io_dat_i[9] ,
    \ccon_0_io_dat_i[8] ,
    \ccon_0_io_dat_i[7] ,
    \ccon_0_io_dat_i[6] ,
    \ccon_0_io_dat_i[5] ,
    \ccon_0_io_dat_i[4] ,
    \ccon_0_io_dat_i[3] ,
    \ccon_0_io_dat_i[2] ,
    \ccon_0_io_dat_i[1] ,
    \ccon_0_io_dat_i[0] }),
    .io_dat_o({\ccon_3_io_dat_o[31] ,
    \ccon_3_io_dat_o[30] ,
    \ccon_3_io_dat_o[29] ,
    \ccon_3_io_dat_o[28] ,
    \ccon_3_io_dat_o[27] ,
    \ccon_3_io_dat_o[26] ,
    \ccon_3_io_dat_o[25] ,
    \ccon_3_io_dat_o[24] ,
    \ccon_3_io_dat_o[23] ,
    \ccon_3_io_dat_o[22] ,
    \ccon_3_io_dat_o[21] ,
    \ccon_3_io_dat_o[20] ,
    \ccon_3_io_dat_o[19] ,
    \ccon_3_io_dat_o[18] ,
    \ccon_3_io_dat_o[17] ,
    \ccon_3_io_dat_o[16] ,
    \ccon_3_io_dat_o[15] ,
    \ccon_3_io_dat_o[14] ,
    \ccon_3_io_dat_o[13] ,
    \ccon_3_io_dat_o[12] ,
    \ccon_3_io_dat_o[11] ,
    \ccon_3_io_dat_o[10] ,
    \ccon_3_io_dat_o[9] ,
    \ccon_3_io_dat_o[8] ,
    \ccon_3_io_dat_o[7] ,
    \ccon_3_io_dat_o[6] ,
    \ccon_3_io_dat_o[5] ,
    \ccon_3_io_dat_o[4] ,
    \ccon_3_io_dat_o[3] ,
    \ccon_3_io_dat_o[2] ,
    \ccon_3_io_dat_o[1] ,
    \ccon_3_io_dat_o[0] }),
    .io_dataLastBlock({\cb_3_0_io_wo[63] ,
    \cb_3_0_io_wo[62] ,
    \cb_3_0_io_wo[61] ,
    \cb_3_0_io_wo[60] ,
    \cb_3_0_io_wo[59] ,
    \cb_3_0_io_wo[58] ,
    \cb_3_0_io_wo[57] ,
    \cb_3_0_io_wo[56] ,
    \cb_3_0_io_wo[55] ,
    \cb_3_0_io_wo[54] ,
    \cb_3_0_io_wo[53] ,
    \cb_3_0_io_wo[52] ,
    \cb_3_0_io_wo[51] ,
    \cb_3_0_io_wo[50] ,
    \cb_3_0_io_wo[49] ,
    \cb_3_0_io_wo[48] ,
    \cb_3_0_io_wo[47] ,
    \cb_3_0_io_wo[46] ,
    \cb_3_0_io_wo[45] ,
    \cb_3_0_io_wo[44] ,
    \cb_3_0_io_wo[43] ,
    \cb_3_0_io_wo[42] ,
    \cb_3_0_io_wo[41] ,
    \cb_3_0_io_wo[40] ,
    \cb_3_0_io_wo[39] ,
    \cb_3_0_io_wo[38] ,
    \cb_3_0_io_wo[37] ,
    \cb_3_0_io_wo[36] ,
    \cb_3_0_io_wo[35] ,
    \cb_3_0_io_wo[34] ,
    \cb_3_0_io_wo[33] ,
    \cb_3_0_io_wo[32] ,
    \cb_3_0_io_wo[31] ,
    \cb_3_0_io_wo[30] ,
    \cb_3_0_io_wo[29] ,
    \cb_3_0_io_wo[28] ,
    \cb_3_0_io_wo[27] ,
    \cb_3_0_io_wo[26] ,
    \cb_3_0_io_wo[25] ,
    \cb_3_0_io_wo[24] ,
    \cb_3_0_io_wo[23] ,
    \cb_3_0_io_wo[22] ,
    \cb_3_0_io_wo[21] ,
    \cb_3_0_io_wo[20] ,
    \cb_3_0_io_wo[19] ,
    \cb_3_0_io_wo[18] ,
    \cb_3_0_io_wo[17] ,
    \cb_3_0_io_wo[16] ,
    \cb_3_0_io_wo[15] ,
    \cb_3_0_io_wo[14] ,
    \cb_3_0_io_wo[13] ,
    \cb_3_0_io_wo[12] ,
    \cb_3_0_io_wo[11] ,
    \cb_3_0_io_wo[10] ,
    \cb_3_0_io_wo[9] ,
    \cb_3_0_io_wo[8] ,
    \cb_3_0_io_wo[7] ,
    \cb_3_0_io_wo[6] ,
    \cb_3_0_io_wo[5] ,
    \cb_3_0_io_wo[4] ,
    \cb_3_0_io_wo[3] ,
    \cb_3_0_io_wo[2] ,
    \cb_3_0_io_wo[1] ,
    \cb_3_0_io_wo[0] }),
    .io_dsi_in({\ccon_0_io_dsi_in[7] ,
    \ccon_0_io_dsi_in[6] ,
    \ccon_0_io_dsi_in[5] ,
    \ccon_0_io_dsi_in[4] ,
    \ccon_0_io_dsi_in[3] ,
    \ccon_0_io_dsi_in[2] ,
    \ccon_0_io_dsi_in[1] ,
    \ccon_0_io_dsi_in[0] }),
    .io_vout({cb_3_10_io_vi,
    cb_3_9_io_vi,
    cb_3_8_io_vi,
    cb_3_7_io_vi,
    cb_3_6_io_vi,
    cb_3_5_io_vi,
    cb_3_4_io_vi,
    cb_3_3_io_vi,
    cb_3_2_io_vi,
    cb_3_1_io_vi,
    cb_3_0_io_vi}));
 cic_con ccon_4 (.io_ack_o(\_T_172[2] ),
    .io_b_cs_i_0(cb_4_0_io_cs_i),
    .io_b_cs_i_1(cb_4_1_io_cs_i),
    .io_b_cs_i_10(cb_4_10_io_cs_i),
    .io_b_cs_i_2(cb_4_2_io_cs_i),
    .io_b_cs_i_3(cb_4_3_io_cs_i),
    .io_b_cs_i_4(cb_4_4_io_cs_i),
    .io_b_cs_i_5(cb_4_5_io_cs_i),
    .io_b_cs_i_6(cb_4_6_io_cs_i),
    .io_b_cs_i_7(cb_4_7_io_cs_i),
    .io_b_cs_i_8(cb_4_8_io_cs_i),
    .io_b_cs_i_9(cb_4_9_io_cs_i),
    .io_b_we_i(cb_4_0_io_we_i),
    .io_cs_i(ccon_4_io_cs_i),
    .io_dsi_o(cb_4_0_io_i_0_ci),
    .io_irq(\_T_183[2] ),
    .io_we_i(ccon_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\ccon_0_io_adr_i[11] ,
    \ccon_0_io_adr_i[10] ,
    \ccon_0_io_adr_i[9] ,
    \ccon_0_io_adr_i[8] ,
    \ccon_0_io_adr_i[7] ,
    \ccon_0_io_adr_i[6] ,
    \ccon_0_io_adr_i[5] ,
    \ccon_0_io_adr_i[4] ,
    \ccon_0_io_adr_i[3] ,
    \ccon_0_io_adr_i[2] ,
    \ccon_0_io_adr_i[1] ,
    \ccon_0_io_adr_i[0] }),
    .io_b_adr_i({\cb_4_0_io_adr_i[1] ,
    \cb_4_0_io_adr_i[0] }),
    .io_b_dat_i({\cb_4_0_io_dat_i[15] ,
    \cb_4_0_io_dat_i[14] ,
    \cb_4_0_io_dat_i[13] ,
    \cb_4_0_io_dat_i[12] ,
    \cb_4_0_io_dat_i[11] ,
    \cb_4_0_io_dat_i[10] ,
    \cb_4_0_io_dat_i[9] ,
    \cb_4_0_io_dat_i[8] ,
    \cb_4_0_io_dat_i[7] ,
    \cb_4_0_io_dat_i[6] ,
    \cb_4_0_io_dat_i[5] ,
    \cb_4_0_io_dat_i[4] ,
    \cb_4_0_io_dat_i[3] ,
    \cb_4_0_io_dat_i[2] ,
    \cb_4_0_io_dat_i[1] ,
    \cb_4_0_io_dat_i[0] }),
    .io_b_dat_o_0({\cb_4_0_io_dat_o[15] ,
    \cb_4_0_io_dat_o[14] ,
    \cb_4_0_io_dat_o[13] ,
    \cb_4_0_io_dat_o[12] ,
    \cb_4_0_io_dat_o[11] ,
    \cb_4_0_io_dat_o[10] ,
    \cb_4_0_io_dat_o[9] ,
    \cb_4_0_io_dat_o[8] ,
    \cb_4_0_io_dat_o[7] ,
    \cb_4_0_io_dat_o[6] ,
    \cb_4_0_io_dat_o[5] ,
    \cb_4_0_io_dat_o[4] ,
    \cb_4_0_io_dat_o[3] ,
    \cb_4_0_io_dat_o[2] ,
    \cb_4_0_io_dat_o[1] ,
    \cb_4_0_io_dat_o[0] }),
    .io_b_dat_o_1({\cb_4_1_io_dat_o[15] ,
    \cb_4_1_io_dat_o[14] ,
    \cb_4_1_io_dat_o[13] ,
    \cb_4_1_io_dat_o[12] ,
    \cb_4_1_io_dat_o[11] ,
    \cb_4_1_io_dat_o[10] ,
    \cb_4_1_io_dat_o[9] ,
    \cb_4_1_io_dat_o[8] ,
    \cb_4_1_io_dat_o[7] ,
    \cb_4_1_io_dat_o[6] ,
    \cb_4_1_io_dat_o[5] ,
    \cb_4_1_io_dat_o[4] ,
    \cb_4_1_io_dat_o[3] ,
    \cb_4_1_io_dat_o[2] ,
    \cb_4_1_io_dat_o[1] ,
    \cb_4_1_io_dat_o[0] }),
    .io_b_dat_o_10({\cb_4_10_io_dat_o[15] ,
    \cb_4_10_io_dat_o[14] ,
    \cb_4_10_io_dat_o[13] ,
    \cb_4_10_io_dat_o[12] ,
    \cb_4_10_io_dat_o[11] ,
    \cb_4_10_io_dat_o[10] ,
    \cb_4_10_io_dat_o[9] ,
    \cb_4_10_io_dat_o[8] ,
    \cb_4_10_io_dat_o[7] ,
    \cb_4_10_io_dat_o[6] ,
    \cb_4_10_io_dat_o[5] ,
    \cb_4_10_io_dat_o[4] ,
    \cb_4_10_io_dat_o[3] ,
    \cb_4_10_io_dat_o[2] ,
    \cb_4_10_io_dat_o[1] ,
    \cb_4_10_io_dat_o[0] }),
    .io_b_dat_o_2({\cb_4_2_io_dat_o[15] ,
    \cb_4_2_io_dat_o[14] ,
    \cb_4_2_io_dat_o[13] ,
    \cb_4_2_io_dat_o[12] ,
    \cb_4_2_io_dat_o[11] ,
    \cb_4_2_io_dat_o[10] ,
    \cb_4_2_io_dat_o[9] ,
    \cb_4_2_io_dat_o[8] ,
    \cb_4_2_io_dat_o[7] ,
    \cb_4_2_io_dat_o[6] ,
    \cb_4_2_io_dat_o[5] ,
    \cb_4_2_io_dat_o[4] ,
    \cb_4_2_io_dat_o[3] ,
    \cb_4_2_io_dat_o[2] ,
    \cb_4_2_io_dat_o[1] ,
    \cb_4_2_io_dat_o[0] }),
    .io_b_dat_o_3({\cb_4_3_io_dat_o[15] ,
    \cb_4_3_io_dat_o[14] ,
    \cb_4_3_io_dat_o[13] ,
    \cb_4_3_io_dat_o[12] ,
    \cb_4_3_io_dat_o[11] ,
    \cb_4_3_io_dat_o[10] ,
    \cb_4_3_io_dat_o[9] ,
    \cb_4_3_io_dat_o[8] ,
    \cb_4_3_io_dat_o[7] ,
    \cb_4_3_io_dat_o[6] ,
    \cb_4_3_io_dat_o[5] ,
    \cb_4_3_io_dat_o[4] ,
    \cb_4_3_io_dat_o[3] ,
    \cb_4_3_io_dat_o[2] ,
    \cb_4_3_io_dat_o[1] ,
    \cb_4_3_io_dat_o[0] }),
    .io_b_dat_o_4({\cb_4_4_io_dat_o[15] ,
    \cb_4_4_io_dat_o[14] ,
    \cb_4_4_io_dat_o[13] ,
    \cb_4_4_io_dat_o[12] ,
    \cb_4_4_io_dat_o[11] ,
    \cb_4_4_io_dat_o[10] ,
    \cb_4_4_io_dat_o[9] ,
    \cb_4_4_io_dat_o[8] ,
    \cb_4_4_io_dat_o[7] ,
    \cb_4_4_io_dat_o[6] ,
    \cb_4_4_io_dat_o[5] ,
    \cb_4_4_io_dat_o[4] ,
    \cb_4_4_io_dat_o[3] ,
    \cb_4_4_io_dat_o[2] ,
    \cb_4_4_io_dat_o[1] ,
    \cb_4_4_io_dat_o[0] }),
    .io_b_dat_o_5({\cb_4_5_io_dat_o[15] ,
    \cb_4_5_io_dat_o[14] ,
    \cb_4_5_io_dat_o[13] ,
    \cb_4_5_io_dat_o[12] ,
    \cb_4_5_io_dat_o[11] ,
    \cb_4_5_io_dat_o[10] ,
    \cb_4_5_io_dat_o[9] ,
    \cb_4_5_io_dat_o[8] ,
    \cb_4_5_io_dat_o[7] ,
    \cb_4_5_io_dat_o[6] ,
    \cb_4_5_io_dat_o[5] ,
    \cb_4_5_io_dat_o[4] ,
    \cb_4_5_io_dat_o[3] ,
    \cb_4_5_io_dat_o[2] ,
    \cb_4_5_io_dat_o[1] ,
    \cb_4_5_io_dat_o[0] }),
    .io_b_dat_o_6({\cb_4_6_io_dat_o[15] ,
    \cb_4_6_io_dat_o[14] ,
    \cb_4_6_io_dat_o[13] ,
    \cb_4_6_io_dat_o[12] ,
    \cb_4_6_io_dat_o[11] ,
    \cb_4_6_io_dat_o[10] ,
    \cb_4_6_io_dat_o[9] ,
    \cb_4_6_io_dat_o[8] ,
    \cb_4_6_io_dat_o[7] ,
    \cb_4_6_io_dat_o[6] ,
    \cb_4_6_io_dat_o[5] ,
    \cb_4_6_io_dat_o[4] ,
    \cb_4_6_io_dat_o[3] ,
    \cb_4_6_io_dat_o[2] ,
    \cb_4_6_io_dat_o[1] ,
    \cb_4_6_io_dat_o[0] }),
    .io_b_dat_o_7({\cb_4_7_io_dat_o[15] ,
    \cb_4_7_io_dat_o[14] ,
    \cb_4_7_io_dat_o[13] ,
    \cb_4_7_io_dat_o[12] ,
    \cb_4_7_io_dat_o[11] ,
    \cb_4_7_io_dat_o[10] ,
    \cb_4_7_io_dat_o[9] ,
    \cb_4_7_io_dat_o[8] ,
    \cb_4_7_io_dat_o[7] ,
    \cb_4_7_io_dat_o[6] ,
    \cb_4_7_io_dat_o[5] ,
    \cb_4_7_io_dat_o[4] ,
    \cb_4_7_io_dat_o[3] ,
    \cb_4_7_io_dat_o[2] ,
    \cb_4_7_io_dat_o[1] ,
    \cb_4_7_io_dat_o[0] }),
    .io_b_dat_o_8({\cb_4_8_io_dat_o[15] ,
    \cb_4_8_io_dat_o[14] ,
    \cb_4_8_io_dat_o[13] ,
    \cb_4_8_io_dat_o[12] ,
    \cb_4_8_io_dat_o[11] ,
    \cb_4_8_io_dat_o[10] ,
    \cb_4_8_io_dat_o[9] ,
    \cb_4_8_io_dat_o[8] ,
    \cb_4_8_io_dat_o[7] ,
    \cb_4_8_io_dat_o[6] ,
    \cb_4_8_io_dat_o[5] ,
    \cb_4_8_io_dat_o[4] ,
    \cb_4_8_io_dat_o[3] ,
    \cb_4_8_io_dat_o[2] ,
    \cb_4_8_io_dat_o[1] ,
    \cb_4_8_io_dat_o[0] }),
    .io_b_dat_o_9({\cb_4_9_io_dat_o[15] ,
    \cb_4_9_io_dat_o[14] ,
    \cb_4_9_io_dat_o[13] ,
    \cb_4_9_io_dat_o[12] ,
    \cb_4_9_io_dat_o[11] ,
    \cb_4_9_io_dat_o[10] ,
    \cb_4_9_io_dat_o[9] ,
    \cb_4_9_io_dat_o[8] ,
    \cb_4_9_io_dat_o[7] ,
    \cb_4_9_io_dat_o[6] ,
    \cb_4_9_io_dat_o[5] ,
    \cb_4_9_io_dat_o[4] ,
    \cb_4_9_io_dat_o[3] ,
    \cb_4_9_io_dat_o[2] ,
    \cb_4_9_io_dat_o[1] ,
    \cb_4_9_io_dat_o[0] }),
    .io_dat_i({\ccon_0_io_dat_i[31] ,
    \ccon_0_io_dat_i[30] ,
    \ccon_0_io_dat_i[29] ,
    \ccon_0_io_dat_i[28] ,
    \ccon_0_io_dat_i[27] ,
    \ccon_0_io_dat_i[26] ,
    \ccon_0_io_dat_i[25] ,
    \ccon_0_io_dat_i[24] ,
    \ccon_0_io_dat_i[23] ,
    \ccon_0_io_dat_i[22] ,
    \ccon_0_io_dat_i[21] ,
    \ccon_0_io_dat_i[20] ,
    \ccon_0_io_dat_i[19] ,
    \ccon_0_io_dat_i[18] ,
    \ccon_0_io_dat_i[17] ,
    \ccon_0_io_dat_i[16] ,
    \ccon_0_io_dat_i[15] ,
    \ccon_0_io_dat_i[14] ,
    \ccon_0_io_dat_i[13] ,
    \ccon_0_io_dat_i[12] ,
    \ccon_0_io_dat_i[11] ,
    \ccon_0_io_dat_i[10] ,
    \ccon_0_io_dat_i[9] ,
    \ccon_0_io_dat_i[8] ,
    \ccon_0_io_dat_i[7] ,
    \ccon_0_io_dat_i[6] ,
    \ccon_0_io_dat_i[5] ,
    \ccon_0_io_dat_i[4] ,
    \ccon_0_io_dat_i[3] ,
    \ccon_0_io_dat_i[2] ,
    \ccon_0_io_dat_i[1] ,
    \ccon_0_io_dat_i[0] }),
    .io_dat_o({\ccon_4_io_dat_o[31] ,
    \ccon_4_io_dat_o[30] ,
    \ccon_4_io_dat_o[29] ,
    \ccon_4_io_dat_o[28] ,
    \ccon_4_io_dat_o[27] ,
    \ccon_4_io_dat_o[26] ,
    \ccon_4_io_dat_o[25] ,
    \ccon_4_io_dat_o[24] ,
    \ccon_4_io_dat_o[23] ,
    \ccon_4_io_dat_o[22] ,
    \ccon_4_io_dat_o[21] ,
    \ccon_4_io_dat_o[20] ,
    \ccon_4_io_dat_o[19] ,
    \ccon_4_io_dat_o[18] ,
    \ccon_4_io_dat_o[17] ,
    \ccon_4_io_dat_o[16] ,
    \ccon_4_io_dat_o[15] ,
    \ccon_4_io_dat_o[14] ,
    \ccon_4_io_dat_o[13] ,
    \ccon_4_io_dat_o[12] ,
    \ccon_4_io_dat_o[11] ,
    \ccon_4_io_dat_o[10] ,
    \ccon_4_io_dat_o[9] ,
    \ccon_4_io_dat_o[8] ,
    \ccon_4_io_dat_o[7] ,
    \ccon_4_io_dat_o[6] ,
    \ccon_4_io_dat_o[5] ,
    \ccon_4_io_dat_o[4] ,
    \ccon_4_io_dat_o[3] ,
    \ccon_4_io_dat_o[2] ,
    \ccon_4_io_dat_o[1] ,
    \ccon_4_io_dat_o[0] }),
    .io_dataLastBlock({\cb_4_0_io_wo[63] ,
    \cb_4_0_io_wo[62] ,
    \cb_4_0_io_wo[61] ,
    \cb_4_0_io_wo[60] ,
    \cb_4_0_io_wo[59] ,
    \cb_4_0_io_wo[58] ,
    \cb_4_0_io_wo[57] ,
    \cb_4_0_io_wo[56] ,
    \cb_4_0_io_wo[55] ,
    \cb_4_0_io_wo[54] ,
    \cb_4_0_io_wo[53] ,
    \cb_4_0_io_wo[52] ,
    \cb_4_0_io_wo[51] ,
    \cb_4_0_io_wo[50] ,
    \cb_4_0_io_wo[49] ,
    \cb_4_0_io_wo[48] ,
    \cb_4_0_io_wo[47] ,
    \cb_4_0_io_wo[46] ,
    \cb_4_0_io_wo[45] ,
    \cb_4_0_io_wo[44] ,
    \cb_4_0_io_wo[43] ,
    \cb_4_0_io_wo[42] ,
    \cb_4_0_io_wo[41] ,
    \cb_4_0_io_wo[40] ,
    \cb_4_0_io_wo[39] ,
    \cb_4_0_io_wo[38] ,
    \cb_4_0_io_wo[37] ,
    \cb_4_0_io_wo[36] ,
    \cb_4_0_io_wo[35] ,
    \cb_4_0_io_wo[34] ,
    \cb_4_0_io_wo[33] ,
    \cb_4_0_io_wo[32] ,
    \cb_4_0_io_wo[31] ,
    \cb_4_0_io_wo[30] ,
    \cb_4_0_io_wo[29] ,
    \cb_4_0_io_wo[28] ,
    \cb_4_0_io_wo[27] ,
    \cb_4_0_io_wo[26] ,
    \cb_4_0_io_wo[25] ,
    \cb_4_0_io_wo[24] ,
    \cb_4_0_io_wo[23] ,
    \cb_4_0_io_wo[22] ,
    \cb_4_0_io_wo[21] ,
    \cb_4_0_io_wo[20] ,
    \cb_4_0_io_wo[19] ,
    \cb_4_0_io_wo[18] ,
    \cb_4_0_io_wo[17] ,
    \cb_4_0_io_wo[16] ,
    \cb_4_0_io_wo[15] ,
    \cb_4_0_io_wo[14] ,
    \cb_4_0_io_wo[13] ,
    \cb_4_0_io_wo[12] ,
    \cb_4_0_io_wo[11] ,
    \cb_4_0_io_wo[10] ,
    \cb_4_0_io_wo[9] ,
    \cb_4_0_io_wo[8] ,
    \cb_4_0_io_wo[7] ,
    \cb_4_0_io_wo[6] ,
    \cb_4_0_io_wo[5] ,
    \cb_4_0_io_wo[4] ,
    \cb_4_0_io_wo[3] ,
    \cb_4_0_io_wo[2] ,
    \cb_4_0_io_wo[1] ,
    \cb_4_0_io_wo[0] }),
    .io_dsi_in({\ccon_0_io_dsi_in[7] ,
    \ccon_0_io_dsi_in[6] ,
    \ccon_0_io_dsi_in[5] ,
    \ccon_0_io_dsi_in[4] ,
    \ccon_0_io_dsi_in[3] ,
    \ccon_0_io_dsi_in[2] ,
    \ccon_0_io_dsi_in[1] ,
    \ccon_0_io_dsi_in[0] }),
    .io_vout({cb_4_10_io_vi,
    cb_4_9_io_vi,
    cb_4_8_io_vi,
    cb_4_7_io_vi,
    cb_4_6_io_vi,
    cb_4_5_io_vi,
    cb_4_4_io_vi,
    cb_4_3_io_vi,
    cb_4_2_io_vi,
    cb_4_1_io_vi,
    cb_4_0_io_vi}));
 cic_con ccon_5 (.io_ack_o(\_T_172[3] ),
    .io_b_cs_i_0(cb_5_0_io_cs_i),
    .io_b_cs_i_1(cb_5_1_io_cs_i),
    .io_b_cs_i_10(cb_5_10_io_cs_i),
    .io_b_cs_i_2(cb_5_2_io_cs_i),
    .io_b_cs_i_3(cb_5_3_io_cs_i),
    .io_b_cs_i_4(cb_5_4_io_cs_i),
    .io_b_cs_i_5(cb_5_5_io_cs_i),
    .io_b_cs_i_6(cb_5_6_io_cs_i),
    .io_b_cs_i_7(cb_5_7_io_cs_i),
    .io_b_cs_i_8(cb_5_8_io_cs_i),
    .io_b_cs_i_9(cb_5_9_io_cs_i),
    .io_b_we_i(cb_5_0_io_we_i),
    .io_cs_i(ccon_5_io_cs_i),
    .io_dsi_o(cb_5_0_io_i_0_ci),
    .io_irq(\_T_183[3] ),
    .io_we_i(ccon_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\ccon_0_io_adr_i[11] ,
    \ccon_0_io_adr_i[10] ,
    \ccon_0_io_adr_i[9] ,
    \ccon_0_io_adr_i[8] ,
    \ccon_0_io_adr_i[7] ,
    \ccon_0_io_adr_i[6] ,
    \ccon_0_io_adr_i[5] ,
    \ccon_0_io_adr_i[4] ,
    \ccon_0_io_adr_i[3] ,
    \ccon_0_io_adr_i[2] ,
    \ccon_0_io_adr_i[1] ,
    \ccon_0_io_adr_i[0] }),
    .io_b_adr_i({\cb_5_0_io_adr_i[1] ,
    \cb_5_0_io_adr_i[0] }),
    .io_b_dat_i({\cb_5_0_io_dat_i[15] ,
    \cb_5_0_io_dat_i[14] ,
    \cb_5_0_io_dat_i[13] ,
    \cb_5_0_io_dat_i[12] ,
    \cb_5_0_io_dat_i[11] ,
    \cb_5_0_io_dat_i[10] ,
    \cb_5_0_io_dat_i[9] ,
    \cb_5_0_io_dat_i[8] ,
    \cb_5_0_io_dat_i[7] ,
    \cb_5_0_io_dat_i[6] ,
    \cb_5_0_io_dat_i[5] ,
    \cb_5_0_io_dat_i[4] ,
    \cb_5_0_io_dat_i[3] ,
    \cb_5_0_io_dat_i[2] ,
    \cb_5_0_io_dat_i[1] ,
    \cb_5_0_io_dat_i[0] }),
    .io_b_dat_o_0({\cb_5_0_io_dat_o[15] ,
    \cb_5_0_io_dat_o[14] ,
    \cb_5_0_io_dat_o[13] ,
    \cb_5_0_io_dat_o[12] ,
    \cb_5_0_io_dat_o[11] ,
    \cb_5_0_io_dat_o[10] ,
    \cb_5_0_io_dat_o[9] ,
    \cb_5_0_io_dat_o[8] ,
    \cb_5_0_io_dat_o[7] ,
    \cb_5_0_io_dat_o[6] ,
    \cb_5_0_io_dat_o[5] ,
    \cb_5_0_io_dat_o[4] ,
    \cb_5_0_io_dat_o[3] ,
    \cb_5_0_io_dat_o[2] ,
    \cb_5_0_io_dat_o[1] ,
    \cb_5_0_io_dat_o[0] }),
    .io_b_dat_o_1({\cb_5_1_io_dat_o[15] ,
    \cb_5_1_io_dat_o[14] ,
    \cb_5_1_io_dat_o[13] ,
    \cb_5_1_io_dat_o[12] ,
    \cb_5_1_io_dat_o[11] ,
    \cb_5_1_io_dat_o[10] ,
    \cb_5_1_io_dat_o[9] ,
    \cb_5_1_io_dat_o[8] ,
    \cb_5_1_io_dat_o[7] ,
    \cb_5_1_io_dat_o[6] ,
    \cb_5_1_io_dat_o[5] ,
    \cb_5_1_io_dat_o[4] ,
    \cb_5_1_io_dat_o[3] ,
    \cb_5_1_io_dat_o[2] ,
    \cb_5_1_io_dat_o[1] ,
    \cb_5_1_io_dat_o[0] }),
    .io_b_dat_o_10({\cb_5_10_io_dat_o[15] ,
    \cb_5_10_io_dat_o[14] ,
    \cb_5_10_io_dat_o[13] ,
    \cb_5_10_io_dat_o[12] ,
    \cb_5_10_io_dat_o[11] ,
    \cb_5_10_io_dat_o[10] ,
    \cb_5_10_io_dat_o[9] ,
    \cb_5_10_io_dat_o[8] ,
    \cb_5_10_io_dat_o[7] ,
    \cb_5_10_io_dat_o[6] ,
    \cb_5_10_io_dat_o[5] ,
    \cb_5_10_io_dat_o[4] ,
    \cb_5_10_io_dat_o[3] ,
    \cb_5_10_io_dat_o[2] ,
    \cb_5_10_io_dat_o[1] ,
    \cb_5_10_io_dat_o[0] }),
    .io_b_dat_o_2({\cb_5_2_io_dat_o[15] ,
    \cb_5_2_io_dat_o[14] ,
    \cb_5_2_io_dat_o[13] ,
    \cb_5_2_io_dat_o[12] ,
    \cb_5_2_io_dat_o[11] ,
    \cb_5_2_io_dat_o[10] ,
    \cb_5_2_io_dat_o[9] ,
    \cb_5_2_io_dat_o[8] ,
    \cb_5_2_io_dat_o[7] ,
    \cb_5_2_io_dat_o[6] ,
    \cb_5_2_io_dat_o[5] ,
    \cb_5_2_io_dat_o[4] ,
    \cb_5_2_io_dat_o[3] ,
    \cb_5_2_io_dat_o[2] ,
    \cb_5_2_io_dat_o[1] ,
    \cb_5_2_io_dat_o[0] }),
    .io_b_dat_o_3({\cb_5_3_io_dat_o[15] ,
    \cb_5_3_io_dat_o[14] ,
    \cb_5_3_io_dat_o[13] ,
    \cb_5_3_io_dat_o[12] ,
    \cb_5_3_io_dat_o[11] ,
    \cb_5_3_io_dat_o[10] ,
    \cb_5_3_io_dat_o[9] ,
    \cb_5_3_io_dat_o[8] ,
    \cb_5_3_io_dat_o[7] ,
    \cb_5_3_io_dat_o[6] ,
    \cb_5_3_io_dat_o[5] ,
    \cb_5_3_io_dat_o[4] ,
    \cb_5_3_io_dat_o[3] ,
    \cb_5_3_io_dat_o[2] ,
    \cb_5_3_io_dat_o[1] ,
    \cb_5_3_io_dat_o[0] }),
    .io_b_dat_o_4({\cb_5_4_io_dat_o[15] ,
    \cb_5_4_io_dat_o[14] ,
    \cb_5_4_io_dat_o[13] ,
    \cb_5_4_io_dat_o[12] ,
    \cb_5_4_io_dat_o[11] ,
    \cb_5_4_io_dat_o[10] ,
    \cb_5_4_io_dat_o[9] ,
    \cb_5_4_io_dat_o[8] ,
    \cb_5_4_io_dat_o[7] ,
    \cb_5_4_io_dat_o[6] ,
    \cb_5_4_io_dat_o[5] ,
    \cb_5_4_io_dat_o[4] ,
    \cb_5_4_io_dat_o[3] ,
    \cb_5_4_io_dat_o[2] ,
    \cb_5_4_io_dat_o[1] ,
    \cb_5_4_io_dat_o[0] }),
    .io_b_dat_o_5({\cb_5_5_io_dat_o[15] ,
    \cb_5_5_io_dat_o[14] ,
    \cb_5_5_io_dat_o[13] ,
    \cb_5_5_io_dat_o[12] ,
    \cb_5_5_io_dat_o[11] ,
    \cb_5_5_io_dat_o[10] ,
    \cb_5_5_io_dat_o[9] ,
    \cb_5_5_io_dat_o[8] ,
    \cb_5_5_io_dat_o[7] ,
    \cb_5_5_io_dat_o[6] ,
    \cb_5_5_io_dat_o[5] ,
    \cb_5_5_io_dat_o[4] ,
    \cb_5_5_io_dat_o[3] ,
    \cb_5_5_io_dat_o[2] ,
    \cb_5_5_io_dat_o[1] ,
    \cb_5_5_io_dat_o[0] }),
    .io_b_dat_o_6({\cb_5_6_io_dat_o[15] ,
    \cb_5_6_io_dat_o[14] ,
    \cb_5_6_io_dat_o[13] ,
    \cb_5_6_io_dat_o[12] ,
    \cb_5_6_io_dat_o[11] ,
    \cb_5_6_io_dat_o[10] ,
    \cb_5_6_io_dat_o[9] ,
    \cb_5_6_io_dat_o[8] ,
    \cb_5_6_io_dat_o[7] ,
    \cb_5_6_io_dat_o[6] ,
    \cb_5_6_io_dat_o[5] ,
    \cb_5_6_io_dat_o[4] ,
    \cb_5_6_io_dat_o[3] ,
    \cb_5_6_io_dat_o[2] ,
    \cb_5_6_io_dat_o[1] ,
    \cb_5_6_io_dat_o[0] }),
    .io_b_dat_o_7({\cb_5_7_io_dat_o[15] ,
    \cb_5_7_io_dat_o[14] ,
    \cb_5_7_io_dat_o[13] ,
    \cb_5_7_io_dat_o[12] ,
    \cb_5_7_io_dat_o[11] ,
    \cb_5_7_io_dat_o[10] ,
    \cb_5_7_io_dat_o[9] ,
    \cb_5_7_io_dat_o[8] ,
    \cb_5_7_io_dat_o[7] ,
    \cb_5_7_io_dat_o[6] ,
    \cb_5_7_io_dat_o[5] ,
    \cb_5_7_io_dat_o[4] ,
    \cb_5_7_io_dat_o[3] ,
    \cb_5_7_io_dat_o[2] ,
    \cb_5_7_io_dat_o[1] ,
    \cb_5_7_io_dat_o[0] }),
    .io_b_dat_o_8({\cb_5_8_io_dat_o[15] ,
    \cb_5_8_io_dat_o[14] ,
    \cb_5_8_io_dat_o[13] ,
    \cb_5_8_io_dat_o[12] ,
    \cb_5_8_io_dat_o[11] ,
    \cb_5_8_io_dat_o[10] ,
    \cb_5_8_io_dat_o[9] ,
    \cb_5_8_io_dat_o[8] ,
    \cb_5_8_io_dat_o[7] ,
    \cb_5_8_io_dat_o[6] ,
    \cb_5_8_io_dat_o[5] ,
    \cb_5_8_io_dat_o[4] ,
    \cb_5_8_io_dat_o[3] ,
    \cb_5_8_io_dat_o[2] ,
    \cb_5_8_io_dat_o[1] ,
    \cb_5_8_io_dat_o[0] }),
    .io_b_dat_o_9({\cb_5_9_io_dat_o[15] ,
    \cb_5_9_io_dat_o[14] ,
    \cb_5_9_io_dat_o[13] ,
    \cb_5_9_io_dat_o[12] ,
    \cb_5_9_io_dat_o[11] ,
    \cb_5_9_io_dat_o[10] ,
    \cb_5_9_io_dat_o[9] ,
    \cb_5_9_io_dat_o[8] ,
    \cb_5_9_io_dat_o[7] ,
    \cb_5_9_io_dat_o[6] ,
    \cb_5_9_io_dat_o[5] ,
    \cb_5_9_io_dat_o[4] ,
    \cb_5_9_io_dat_o[3] ,
    \cb_5_9_io_dat_o[2] ,
    \cb_5_9_io_dat_o[1] ,
    \cb_5_9_io_dat_o[0] }),
    .io_dat_i({\ccon_0_io_dat_i[31] ,
    \ccon_0_io_dat_i[30] ,
    \ccon_0_io_dat_i[29] ,
    \ccon_0_io_dat_i[28] ,
    \ccon_0_io_dat_i[27] ,
    \ccon_0_io_dat_i[26] ,
    \ccon_0_io_dat_i[25] ,
    \ccon_0_io_dat_i[24] ,
    \ccon_0_io_dat_i[23] ,
    \ccon_0_io_dat_i[22] ,
    \ccon_0_io_dat_i[21] ,
    \ccon_0_io_dat_i[20] ,
    \ccon_0_io_dat_i[19] ,
    \ccon_0_io_dat_i[18] ,
    \ccon_0_io_dat_i[17] ,
    \ccon_0_io_dat_i[16] ,
    \ccon_0_io_dat_i[15] ,
    \ccon_0_io_dat_i[14] ,
    \ccon_0_io_dat_i[13] ,
    \ccon_0_io_dat_i[12] ,
    \ccon_0_io_dat_i[11] ,
    \ccon_0_io_dat_i[10] ,
    \ccon_0_io_dat_i[9] ,
    \ccon_0_io_dat_i[8] ,
    \ccon_0_io_dat_i[7] ,
    \ccon_0_io_dat_i[6] ,
    \ccon_0_io_dat_i[5] ,
    \ccon_0_io_dat_i[4] ,
    \ccon_0_io_dat_i[3] ,
    \ccon_0_io_dat_i[2] ,
    \ccon_0_io_dat_i[1] ,
    \ccon_0_io_dat_i[0] }),
    .io_dat_o({\ccon_5_io_dat_o[31] ,
    \ccon_5_io_dat_o[30] ,
    \ccon_5_io_dat_o[29] ,
    \ccon_5_io_dat_o[28] ,
    \ccon_5_io_dat_o[27] ,
    \ccon_5_io_dat_o[26] ,
    \ccon_5_io_dat_o[25] ,
    \ccon_5_io_dat_o[24] ,
    \ccon_5_io_dat_o[23] ,
    \ccon_5_io_dat_o[22] ,
    \ccon_5_io_dat_o[21] ,
    \ccon_5_io_dat_o[20] ,
    \ccon_5_io_dat_o[19] ,
    \ccon_5_io_dat_o[18] ,
    \ccon_5_io_dat_o[17] ,
    \ccon_5_io_dat_o[16] ,
    \ccon_5_io_dat_o[15] ,
    \ccon_5_io_dat_o[14] ,
    \ccon_5_io_dat_o[13] ,
    \ccon_5_io_dat_o[12] ,
    \ccon_5_io_dat_o[11] ,
    \ccon_5_io_dat_o[10] ,
    \ccon_5_io_dat_o[9] ,
    \ccon_5_io_dat_o[8] ,
    \ccon_5_io_dat_o[7] ,
    \ccon_5_io_dat_o[6] ,
    \ccon_5_io_dat_o[5] ,
    \ccon_5_io_dat_o[4] ,
    \ccon_5_io_dat_o[3] ,
    \ccon_5_io_dat_o[2] ,
    \ccon_5_io_dat_o[1] ,
    \ccon_5_io_dat_o[0] }),
    .io_dataLastBlock({\cb_5_0_io_wo[63] ,
    \cb_5_0_io_wo[62] ,
    \cb_5_0_io_wo[61] ,
    \cb_5_0_io_wo[60] ,
    \cb_5_0_io_wo[59] ,
    \cb_5_0_io_wo[58] ,
    \cb_5_0_io_wo[57] ,
    \cb_5_0_io_wo[56] ,
    \cb_5_0_io_wo[55] ,
    \cb_5_0_io_wo[54] ,
    \cb_5_0_io_wo[53] ,
    \cb_5_0_io_wo[52] ,
    \cb_5_0_io_wo[51] ,
    \cb_5_0_io_wo[50] ,
    \cb_5_0_io_wo[49] ,
    \cb_5_0_io_wo[48] ,
    \cb_5_0_io_wo[47] ,
    \cb_5_0_io_wo[46] ,
    \cb_5_0_io_wo[45] ,
    \cb_5_0_io_wo[44] ,
    \cb_5_0_io_wo[43] ,
    \cb_5_0_io_wo[42] ,
    \cb_5_0_io_wo[41] ,
    \cb_5_0_io_wo[40] ,
    \cb_5_0_io_wo[39] ,
    \cb_5_0_io_wo[38] ,
    \cb_5_0_io_wo[37] ,
    \cb_5_0_io_wo[36] ,
    \cb_5_0_io_wo[35] ,
    \cb_5_0_io_wo[34] ,
    \cb_5_0_io_wo[33] ,
    \cb_5_0_io_wo[32] ,
    \cb_5_0_io_wo[31] ,
    \cb_5_0_io_wo[30] ,
    \cb_5_0_io_wo[29] ,
    \cb_5_0_io_wo[28] ,
    \cb_5_0_io_wo[27] ,
    \cb_5_0_io_wo[26] ,
    \cb_5_0_io_wo[25] ,
    \cb_5_0_io_wo[24] ,
    \cb_5_0_io_wo[23] ,
    \cb_5_0_io_wo[22] ,
    \cb_5_0_io_wo[21] ,
    \cb_5_0_io_wo[20] ,
    \cb_5_0_io_wo[19] ,
    \cb_5_0_io_wo[18] ,
    \cb_5_0_io_wo[17] ,
    \cb_5_0_io_wo[16] ,
    \cb_5_0_io_wo[15] ,
    \cb_5_0_io_wo[14] ,
    \cb_5_0_io_wo[13] ,
    \cb_5_0_io_wo[12] ,
    \cb_5_0_io_wo[11] ,
    \cb_5_0_io_wo[10] ,
    \cb_5_0_io_wo[9] ,
    \cb_5_0_io_wo[8] ,
    \cb_5_0_io_wo[7] ,
    \cb_5_0_io_wo[6] ,
    \cb_5_0_io_wo[5] ,
    \cb_5_0_io_wo[4] ,
    \cb_5_0_io_wo[3] ,
    \cb_5_0_io_wo[2] ,
    \cb_5_0_io_wo[1] ,
    \cb_5_0_io_wo[0] }),
    .io_dsi_in({\ccon_0_io_dsi_in[7] ,
    \ccon_0_io_dsi_in[6] ,
    \ccon_0_io_dsi_in[5] ,
    \ccon_0_io_dsi_in[4] ,
    \ccon_0_io_dsi_in[3] ,
    \ccon_0_io_dsi_in[2] ,
    \ccon_0_io_dsi_in[1] ,
    \ccon_0_io_dsi_in[0] }),
    .io_vout({cb_5_10_io_vi,
    cb_5_9_io_vi,
    cb_5_8_io_vi,
    cb_5_7_io_vi,
    cb_5_6_io_vi,
    cb_5_5_io_vi,
    cb_5_4_io_vi,
    cb_5_3_io_vi,
    cb_5_2_io_vi,
    cb_5_1_io_vi,
    cb_5_0_io_vi}));
 cic_con ccon_6 (.io_ack_o(\_T_172[4] ),
    .io_b_cs_i_0(cb_6_0_io_cs_i),
    .io_b_cs_i_1(cb_6_1_io_cs_i),
    .io_b_cs_i_10(cb_6_10_io_cs_i),
    .io_b_cs_i_2(cb_6_2_io_cs_i),
    .io_b_cs_i_3(cb_6_3_io_cs_i),
    .io_b_cs_i_4(cb_6_4_io_cs_i),
    .io_b_cs_i_5(cb_6_5_io_cs_i),
    .io_b_cs_i_6(cb_6_6_io_cs_i),
    .io_b_cs_i_7(cb_6_7_io_cs_i),
    .io_b_cs_i_8(cb_6_8_io_cs_i),
    .io_b_cs_i_9(cb_6_9_io_cs_i),
    .io_b_we_i(cb_6_0_io_we_i),
    .io_cs_i(ccon_6_io_cs_i),
    .io_dsi_o(cb_6_0_io_i_0_ci),
    .io_irq(\_T_183[4] ),
    .io_we_i(ccon_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\ccon_0_io_adr_i[11] ,
    \ccon_0_io_adr_i[10] ,
    \ccon_0_io_adr_i[9] ,
    \ccon_0_io_adr_i[8] ,
    \ccon_0_io_adr_i[7] ,
    \ccon_0_io_adr_i[6] ,
    \ccon_0_io_adr_i[5] ,
    \ccon_0_io_adr_i[4] ,
    \ccon_0_io_adr_i[3] ,
    \ccon_0_io_adr_i[2] ,
    \ccon_0_io_adr_i[1] ,
    \ccon_0_io_adr_i[0] }),
    .io_b_adr_i({\cb_6_0_io_adr_i[1] ,
    \cb_6_0_io_adr_i[0] }),
    .io_b_dat_i({\cb_6_0_io_dat_i[15] ,
    \cb_6_0_io_dat_i[14] ,
    \cb_6_0_io_dat_i[13] ,
    \cb_6_0_io_dat_i[12] ,
    \cb_6_0_io_dat_i[11] ,
    \cb_6_0_io_dat_i[10] ,
    \cb_6_0_io_dat_i[9] ,
    \cb_6_0_io_dat_i[8] ,
    \cb_6_0_io_dat_i[7] ,
    \cb_6_0_io_dat_i[6] ,
    \cb_6_0_io_dat_i[5] ,
    \cb_6_0_io_dat_i[4] ,
    \cb_6_0_io_dat_i[3] ,
    \cb_6_0_io_dat_i[2] ,
    \cb_6_0_io_dat_i[1] ,
    \cb_6_0_io_dat_i[0] }),
    .io_b_dat_o_0({\cb_6_0_io_dat_o[15] ,
    \cb_6_0_io_dat_o[14] ,
    \cb_6_0_io_dat_o[13] ,
    \cb_6_0_io_dat_o[12] ,
    \cb_6_0_io_dat_o[11] ,
    \cb_6_0_io_dat_o[10] ,
    \cb_6_0_io_dat_o[9] ,
    \cb_6_0_io_dat_o[8] ,
    \cb_6_0_io_dat_o[7] ,
    \cb_6_0_io_dat_o[6] ,
    \cb_6_0_io_dat_o[5] ,
    \cb_6_0_io_dat_o[4] ,
    \cb_6_0_io_dat_o[3] ,
    \cb_6_0_io_dat_o[2] ,
    \cb_6_0_io_dat_o[1] ,
    \cb_6_0_io_dat_o[0] }),
    .io_b_dat_o_1({\cb_6_1_io_dat_o[15] ,
    \cb_6_1_io_dat_o[14] ,
    \cb_6_1_io_dat_o[13] ,
    \cb_6_1_io_dat_o[12] ,
    \cb_6_1_io_dat_o[11] ,
    \cb_6_1_io_dat_o[10] ,
    \cb_6_1_io_dat_o[9] ,
    \cb_6_1_io_dat_o[8] ,
    \cb_6_1_io_dat_o[7] ,
    \cb_6_1_io_dat_o[6] ,
    \cb_6_1_io_dat_o[5] ,
    \cb_6_1_io_dat_o[4] ,
    \cb_6_1_io_dat_o[3] ,
    \cb_6_1_io_dat_o[2] ,
    \cb_6_1_io_dat_o[1] ,
    \cb_6_1_io_dat_o[0] }),
    .io_b_dat_o_10({\cb_6_10_io_dat_o[15] ,
    \cb_6_10_io_dat_o[14] ,
    \cb_6_10_io_dat_o[13] ,
    \cb_6_10_io_dat_o[12] ,
    \cb_6_10_io_dat_o[11] ,
    \cb_6_10_io_dat_o[10] ,
    \cb_6_10_io_dat_o[9] ,
    \cb_6_10_io_dat_o[8] ,
    \cb_6_10_io_dat_o[7] ,
    \cb_6_10_io_dat_o[6] ,
    \cb_6_10_io_dat_o[5] ,
    \cb_6_10_io_dat_o[4] ,
    \cb_6_10_io_dat_o[3] ,
    \cb_6_10_io_dat_o[2] ,
    \cb_6_10_io_dat_o[1] ,
    \cb_6_10_io_dat_o[0] }),
    .io_b_dat_o_2({\cb_6_2_io_dat_o[15] ,
    \cb_6_2_io_dat_o[14] ,
    \cb_6_2_io_dat_o[13] ,
    \cb_6_2_io_dat_o[12] ,
    \cb_6_2_io_dat_o[11] ,
    \cb_6_2_io_dat_o[10] ,
    \cb_6_2_io_dat_o[9] ,
    \cb_6_2_io_dat_o[8] ,
    \cb_6_2_io_dat_o[7] ,
    \cb_6_2_io_dat_o[6] ,
    \cb_6_2_io_dat_o[5] ,
    \cb_6_2_io_dat_o[4] ,
    \cb_6_2_io_dat_o[3] ,
    \cb_6_2_io_dat_o[2] ,
    \cb_6_2_io_dat_o[1] ,
    \cb_6_2_io_dat_o[0] }),
    .io_b_dat_o_3({\cb_6_3_io_dat_o[15] ,
    \cb_6_3_io_dat_o[14] ,
    \cb_6_3_io_dat_o[13] ,
    \cb_6_3_io_dat_o[12] ,
    \cb_6_3_io_dat_o[11] ,
    \cb_6_3_io_dat_o[10] ,
    \cb_6_3_io_dat_o[9] ,
    \cb_6_3_io_dat_o[8] ,
    \cb_6_3_io_dat_o[7] ,
    \cb_6_3_io_dat_o[6] ,
    \cb_6_3_io_dat_o[5] ,
    \cb_6_3_io_dat_o[4] ,
    \cb_6_3_io_dat_o[3] ,
    \cb_6_3_io_dat_o[2] ,
    \cb_6_3_io_dat_o[1] ,
    \cb_6_3_io_dat_o[0] }),
    .io_b_dat_o_4({\cb_6_4_io_dat_o[15] ,
    \cb_6_4_io_dat_o[14] ,
    \cb_6_4_io_dat_o[13] ,
    \cb_6_4_io_dat_o[12] ,
    \cb_6_4_io_dat_o[11] ,
    \cb_6_4_io_dat_o[10] ,
    \cb_6_4_io_dat_o[9] ,
    \cb_6_4_io_dat_o[8] ,
    \cb_6_4_io_dat_o[7] ,
    \cb_6_4_io_dat_o[6] ,
    \cb_6_4_io_dat_o[5] ,
    \cb_6_4_io_dat_o[4] ,
    \cb_6_4_io_dat_o[3] ,
    \cb_6_4_io_dat_o[2] ,
    \cb_6_4_io_dat_o[1] ,
    \cb_6_4_io_dat_o[0] }),
    .io_b_dat_o_5({\cb_6_5_io_dat_o[15] ,
    \cb_6_5_io_dat_o[14] ,
    \cb_6_5_io_dat_o[13] ,
    \cb_6_5_io_dat_o[12] ,
    \cb_6_5_io_dat_o[11] ,
    \cb_6_5_io_dat_o[10] ,
    \cb_6_5_io_dat_o[9] ,
    \cb_6_5_io_dat_o[8] ,
    \cb_6_5_io_dat_o[7] ,
    \cb_6_5_io_dat_o[6] ,
    \cb_6_5_io_dat_o[5] ,
    \cb_6_5_io_dat_o[4] ,
    \cb_6_5_io_dat_o[3] ,
    \cb_6_5_io_dat_o[2] ,
    \cb_6_5_io_dat_o[1] ,
    \cb_6_5_io_dat_o[0] }),
    .io_b_dat_o_6({\cb_6_6_io_dat_o[15] ,
    \cb_6_6_io_dat_o[14] ,
    \cb_6_6_io_dat_o[13] ,
    \cb_6_6_io_dat_o[12] ,
    \cb_6_6_io_dat_o[11] ,
    \cb_6_6_io_dat_o[10] ,
    \cb_6_6_io_dat_o[9] ,
    \cb_6_6_io_dat_o[8] ,
    \cb_6_6_io_dat_o[7] ,
    \cb_6_6_io_dat_o[6] ,
    \cb_6_6_io_dat_o[5] ,
    \cb_6_6_io_dat_o[4] ,
    \cb_6_6_io_dat_o[3] ,
    \cb_6_6_io_dat_o[2] ,
    \cb_6_6_io_dat_o[1] ,
    \cb_6_6_io_dat_o[0] }),
    .io_b_dat_o_7({\cb_6_7_io_dat_o[15] ,
    \cb_6_7_io_dat_o[14] ,
    \cb_6_7_io_dat_o[13] ,
    \cb_6_7_io_dat_o[12] ,
    \cb_6_7_io_dat_o[11] ,
    \cb_6_7_io_dat_o[10] ,
    \cb_6_7_io_dat_o[9] ,
    \cb_6_7_io_dat_o[8] ,
    \cb_6_7_io_dat_o[7] ,
    \cb_6_7_io_dat_o[6] ,
    \cb_6_7_io_dat_o[5] ,
    \cb_6_7_io_dat_o[4] ,
    \cb_6_7_io_dat_o[3] ,
    \cb_6_7_io_dat_o[2] ,
    \cb_6_7_io_dat_o[1] ,
    \cb_6_7_io_dat_o[0] }),
    .io_b_dat_o_8({\cb_6_8_io_dat_o[15] ,
    \cb_6_8_io_dat_o[14] ,
    \cb_6_8_io_dat_o[13] ,
    \cb_6_8_io_dat_o[12] ,
    \cb_6_8_io_dat_o[11] ,
    \cb_6_8_io_dat_o[10] ,
    \cb_6_8_io_dat_o[9] ,
    \cb_6_8_io_dat_o[8] ,
    \cb_6_8_io_dat_o[7] ,
    \cb_6_8_io_dat_o[6] ,
    \cb_6_8_io_dat_o[5] ,
    \cb_6_8_io_dat_o[4] ,
    \cb_6_8_io_dat_o[3] ,
    \cb_6_8_io_dat_o[2] ,
    \cb_6_8_io_dat_o[1] ,
    \cb_6_8_io_dat_o[0] }),
    .io_b_dat_o_9({\cb_6_9_io_dat_o[15] ,
    \cb_6_9_io_dat_o[14] ,
    \cb_6_9_io_dat_o[13] ,
    \cb_6_9_io_dat_o[12] ,
    \cb_6_9_io_dat_o[11] ,
    \cb_6_9_io_dat_o[10] ,
    \cb_6_9_io_dat_o[9] ,
    \cb_6_9_io_dat_o[8] ,
    \cb_6_9_io_dat_o[7] ,
    \cb_6_9_io_dat_o[6] ,
    \cb_6_9_io_dat_o[5] ,
    \cb_6_9_io_dat_o[4] ,
    \cb_6_9_io_dat_o[3] ,
    \cb_6_9_io_dat_o[2] ,
    \cb_6_9_io_dat_o[1] ,
    \cb_6_9_io_dat_o[0] }),
    .io_dat_i({\ccon_0_io_dat_i[31] ,
    \ccon_0_io_dat_i[30] ,
    \ccon_0_io_dat_i[29] ,
    \ccon_0_io_dat_i[28] ,
    \ccon_0_io_dat_i[27] ,
    \ccon_0_io_dat_i[26] ,
    \ccon_0_io_dat_i[25] ,
    \ccon_0_io_dat_i[24] ,
    \ccon_0_io_dat_i[23] ,
    \ccon_0_io_dat_i[22] ,
    \ccon_0_io_dat_i[21] ,
    \ccon_0_io_dat_i[20] ,
    \ccon_0_io_dat_i[19] ,
    \ccon_0_io_dat_i[18] ,
    \ccon_0_io_dat_i[17] ,
    \ccon_0_io_dat_i[16] ,
    \ccon_0_io_dat_i[15] ,
    \ccon_0_io_dat_i[14] ,
    \ccon_0_io_dat_i[13] ,
    \ccon_0_io_dat_i[12] ,
    \ccon_0_io_dat_i[11] ,
    \ccon_0_io_dat_i[10] ,
    \ccon_0_io_dat_i[9] ,
    \ccon_0_io_dat_i[8] ,
    \ccon_0_io_dat_i[7] ,
    \ccon_0_io_dat_i[6] ,
    \ccon_0_io_dat_i[5] ,
    \ccon_0_io_dat_i[4] ,
    \ccon_0_io_dat_i[3] ,
    \ccon_0_io_dat_i[2] ,
    \ccon_0_io_dat_i[1] ,
    \ccon_0_io_dat_i[0] }),
    .io_dat_o({\ccon_6_io_dat_o[31] ,
    \ccon_6_io_dat_o[30] ,
    \ccon_6_io_dat_o[29] ,
    \ccon_6_io_dat_o[28] ,
    \ccon_6_io_dat_o[27] ,
    \ccon_6_io_dat_o[26] ,
    \ccon_6_io_dat_o[25] ,
    \ccon_6_io_dat_o[24] ,
    \ccon_6_io_dat_o[23] ,
    \ccon_6_io_dat_o[22] ,
    \ccon_6_io_dat_o[21] ,
    \ccon_6_io_dat_o[20] ,
    \ccon_6_io_dat_o[19] ,
    \ccon_6_io_dat_o[18] ,
    \ccon_6_io_dat_o[17] ,
    \ccon_6_io_dat_o[16] ,
    \ccon_6_io_dat_o[15] ,
    \ccon_6_io_dat_o[14] ,
    \ccon_6_io_dat_o[13] ,
    \ccon_6_io_dat_o[12] ,
    \ccon_6_io_dat_o[11] ,
    \ccon_6_io_dat_o[10] ,
    \ccon_6_io_dat_o[9] ,
    \ccon_6_io_dat_o[8] ,
    \ccon_6_io_dat_o[7] ,
    \ccon_6_io_dat_o[6] ,
    \ccon_6_io_dat_o[5] ,
    \ccon_6_io_dat_o[4] ,
    \ccon_6_io_dat_o[3] ,
    \ccon_6_io_dat_o[2] ,
    \ccon_6_io_dat_o[1] ,
    \ccon_6_io_dat_o[0] }),
    .io_dataLastBlock({\cb_6_0_io_wo[63] ,
    \cb_6_0_io_wo[62] ,
    \cb_6_0_io_wo[61] ,
    \cb_6_0_io_wo[60] ,
    \cb_6_0_io_wo[59] ,
    \cb_6_0_io_wo[58] ,
    \cb_6_0_io_wo[57] ,
    \cb_6_0_io_wo[56] ,
    \cb_6_0_io_wo[55] ,
    \cb_6_0_io_wo[54] ,
    \cb_6_0_io_wo[53] ,
    \cb_6_0_io_wo[52] ,
    \cb_6_0_io_wo[51] ,
    \cb_6_0_io_wo[50] ,
    \cb_6_0_io_wo[49] ,
    \cb_6_0_io_wo[48] ,
    \cb_6_0_io_wo[47] ,
    \cb_6_0_io_wo[46] ,
    \cb_6_0_io_wo[45] ,
    \cb_6_0_io_wo[44] ,
    \cb_6_0_io_wo[43] ,
    \cb_6_0_io_wo[42] ,
    \cb_6_0_io_wo[41] ,
    \cb_6_0_io_wo[40] ,
    \cb_6_0_io_wo[39] ,
    \cb_6_0_io_wo[38] ,
    \cb_6_0_io_wo[37] ,
    \cb_6_0_io_wo[36] ,
    \cb_6_0_io_wo[35] ,
    \cb_6_0_io_wo[34] ,
    \cb_6_0_io_wo[33] ,
    \cb_6_0_io_wo[32] ,
    \cb_6_0_io_wo[31] ,
    \cb_6_0_io_wo[30] ,
    \cb_6_0_io_wo[29] ,
    \cb_6_0_io_wo[28] ,
    \cb_6_0_io_wo[27] ,
    \cb_6_0_io_wo[26] ,
    \cb_6_0_io_wo[25] ,
    \cb_6_0_io_wo[24] ,
    \cb_6_0_io_wo[23] ,
    \cb_6_0_io_wo[22] ,
    \cb_6_0_io_wo[21] ,
    \cb_6_0_io_wo[20] ,
    \cb_6_0_io_wo[19] ,
    \cb_6_0_io_wo[18] ,
    \cb_6_0_io_wo[17] ,
    \cb_6_0_io_wo[16] ,
    \cb_6_0_io_wo[15] ,
    \cb_6_0_io_wo[14] ,
    \cb_6_0_io_wo[13] ,
    \cb_6_0_io_wo[12] ,
    \cb_6_0_io_wo[11] ,
    \cb_6_0_io_wo[10] ,
    \cb_6_0_io_wo[9] ,
    \cb_6_0_io_wo[8] ,
    \cb_6_0_io_wo[7] ,
    \cb_6_0_io_wo[6] ,
    \cb_6_0_io_wo[5] ,
    \cb_6_0_io_wo[4] ,
    \cb_6_0_io_wo[3] ,
    \cb_6_0_io_wo[2] ,
    \cb_6_0_io_wo[1] ,
    \cb_6_0_io_wo[0] }),
    .io_dsi_in({\ccon_0_io_dsi_in[7] ,
    \ccon_0_io_dsi_in[6] ,
    \ccon_0_io_dsi_in[5] ,
    \ccon_0_io_dsi_in[4] ,
    \ccon_0_io_dsi_in[3] ,
    \ccon_0_io_dsi_in[2] ,
    \ccon_0_io_dsi_in[1] ,
    \ccon_0_io_dsi_in[0] }),
    .io_vout({cb_6_10_io_vi,
    cb_6_9_io_vi,
    cb_6_8_io_vi,
    cb_6_7_io_vi,
    cb_6_6_io_vi,
    cb_6_5_io_vi,
    cb_6_4_io_vi,
    cb_6_3_io_vi,
    cb_6_2_io_vi,
    cb_6_1_io_vi,
    cb_6_0_io_vi}));
 cic_con ccon_7 (.io_ack_o(\_T_172[5] ),
    .io_b_cs_i_0(cb_7_0_io_cs_i),
    .io_b_cs_i_1(cb_7_1_io_cs_i),
    .io_b_cs_i_10(cb_7_10_io_cs_i),
    .io_b_cs_i_2(cb_7_2_io_cs_i),
    .io_b_cs_i_3(cb_7_3_io_cs_i),
    .io_b_cs_i_4(cb_7_4_io_cs_i),
    .io_b_cs_i_5(cb_7_5_io_cs_i),
    .io_b_cs_i_6(cb_7_6_io_cs_i),
    .io_b_cs_i_7(cb_7_7_io_cs_i),
    .io_b_cs_i_8(cb_7_8_io_cs_i),
    .io_b_cs_i_9(cb_7_9_io_cs_i),
    .io_b_we_i(cb_7_0_io_we_i),
    .io_cs_i(ccon_7_io_cs_i),
    .io_dsi_o(cb_7_0_io_i_0_ci),
    .io_irq(\_T_183[5] ),
    .io_we_i(ccon_0_io_we_i),
    .wb_clk_i(cb_0_0_wb_clk_i),
    .wb_rst_i(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_adr_i({\ccon_0_io_adr_i[11] ,
    \ccon_0_io_adr_i[10] ,
    \ccon_0_io_adr_i[9] ,
    \ccon_0_io_adr_i[8] ,
    \ccon_0_io_adr_i[7] ,
    \ccon_0_io_adr_i[6] ,
    \ccon_0_io_adr_i[5] ,
    \ccon_0_io_adr_i[4] ,
    \ccon_0_io_adr_i[3] ,
    \ccon_0_io_adr_i[2] ,
    \ccon_0_io_adr_i[1] ,
    \ccon_0_io_adr_i[0] }),
    .io_b_adr_i({\cb_7_0_io_adr_i[1] ,
    \cb_7_0_io_adr_i[0] }),
    .io_b_dat_i({\cb_7_0_io_dat_i[15] ,
    \cb_7_0_io_dat_i[14] ,
    \cb_7_0_io_dat_i[13] ,
    \cb_7_0_io_dat_i[12] ,
    \cb_7_0_io_dat_i[11] ,
    \cb_7_0_io_dat_i[10] ,
    \cb_7_0_io_dat_i[9] ,
    \cb_7_0_io_dat_i[8] ,
    \cb_7_0_io_dat_i[7] ,
    \cb_7_0_io_dat_i[6] ,
    \cb_7_0_io_dat_i[5] ,
    \cb_7_0_io_dat_i[4] ,
    \cb_7_0_io_dat_i[3] ,
    \cb_7_0_io_dat_i[2] ,
    \cb_7_0_io_dat_i[1] ,
    \cb_7_0_io_dat_i[0] }),
    .io_b_dat_o_0({\cb_7_0_io_dat_o[15] ,
    \cb_7_0_io_dat_o[14] ,
    \cb_7_0_io_dat_o[13] ,
    \cb_7_0_io_dat_o[12] ,
    \cb_7_0_io_dat_o[11] ,
    \cb_7_0_io_dat_o[10] ,
    \cb_7_0_io_dat_o[9] ,
    \cb_7_0_io_dat_o[8] ,
    \cb_7_0_io_dat_o[7] ,
    \cb_7_0_io_dat_o[6] ,
    \cb_7_0_io_dat_o[5] ,
    \cb_7_0_io_dat_o[4] ,
    \cb_7_0_io_dat_o[3] ,
    \cb_7_0_io_dat_o[2] ,
    \cb_7_0_io_dat_o[1] ,
    \cb_7_0_io_dat_o[0] }),
    .io_b_dat_o_1({\cb_7_1_io_dat_o[15] ,
    \cb_7_1_io_dat_o[14] ,
    \cb_7_1_io_dat_o[13] ,
    \cb_7_1_io_dat_o[12] ,
    \cb_7_1_io_dat_o[11] ,
    \cb_7_1_io_dat_o[10] ,
    \cb_7_1_io_dat_o[9] ,
    \cb_7_1_io_dat_o[8] ,
    \cb_7_1_io_dat_o[7] ,
    \cb_7_1_io_dat_o[6] ,
    \cb_7_1_io_dat_o[5] ,
    \cb_7_1_io_dat_o[4] ,
    \cb_7_1_io_dat_o[3] ,
    \cb_7_1_io_dat_o[2] ,
    \cb_7_1_io_dat_o[1] ,
    \cb_7_1_io_dat_o[0] }),
    .io_b_dat_o_10({\cb_7_10_io_dat_o[15] ,
    \cb_7_10_io_dat_o[14] ,
    \cb_7_10_io_dat_o[13] ,
    \cb_7_10_io_dat_o[12] ,
    \cb_7_10_io_dat_o[11] ,
    \cb_7_10_io_dat_o[10] ,
    \cb_7_10_io_dat_o[9] ,
    \cb_7_10_io_dat_o[8] ,
    \cb_7_10_io_dat_o[7] ,
    \cb_7_10_io_dat_o[6] ,
    \cb_7_10_io_dat_o[5] ,
    \cb_7_10_io_dat_o[4] ,
    \cb_7_10_io_dat_o[3] ,
    \cb_7_10_io_dat_o[2] ,
    \cb_7_10_io_dat_o[1] ,
    \cb_7_10_io_dat_o[0] }),
    .io_b_dat_o_2({\cb_7_2_io_dat_o[15] ,
    \cb_7_2_io_dat_o[14] ,
    \cb_7_2_io_dat_o[13] ,
    \cb_7_2_io_dat_o[12] ,
    \cb_7_2_io_dat_o[11] ,
    \cb_7_2_io_dat_o[10] ,
    \cb_7_2_io_dat_o[9] ,
    \cb_7_2_io_dat_o[8] ,
    \cb_7_2_io_dat_o[7] ,
    \cb_7_2_io_dat_o[6] ,
    \cb_7_2_io_dat_o[5] ,
    \cb_7_2_io_dat_o[4] ,
    \cb_7_2_io_dat_o[3] ,
    \cb_7_2_io_dat_o[2] ,
    \cb_7_2_io_dat_o[1] ,
    \cb_7_2_io_dat_o[0] }),
    .io_b_dat_o_3({\cb_7_3_io_dat_o[15] ,
    \cb_7_3_io_dat_o[14] ,
    \cb_7_3_io_dat_o[13] ,
    \cb_7_3_io_dat_o[12] ,
    \cb_7_3_io_dat_o[11] ,
    \cb_7_3_io_dat_o[10] ,
    \cb_7_3_io_dat_o[9] ,
    \cb_7_3_io_dat_o[8] ,
    \cb_7_3_io_dat_o[7] ,
    \cb_7_3_io_dat_o[6] ,
    \cb_7_3_io_dat_o[5] ,
    \cb_7_3_io_dat_o[4] ,
    \cb_7_3_io_dat_o[3] ,
    \cb_7_3_io_dat_o[2] ,
    \cb_7_3_io_dat_o[1] ,
    \cb_7_3_io_dat_o[0] }),
    .io_b_dat_o_4({\cb_7_4_io_dat_o[15] ,
    \cb_7_4_io_dat_o[14] ,
    \cb_7_4_io_dat_o[13] ,
    \cb_7_4_io_dat_o[12] ,
    \cb_7_4_io_dat_o[11] ,
    \cb_7_4_io_dat_o[10] ,
    \cb_7_4_io_dat_o[9] ,
    \cb_7_4_io_dat_o[8] ,
    \cb_7_4_io_dat_o[7] ,
    \cb_7_4_io_dat_o[6] ,
    \cb_7_4_io_dat_o[5] ,
    \cb_7_4_io_dat_o[4] ,
    \cb_7_4_io_dat_o[3] ,
    \cb_7_4_io_dat_o[2] ,
    \cb_7_4_io_dat_o[1] ,
    \cb_7_4_io_dat_o[0] }),
    .io_b_dat_o_5({\cb_7_5_io_dat_o[15] ,
    \cb_7_5_io_dat_o[14] ,
    \cb_7_5_io_dat_o[13] ,
    \cb_7_5_io_dat_o[12] ,
    \cb_7_5_io_dat_o[11] ,
    \cb_7_5_io_dat_o[10] ,
    \cb_7_5_io_dat_o[9] ,
    \cb_7_5_io_dat_o[8] ,
    \cb_7_5_io_dat_o[7] ,
    \cb_7_5_io_dat_o[6] ,
    \cb_7_5_io_dat_o[5] ,
    \cb_7_5_io_dat_o[4] ,
    \cb_7_5_io_dat_o[3] ,
    \cb_7_5_io_dat_o[2] ,
    \cb_7_5_io_dat_o[1] ,
    \cb_7_5_io_dat_o[0] }),
    .io_b_dat_o_6({\cb_7_6_io_dat_o[15] ,
    \cb_7_6_io_dat_o[14] ,
    \cb_7_6_io_dat_o[13] ,
    \cb_7_6_io_dat_o[12] ,
    \cb_7_6_io_dat_o[11] ,
    \cb_7_6_io_dat_o[10] ,
    \cb_7_6_io_dat_o[9] ,
    \cb_7_6_io_dat_o[8] ,
    \cb_7_6_io_dat_o[7] ,
    \cb_7_6_io_dat_o[6] ,
    \cb_7_6_io_dat_o[5] ,
    \cb_7_6_io_dat_o[4] ,
    \cb_7_6_io_dat_o[3] ,
    \cb_7_6_io_dat_o[2] ,
    \cb_7_6_io_dat_o[1] ,
    \cb_7_6_io_dat_o[0] }),
    .io_b_dat_o_7({\cb_7_7_io_dat_o[15] ,
    \cb_7_7_io_dat_o[14] ,
    \cb_7_7_io_dat_o[13] ,
    \cb_7_7_io_dat_o[12] ,
    \cb_7_7_io_dat_o[11] ,
    \cb_7_7_io_dat_o[10] ,
    \cb_7_7_io_dat_o[9] ,
    \cb_7_7_io_dat_o[8] ,
    \cb_7_7_io_dat_o[7] ,
    \cb_7_7_io_dat_o[6] ,
    \cb_7_7_io_dat_o[5] ,
    \cb_7_7_io_dat_o[4] ,
    \cb_7_7_io_dat_o[3] ,
    \cb_7_7_io_dat_o[2] ,
    \cb_7_7_io_dat_o[1] ,
    \cb_7_7_io_dat_o[0] }),
    .io_b_dat_o_8({\cb_7_8_io_dat_o[15] ,
    \cb_7_8_io_dat_o[14] ,
    \cb_7_8_io_dat_o[13] ,
    \cb_7_8_io_dat_o[12] ,
    \cb_7_8_io_dat_o[11] ,
    \cb_7_8_io_dat_o[10] ,
    \cb_7_8_io_dat_o[9] ,
    \cb_7_8_io_dat_o[8] ,
    \cb_7_8_io_dat_o[7] ,
    \cb_7_8_io_dat_o[6] ,
    \cb_7_8_io_dat_o[5] ,
    \cb_7_8_io_dat_o[4] ,
    \cb_7_8_io_dat_o[3] ,
    \cb_7_8_io_dat_o[2] ,
    \cb_7_8_io_dat_o[1] ,
    \cb_7_8_io_dat_o[0] }),
    .io_b_dat_o_9({\cb_7_9_io_dat_o[15] ,
    \cb_7_9_io_dat_o[14] ,
    \cb_7_9_io_dat_o[13] ,
    \cb_7_9_io_dat_o[12] ,
    \cb_7_9_io_dat_o[11] ,
    \cb_7_9_io_dat_o[10] ,
    \cb_7_9_io_dat_o[9] ,
    \cb_7_9_io_dat_o[8] ,
    \cb_7_9_io_dat_o[7] ,
    \cb_7_9_io_dat_o[6] ,
    \cb_7_9_io_dat_o[5] ,
    \cb_7_9_io_dat_o[4] ,
    \cb_7_9_io_dat_o[3] ,
    \cb_7_9_io_dat_o[2] ,
    \cb_7_9_io_dat_o[1] ,
    \cb_7_9_io_dat_o[0] }),
    .io_dat_i({\ccon_0_io_dat_i[31] ,
    \ccon_0_io_dat_i[30] ,
    \ccon_0_io_dat_i[29] ,
    \ccon_0_io_dat_i[28] ,
    \ccon_0_io_dat_i[27] ,
    \ccon_0_io_dat_i[26] ,
    \ccon_0_io_dat_i[25] ,
    \ccon_0_io_dat_i[24] ,
    \ccon_0_io_dat_i[23] ,
    \ccon_0_io_dat_i[22] ,
    \ccon_0_io_dat_i[21] ,
    \ccon_0_io_dat_i[20] ,
    \ccon_0_io_dat_i[19] ,
    \ccon_0_io_dat_i[18] ,
    \ccon_0_io_dat_i[17] ,
    \ccon_0_io_dat_i[16] ,
    \ccon_0_io_dat_i[15] ,
    \ccon_0_io_dat_i[14] ,
    \ccon_0_io_dat_i[13] ,
    \ccon_0_io_dat_i[12] ,
    \ccon_0_io_dat_i[11] ,
    \ccon_0_io_dat_i[10] ,
    \ccon_0_io_dat_i[9] ,
    \ccon_0_io_dat_i[8] ,
    \ccon_0_io_dat_i[7] ,
    \ccon_0_io_dat_i[6] ,
    \ccon_0_io_dat_i[5] ,
    \ccon_0_io_dat_i[4] ,
    \ccon_0_io_dat_i[3] ,
    \ccon_0_io_dat_i[2] ,
    \ccon_0_io_dat_i[1] ,
    \ccon_0_io_dat_i[0] }),
    .io_dat_o({\ccon_7_io_dat_o[31] ,
    \ccon_7_io_dat_o[30] ,
    \ccon_7_io_dat_o[29] ,
    \ccon_7_io_dat_o[28] ,
    \ccon_7_io_dat_o[27] ,
    \ccon_7_io_dat_o[26] ,
    \ccon_7_io_dat_o[25] ,
    \ccon_7_io_dat_o[24] ,
    \ccon_7_io_dat_o[23] ,
    \ccon_7_io_dat_o[22] ,
    \ccon_7_io_dat_o[21] ,
    \ccon_7_io_dat_o[20] ,
    \ccon_7_io_dat_o[19] ,
    \ccon_7_io_dat_o[18] ,
    \ccon_7_io_dat_o[17] ,
    \ccon_7_io_dat_o[16] ,
    \ccon_7_io_dat_o[15] ,
    \ccon_7_io_dat_o[14] ,
    \ccon_7_io_dat_o[13] ,
    \ccon_7_io_dat_o[12] ,
    \ccon_7_io_dat_o[11] ,
    \ccon_7_io_dat_o[10] ,
    \ccon_7_io_dat_o[9] ,
    \ccon_7_io_dat_o[8] ,
    \ccon_7_io_dat_o[7] ,
    \ccon_7_io_dat_o[6] ,
    \ccon_7_io_dat_o[5] ,
    \ccon_7_io_dat_o[4] ,
    \ccon_7_io_dat_o[3] ,
    \ccon_7_io_dat_o[2] ,
    \ccon_7_io_dat_o[1] ,
    \ccon_7_io_dat_o[0] }),
    .io_dataLastBlock({\cb_7_0_io_wo[63] ,
    \cb_7_0_io_wo[62] ,
    \cb_7_0_io_wo[61] ,
    \cb_7_0_io_wo[60] ,
    \cb_7_0_io_wo[59] ,
    \cb_7_0_io_wo[58] ,
    \cb_7_0_io_wo[57] ,
    \cb_7_0_io_wo[56] ,
    \cb_7_0_io_wo[55] ,
    \cb_7_0_io_wo[54] ,
    \cb_7_0_io_wo[53] ,
    \cb_7_0_io_wo[52] ,
    \cb_7_0_io_wo[51] ,
    \cb_7_0_io_wo[50] ,
    \cb_7_0_io_wo[49] ,
    \cb_7_0_io_wo[48] ,
    \cb_7_0_io_wo[47] ,
    \cb_7_0_io_wo[46] ,
    \cb_7_0_io_wo[45] ,
    \cb_7_0_io_wo[44] ,
    \cb_7_0_io_wo[43] ,
    \cb_7_0_io_wo[42] ,
    \cb_7_0_io_wo[41] ,
    \cb_7_0_io_wo[40] ,
    \cb_7_0_io_wo[39] ,
    \cb_7_0_io_wo[38] ,
    \cb_7_0_io_wo[37] ,
    \cb_7_0_io_wo[36] ,
    \cb_7_0_io_wo[35] ,
    \cb_7_0_io_wo[34] ,
    \cb_7_0_io_wo[33] ,
    \cb_7_0_io_wo[32] ,
    \cb_7_0_io_wo[31] ,
    \cb_7_0_io_wo[30] ,
    \cb_7_0_io_wo[29] ,
    \cb_7_0_io_wo[28] ,
    \cb_7_0_io_wo[27] ,
    \cb_7_0_io_wo[26] ,
    \cb_7_0_io_wo[25] ,
    \cb_7_0_io_wo[24] ,
    \cb_7_0_io_wo[23] ,
    \cb_7_0_io_wo[22] ,
    \cb_7_0_io_wo[21] ,
    \cb_7_0_io_wo[20] ,
    \cb_7_0_io_wo[19] ,
    \cb_7_0_io_wo[18] ,
    \cb_7_0_io_wo[17] ,
    \cb_7_0_io_wo[16] ,
    \cb_7_0_io_wo[15] ,
    \cb_7_0_io_wo[14] ,
    \cb_7_0_io_wo[13] ,
    \cb_7_0_io_wo[12] ,
    \cb_7_0_io_wo[11] ,
    \cb_7_0_io_wo[10] ,
    \cb_7_0_io_wo[9] ,
    \cb_7_0_io_wo[8] ,
    \cb_7_0_io_wo[7] ,
    \cb_7_0_io_wo[6] ,
    \cb_7_0_io_wo[5] ,
    \cb_7_0_io_wo[4] ,
    \cb_7_0_io_wo[3] ,
    \cb_7_0_io_wo[2] ,
    \cb_7_0_io_wo[1] ,
    \cb_7_0_io_wo[0] }),
    .io_dsi_in({\ccon_0_io_dsi_in[7] ,
    \ccon_0_io_dsi_in[6] ,
    \ccon_0_io_dsi_in[5] ,
    \ccon_0_io_dsi_in[4] ,
    \ccon_0_io_dsi_in[3] ,
    \ccon_0_io_dsi_in[2] ,
    \ccon_0_io_dsi_in[1] ,
    \ccon_0_io_dsi_in[0] }),
    .io_vout({cb_7_10_io_vi,
    cb_7_9_io_vi,
    cb_7_8_io_vi,
    cb_7_7_io_vi,
    cb_7_6_io_vi,
    cb_7_5_io_vi,
    cb_7_4_io_vi,
    cb_7_3_io_vi,
    cb_7_2_io_vi,
    cb_7_1_io_vi,
    cb_7_0_io_vi}));
 sin3 cordic (.vccd1(vccd1),
    .vssd1(vssd1),
    .ao_reg({_NC513,
    _NC514,
    _NC515,
    _NC516,
    _NC517,
    _NC518,
    _NC519,
    _NC520,
    _NC521,
    _NC522,
    _NC523,
    _NC524,
    _NC525,
    _NC526,
    _NC527,
    _NC528,
    _NC529,
    _NC530,
    _NC531,
    _NC532,
    _NC533,
    _NC534,
    _NC535,
    _NC536,
    _NC537,
    _NC538,
    _NC539,
    _NC540,
    _NC541,
    _NC542,
    _NC543,
    _NC544}),
    .bo_reg({_NC545,
    _NC546,
    _NC547,
    _NC548,
    _NC549,
    _NC550,
    _NC551,
    _NC552,
    _NC553,
    _NC554,
    _NC555,
    _NC556,
    _NC557,
    _NC558,
    _NC559,
    _NC560,
    _NC561,
    _NC562,
    _NC563,
    _NC564,
    _NC565,
    _NC566,
    _NC567,
    _NC568,
    _NC569,
    _NC570,
    _NC571,
    _NC572,
    _NC573,
    _NC574,
    _NC575,
    _NC576}),
    .e_i({la_data_in[127],
    la_data_in[126],
    la_data_in[125],
    la_data_in[124],
    la_data_in[123],
    la_data_in[122],
    la_data_in[121],
    la_data_in[120],
    la_data_in[119],
    la_data_in[118],
    la_data_in[117],
    la_data_in[116],
    la_data_in[115],
    la_data_in[114],
    la_data_in[113],
    la_data_in[112],
    la_data_in[111],
    la_data_in[110],
    la_data_in[109],
    la_data_in[108],
    la_data_in[107],
    la_data_in[106],
    la_data_in[105],
    la_data_in[104],
    la_data_in[103],
    la_data_in[102],
    la_data_in[101],
    la_data_in[100],
    la_data_in[99],
    la_data_in[98],
    la_data_in[97],
    la_data_in[96]}),
    .e_o({la_data_out[127],
    la_data_out[126],
    la_data_out[125],
    la_data_out[124],
    la_data_out[123],
    la_data_out[122],
    la_data_out[121],
    la_data_out[120],
    la_data_out[119],
    la_data_out[118],
    la_data_out[117],
    la_data_out[116],
    la_data_out[115],
    la_data_out[114],
    la_data_out[113],
    la_data_out[112],
    la_data_out[111],
    la_data_out[110],
    la_data_out[109],
    la_data_out[108],
    la_data_out[107],
    la_data_out[106],
    la_data_out[105],
    la_data_out[104],
    la_data_out[103],
    la_data_out[102],
    la_data_out[101],
    la_data_out[100],
    la_data_out[99],
    la_data_out[98],
    la_data_out[97],
    la_data_out[96]}),
    .se_i({la_data_in[95],
    la_data_in[94],
    la_data_in[93],
    la_data_in[92],
    la_data_in[91],
    la_data_in[90],
    la_data_in[89],
    la_data_in[88],
    la_data_in[87],
    la_data_in[86],
    la_data_in[85],
    la_data_in[84],
    la_data_in[83],
    la_data_in[82],
    la_data_in[81],
    la_data_in[80],
    la_data_in[79],
    la_data_in[78],
    la_data_in[77],
    la_data_in[76],
    la_data_in[75],
    la_data_in[74],
    la_data_in[73],
    la_data_in[72],
    la_data_in[71],
    la_data_in[70],
    la_data_in[69],
    la_data_in[68],
    la_data_in[67],
    la_data_in[66],
    la_data_in[65],
    la_data_in[64]}),
    .se_o({la_data_out[95],
    la_data_out[94],
    la_data_out[93],
    la_data_out[92],
    la_data_out[91],
    la_data_out[90],
    la_data_out[89],
    la_data_out[88],
    la_data_out[87],
    la_data_out[86],
    la_data_out[85],
    la_data_out[84],
    la_data_out[83],
    la_data_out[82],
    la_data_out[81],
    la_data_out[80],
    la_data_out[79],
    la_data_out[78],
    la_data_out[77],
    la_data_out[76],
    la_data_out[75],
    la_data_out[74],
    la_data_out[73],
    la_data_out[72],
    la_data_out[71],
    la_data_out[70],
    la_data_out[69],
    la_data_out[68],
    la_data_out[67],
    la_data_out[66],
    la_data_out[65],
    la_data_out[64]}),
    .sw_i({la_data_in[63],
    la_data_in[62],
    la_data_in[61],
    la_data_in[60],
    la_data_in[59],
    la_data_in[58],
    la_data_in[57],
    la_data_in[56],
    la_data_in[55],
    la_data_in[54],
    la_data_in[53],
    la_data_in[52],
    la_data_in[51],
    la_data_in[50],
    la_data_in[49],
    la_data_in[48],
    la_data_in[47],
    la_data_in[46],
    la_data_in[45],
    la_data_in[44],
    la_data_in[43],
    la_data_in[42],
    la_data_in[41],
    la_data_in[40],
    la_data_in[39],
    la_data_in[38],
    la_data_in[37],
    la_data_in[36],
    la_data_in[35],
    la_data_in[34],
    la_data_in[33],
    la_data_in[32]}),
    .sw_o({la_data_out[63],
    la_data_out[62],
    la_data_out[61],
    la_data_out[60],
    la_data_out[59],
    la_data_out[58],
    la_data_out[57],
    la_data_out[56],
    la_data_out[55],
    la_data_out[54],
    la_data_out[53],
    la_data_out[52],
    la_data_out[51],
    la_data_out[50],
    la_data_out[49],
    la_data_out[48],
    la_data_out[47],
    la_data_out[46],
    la_data_out[45],
    la_data_out[44],
    la_data_out[43],
    la_data_out[42],
    la_data_out[41],
    la_data_out[40],
    la_data_out[39],
    la_data_out[38],
    la_data_out[37],
    la_data_out[36],
    la_data_out[35],
    la_data_out[34],
    la_data_out[33],
    la_data_out[32]}),
    .w_i({la_data_in[31],
    la_data_in[30],
    la_data_in[29],
    la_data_in[28],
    la_data_in[27],
    la_data_in[26],
    la_data_in[25],
    la_data_in[24],
    la_data_in[23],
    la_data_in[22],
    la_data_in[21],
    la_data_in[20],
    la_data_in[19],
    la_data_in[18],
    la_data_in[17],
    la_data_in[16],
    la_data_in[15],
    la_data_in[14],
    la_data_in[13],
    la_data_in[12],
    la_data_in[11],
    la_data_in[10],
    la_data_in[9],
    la_data_in[8],
    la_data_in[7],
    la_data_in[6],
    la_data_in[5],
    la_data_in[4],
    la_data_in[3],
    la_data_in[2],
    la_data_in[1],
    la_data_in[0]}),
    .w_o({la_data_out[31],
    la_data_out[30],
    la_data_out[29],
    la_data_out[28],
    la_data_out[27],
    la_data_out[26],
    la_data_out[25],
    la_data_out[24],
    la_data_out[23],
    la_data_out[22],
    la_data_out[21],
    la_data_out[20],
    la_data_out[19],
    la_data_out[18],
    la_data_out[17],
    la_data_out[16],
    la_data_out[15],
    la_data_out[14],
    la_data_out[13],
    la_data_out[12],
    la_data_out[11],
    la_data_out[10],
    la_data_out[9],
    la_data_out[8],
    la_data_out[7],
    la_data_out[6],
    la_data_out[5],
    la_data_out[4],
    la_data_out[3],
    la_data_out[2],
    la_data_out[1],
    la_data_out[0]}));
 wb_local icon (.m_wb_clk_i(cb_0_0_wb_clk_i),
    .m_wb_rst_i(cb_0_0_wb_rst_i),
    .m_wbs_we_i(ccon_0_io_we_i),
    .mt_QEI_ChA_0(icon_mt_QEI_ChA_0),
    .mt_QEI_ChA_1(icon_mt_QEI_ChA_1),
    .mt_QEI_ChA_2(icon_mt_QEI_ChA_2),
    .mt_QEI_ChA_3(icon_mt_QEI_ChA_3),
    .mt_QEI_ChB_0(icon_mt_QEI_ChB_0),
    .mt_QEI_ChB_1(icon_mt_QEI_ChB_1),
    .mt_QEI_ChB_2(icon_mt_QEI_ChB_2),
    .mt_QEI_ChB_3(icon_mt_QEI_ChB_3),
    .mt_pwm_h_0(icon_mt_pwm_h_0),
    .mt_pwm_h_1(icon_mt_pwm_h_1),
    .mt_pwm_h_2(icon_mt_pwm_h_2),
    .mt_pwm_h_3(icon_mt_pwm_h_3),
    .mt_pwm_l_0(icon_mt_pwm_l_0),
    .mt_pwm_l_1(icon_mt_pwm_l_1),
    .mt_pwm_l_2(icon_mt_pwm_l_2),
    .mt_pwm_l_3(icon_mt_pwm_l_3),
    .wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),
    .wbs_ack_o(wbs_ack_o),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(wbs_stb_i),
    .wbs_we_i(wbs_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .dsi({\ccon_0_io_dsi_in[7] ,
    \ccon_0_io_dsi_in[6] ,
    \ccon_0_io_dsi_in[5] ,
    \ccon_0_io_dsi_in[4] ,
    \ccon_0_io_dsi_in[3] ,
    \ccon_0_io_dsi_in[2] ,
    \ccon_0_io_dsi_in[1] ,
    \ccon_0_io_dsi_in[0] }),
    .io_in({io_in[37],
    io_in[36],
    io_in[35],
    io_in[34],
    io_in[33],
    io_in[32],
    io_in[31],
    io_in[30],
    io_in[29],
    io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24],
    io_in[23],
    io_in[22],
    io_in[21],
    io_in[20],
    io_in[19],
    io_in[18],
    io_in[17],
    io_in[16],
    io_in[15],
    io_in[14],
    io_in[13],
    io_in[12],
    io_in[11],
    io_in[10],
    io_in[9],
    io_in[8],
    io_in[7],
    io_in[6],
    io_in[5],
    io_in[4],
    io_in[3],
    io_in[2],
    io_in[1],
    io_in[0]}),
    .io_oeb({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21],
    io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13],
    io_oeb[12],
    io_oeb[11],
    io_oeb[10],
    io_oeb[9],
    io_oeb[8],
    io_oeb[7],
    io_oeb[6],
    io_oeb[5],
    io_oeb[4],
    io_oeb[3],
    io_oeb[2],
    io_oeb[1],
    io_oeb[0]}),
    .io_out({io_out[37],
    io_out[36],
    io_out[35],
    io_out[34],
    io_out[33],
    io_out[32],
    io_out[31],
    io_out[30],
    io_out[29],
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24],
    io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16],
    io_out[15],
    io_out[14],
    io_out[13],
    io_out[12],
    io_out[11],
    io_out[10],
    io_out[9],
    io_out[8],
    io_out[7],
    io_out[6],
    io_out[5],
    io_out[4],
    io_out[3],
    io_out[2],
    io_out[1],
    io_out[0]}),
    .irq({user_irq[2],
    user_irq[1],
    user_irq[0]}),
    .m_irqs({\_T_183[5] ,
    \_T_183[4] ,
    \_T_183[3] ,
    \_T_183[2] ,
    \_T_183[1] ,
    \_T_183[0] ,
    \_T_178[5] ,
    \_T_178[4] ,
    \_T_178[3] ,
    \_T_178[2] ,
    \_T_178[1] ,
    \_T_178[0] }),
    .m_wbs_ack_o({\_T_172[5] ,
    \_T_172[4] ,
    \_T_172[3] ,
    \_T_172[2] ,
    \_T_172[1] ,
    \_T_172[0] ,
    \_T_167[5] ,
    \_T_167[4] ,
    \_T_167[3] ,
    \_T_167[2] ,
    \_T_167[1] ,
    \_T_167[0] }),
    .m_wbs_adr_i({\ccon_0_io_adr_i[11] ,
    \ccon_0_io_adr_i[10] ,
    \ccon_0_io_adr_i[9] ,
    \ccon_0_io_adr_i[8] ,
    \ccon_0_io_adr_i[7] ,
    \ccon_0_io_adr_i[6] ,
    \ccon_0_io_adr_i[5] ,
    \ccon_0_io_adr_i[4] ,
    \ccon_0_io_adr_i[3] ,
    \ccon_0_io_adr_i[2] ,
    \ccon_0_io_adr_i[1] ,
    \ccon_0_io_adr_i[0] }),
    .m_wbs_cs_i({ccon_7_io_cs_i,
    ccon_6_io_cs_i,
    ccon_5_io_cs_i,
    ccon_4_io_cs_i,
    ccon_3_io_cs_i,
    ccon_2_io_cs_i,
    ccon_1_io_cs_i,
    ccon_0_io_cs_i,
    \icon_m_wbs_cs_i[3] ,
    \icon_m_wbs_cs_i[2] ,
    \icon_m_wbs_cs_i[1] ,
    \icon_m_wbs_cs_i[0] }),
    .m_wbs_dat_i({\ccon_0_io_dat_i[31] ,
    \ccon_0_io_dat_i[30] ,
    \ccon_0_io_dat_i[29] ,
    \ccon_0_io_dat_i[28] ,
    \ccon_0_io_dat_i[27] ,
    \ccon_0_io_dat_i[26] ,
    \ccon_0_io_dat_i[25] ,
    \ccon_0_io_dat_i[24] ,
    \ccon_0_io_dat_i[23] ,
    \ccon_0_io_dat_i[22] ,
    \ccon_0_io_dat_i[21] ,
    \ccon_0_io_dat_i[20] ,
    \ccon_0_io_dat_i[19] ,
    \ccon_0_io_dat_i[18] ,
    \ccon_0_io_dat_i[17] ,
    \ccon_0_io_dat_i[16] ,
    \ccon_0_io_dat_i[15] ,
    \ccon_0_io_dat_i[14] ,
    \ccon_0_io_dat_i[13] ,
    \ccon_0_io_dat_i[12] ,
    \ccon_0_io_dat_i[11] ,
    \ccon_0_io_dat_i[10] ,
    \ccon_0_io_dat_i[9] ,
    \ccon_0_io_dat_i[8] ,
    \ccon_0_io_dat_i[7] ,
    \ccon_0_io_dat_i[6] ,
    \ccon_0_io_dat_i[5] ,
    \ccon_0_io_dat_i[4] ,
    \ccon_0_io_dat_i[3] ,
    \ccon_0_io_dat_i[2] ,
    \ccon_0_io_dat_i[1] ,
    \ccon_0_io_dat_i[0] }),
    .m_wbs_dat_o_0({\icon_m_wbs_dat_o_0[31] ,
    \icon_m_wbs_dat_o_0[30] ,
    \icon_m_wbs_dat_o_0[29] ,
    \icon_m_wbs_dat_o_0[28] ,
    \icon_m_wbs_dat_o_0[27] ,
    \icon_m_wbs_dat_o_0[26] ,
    \icon_m_wbs_dat_o_0[25] ,
    \icon_m_wbs_dat_o_0[24] ,
    \icon_m_wbs_dat_o_0[23] ,
    \icon_m_wbs_dat_o_0[22] ,
    \icon_m_wbs_dat_o_0[21] ,
    \icon_m_wbs_dat_o_0[20] ,
    \icon_m_wbs_dat_o_0[19] ,
    \icon_m_wbs_dat_o_0[18] ,
    \icon_m_wbs_dat_o_0[17] ,
    \icon_m_wbs_dat_o_0[16] ,
    \icon_m_wbs_dat_o_0[15] ,
    \icon_m_wbs_dat_o_0[14] ,
    \icon_m_wbs_dat_o_0[13] ,
    \icon_m_wbs_dat_o_0[12] ,
    \icon_m_wbs_dat_o_0[11] ,
    \icon_m_wbs_dat_o_0[10] ,
    \icon_m_wbs_dat_o_0[9] ,
    \icon_m_wbs_dat_o_0[8] ,
    \icon_m_wbs_dat_o_0[7] ,
    \icon_m_wbs_dat_o_0[6] ,
    \icon_m_wbs_dat_o_0[5] ,
    \icon_m_wbs_dat_o_0[4] ,
    \icon_m_wbs_dat_o_0[3] ,
    \icon_m_wbs_dat_o_0[2] ,
    \icon_m_wbs_dat_o_0[1] ,
    \icon_m_wbs_dat_o_0[0] }),
    .m_wbs_dat_o_1({\icon_m_wbs_dat_o_1[31] ,
    \icon_m_wbs_dat_o_1[30] ,
    \icon_m_wbs_dat_o_1[29] ,
    \icon_m_wbs_dat_o_1[28] ,
    \icon_m_wbs_dat_o_1[27] ,
    \icon_m_wbs_dat_o_1[26] ,
    \icon_m_wbs_dat_o_1[25] ,
    \icon_m_wbs_dat_o_1[24] ,
    \icon_m_wbs_dat_o_1[23] ,
    \icon_m_wbs_dat_o_1[22] ,
    \icon_m_wbs_dat_o_1[21] ,
    \icon_m_wbs_dat_o_1[20] ,
    \icon_m_wbs_dat_o_1[19] ,
    \icon_m_wbs_dat_o_1[18] ,
    \icon_m_wbs_dat_o_1[17] ,
    \icon_m_wbs_dat_o_1[16] ,
    \icon_m_wbs_dat_o_1[15] ,
    \icon_m_wbs_dat_o_1[14] ,
    \icon_m_wbs_dat_o_1[13] ,
    \icon_m_wbs_dat_o_1[12] ,
    \icon_m_wbs_dat_o_1[11] ,
    \icon_m_wbs_dat_o_1[10] ,
    \icon_m_wbs_dat_o_1[9] ,
    \icon_m_wbs_dat_o_1[8] ,
    \icon_m_wbs_dat_o_1[7] ,
    \icon_m_wbs_dat_o_1[6] ,
    \icon_m_wbs_dat_o_1[5] ,
    \icon_m_wbs_dat_o_1[4] ,
    \icon_m_wbs_dat_o_1[3] ,
    \icon_m_wbs_dat_o_1[2] ,
    \icon_m_wbs_dat_o_1[1] ,
    \icon_m_wbs_dat_o_1[0] }),
    .m_wbs_dat_o_10({\ccon_6_io_dat_o[31] ,
    \ccon_6_io_dat_o[30] ,
    \ccon_6_io_dat_o[29] ,
    \ccon_6_io_dat_o[28] ,
    \ccon_6_io_dat_o[27] ,
    \ccon_6_io_dat_o[26] ,
    \ccon_6_io_dat_o[25] ,
    \ccon_6_io_dat_o[24] ,
    \ccon_6_io_dat_o[23] ,
    \ccon_6_io_dat_o[22] ,
    \ccon_6_io_dat_o[21] ,
    \ccon_6_io_dat_o[20] ,
    \ccon_6_io_dat_o[19] ,
    \ccon_6_io_dat_o[18] ,
    \ccon_6_io_dat_o[17] ,
    \ccon_6_io_dat_o[16] ,
    \ccon_6_io_dat_o[15] ,
    \ccon_6_io_dat_o[14] ,
    \ccon_6_io_dat_o[13] ,
    \ccon_6_io_dat_o[12] ,
    \ccon_6_io_dat_o[11] ,
    \ccon_6_io_dat_o[10] ,
    \ccon_6_io_dat_o[9] ,
    \ccon_6_io_dat_o[8] ,
    \ccon_6_io_dat_o[7] ,
    \ccon_6_io_dat_o[6] ,
    \ccon_6_io_dat_o[5] ,
    \ccon_6_io_dat_o[4] ,
    \ccon_6_io_dat_o[3] ,
    \ccon_6_io_dat_o[2] ,
    \ccon_6_io_dat_o[1] ,
    \ccon_6_io_dat_o[0] }),
    .m_wbs_dat_o_11({\ccon_7_io_dat_o[31] ,
    \ccon_7_io_dat_o[30] ,
    \ccon_7_io_dat_o[29] ,
    \ccon_7_io_dat_o[28] ,
    \ccon_7_io_dat_o[27] ,
    \ccon_7_io_dat_o[26] ,
    \ccon_7_io_dat_o[25] ,
    \ccon_7_io_dat_o[24] ,
    \ccon_7_io_dat_o[23] ,
    \ccon_7_io_dat_o[22] ,
    \ccon_7_io_dat_o[21] ,
    \ccon_7_io_dat_o[20] ,
    \ccon_7_io_dat_o[19] ,
    \ccon_7_io_dat_o[18] ,
    \ccon_7_io_dat_o[17] ,
    \ccon_7_io_dat_o[16] ,
    \ccon_7_io_dat_o[15] ,
    \ccon_7_io_dat_o[14] ,
    \ccon_7_io_dat_o[13] ,
    \ccon_7_io_dat_o[12] ,
    \ccon_7_io_dat_o[11] ,
    \ccon_7_io_dat_o[10] ,
    \ccon_7_io_dat_o[9] ,
    \ccon_7_io_dat_o[8] ,
    \ccon_7_io_dat_o[7] ,
    \ccon_7_io_dat_o[6] ,
    \ccon_7_io_dat_o[5] ,
    \ccon_7_io_dat_o[4] ,
    \ccon_7_io_dat_o[3] ,
    \ccon_7_io_dat_o[2] ,
    \ccon_7_io_dat_o[1] ,
    \ccon_7_io_dat_o[0] }),
    .m_wbs_dat_o_2({\icon_m_wbs_dat_o_2[31] ,
    \icon_m_wbs_dat_o_2[30] ,
    \icon_m_wbs_dat_o_2[29] ,
    \icon_m_wbs_dat_o_2[28] ,
    \icon_m_wbs_dat_o_2[27] ,
    \icon_m_wbs_dat_o_2[26] ,
    \icon_m_wbs_dat_o_2[25] ,
    \icon_m_wbs_dat_o_2[24] ,
    \icon_m_wbs_dat_o_2[23] ,
    \icon_m_wbs_dat_o_2[22] ,
    \icon_m_wbs_dat_o_2[21] ,
    \icon_m_wbs_dat_o_2[20] ,
    \icon_m_wbs_dat_o_2[19] ,
    \icon_m_wbs_dat_o_2[18] ,
    \icon_m_wbs_dat_o_2[17] ,
    \icon_m_wbs_dat_o_2[16] ,
    \icon_m_wbs_dat_o_2[15] ,
    \icon_m_wbs_dat_o_2[14] ,
    \icon_m_wbs_dat_o_2[13] ,
    \icon_m_wbs_dat_o_2[12] ,
    \icon_m_wbs_dat_o_2[11] ,
    \icon_m_wbs_dat_o_2[10] ,
    \icon_m_wbs_dat_o_2[9] ,
    \icon_m_wbs_dat_o_2[8] ,
    \icon_m_wbs_dat_o_2[7] ,
    \icon_m_wbs_dat_o_2[6] ,
    \icon_m_wbs_dat_o_2[5] ,
    \icon_m_wbs_dat_o_2[4] ,
    \icon_m_wbs_dat_o_2[3] ,
    \icon_m_wbs_dat_o_2[2] ,
    \icon_m_wbs_dat_o_2[1] ,
    \icon_m_wbs_dat_o_2[0] }),
    .m_wbs_dat_o_3({\icon_m_wbs_dat_o_3[31] ,
    \icon_m_wbs_dat_o_3[30] ,
    \icon_m_wbs_dat_o_3[29] ,
    \icon_m_wbs_dat_o_3[28] ,
    \icon_m_wbs_dat_o_3[27] ,
    \icon_m_wbs_dat_o_3[26] ,
    \icon_m_wbs_dat_o_3[25] ,
    \icon_m_wbs_dat_o_3[24] ,
    \icon_m_wbs_dat_o_3[23] ,
    \icon_m_wbs_dat_o_3[22] ,
    \icon_m_wbs_dat_o_3[21] ,
    \icon_m_wbs_dat_o_3[20] ,
    \icon_m_wbs_dat_o_3[19] ,
    \icon_m_wbs_dat_o_3[18] ,
    \icon_m_wbs_dat_o_3[17] ,
    \icon_m_wbs_dat_o_3[16] ,
    \icon_m_wbs_dat_o_3[15] ,
    \icon_m_wbs_dat_o_3[14] ,
    \icon_m_wbs_dat_o_3[13] ,
    \icon_m_wbs_dat_o_3[12] ,
    \icon_m_wbs_dat_o_3[11] ,
    \icon_m_wbs_dat_o_3[10] ,
    \icon_m_wbs_dat_o_3[9] ,
    \icon_m_wbs_dat_o_3[8] ,
    \icon_m_wbs_dat_o_3[7] ,
    \icon_m_wbs_dat_o_3[6] ,
    \icon_m_wbs_dat_o_3[5] ,
    \icon_m_wbs_dat_o_3[4] ,
    \icon_m_wbs_dat_o_3[3] ,
    \icon_m_wbs_dat_o_3[2] ,
    \icon_m_wbs_dat_o_3[1] ,
    \icon_m_wbs_dat_o_3[0] }),
    .m_wbs_dat_o_4({\ccon_0_io_dat_o[31] ,
    \ccon_0_io_dat_o[30] ,
    \ccon_0_io_dat_o[29] ,
    \ccon_0_io_dat_o[28] ,
    \ccon_0_io_dat_o[27] ,
    \ccon_0_io_dat_o[26] ,
    \ccon_0_io_dat_o[25] ,
    \ccon_0_io_dat_o[24] ,
    \ccon_0_io_dat_o[23] ,
    \ccon_0_io_dat_o[22] ,
    \ccon_0_io_dat_o[21] ,
    \ccon_0_io_dat_o[20] ,
    \ccon_0_io_dat_o[19] ,
    \ccon_0_io_dat_o[18] ,
    \ccon_0_io_dat_o[17] ,
    \ccon_0_io_dat_o[16] ,
    \ccon_0_io_dat_o[15] ,
    \ccon_0_io_dat_o[14] ,
    \ccon_0_io_dat_o[13] ,
    \ccon_0_io_dat_o[12] ,
    \ccon_0_io_dat_o[11] ,
    \ccon_0_io_dat_o[10] ,
    \ccon_0_io_dat_o[9] ,
    \ccon_0_io_dat_o[8] ,
    \ccon_0_io_dat_o[7] ,
    \ccon_0_io_dat_o[6] ,
    \ccon_0_io_dat_o[5] ,
    \ccon_0_io_dat_o[4] ,
    \ccon_0_io_dat_o[3] ,
    \ccon_0_io_dat_o[2] ,
    \ccon_0_io_dat_o[1] ,
    \ccon_0_io_dat_o[0] }),
    .m_wbs_dat_o_5({\ccon_1_io_dat_o[31] ,
    \ccon_1_io_dat_o[30] ,
    \ccon_1_io_dat_o[29] ,
    \ccon_1_io_dat_o[28] ,
    \ccon_1_io_dat_o[27] ,
    \ccon_1_io_dat_o[26] ,
    \ccon_1_io_dat_o[25] ,
    \ccon_1_io_dat_o[24] ,
    \ccon_1_io_dat_o[23] ,
    \ccon_1_io_dat_o[22] ,
    \ccon_1_io_dat_o[21] ,
    \ccon_1_io_dat_o[20] ,
    \ccon_1_io_dat_o[19] ,
    \ccon_1_io_dat_o[18] ,
    \ccon_1_io_dat_o[17] ,
    \ccon_1_io_dat_o[16] ,
    \ccon_1_io_dat_o[15] ,
    \ccon_1_io_dat_o[14] ,
    \ccon_1_io_dat_o[13] ,
    \ccon_1_io_dat_o[12] ,
    \ccon_1_io_dat_o[11] ,
    \ccon_1_io_dat_o[10] ,
    \ccon_1_io_dat_o[9] ,
    \ccon_1_io_dat_o[8] ,
    \ccon_1_io_dat_o[7] ,
    \ccon_1_io_dat_o[6] ,
    \ccon_1_io_dat_o[5] ,
    \ccon_1_io_dat_o[4] ,
    \ccon_1_io_dat_o[3] ,
    \ccon_1_io_dat_o[2] ,
    \ccon_1_io_dat_o[1] ,
    \ccon_1_io_dat_o[0] }),
    .m_wbs_dat_o_6({\ccon_2_io_dat_o[31] ,
    \ccon_2_io_dat_o[30] ,
    \ccon_2_io_dat_o[29] ,
    \ccon_2_io_dat_o[28] ,
    \ccon_2_io_dat_o[27] ,
    \ccon_2_io_dat_o[26] ,
    \ccon_2_io_dat_o[25] ,
    \ccon_2_io_dat_o[24] ,
    \ccon_2_io_dat_o[23] ,
    \ccon_2_io_dat_o[22] ,
    \ccon_2_io_dat_o[21] ,
    \ccon_2_io_dat_o[20] ,
    \ccon_2_io_dat_o[19] ,
    \ccon_2_io_dat_o[18] ,
    \ccon_2_io_dat_o[17] ,
    \ccon_2_io_dat_o[16] ,
    \ccon_2_io_dat_o[15] ,
    \ccon_2_io_dat_o[14] ,
    \ccon_2_io_dat_o[13] ,
    \ccon_2_io_dat_o[12] ,
    \ccon_2_io_dat_o[11] ,
    \ccon_2_io_dat_o[10] ,
    \ccon_2_io_dat_o[9] ,
    \ccon_2_io_dat_o[8] ,
    \ccon_2_io_dat_o[7] ,
    \ccon_2_io_dat_o[6] ,
    \ccon_2_io_dat_o[5] ,
    \ccon_2_io_dat_o[4] ,
    \ccon_2_io_dat_o[3] ,
    \ccon_2_io_dat_o[2] ,
    \ccon_2_io_dat_o[1] ,
    \ccon_2_io_dat_o[0] }),
    .m_wbs_dat_o_7({\ccon_3_io_dat_o[31] ,
    \ccon_3_io_dat_o[30] ,
    \ccon_3_io_dat_o[29] ,
    \ccon_3_io_dat_o[28] ,
    \ccon_3_io_dat_o[27] ,
    \ccon_3_io_dat_o[26] ,
    \ccon_3_io_dat_o[25] ,
    \ccon_3_io_dat_o[24] ,
    \ccon_3_io_dat_o[23] ,
    \ccon_3_io_dat_o[22] ,
    \ccon_3_io_dat_o[21] ,
    \ccon_3_io_dat_o[20] ,
    \ccon_3_io_dat_o[19] ,
    \ccon_3_io_dat_o[18] ,
    \ccon_3_io_dat_o[17] ,
    \ccon_3_io_dat_o[16] ,
    \ccon_3_io_dat_o[15] ,
    \ccon_3_io_dat_o[14] ,
    \ccon_3_io_dat_o[13] ,
    \ccon_3_io_dat_o[12] ,
    \ccon_3_io_dat_o[11] ,
    \ccon_3_io_dat_o[10] ,
    \ccon_3_io_dat_o[9] ,
    \ccon_3_io_dat_o[8] ,
    \ccon_3_io_dat_o[7] ,
    \ccon_3_io_dat_o[6] ,
    \ccon_3_io_dat_o[5] ,
    \ccon_3_io_dat_o[4] ,
    \ccon_3_io_dat_o[3] ,
    \ccon_3_io_dat_o[2] ,
    \ccon_3_io_dat_o[1] ,
    \ccon_3_io_dat_o[0] }),
    .m_wbs_dat_o_8({\ccon_4_io_dat_o[31] ,
    \ccon_4_io_dat_o[30] ,
    \ccon_4_io_dat_o[29] ,
    \ccon_4_io_dat_o[28] ,
    \ccon_4_io_dat_o[27] ,
    \ccon_4_io_dat_o[26] ,
    \ccon_4_io_dat_o[25] ,
    \ccon_4_io_dat_o[24] ,
    \ccon_4_io_dat_o[23] ,
    \ccon_4_io_dat_o[22] ,
    \ccon_4_io_dat_o[21] ,
    \ccon_4_io_dat_o[20] ,
    \ccon_4_io_dat_o[19] ,
    \ccon_4_io_dat_o[18] ,
    \ccon_4_io_dat_o[17] ,
    \ccon_4_io_dat_o[16] ,
    \ccon_4_io_dat_o[15] ,
    \ccon_4_io_dat_o[14] ,
    \ccon_4_io_dat_o[13] ,
    \ccon_4_io_dat_o[12] ,
    \ccon_4_io_dat_o[11] ,
    \ccon_4_io_dat_o[10] ,
    \ccon_4_io_dat_o[9] ,
    \ccon_4_io_dat_o[8] ,
    \ccon_4_io_dat_o[7] ,
    \ccon_4_io_dat_o[6] ,
    \ccon_4_io_dat_o[5] ,
    \ccon_4_io_dat_o[4] ,
    \ccon_4_io_dat_o[3] ,
    \ccon_4_io_dat_o[2] ,
    \ccon_4_io_dat_o[1] ,
    \ccon_4_io_dat_o[0] }),
    .m_wbs_dat_o_9({\ccon_5_io_dat_o[31] ,
    \ccon_5_io_dat_o[30] ,
    \ccon_5_io_dat_o[29] ,
    \ccon_5_io_dat_o[28] ,
    \ccon_5_io_dat_o[27] ,
    \ccon_5_io_dat_o[26] ,
    \ccon_5_io_dat_o[25] ,
    \ccon_5_io_dat_o[24] ,
    \ccon_5_io_dat_o[23] ,
    \ccon_5_io_dat_o[22] ,
    \ccon_5_io_dat_o[21] ,
    \ccon_5_io_dat_o[20] ,
    \ccon_5_io_dat_o[19] ,
    \ccon_5_io_dat_o[18] ,
    \ccon_5_io_dat_o[17] ,
    \ccon_5_io_dat_o[16] ,
    \ccon_5_io_dat_o[15] ,
    \ccon_5_io_dat_o[14] ,
    \ccon_5_io_dat_o[13] ,
    \ccon_5_io_dat_o[12] ,
    \ccon_5_io_dat_o[11] ,
    \ccon_5_io_dat_o[10] ,
    \ccon_5_io_dat_o[9] ,
    \ccon_5_io_dat_o[8] ,
    \ccon_5_io_dat_o[7] ,
    \ccon_5_io_dat_o[6] ,
    \ccon_5_io_dat_o[5] ,
    \ccon_5_io_dat_o[4] ,
    \ccon_5_io_dat_o[3] ,
    \ccon_5_io_dat_o[2] ,
    \ccon_5_io_dat_o[1] ,
    \ccon_5_io_dat_o[0] }),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({wbs_dat_o[31],
    wbs_dat_o[30],
    wbs_dat_o[29],
    wbs_dat_o[28],
    wbs_dat_o[27],
    wbs_dat_o[26],
    wbs_dat_o[25],
    wbs_dat_o[24],
    wbs_dat_o[23],
    wbs_dat_o[22],
    wbs_dat_o[21],
    wbs_dat_o[20],
    wbs_dat_o[19],
    wbs_dat_o[18],
    wbs_dat_o[17],
    wbs_dat_o[16],
    wbs_dat_o[15],
    wbs_dat_o[14],
    wbs_dat_o[13],
    wbs_dat_o[12],
    wbs_dat_o[11],
    wbs_dat_o[10],
    wbs_dat_o[9],
    wbs_dat_o[8],
    wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 motor_top mcons_0 (.clock(cb_0_0_wb_clk_i),
    .io_QEI_ChA(icon_mt_QEI_ChA_0),
    .io_QEI_ChB(icon_mt_QEI_ChB_0),
    .io_irq(\_T_178[0] ),
    .io_pwm_h(icon_mt_pwm_h_0),
    .io_pwm_l(icon_mt_pwm_l_0),
    .io_wb_ack_o(\_T_167[0] ),
    .io_wb_cs_i(\icon_m_wbs_cs_i[0] ),
    .io_wb_we_i(ccon_0_io_we_i),
    .reset(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_wb_adr_i({\ccon_0_io_adr_i[11] ,
    \ccon_0_io_adr_i[10] ,
    \ccon_0_io_adr_i[9] ,
    \ccon_0_io_adr_i[8] ,
    \ccon_0_io_adr_i[7] ,
    \ccon_0_io_adr_i[6] ,
    \ccon_0_io_adr_i[5] ,
    \ccon_0_io_adr_i[4] ,
    \ccon_0_io_adr_i[3] ,
    \ccon_0_io_adr_i[2] ,
    \ccon_0_io_adr_i[1] ,
    \ccon_0_io_adr_i[0] }),
    .io_wb_dat_i({\ccon_0_io_dat_i[31] ,
    \ccon_0_io_dat_i[30] ,
    \ccon_0_io_dat_i[29] ,
    \ccon_0_io_dat_i[28] ,
    \ccon_0_io_dat_i[27] ,
    \ccon_0_io_dat_i[26] ,
    \ccon_0_io_dat_i[25] ,
    \ccon_0_io_dat_i[24] ,
    \ccon_0_io_dat_i[23] ,
    \ccon_0_io_dat_i[22] ,
    \ccon_0_io_dat_i[21] ,
    \ccon_0_io_dat_i[20] ,
    \ccon_0_io_dat_i[19] ,
    \ccon_0_io_dat_i[18] ,
    \ccon_0_io_dat_i[17] ,
    \ccon_0_io_dat_i[16] ,
    \ccon_0_io_dat_i[15] ,
    \ccon_0_io_dat_i[14] ,
    \ccon_0_io_dat_i[13] ,
    \ccon_0_io_dat_i[12] ,
    \ccon_0_io_dat_i[11] ,
    \ccon_0_io_dat_i[10] ,
    \ccon_0_io_dat_i[9] ,
    \ccon_0_io_dat_i[8] ,
    \ccon_0_io_dat_i[7] ,
    \ccon_0_io_dat_i[6] ,
    \ccon_0_io_dat_i[5] ,
    \ccon_0_io_dat_i[4] ,
    \ccon_0_io_dat_i[3] ,
    \ccon_0_io_dat_i[2] ,
    \ccon_0_io_dat_i[1] ,
    \ccon_0_io_dat_i[0] }),
    .io_wb_dat_o({\icon_m_wbs_dat_o_0[31] ,
    \icon_m_wbs_dat_o_0[30] ,
    \icon_m_wbs_dat_o_0[29] ,
    \icon_m_wbs_dat_o_0[28] ,
    \icon_m_wbs_dat_o_0[27] ,
    \icon_m_wbs_dat_o_0[26] ,
    \icon_m_wbs_dat_o_0[25] ,
    \icon_m_wbs_dat_o_0[24] ,
    \icon_m_wbs_dat_o_0[23] ,
    \icon_m_wbs_dat_o_0[22] ,
    \icon_m_wbs_dat_o_0[21] ,
    \icon_m_wbs_dat_o_0[20] ,
    \icon_m_wbs_dat_o_0[19] ,
    \icon_m_wbs_dat_o_0[18] ,
    \icon_m_wbs_dat_o_0[17] ,
    \icon_m_wbs_dat_o_0[16] ,
    \icon_m_wbs_dat_o_0[15] ,
    \icon_m_wbs_dat_o_0[14] ,
    \icon_m_wbs_dat_o_0[13] ,
    \icon_m_wbs_dat_o_0[12] ,
    \icon_m_wbs_dat_o_0[11] ,
    \icon_m_wbs_dat_o_0[10] ,
    \icon_m_wbs_dat_o_0[9] ,
    \icon_m_wbs_dat_o_0[8] ,
    \icon_m_wbs_dat_o_0[7] ,
    \icon_m_wbs_dat_o_0[6] ,
    \icon_m_wbs_dat_o_0[5] ,
    \icon_m_wbs_dat_o_0[4] ,
    \icon_m_wbs_dat_o_0[3] ,
    \icon_m_wbs_dat_o_0[2] ,
    \icon_m_wbs_dat_o_0[1] ,
    \icon_m_wbs_dat_o_0[0] }));
 motor_top mcons_1 (.clock(cb_0_0_wb_clk_i),
    .io_QEI_ChA(icon_mt_QEI_ChA_1),
    .io_QEI_ChB(icon_mt_QEI_ChB_1),
    .io_irq(\_T_178[1] ),
    .io_pwm_h(icon_mt_pwm_h_1),
    .io_pwm_l(icon_mt_pwm_l_1),
    .io_wb_ack_o(\_T_167[1] ),
    .io_wb_cs_i(\icon_m_wbs_cs_i[1] ),
    .io_wb_we_i(ccon_0_io_we_i),
    .reset(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_wb_adr_i({\ccon_0_io_adr_i[11] ,
    \ccon_0_io_adr_i[10] ,
    \ccon_0_io_adr_i[9] ,
    \ccon_0_io_adr_i[8] ,
    \ccon_0_io_adr_i[7] ,
    \ccon_0_io_adr_i[6] ,
    \ccon_0_io_adr_i[5] ,
    \ccon_0_io_adr_i[4] ,
    \ccon_0_io_adr_i[3] ,
    \ccon_0_io_adr_i[2] ,
    \ccon_0_io_adr_i[1] ,
    \ccon_0_io_adr_i[0] }),
    .io_wb_dat_i({\ccon_0_io_dat_i[31] ,
    \ccon_0_io_dat_i[30] ,
    \ccon_0_io_dat_i[29] ,
    \ccon_0_io_dat_i[28] ,
    \ccon_0_io_dat_i[27] ,
    \ccon_0_io_dat_i[26] ,
    \ccon_0_io_dat_i[25] ,
    \ccon_0_io_dat_i[24] ,
    \ccon_0_io_dat_i[23] ,
    \ccon_0_io_dat_i[22] ,
    \ccon_0_io_dat_i[21] ,
    \ccon_0_io_dat_i[20] ,
    \ccon_0_io_dat_i[19] ,
    \ccon_0_io_dat_i[18] ,
    \ccon_0_io_dat_i[17] ,
    \ccon_0_io_dat_i[16] ,
    \ccon_0_io_dat_i[15] ,
    \ccon_0_io_dat_i[14] ,
    \ccon_0_io_dat_i[13] ,
    \ccon_0_io_dat_i[12] ,
    \ccon_0_io_dat_i[11] ,
    \ccon_0_io_dat_i[10] ,
    \ccon_0_io_dat_i[9] ,
    \ccon_0_io_dat_i[8] ,
    \ccon_0_io_dat_i[7] ,
    \ccon_0_io_dat_i[6] ,
    \ccon_0_io_dat_i[5] ,
    \ccon_0_io_dat_i[4] ,
    \ccon_0_io_dat_i[3] ,
    \ccon_0_io_dat_i[2] ,
    \ccon_0_io_dat_i[1] ,
    \ccon_0_io_dat_i[0] }),
    .io_wb_dat_o({\icon_m_wbs_dat_o_1[31] ,
    \icon_m_wbs_dat_o_1[30] ,
    \icon_m_wbs_dat_o_1[29] ,
    \icon_m_wbs_dat_o_1[28] ,
    \icon_m_wbs_dat_o_1[27] ,
    \icon_m_wbs_dat_o_1[26] ,
    \icon_m_wbs_dat_o_1[25] ,
    \icon_m_wbs_dat_o_1[24] ,
    \icon_m_wbs_dat_o_1[23] ,
    \icon_m_wbs_dat_o_1[22] ,
    \icon_m_wbs_dat_o_1[21] ,
    \icon_m_wbs_dat_o_1[20] ,
    \icon_m_wbs_dat_o_1[19] ,
    \icon_m_wbs_dat_o_1[18] ,
    \icon_m_wbs_dat_o_1[17] ,
    \icon_m_wbs_dat_o_1[16] ,
    \icon_m_wbs_dat_o_1[15] ,
    \icon_m_wbs_dat_o_1[14] ,
    \icon_m_wbs_dat_o_1[13] ,
    \icon_m_wbs_dat_o_1[12] ,
    \icon_m_wbs_dat_o_1[11] ,
    \icon_m_wbs_dat_o_1[10] ,
    \icon_m_wbs_dat_o_1[9] ,
    \icon_m_wbs_dat_o_1[8] ,
    \icon_m_wbs_dat_o_1[7] ,
    \icon_m_wbs_dat_o_1[6] ,
    \icon_m_wbs_dat_o_1[5] ,
    \icon_m_wbs_dat_o_1[4] ,
    \icon_m_wbs_dat_o_1[3] ,
    \icon_m_wbs_dat_o_1[2] ,
    \icon_m_wbs_dat_o_1[1] ,
    \icon_m_wbs_dat_o_1[0] }));
 motor_top mcons_2 (.clock(cb_0_0_wb_clk_i),
    .io_QEI_ChA(icon_mt_QEI_ChA_2),
    .io_QEI_ChB(icon_mt_QEI_ChB_2),
    .io_irq(\_T_178[2] ),
    .io_pwm_h(icon_mt_pwm_h_2),
    .io_pwm_l(icon_mt_pwm_l_2),
    .io_wb_ack_o(\_T_167[2] ),
    .io_wb_cs_i(\icon_m_wbs_cs_i[2] ),
    .io_wb_we_i(ccon_0_io_we_i),
    .reset(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_wb_adr_i({\ccon_0_io_adr_i[11] ,
    \ccon_0_io_adr_i[10] ,
    \ccon_0_io_adr_i[9] ,
    \ccon_0_io_adr_i[8] ,
    \ccon_0_io_adr_i[7] ,
    \ccon_0_io_adr_i[6] ,
    \ccon_0_io_adr_i[5] ,
    \ccon_0_io_adr_i[4] ,
    \ccon_0_io_adr_i[3] ,
    \ccon_0_io_adr_i[2] ,
    \ccon_0_io_adr_i[1] ,
    \ccon_0_io_adr_i[0] }),
    .io_wb_dat_i({\ccon_0_io_dat_i[31] ,
    \ccon_0_io_dat_i[30] ,
    \ccon_0_io_dat_i[29] ,
    \ccon_0_io_dat_i[28] ,
    \ccon_0_io_dat_i[27] ,
    \ccon_0_io_dat_i[26] ,
    \ccon_0_io_dat_i[25] ,
    \ccon_0_io_dat_i[24] ,
    \ccon_0_io_dat_i[23] ,
    \ccon_0_io_dat_i[22] ,
    \ccon_0_io_dat_i[21] ,
    \ccon_0_io_dat_i[20] ,
    \ccon_0_io_dat_i[19] ,
    \ccon_0_io_dat_i[18] ,
    \ccon_0_io_dat_i[17] ,
    \ccon_0_io_dat_i[16] ,
    \ccon_0_io_dat_i[15] ,
    \ccon_0_io_dat_i[14] ,
    \ccon_0_io_dat_i[13] ,
    \ccon_0_io_dat_i[12] ,
    \ccon_0_io_dat_i[11] ,
    \ccon_0_io_dat_i[10] ,
    \ccon_0_io_dat_i[9] ,
    \ccon_0_io_dat_i[8] ,
    \ccon_0_io_dat_i[7] ,
    \ccon_0_io_dat_i[6] ,
    \ccon_0_io_dat_i[5] ,
    \ccon_0_io_dat_i[4] ,
    \ccon_0_io_dat_i[3] ,
    \ccon_0_io_dat_i[2] ,
    \ccon_0_io_dat_i[1] ,
    \ccon_0_io_dat_i[0] }),
    .io_wb_dat_o({\icon_m_wbs_dat_o_2[31] ,
    \icon_m_wbs_dat_o_2[30] ,
    \icon_m_wbs_dat_o_2[29] ,
    \icon_m_wbs_dat_o_2[28] ,
    \icon_m_wbs_dat_o_2[27] ,
    \icon_m_wbs_dat_o_2[26] ,
    \icon_m_wbs_dat_o_2[25] ,
    \icon_m_wbs_dat_o_2[24] ,
    \icon_m_wbs_dat_o_2[23] ,
    \icon_m_wbs_dat_o_2[22] ,
    \icon_m_wbs_dat_o_2[21] ,
    \icon_m_wbs_dat_o_2[20] ,
    \icon_m_wbs_dat_o_2[19] ,
    \icon_m_wbs_dat_o_2[18] ,
    \icon_m_wbs_dat_o_2[17] ,
    \icon_m_wbs_dat_o_2[16] ,
    \icon_m_wbs_dat_o_2[15] ,
    \icon_m_wbs_dat_o_2[14] ,
    \icon_m_wbs_dat_o_2[13] ,
    \icon_m_wbs_dat_o_2[12] ,
    \icon_m_wbs_dat_o_2[11] ,
    \icon_m_wbs_dat_o_2[10] ,
    \icon_m_wbs_dat_o_2[9] ,
    \icon_m_wbs_dat_o_2[8] ,
    \icon_m_wbs_dat_o_2[7] ,
    \icon_m_wbs_dat_o_2[6] ,
    \icon_m_wbs_dat_o_2[5] ,
    \icon_m_wbs_dat_o_2[4] ,
    \icon_m_wbs_dat_o_2[3] ,
    \icon_m_wbs_dat_o_2[2] ,
    \icon_m_wbs_dat_o_2[1] ,
    \icon_m_wbs_dat_o_2[0] }));
 motor_top mcons_3 (.clock(cb_0_0_wb_clk_i),
    .io_QEI_ChA(icon_mt_QEI_ChA_3),
    .io_QEI_ChB(icon_mt_QEI_ChB_3),
    .io_irq(\_T_178[3] ),
    .io_pwm_h(icon_mt_pwm_h_3),
    .io_pwm_l(icon_mt_pwm_l_3),
    .io_wb_ack_o(\_T_167[3] ),
    .io_wb_cs_i(\icon_m_wbs_cs_i[3] ),
    .io_wb_we_i(ccon_0_io_we_i),
    .reset(cb_0_0_wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_wb_adr_i({\ccon_0_io_adr_i[11] ,
    \ccon_0_io_adr_i[10] ,
    \ccon_0_io_adr_i[9] ,
    \ccon_0_io_adr_i[8] ,
    \ccon_0_io_adr_i[7] ,
    \ccon_0_io_adr_i[6] ,
    \ccon_0_io_adr_i[5] ,
    \ccon_0_io_adr_i[4] ,
    \ccon_0_io_adr_i[3] ,
    \ccon_0_io_adr_i[2] ,
    \ccon_0_io_adr_i[1] ,
    \ccon_0_io_adr_i[0] }),
    .io_wb_dat_i({\ccon_0_io_dat_i[31] ,
    \ccon_0_io_dat_i[30] ,
    \ccon_0_io_dat_i[29] ,
    \ccon_0_io_dat_i[28] ,
    \ccon_0_io_dat_i[27] ,
    \ccon_0_io_dat_i[26] ,
    \ccon_0_io_dat_i[25] ,
    \ccon_0_io_dat_i[24] ,
    \ccon_0_io_dat_i[23] ,
    \ccon_0_io_dat_i[22] ,
    \ccon_0_io_dat_i[21] ,
    \ccon_0_io_dat_i[20] ,
    \ccon_0_io_dat_i[19] ,
    \ccon_0_io_dat_i[18] ,
    \ccon_0_io_dat_i[17] ,
    \ccon_0_io_dat_i[16] ,
    \ccon_0_io_dat_i[15] ,
    \ccon_0_io_dat_i[14] ,
    \ccon_0_io_dat_i[13] ,
    \ccon_0_io_dat_i[12] ,
    \ccon_0_io_dat_i[11] ,
    \ccon_0_io_dat_i[10] ,
    \ccon_0_io_dat_i[9] ,
    \ccon_0_io_dat_i[8] ,
    \ccon_0_io_dat_i[7] ,
    \ccon_0_io_dat_i[6] ,
    \ccon_0_io_dat_i[5] ,
    \ccon_0_io_dat_i[4] ,
    \ccon_0_io_dat_i[3] ,
    \ccon_0_io_dat_i[2] ,
    \ccon_0_io_dat_i[1] ,
    \ccon_0_io_dat_i[0] }),
    .io_wb_dat_o({\icon_m_wbs_dat_o_3[31] ,
    \icon_m_wbs_dat_o_3[30] ,
    \icon_m_wbs_dat_o_3[29] ,
    \icon_m_wbs_dat_o_3[28] ,
    \icon_m_wbs_dat_o_3[27] ,
    \icon_m_wbs_dat_o_3[26] ,
    \icon_m_wbs_dat_o_3[25] ,
    \icon_m_wbs_dat_o_3[24] ,
    \icon_m_wbs_dat_o_3[23] ,
    \icon_m_wbs_dat_o_3[22] ,
    \icon_m_wbs_dat_o_3[21] ,
    \icon_m_wbs_dat_o_3[20] ,
    \icon_m_wbs_dat_o_3[19] ,
    \icon_m_wbs_dat_o_3[18] ,
    \icon_m_wbs_dat_o_3[17] ,
    \icon_m_wbs_dat_o_3[16] ,
    \icon_m_wbs_dat_o_3[15] ,
    \icon_m_wbs_dat_o_3[14] ,
    \icon_m_wbs_dat_o_3[13] ,
    \icon_m_wbs_dat_o_3[12] ,
    \icon_m_wbs_dat_o_3[11] ,
    \icon_m_wbs_dat_o_3[10] ,
    \icon_m_wbs_dat_o_3[9] ,
    \icon_m_wbs_dat_o_3[8] ,
    \icon_m_wbs_dat_o_3[7] ,
    \icon_m_wbs_dat_o_3[6] ,
    \icon_m_wbs_dat_o_3[5] ,
    \icon_m_wbs_dat_o_3[4] ,
    \icon_m_wbs_dat_o_3[3] ,
    \icon_m_wbs_dat_o_3[2] ,
    \icon_m_wbs_dat_o_3[1] ,
    \icon_m_wbs_dat_o_3[0] }));
endmodule
