magic
tech sky130A
magscale 1 2
timestamp 1623893289
<< locali >>
rect 2973 115447 3007 115549
rect 35173 112795 35207 113033
rect 37105 87227 37139 87465
rect 32137 80631 32171 80801
rect 38945 71791 38979 72573
rect 39221 69207 39255 75089
rect 39313 70363 39347 74885
rect 39405 67167 39439 75021
rect 39773 67167 39807 69649
rect 29285 18615 29319 18921
rect 38945 11067 38979 11645
rect 38945 5559 38979 6205
rect 34437 2975 34471 3077
rect 35633 2431 35667 2601
<< viali >>
rect 2697 117385 2731 117419
rect 12449 117385 12483 117419
rect 27261 117385 27295 117419
rect 34989 117385 35023 117419
rect 7205 117317 7239 117351
rect 2053 117249 2087 117283
rect 4537 117249 4571 117283
rect 6009 117249 6043 117283
rect 7941 117249 7975 117283
rect 9873 117249 9907 117283
rect 11345 117249 11379 117283
rect 13277 117249 13311 117283
rect 15209 117249 15243 117283
rect 18613 117249 18647 117283
rect 19349 117249 19383 117283
rect 21281 117249 21315 117283
rect 24685 117249 24719 117283
rect 26617 117249 26651 117283
rect 32689 117249 32723 117283
rect 33885 117249 33919 117283
rect 5273 117181 5307 117215
rect 8493 117181 8527 117215
rect 10609 117181 10643 117215
rect 15945 117181 15979 117215
rect 18429 117181 18463 117215
rect 25881 117181 25915 117215
rect 32505 117181 32539 117215
rect 36369 117181 36403 117215
rect 37197 117181 37231 117215
rect 1869 117113 1903 117147
rect 2605 117113 2639 117147
rect 4353 117113 4387 117147
rect 5089 117113 5123 117147
rect 5825 117113 5859 117147
rect 7021 117113 7055 117147
rect 7757 117113 7791 117147
rect 9689 117113 9723 117147
rect 10425 117113 10459 117147
rect 11161 117113 11195 117147
rect 12357 117113 12391 117147
rect 13093 117113 13127 117147
rect 13829 117113 13863 117147
rect 15025 117113 15059 117147
rect 15761 117113 15795 117147
rect 16497 117113 16531 117147
rect 17693 117113 17727 117147
rect 19165 117113 19199 117147
rect 20361 117113 20395 117147
rect 21097 117113 21131 117147
rect 21833 117113 21867 117147
rect 23029 117113 23063 117147
rect 23765 117113 23799 117147
rect 24501 117113 24535 117147
rect 25697 117113 25731 117147
rect 26433 117113 26467 117147
rect 27169 117113 27203 117147
rect 28365 117113 28399 117147
rect 29101 117113 29135 117147
rect 29837 117113 29871 117147
rect 31033 117113 31067 117147
rect 31769 117113 31803 117147
rect 33701 117113 33735 117147
rect 34897 117113 34931 117147
rect 37473 117113 37507 117147
rect 8585 117045 8619 117079
rect 13921 117045 13955 117079
rect 16589 117045 16623 117079
rect 17785 117045 17819 117079
rect 20453 117045 20487 117079
rect 21925 117045 21959 117079
rect 23121 117045 23155 117079
rect 23857 117045 23891 117079
rect 28457 117045 28491 117079
rect 29193 117045 29227 117079
rect 29929 117045 29963 117079
rect 31125 117045 31159 117079
rect 31861 117045 31895 117079
rect 36461 117045 36495 117079
rect 1961 116841 1995 116875
rect 5181 116841 5215 116875
rect 7021 116841 7055 116875
rect 7757 116841 7791 116875
rect 9229 116841 9263 116875
rect 9965 116841 9999 116875
rect 10701 116841 10735 116875
rect 12265 116841 12299 116875
rect 13737 116841 13771 116875
rect 15209 116841 15243 116875
rect 15945 116841 15979 116875
rect 17509 116841 17543 116875
rect 18245 116841 18279 116875
rect 18981 116841 19015 116875
rect 19717 116841 19751 116875
rect 21189 116841 21223 116875
rect 22753 116841 22787 116875
rect 24225 116841 24259 116875
rect 24961 116841 24995 116875
rect 25697 116841 25731 116875
rect 26433 116841 26467 116875
rect 27997 116841 28031 116875
rect 28733 116841 28767 116875
rect 33609 116841 33643 116875
rect 37289 116841 37323 116875
rect 2789 116773 2823 116807
rect 4537 116773 4571 116807
rect 13093 116773 13127 116807
rect 14565 116773 14599 116807
rect 20545 116773 20579 116807
rect 23581 116773 23615 116807
rect 29561 116773 29595 116807
rect 31401 116773 31435 116807
rect 35173 116773 35207 116807
rect 35909 116773 35943 116807
rect 1869 116705 1903 116739
rect 2605 116705 2639 116739
rect 3341 116705 3375 116739
rect 4353 116705 4387 116739
rect 5089 116705 5123 116739
rect 6929 116705 6963 116739
rect 7665 116705 7699 116739
rect 8401 116705 8435 116739
rect 9137 116705 9171 116739
rect 9873 116705 9907 116739
rect 10609 116705 10643 116739
rect 12173 116705 12207 116739
rect 12909 116705 12943 116739
rect 13645 116705 13679 116739
rect 14381 116705 14415 116739
rect 15117 116705 15151 116739
rect 15853 116705 15887 116739
rect 17417 116705 17451 116739
rect 18153 116705 18187 116739
rect 18889 116705 18923 116739
rect 19625 116705 19659 116739
rect 20361 116705 20395 116739
rect 21097 116705 21131 116739
rect 22661 116705 22695 116739
rect 23397 116705 23431 116739
rect 24133 116705 24167 116739
rect 24869 116705 24903 116739
rect 25605 116705 25639 116739
rect 26341 116705 26375 116739
rect 27905 116705 27939 116739
rect 28641 116705 28675 116739
rect 29377 116705 29411 116739
rect 30481 116705 30515 116739
rect 31217 116705 31251 116739
rect 31953 116705 31987 116739
rect 33517 116705 33551 116739
rect 34253 116705 34287 116739
rect 34989 116705 35023 116739
rect 35725 116705 35759 116739
rect 36369 116705 36403 116739
rect 37197 116705 37231 116739
rect 30665 116569 30699 116603
rect 34437 116569 34471 116603
rect 3433 116501 3467 116535
rect 5917 116501 5951 116535
rect 8493 116501 8527 116535
rect 32045 116501 32079 116535
rect 36553 116501 36587 116535
rect 3249 116297 3283 116331
rect 4445 116297 4479 116331
rect 5181 116297 5215 116331
rect 5825 116297 5859 116331
rect 6561 116297 6595 116331
rect 7297 116297 7331 116331
rect 9689 116297 9723 116331
rect 10885 116297 10919 116331
rect 11621 116297 11655 116331
rect 12265 116297 12299 116331
rect 13553 116297 13587 116331
rect 15025 116297 15059 116331
rect 15761 116297 15795 116331
rect 17877 116297 17911 116331
rect 21281 116297 21315 116331
rect 24041 116297 24075 116331
rect 26893 116297 26927 116331
rect 27629 116297 27663 116331
rect 28457 116297 28491 116331
rect 29193 116297 29227 116331
rect 32689 116297 32723 116331
rect 35909 116297 35943 116331
rect 8125 116229 8159 116263
rect 12909 116229 12943 116263
rect 16589 116229 16623 116263
rect 17233 116229 17267 116263
rect 20177 116229 20211 116263
rect 31309 116229 31343 116263
rect 31677 116229 31711 116263
rect 32505 116229 32539 116263
rect 33701 116229 33735 116263
rect 37105 116229 37139 116263
rect 2053 116161 2087 116195
rect 18521 116161 18555 116195
rect 21833 116161 21867 116195
rect 22477 116161 22511 116195
rect 25237 116161 25271 116195
rect 31401 116161 31435 116195
rect 32376 116161 32410 116195
rect 32597 116161 32631 116195
rect 33572 116161 33606 116195
rect 33793 116161 33827 116195
rect 37749 116161 37783 116195
rect 5733 116093 5767 116127
rect 23121 116093 23155 116127
rect 29101 116093 29135 116127
rect 31180 116093 31214 116127
rect 34805 116093 34839 116127
rect 37565 116093 37599 116127
rect 1869 116025 1903 116059
rect 3157 116025 3191 116059
rect 4353 116025 4387 116059
rect 6469 116025 6503 116059
rect 7205 116025 7239 116059
rect 7941 116025 7975 116059
rect 9597 116025 9631 116059
rect 10793 116025 10827 116059
rect 14933 116025 14967 116059
rect 16405 116025 16439 116059
rect 21189 116025 21223 116059
rect 23949 116025 23983 116059
rect 26801 116025 26835 116059
rect 28365 116025 28399 116059
rect 31033 116025 31067 116059
rect 32229 116025 32263 116059
rect 33425 116025 33459 116059
rect 35817 116025 35851 116059
rect 36921 116025 36955 116059
rect 25881 115957 25915 115991
rect 34069 115957 34103 115991
rect 34621 115957 34655 115991
rect 3249 115753 3283 115787
rect 5365 115753 5399 115787
rect 8125 115753 8159 115787
rect 8677 115753 8711 115787
rect 22569 115753 22603 115787
rect 23581 115753 23615 115787
rect 24961 115753 24995 115787
rect 29929 115753 29963 115787
rect 31217 115753 31251 115787
rect 34345 115753 34379 115787
rect 4721 115685 4755 115719
rect 7297 115685 7331 115719
rect 29101 115685 29135 115719
rect 30757 115685 30791 115719
rect 32137 115685 32171 115719
rect 35909 115685 35943 115719
rect 1869 115617 1903 115651
rect 3157 115617 3191 115651
rect 4537 115617 4571 115651
rect 5273 115617 5307 115651
rect 8033 115617 8067 115651
rect 9505 115617 9539 115651
rect 10149 115617 10183 115651
rect 10793 115617 10827 115651
rect 12265 115617 12299 115651
rect 12909 115617 12943 115651
rect 15301 115617 15335 115651
rect 16037 115617 16071 115651
rect 17509 115617 17543 115651
rect 18153 115617 18187 115651
rect 19441 115617 19475 115651
rect 20177 115617 20211 115651
rect 21557 115617 21591 115651
rect 22753 115617 22787 115651
rect 25145 115617 25179 115651
rect 25881 115617 25915 115651
rect 27997 115617 28031 115651
rect 29837 115617 29871 115651
rect 30573 115617 30607 115651
rect 31401 115617 31435 115651
rect 31953 115617 31987 115651
rect 33517 115617 33551 115651
rect 34253 115617 34287 115651
rect 34989 115617 35023 115651
rect 35725 115617 35759 115651
rect 36461 115617 36495 115651
rect 37197 115617 37231 115651
rect 2973 115549 3007 115583
rect 3985 115549 4019 115583
rect 13921 115549 13955 115583
rect 18797 115549 18831 115583
rect 20913 115549 20947 115583
rect 24317 115549 24351 115583
rect 26341 115549 26375 115583
rect 29285 115549 29319 115583
rect 33701 115549 33735 115583
rect 35173 115549 35207 115583
rect 14657 115481 14691 115515
rect 25697 115481 25731 115515
rect 37381 115481 37415 115515
rect 1961 115413 1995 115447
rect 2973 115413 3007 115447
rect 36553 115413 36587 115447
rect 1961 115209 1995 115243
rect 5733 115209 5767 115243
rect 6377 115209 6411 115243
rect 7021 115209 7055 115243
rect 7665 115209 7699 115243
rect 8309 115209 8343 115243
rect 9689 115209 9723 115243
rect 10333 115209 10367 115243
rect 10977 115209 11011 115243
rect 12817 115209 12851 115243
rect 13461 115209 13495 115243
rect 14933 115209 14967 115243
rect 15577 115209 15611 115243
rect 16313 115209 16347 115243
rect 18337 115209 18371 115243
rect 20177 115209 20211 115243
rect 20821 115209 20855 115243
rect 26249 115209 26283 115243
rect 28089 115209 28123 115243
rect 29193 115209 29227 115243
rect 30665 115209 30699 115243
rect 31309 115209 31343 115243
rect 31953 115209 31987 115243
rect 33977 115209 34011 115243
rect 2789 115141 2823 115175
rect 4445 115141 4479 115175
rect 11437 115141 11471 115175
rect 18797 115141 18831 115175
rect 22753 115141 22787 115175
rect 24133 115141 24167 115175
rect 25237 115141 25271 115175
rect 33333 115141 33367 115175
rect 34805 115141 34839 115175
rect 5089 115073 5123 115107
rect 27353 115073 27387 115107
rect 2605 115005 2639 115039
rect 11621 115005 11655 115039
rect 16957 115005 16991 115039
rect 17601 115005 17635 115039
rect 18981 115005 19015 115039
rect 21465 115005 21499 115039
rect 21925 115005 21959 115039
rect 22937 115005 22971 115039
rect 23673 115005 23707 115039
rect 24317 115005 24351 115039
rect 25429 115005 25463 115039
rect 26433 115005 26467 115039
rect 28733 115005 28767 115039
rect 29377 115005 29411 115039
rect 31493 115005 31527 115039
rect 32137 115005 32171 115039
rect 33885 115005 33919 115039
rect 35725 115005 35759 115039
rect 36185 115005 36219 115039
rect 36553 115005 36587 115039
rect 1869 114937 1903 114971
rect 30573 114937 30607 114971
rect 33149 114937 33183 114971
rect 34621 114937 34655 114971
rect 37933 114937 37967 114971
rect 16773 114869 16807 114903
rect 17417 114869 17451 114903
rect 21281 114869 21315 114903
rect 23489 114869 23523 114903
rect 28549 114869 28583 114903
rect 35817 114869 35851 114903
rect 38025 114869 38059 114903
rect 3433 114665 3467 114699
rect 8125 114665 8159 114699
rect 12081 114665 12115 114699
rect 13369 114665 13403 114699
rect 14013 114665 14047 114699
rect 15301 114665 15335 114699
rect 15945 114665 15979 114699
rect 17877 114665 17911 114699
rect 22661 114665 22695 114699
rect 27813 114665 27847 114699
rect 28457 114665 28491 114699
rect 29101 114665 29135 114699
rect 30113 114665 30147 114699
rect 30665 114665 30699 114699
rect 31309 114665 31343 114699
rect 31953 114665 31987 114699
rect 36277 114665 36311 114699
rect 1869 114597 1903 114631
rect 2605 114529 2639 114563
rect 3341 114529 3375 114563
rect 5457 114529 5491 114563
rect 7665 114529 7699 114563
rect 8309 114529 8343 114563
rect 8769 114529 8803 114563
rect 9413 114529 9447 114563
rect 10057 114529 10091 114563
rect 10885 114529 10919 114563
rect 12265 114529 12299 114563
rect 12909 114529 12943 114563
rect 13553 114529 13587 114563
rect 14197 114529 14231 114563
rect 14841 114529 14875 114563
rect 15485 114529 15519 114563
rect 16129 114529 16163 114563
rect 18061 114529 18095 114563
rect 19441 114529 19475 114563
rect 20177 114529 20211 114563
rect 22845 114529 22879 114563
rect 23305 114529 23339 114563
rect 24501 114529 24535 114563
rect 24961 114529 24995 114563
rect 25605 114529 25639 114563
rect 26249 114529 26283 114563
rect 27997 114529 28031 114563
rect 28641 114529 28675 114563
rect 29285 114529 29319 114563
rect 30021 114529 30055 114563
rect 30849 114529 30883 114563
rect 31493 114529 31527 114563
rect 32137 114529 32171 114563
rect 33241 114529 33275 114563
rect 33977 114529 34011 114563
rect 34805 114529 34839 114563
rect 35449 114529 35483 114563
rect 35725 114529 35759 114563
rect 36185 114529 36219 114563
rect 37013 114529 37047 114563
rect 2053 114461 2087 114495
rect 2789 114461 2823 114495
rect 4169 114461 4203 114495
rect 4813 114461 4847 114495
rect 7021 114461 7055 114495
rect 33425 114461 33459 114495
rect 35357 114461 35391 114495
rect 36921 114461 36955 114495
rect 7481 114393 7515 114427
rect 8953 114393 8987 114427
rect 10701 114393 10735 114427
rect 19257 114393 19291 114427
rect 19993 114393 20027 114427
rect 24317 114393 24351 114427
rect 12725 114325 12759 114359
rect 14657 114325 14691 114359
rect 34069 114325 34103 114359
rect 3065 114121 3099 114155
rect 4445 114121 4479 114155
rect 4997 114121 5031 114155
rect 5825 114121 5859 114155
rect 8217 114121 8251 114155
rect 30481 114121 30515 114155
rect 31861 114121 31895 114155
rect 33149 114121 33183 114155
rect 33885 114121 33919 114155
rect 6929 114053 6963 114087
rect 31125 114053 31159 114087
rect 32505 114053 32539 114087
rect 34805 114053 34839 114087
rect 5181 113917 5215 113951
rect 6469 113917 6503 113951
rect 7113 113917 7147 113951
rect 7757 113917 7791 113951
rect 8401 113917 8435 113951
rect 22017 113917 22051 113951
rect 23397 113917 23431 113951
rect 26249 113917 26283 113951
rect 26893 113917 26927 113951
rect 27629 113917 27663 113951
rect 30665 113917 30699 113951
rect 31309 113917 31343 113951
rect 32045 113917 32079 113951
rect 32689 113917 32723 113951
rect 33333 113917 33367 113951
rect 34069 113917 34103 113951
rect 36001 113917 36035 113951
rect 36277 113917 36311 113951
rect 36553 113917 36587 113951
rect 1869 113849 1903 113883
rect 2053 113849 2087 113883
rect 34621 113849 34655 113883
rect 37933 113849 37967 113883
rect 6285 113781 6319 113815
rect 7573 113781 7607 113815
rect 35817 113781 35851 113815
rect 38025 113781 38059 113815
rect 30849 113577 30883 113611
rect 33149 113577 33183 113611
rect 34253 113577 34287 113611
rect 34621 113577 34655 113611
rect 34462 113509 34496 113543
rect 35909 113509 35943 113543
rect 36645 113509 36679 113543
rect 2145 113441 2179 113475
rect 2789 113441 2823 113475
rect 3433 113441 3467 113475
rect 4261 113441 4295 113475
rect 4905 113441 4939 113475
rect 5549 113441 5583 113475
rect 6837 113441 6871 113475
rect 7481 113441 7515 113475
rect 8401 113441 8435 113475
rect 9045 113441 9079 113475
rect 31033 113441 31067 113475
rect 31677 113441 31711 113475
rect 33333 113441 33367 113475
rect 34345 113441 34379 113475
rect 35725 113441 35759 113475
rect 36461 113441 36495 113475
rect 37197 113441 37231 113475
rect 33977 113373 34011 113407
rect 31493 113305 31527 113339
rect 37289 113237 37323 113271
rect 1961 113033 1995 113067
rect 31309 113033 31343 113067
rect 32597 113033 32631 113067
rect 33425 113033 33459 113067
rect 34713 113033 34747 113067
rect 35173 113033 35207 113067
rect 36553 113033 36587 113067
rect 28917 112965 28951 112999
rect 31953 112965 31987 112999
rect 34554 112897 34588 112931
rect 28825 112829 28859 112863
rect 29101 112829 29135 112863
rect 31493 112829 31527 112863
rect 32137 112829 32171 112863
rect 32781 112829 32815 112863
rect 33609 112829 33643 112863
rect 34069 112829 34103 112863
rect 34437 112829 34471 112863
rect 37381 112965 37415 112999
rect 35725 112829 35759 112863
rect 37933 112829 37967 112863
rect 1869 112761 1903 112795
rect 35173 112761 35207 112795
rect 36461 112761 36495 112795
rect 37197 112761 37231 112795
rect 29285 112693 29319 112727
rect 34345 112693 34379 112727
rect 35909 112693 35943 112727
rect 38025 112693 38059 112727
rect 34069 112489 34103 112523
rect 36553 112489 36587 112523
rect 1869 112353 1903 112387
rect 34253 112353 34287 112387
rect 35725 112353 35759 112387
rect 36461 112353 36495 112387
rect 37105 112353 37139 112387
rect 2053 112285 2087 112319
rect 37289 112217 37323 112251
rect 35909 112149 35943 112183
rect 35725 111809 35759 111843
rect 36093 111741 36127 111775
rect 37105 111741 37139 111775
rect 37841 111741 37875 111775
rect 36210 111673 36244 111707
rect 36001 111605 36035 111639
rect 36369 111605 36403 111639
rect 37289 111605 37323 111639
rect 38025 111605 38059 111639
rect 1961 111401 1995 111435
rect 36001 111401 36035 111435
rect 35725 111333 35759 111367
rect 1869 111265 1903 111299
rect 35842 111265 35876 111299
rect 37105 111265 37139 111299
rect 35357 111197 35391 111231
rect 35633 111197 35667 111231
rect 37289 111061 37323 111095
rect 1869 110653 1903 110687
rect 26617 110653 26651 110687
rect 37841 110653 37875 110687
rect 2053 110585 2087 110619
rect 26801 110517 26835 110551
rect 38025 110517 38059 110551
rect 37105 110177 37139 110211
rect 37289 109973 37323 110007
rect 1961 109769 1995 109803
rect 34621 109769 34655 109803
rect 37289 109769 37323 109803
rect 32689 109565 32723 109599
rect 32965 109565 32999 109599
rect 33241 109565 33275 109599
rect 33333 109565 33367 109599
rect 33977 109565 34011 109599
rect 37105 109565 37139 109599
rect 37841 109565 37875 109599
rect 1869 109497 1903 109531
rect 34462 109497 34496 109531
rect 33241 109429 33275 109463
rect 34253 109429 34287 109463
rect 34345 109429 34379 109463
rect 38025 109429 38059 109463
rect 34437 109225 34471 109259
rect 37289 109225 37323 109259
rect 34161 109157 34195 109191
rect 1869 109089 1903 109123
rect 34069 109089 34103 109123
rect 37105 109089 37139 109123
rect 2145 109021 2179 109055
rect 33793 109021 33827 109055
rect 34278 109021 34312 109055
rect 13093 108681 13127 108715
rect 28733 108681 28767 108715
rect 38025 108613 38059 108647
rect 33701 108545 33735 108579
rect 12909 108477 12943 108511
rect 28549 108477 28583 108511
rect 33333 108477 33367 108511
rect 34161 108477 34195 108511
rect 37841 108477 37875 108511
rect 33149 108409 33183 108443
rect 34345 108341 34379 108375
rect 1961 108137 1995 108171
rect 1869 108001 1903 108035
rect 33333 108001 33367 108035
rect 37197 108001 37231 108035
rect 37381 107865 37415 107899
rect 33517 107797 33551 107831
rect 33149 107525 33183 107559
rect 1869 107389 1903 107423
rect 32965 107389 32999 107423
rect 37197 107389 37231 107423
rect 2053 107321 2087 107355
rect 37933 107321 37967 107355
rect 37289 107253 37323 107287
rect 38025 107253 38059 107287
rect 1869 106913 1903 106947
rect 37197 106913 37231 106947
rect 1961 106709 1995 106743
rect 37289 106709 37323 106743
rect 38117 106369 38151 106403
rect 37933 106301 37967 106335
rect 10149 105961 10183 105995
rect 33149 105893 33183 105927
rect 35265 105893 35299 105927
rect 1409 105825 1443 105859
rect 9965 105825 9999 105859
rect 35081 105825 35115 105859
rect 35173 105825 35207 105859
rect 37197 105825 37231 105859
rect 1593 105757 1627 105791
rect 34621 105757 34655 105791
rect 34713 105757 34747 105791
rect 33241 105621 33275 105655
rect 37289 105621 37323 105655
rect 37933 105213 37967 105247
rect 1869 105145 1903 105179
rect 1961 105077 1995 105111
rect 38025 105077 38059 105111
rect 37197 104805 37231 104839
rect 37289 104533 37323 104567
rect 30665 104329 30699 104363
rect 1501 104125 1535 104159
rect 30481 104125 30515 104159
rect 37197 104125 37231 104159
rect 2053 104057 2087 104091
rect 37933 104057 37967 104091
rect 37289 103989 37323 104023
rect 38025 103989 38059 104023
rect 30941 103785 30975 103819
rect 30389 103717 30423 103751
rect 1869 103649 1903 103683
rect 30021 103649 30055 103683
rect 30849 103649 30883 103683
rect 37197 103649 37231 103683
rect 2053 103513 2087 103547
rect 37381 103513 37415 103547
rect 7113 103241 7147 103275
rect 30573 103241 30607 103275
rect 25697 103105 25731 103139
rect 6929 103037 6963 103071
rect 30481 103037 30515 103071
rect 25513 102969 25547 103003
rect 37933 102969 37967 103003
rect 38025 102901 38059 102935
rect 7757 102697 7791 102731
rect 1869 102561 1903 102595
rect 2053 102561 2087 102595
rect 7573 102561 7607 102595
rect 37197 102561 37231 102595
rect 37289 102357 37323 102391
rect 25881 102085 25915 102119
rect 1409 101949 1443 101983
rect 9505 101949 9539 101983
rect 37197 101949 37231 101983
rect 37381 101949 37415 101983
rect 25697 101881 25731 101915
rect 37933 101881 37967 101915
rect 9689 101813 9723 101847
rect 38025 101813 38059 101847
rect 37197 101473 37231 101507
rect 37289 101269 37323 101303
rect 6561 101065 6595 101099
rect 1409 100861 1443 100895
rect 6377 100861 6411 100895
rect 37933 100793 37967 100827
rect 38025 100725 38059 100759
rect 1409 100385 1443 100419
rect 37197 100385 37231 100419
rect 37289 100181 37323 100215
rect 6285 99977 6319 100011
rect 38117 99909 38151 99943
rect 6101 99773 6135 99807
rect 37289 99773 37323 99807
rect 37933 99773 37967 99807
rect 37473 99637 37507 99671
rect 1409 99297 1443 99331
rect 5089 99297 5123 99331
rect 37197 99297 37231 99331
rect 5273 99161 5307 99195
rect 37381 99093 37415 99127
rect 1409 98685 1443 98719
rect 37933 98685 37967 98719
rect 38117 98549 38151 98583
rect 5089 98345 5123 98379
rect 4905 98209 4939 98243
rect 37105 98209 37139 98243
rect 37289 98005 37323 98039
rect 4445 97801 4479 97835
rect 1409 97597 1443 97631
rect 4261 97597 4295 97631
rect 37841 97597 37875 97631
rect 38025 97461 38059 97495
rect 1409 97121 1443 97155
rect 37105 97121 37139 97155
rect 37289 96917 37323 96951
rect 37105 96509 37139 96543
rect 37933 96441 37967 96475
rect 37289 96373 37323 96407
rect 38025 96373 38059 96407
rect 3525 96169 3559 96203
rect 1409 96033 1443 96067
rect 3341 96033 3375 96067
rect 37197 96033 37231 96067
rect 37381 95897 37415 95931
rect 2973 95625 3007 95659
rect 1409 95421 1443 95455
rect 2789 95421 2823 95455
rect 38117 95421 38151 95455
rect 37933 95353 37967 95387
rect 37197 94945 37231 94979
rect 37289 94741 37323 94775
rect 2881 94537 2915 94571
rect 1409 94333 1443 94367
rect 2697 94333 2731 94367
rect 37197 94333 37231 94367
rect 37933 94265 37967 94299
rect 37289 94197 37323 94231
rect 38025 94197 38059 94231
rect 37381 93993 37415 94027
rect 1409 93857 1443 93891
rect 37197 93857 37231 93891
rect 1409 93245 1443 93279
rect 37289 93245 37323 93279
rect 37933 93245 37967 93279
rect 37473 93109 37507 93143
rect 38117 93109 38151 93143
rect 2329 92905 2363 92939
rect 30757 92837 30791 92871
rect 2145 92769 2179 92803
rect 30573 92769 30607 92803
rect 1409 92157 1443 92191
rect 37289 92157 37323 92191
rect 37933 92157 37967 92191
rect 37473 92021 37507 92055
rect 38117 92021 38151 92055
rect 1409 91681 1443 91715
rect 37197 91681 37231 91715
rect 37381 91477 37415 91511
rect 1593 91273 1627 91307
rect 38117 91205 38151 91239
rect 1409 91069 1443 91103
rect 37289 91069 37323 91103
rect 37933 91069 37967 91103
rect 37473 90933 37507 90967
rect 1593 90729 1627 90763
rect 1409 90593 1443 90627
rect 2053 90593 2087 90627
rect 38117 90117 38151 90151
rect 1409 89981 1443 90015
rect 37289 89981 37323 90015
rect 37933 89981 37967 90015
rect 37473 89845 37507 89879
rect 37197 89505 37231 89539
rect 37381 89301 37415 89335
rect 1409 88893 1443 88927
rect 37289 88893 37323 88927
rect 37933 88893 37967 88927
rect 37473 88757 37507 88791
rect 38117 88757 38151 88791
rect 1409 88417 1443 88451
rect 33701 87805 33735 87839
rect 33793 87805 33827 87839
rect 34069 87805 34103 87839
rect 34345 87805 34379 87839
rect 34621 87805 34655 87839
rect 37289 87805 37323 87839
rect 37933 87805 37967 87839
rect 33241 87737 33275 87771
rect 37473 87669 37507 87703
rect 38117 87669 38151 87703
rect 37105 87465 37139 87499
rect 1409 87329 1443 87363
rect 33701 87329 33735 87363
rect 33793 87329 33827 87363
rect 34069 87329 34103 87363
rect 34345 87329 34379 87363
rect 34621 87329 34655 87363
rect 37197 87329 37231 87363
rect 37105 87193 37139 87227
rect 33333 87125 33367 87159
rect 37381 87125 37415 87159
rect 27261 86853 27295 86887
rect 32689 86853 32723 86887
rect 38117 86853 38151 86887
rect 1409 86717 1443 86751
rect 27077 86717 27111 86751
rect 27813 86717 27847 86751
rect 31769 86717 31803 86751
rect 32505 86717 32539 86751
rect 33701 86717 33735 86751
rect 33793 86717 33827 86751
rect 34069 86717 34103 86751
rect 34345 86717 34379 86751
rect 34621 86717 34655 86751
rect 37289 86717 37323 86751
rect 37933 86717 37967 86751
rect 33241 86649 33275 86683
rect 27997 86581 28031 86615
rect 31953 86581 31987 86615
rect 37473 86581 37507 86615
rect 33701 86241 33735 86275
rect 33793 86241 33827 86275
rect 34069 86241 34103 86275
rect 34345 86241 34379 86275
rect 34529 86241 34563 86275
rect 33333 86037 33367 86071
rect 27353 85833 27387 85867
rect 38117 85833 38151 85867
rect 37473 85765 37507 85799
rect 1409 85629 1443 85663
rect 27169 85629 27203 85663
rect 32413 85629 32447 85663
rect 32505 85629 32539 85663
rect 32781 85629 32815 85663
rect 33057 85629 33091 85663
rect 33333 85629 33367 85663
rect 37289 85629 37323 85663
rect 37933 85629 37967 85663
rect 31953 85561 31987 85595
rect 1409 85153 1443 85187
rect 33057 85153 33091 85187
rect 33241 84949 33275 84983
rect 27169 84677 27203 84711
rect 26985 84541 27019 84575
rect 31309 84541 31343 84575
rect 32505 84541 32539 84575
rect 32781 84541 32815 84575
rect 32873 84541 32907 84575
rect 33149 84541 33183 84575
rect 33425 84541 33459 84575
rect 37289 84541 37323 84575
rect 37933 84541 37967 84575
rect 32045 84473 32079 84507
rect 31493 84405 31527 84439
rect 37473 84405 37507 84439
rect 38117 84405 38151 84439
rect 1409 84065 1443 84099
rect 31125 84065 31159 84099
rect 31401 84065 31435 84099
rect 31493 84065 31527 84099
rect 31769 84065 31803 84099
rect 32045 84065 32079 84099
rect 33517 84065 33551 84099
rect 33793 84065 33827 84099
rect 33931 84065 33965 84099
rect 34161 84065 34195 84099
rect 34437 84065 34471 84099
rect 37197 84065 37231 84099
rect 30757 83861 30791 83895
rect 33149 83861 33183 83895
rect 37381 83861 37415 83895
rect 1409 83453 1443 83487
rect 32321 83453 32355 83487
rect 32413 83453 32447 83487
rect 32689 83453 32723 83487
rect 32965 83453 32999 83487
rect 33241 83453 33275 83487
rect 37289 83453 37323 83487
rect 37933 83453 37967 83487
rect 31861 83385 31895 83419
rect 37473 83317 37507 83351
rect 38117 83317 38151 83351
rect 30665 82977 30699 83011
rect 31125 82977 31159 83011
rect 31401 82977 31435 83011
rect 31493 82977 31527 83011
rect 31769 82977 31803 83011
rect 32045 82977 32079 83011
rect 33517 82977 33551 83011
rect 33609 82977 33643 83011
rect 33885 82977 33919 83011
rect 34161 82977 34195 83011
rect 34437 82977 34471 83011
rect 33149 82841 33183 82875
rect 1409 82365 1443 82399
rect 31953 82365 31987 82399
rect 32045 82365 32079 82399
rect 32321 82365 32355 82399
rect 32597 82365 32631 82399
rect 32873 82365 32907 82399
rect 37289 82365 37323 82399
rect 37933 82365 37967 82399
rect 31493 82297 31527 82331
rect 37473 82229 37507 82263
rect 38117 82229 38151 82263
rect 1409 81889 1443 81923
rect 31125 81889 31159 81923
rect 31401 81889 31435 81923
rect 31493 81889 31527 81923
rect 31769 81889 31803 81923
rect 32045 81889 32079 81923
rect 33517 81889 33551 81923
rect 33609 81889 33643 81923
rect 33885 81889 33919 81923
rect 34161 81889 34195 81923
rect 34437 81889 34471 81923
rect 37197 81889 37231 81923
rect 30757 81685 30791 81719
rect 33149 81685 33183 81719
rect 37381 81685 37415 81719
rect 37473 81481 37507 81515
rect 31769 81277 31803 81311
rect 32045 81277 32079 81311
rect 32137 81277 32171 81311
rect 32413 81277 32447 81311
rect 32689 81277 32723 81311
rect 33701 81277 33735 81311
rect 33793 81277 33827 81311
rect 34069 81277 34103 81311
rect 34345 81277 34379 81311
rect 34621 81277 34655 81311
rect 37289 81277 37323 81311
rect 37933 81277 37967 81311
rect 31401 81141 31435 81175
rect 33333 81141 33367 81175
rect 38117 81141 38151 81175
rect 33149 80937 33183 80971
rect 1409 80801 1443 80835
rect 31125 80801 31159 80835
rect 31217 80801 31251 80835
rect 31493 80801 31527 80835
rect 31769 80801 31803 80835
rect 31953 80801 31987 80835
rect 32137 80801 32171 80835
rect 33517 80801 33551 80835
rect 33793 80801 33827 80835
rect 33885 80801 33919 80835
rect 34161 80801 34195 80835
rect 34437 80801 34471 80835
rect 30757 80597 30791 80631
rect 32137 80597 32171 80631
rect 37473 80325 37507 80359
rect 1409 80189 1443 80223
rect 31401 80189 31435 80223
rect 31677 80189 31711 80223
rect 31769 80189 31803 80223
rect 32045 80189 32079 80223
rect 32321 80189 32355 80223
rect 37289 80189 37323 80223
rect 37933 80189 37967 80223
rect 30941 80121 30975 80155
rect 38117 80053 38151 80087
rect 1409 79713 1443 79747
rect 14841 79713 14875 79747
rect 37197 79713 37231 79747
rect 15025 79509 15059 79543
rect 37381 79509 37415 79543
rect 37473 79237 37507 79271
rect 37289 79101 37323 79135
rect 37933 79101 37967 79135
rect 38117 78965 38151 78999
rect 1409 78625 1443 78659
rect 27813 78625 27847 78659
rect 27997 78421 28031 78455
rect 37473 78149 37507 78183
rect 1409 78013 1443 78047
rect 32413 78013 32447 78047
rect 37289 78013 37323 78047
rect 37933 78013 37967 78047
rect 32597 77877 32631 77911
rect 38117 77877 38151 77911
rect 1409 76925 1443 76959
rect 37289 76925 37323 76959
rect 37933 76925 37967 76959
rect 37473 76789 37507 76823
rect 38117 76789 38151 76823
rect 31125 76585 31159 76619
rect 23489 76517 23523 76551
rect 1409 76449 1443 76483
rect 30941 76449 30975 76483
rect 23673 76313 23707 76347
rect 20085 75837 20119 75871
rect 20177 75837 20211 75871
rect 20361 75837 20395 75871
rect 37289 75837 37323 75871
rect 37933 75837 37967 75871
rect 37473 75701 37507 75735
rect 38117 75701 38151 75735
rect 20361 75497 20395 75531
rect 21189 75497 21223 75531
rect 29653 75497 29687 75531
rect 1409 75361 1443 75395
rect 20177 75361 20211 75395
rect 20821 75361 20855 75395
rect 21005 75361 21039 75395
rect 29469 75361 29503 75395
rect 29653 75361 29687 75395
rect 29929 75361 29963 75395
rect 30113 75361 30147 75395
rect 37197 75361 37231 75395
rect 19993 75293 20027 75327
rect 37381 75157 37415 75191
rect 39221 75089 39255 75123
rect 20361 74953 20395 74987
rect 37473 74885 37507 74919
rect 19993 74817 20027 74851
rect 1409 74749 1443 74783
rect 20177 74749 20211 74783
rect 37289 74749 37323 74783
rect 37933 74749 37967 74783
rect 38117 74613 38151 74647
rect 37197 74273 37231 74307
rect 37381 74069 37415 74103
rect 38117 73797 38151 73831
rect 1409 73661 1443 73695
rect 20085 73661 20119 73695
rect 20729 73661 20763 73695
rect 37289 73661 37323 73695
rect 37933 73661 37967 73695
rect 20269 73525 20303 73559
rect 20913 73525 20947 73559
rect 37473 73525 37507 73559
rect 1409 73185 1443 73219
rect 16129 72777 16163 72811
rect 16957 72777 16991 72811
rect 17785 72777 17819 72811
rect 15761 72641 15795 72675
rect 16589 72641 16623 72675
rect 17417 72641 17451 72675
rect 15945 72573 15979 72607
rect 16773 72573 16807 72607
rect 17601 72573 17635 72607
rect 19993 72573 20027 72607
rect 37289 72573 37323 72607
rect 37933 72573 37967 72607
rect 38945 72573 38979 72607
rect 20177 72437 20211 72471
rect 37473 72437 37507 72471
rect 38117 72437 38151 72471
rect 16405 72233 16439 72267
rect 17693 72233 17727 72267
rect 17141 72165 17175 72199
rect 1409 72097 1443 72131
rect 16221 72097 16255 72131
rect 17417 72097 17451 72131
rect 17509 72097 17543 72131
rect 37197 72097 37231 72131
rect 16037 72029 16071 72063
rect 37381 71893 37415 71927
rect 38945 71757 38979 71791
rect 16957 71689 16991 71723
rect 17785 71689 17819 71723
rect 35909 71689 35943 71723
rect 16129 71621 16163 71655
rect 15761 71553 15795 71587
rect 16589 71553 16623 71587
rect 17417 71553 17451 71587
rect 1409 71485 1443 71519
rect 15945 71485 15979 71519
rect 16773 71485 16807 71519
rect 17601 71485 17635 71519
rect 31493 71485 31527 71519
rect 31585 71485 31619 71519
rect 31861 71485 31895 71519
rect 32137 71485 32171 71519
rect 32413 71485 32447 71519
rect 35817 71485 35851 71519
rect 37473 71485 37507 71519
rect 38117 71485 38151 71519
rect 31033 71417 31067 71451
rect 37289 71349 37323 71383
rect 37933 71349 37967 71383
rect 15577 71145 15611 71179
rect 16405 71145 16439 71179
rect 15393 71009 15427 71043
rect 16221 71009 16255 71043
rect 31125 71009 31159 71043
rect 31401 71009 31435 71043
rect 31493 71009 31527 71043
rect 31769 71009 31803 71043
rect 32045 71009 32079 71043
rect 37381 71009 37415 71043
rect 15209 70941 15243 70975
rect 16037 70941 16071 70975
rect 30757 70805 30791 70839
rect 37197 70805 37231 70839
rect 15853 70601 15887 70635
rect 16681 70601 16715 70635
rect 17509 70601 17543 70635
rect 37289 70533 37323 70567
rect 37933 70533 37967 70567
rect 16313 70465 16347 70499
rect 1409 70397 1443 70431
rect 15485 70397 15519 70431
rect 15669 70397 15703 70431
rect 16497 70397 16531 70431
rect 16957 70397 16991 70431
rect 17233 70397 17267 70431
rect 17325 70397 17359 70431
rect 31401 70397 31435 70431
rect 31677 70397 31711 70431
rect 31769 70397 31803 70431
rect 32045 70397 32079 70431
rect 32321 70397 32355 70431
rect 37473 70397 37507 70431
rect 38117 70397 38151 70431
rect 30941 70329 30975 70363
rect 16405 70057 16439 70091
rect 1409 69921 1443 69955
rect 16221 69921 16255 69955
rect 36737 69921 36771 69955
rect 37381 69921 37415 69955
rect 16037 69853 16071 69887
rect 36553 69785 36587 69819
rect 37197 69717 37231 69751
rect 16497 69513 16531 69547
rect 37197 69445 37231 69479
rect 16129 69377 16163 69411
rect 16313 69309 16347 69343
rect 36645 69309 36679 69343
rect 37013 69309 37047 69343
rect 38117 69309 38151 69343
rect 36829 69241 36863 69275
rect 36921 69241 36955 69275
rect 39405 75021 39439 75055
rect 39313 74885 39347 74919
rect 39313 70329 39347 70363
rect 37933 69173 37967 69207
rect 39221 69173 39255 69207
rect 36921 68901 36955 68935
rect 37013 68901 37047 68935
rect 1409 68833 1443 68867
rect 36277 68833 36311 68867
rect 36737 68833 36771 68867
rect 37105 68833 37139 68867
rect 36093 68697 36127 68731
rect 37289 68629 37323 68663
rect 37289 68425 37323 68459
rect 1409 68221 1443 68255
rect 31953 68221 31987 68255
rect 36277 68221 36311 68255
rect 36737 68221 36771 68255
rect 36921 68221 36955 68255
rect 37105 68221 37139 68255
rect 38117 68221 38151 68255
rect 31861 68153 31895 68187
rect 37013 68153 37047 68187
rect 32137 68085 32171 68119
rect 36093 68085 36127 68119
rect 37933 68085 37967 68119
rect 36921 67813 36955 67847
rect 37013 67813 37047 67847
rect 36001 67745 36035 67779
rect 36737 67745 36771 67779
rect 37105 67745 37139 67779
rect 37289 67609 37323 67643
rect 36185 67541 36219 67575
rect 38117 67337 38151 67371
rect 37105 67269 37139 67303
rect 1409 67133 1443 67167
rect 32965 67133 32999 67167
rect 35909 67133 35943 67167
rect 36553 67133 36587 67167
rect 36921 67133 36955 67167
rect 37565 67133 37599 67167
rect 37933 67133 37967 67167
rect 39405 67133 39439 67167
rect 39773 69649 39807 69683
rect 39773 67133 39807 67167
rect 33149 67065 33183 67099
rect 36737 67065 36771 67099
rect 36829 67065 36863 67099
rect 37749 67065 37783 67099
rect 37841 67065 37875 67099
rect 36093 66997 36127 67031
rect 36001 66725 36035 66759
rect 37013 66725 37047 66759
rect 1409 66657 1443 66691
rect 34713 66657 34747 66691
rect 35357 66657 35391 66691
rect 35817 66657 35851 66691
rect 36093 66657 36127 66691
rect 36185 66657 36219 66691
rect 36829 66657 36863 66691
rect 37105 66657 37139 66691
rect 37197 66657 37231 66691
rect 36369 66521 36403 66555
rect 34529 66453 34563 66487
rect 35173 66453 35207 66487
rect 37381 66453 37415 66487
rect 38117 66181 38151 66215
rect 1409 66045 1443 66079
rect 32965 66045 32999 66079
rect 35909 66045 35943 66079
rect 36645 66045 36679 66079
rect 37565 66045 37599 66079
rect 37933 66045 37967 66079
rect 33149 65977 33183 66011
rect 36829 65977 36863 66011
rect 37749 65977 37783 66011
rect 37841 65977 37875 66011
rect 36001 65909 36035 65943
rect 33149 65569 33183 65603
rect 35081 65569 35115 65603
rect 35725 65569 35759 65603
rect 36369 65569 36403 65603
rect 36829 65569 36863 65603
rect 37013 65569 37047 65603
rect 37105 65569 37139 65603
rect 37243 65569 37277 65603
rect 33241 65365 33275 65399
rect 34897 65365 34931 65399
rect 35541 65365 35575 65399
rect 36185 65365 36219 65399
rect 37381 65365 37415 65399
rect 32965 65161 32999 65195
rect 36001 65161 36035 65195
rect 37105 65093 37139 65127
rect 38117 65093 38151 65127
rect 1409 64957 1443 64991
rect 32873 64957 32907 64991
rect 34805 64957 34839 64991
rect 35909 64957 35943 64991
rect 36553 64957 36587 64991
rect 36921 64957 36955 64991
rect 37565 64957 37599 64991
rect 37933 64957 37967 64991
rect 36737 64889 36771 64923
rect 36829 64889 36863 64923
rect 37749 64889 37783 64923
rect 37841 64889 37875 64923
rect 34621 64821 34655 64855
rect 35357 64617 35391 64651
rect 20177 64549 20211 64583
rect 33149 64549 33183 64583
rect 36093 64549 36127 64583
rect 37013 64549 37047 64583
rect 37105 64549 37139 64583
rect 1409 64481 1443 64515
rect 31677 64481 31711 64515
rect 34713 64481 34747 64515
rect 35173 64481 35207 64515
rect 35817 64481 35851 64515
rect 36001 64481 36035 64515
rect 36185 64481 36219 64515
rect 36829 64481 36863 64515
rect 37197 64481 37231 64515
rect 31861 64345 31895 64379
rect 20269 64277 20303 64311
rect 33241 64277 33275 64311
rect 34529 64277 34563 64311
rect 36369 64277 36403 64311
rect 37381 64277 37415 64311
rect 36093 64005 36127 64039
rect 34805 63869 34839 63903
rect 35909 63869 35943 63903
rect 36553 63869 36587 63903
rect 36921 63869 36955 63903
rect 37565 63869 37599 63903
rect 37749 63869 37783 63903
rect 37933 63869 37967 63903
rect 36737 63801 36771 63835
rect 36829 63801 36863 63835
rect 37841 63801 37875 63835
rect 34621 63733 34655 63767
rect 37105 63733 37139 63767
rect 38117 63733 38151 63767
rect 34713 63529 34747 63563
rect 36093 63461 36127 63495
rect 37013 63461 37047 63495
rect 1409 63393 1443 63427
rect 34529 63393 34563 63427
rect 35173 63393 35207 63427
rect 35817 63393 35851 63427
rect 36001 63393 36035 63427
rect 36185 63393 36219 63427
rect 36829 63393 36863 63427
rect 37105 63393 37139 63427
rect 37197 63393 37231 63427
rect 35357 63189 35391 63223
rect 36369 63189 36403 63223
rect 37381 63189 37415 63223
rect 37657 62917 37691 62951
rect 1409 62781 1443 62815
rect 31861 62781 31895 62815
rect 32689 62781 32723 62815
rect 36093 62781 36127 62815
rect 36461 62781 36495 62815
rect 37105 62781 37139 62815
rect 37289 62781 37323 62815
rect 37381 62781 37415 62815
rect 37478 62781 37512 62815
rect 32045 62713 32079 62747
rect 32873 62713 32907 62747
rect 36277 62713 36311 62747
rect 36369 62713 36403 62747
rect 36645 62645 36679 62679
rect 35449 62441 35483 62475
rect 36921 62373 36955 62407
rect 15393 62305 15427 62339
rect 35633 62305 35667 62339
rect 36277 62305 36311 62339
rect 36737 62305 36771 62339
rect 37013 62305 37047 62339
rect 37157 62305 37191 62339
rect 36093 62169 36127 62203
rect 15485 62101 15519 62135
rect 37289 62101 37323 62135
rect 35817 61829 35851 61863
rect 37657 61829 37691 61863
rect 1409 61693 1443 61727
rect 36001 61693 36035 61727
rect 36645 61693 36679 61727
rect 37105 61693 37139 61727
rect 37478 61693 37512 61727
rect 37289 61625 37323 61659
rect 37381 61625 37415 61659
rect 36461 61557 36495 61591
rect 36185 61353 36219 61387
rect 36921 61285 36955 61319
rect 1409 61217 1443 61251
rect 34897 61217 34931 61251
rect 35541 61217 35575 61251
rect 36001 61217 36035 61251
rect 36737 61217 36771 61251
rect 37013 61217 37047 61251
rect 37110 61217 37144 61251
rect 34713 61081 34747 61115
rect 37289 61081 37323 61115
rect 35357 61013 35391 61047
rect 37657 60741 37691 60775
rect 36001 60605 36035 60639
rect 36277 60605 36311 60639
rect 36421 60605 36455 60639
rect 37105 60605 37139 60639
rect 37289 60605 37323 60639
rect 37478 60605 37512 60639
rect 36185 60537 36219 60571
rect 37381 60537 37415 60571
rect 36561 60469 36595 60503
rect 33425 60197 33459 60231
rect 35909 60197 35943 60231
rect 37014 60197 37048 60231
rect 1409 60129 1443 60163
rect 33057 60129 33091 60163
rect 33205 60129 33239 60163
rect 33333 60129 33367 60163
rect 33563 60129 33597 60163
rect 35173 60129 35207 60163
rect 35633 60129 35667 60163
rect 35817 60129 35851 60163
rect 36006 60129 36040 60163
rect 36757 60129 36791 60163
rect 36921 60129 36955 60163
rect 37157 60129 37191 60163
rect 36185 59993 36219 60027
rect 33701 59925 33735 59959
rect 34989 59925 35023 59959
rect 37289 59925 37323 59959
rect 34621 59721 34655 59755
rect 36553 59653 36587 59687
rect 37657 59653 37691 59687
rect 1409 59517 1443 59551
rect 32965 59517 32999 59551
rect 33241 59517 33275 59551
rect 33333 59517 33367 59551
rect 33609 59517 33643 59551
rect 33793 59517 33827 59551
rect 34805 59517 34839 59551
rect 36001 59517 36035 59551
rect 36421 59517 36455 59551
rect 37105 59517 37139 59551
rect 37478 59517 37512 59551
rect 32505 59449 32539 59483
rect 36185 59449 36219 59483
rect 36277 59449 36311 59483
rect 37289 59449 37323 59483
rect 37381 59449 37415 59483
rect 31677 59109 31711 59143
rect 31769 59109 31803 59143
rect 35909 59109 35943 59143
rect 36921 59109 36955 59143
rect 37013 59109 37047 59143
rect 31401 59041 31435 59075
rect 31494 59041 31528 59075
rect 31907 59041 31941 59075
rect 33517 59041 33551 59075
rect 33609 59041 33643 59075
rect 33885 59041 33919 59075
rect 34161 59041 34195 59075
rect 34345 59041 34379 59075
rect 35633 59041 35667 59075
rect 35817 59041 35851 59075
rect 36006 59041 36040 59075
rect 36737 59041 36771 59075
rect 37157 59041 37191 59075
rect 32045 58837 32079 58871
rect 33149 58837 33183 58871
rect 36185 58837 36219 58871
rect 37289 58837 37323 58871
rect 36461 58633 36495 58667
rect 35817 58565 35851 58599
rect 37657 58565 37691 58599
rect 1409 58429 1443 58463
rect 32873 58429 32907 58463
rect 33149 58429 33183 58463
rect 33241 58429 33275 58463
rect 33517 58429 33551 58463
rect 33793 58429 33827 58463
rect 36001 58429 36035 58463
rect 36645 58429 36679 58463
rect 37105 58429 37139 58463
rect 37478 58429 37512 58463
rect 32413 58361 32447 58395
rect 37289 58361 37323 58395
rect 37381 58361 37415 58395
rect 36553 58089 36587 58123
rect 1409 57953 1443 57987
rect 36737 57953 36771 57987
rect 37381 57953 37415 57987
rect 37197 57817 37231 57851
rect 37289 57545 37323 57579
rect 37473 57341 37507 57375
rect 37933 57341 37967 57375
rect 1409 56865 1443 56899
rect 15761 56457 15795 56491
rect 16681 56457 16715 56491
rect 17601 56457 17635 56491
rect 1409 56253 1443 56287
rect 15393 56253 15427 56287
rect 15577 56253 15611 56287
rect 16313 56253 16347 56287
rect 16497 56253 16531 56287
rect 17325 56253 17359 56287
rect 17417 56253 17451 56287
rect 33057 56253 33091 56287
rect 33205 56253 33239 56287
rect 33563 56253 33597 56287
rect 37473 56253 37507 56287
rect 37933 56253 37967 56287
rect 33333 56185 33367 56219
rect 33425 56185 33459 56219
rect 17049 56117 17083 56151
rect 33701 56117 33735 56151
rect 37289 56117 37323 56151
rect 33609 55845 33643 55879
rect 33241 55777 33275 55811
rect 33389 55777 33423 55811
rect 33517 55777 33551 55811
rect 33747 55777 33781 55811
rect 37197 55777 37231 55811
rect 33885 55641 33919 55675
rect 1409 55165 1443 55199
rect 32045 55165 32079 55199
rect 32193 55165 32227 55199
rect 32321 55165 32355 55199
rect 32551 55165 32585 55199
rect 33241 55165 33275 55199
rect 33389 55165 33423 55199
rect 33609 55165 33643 55199
rect 33747 55165 33781 55199
rect 37473 55165 37507 55199
rect 37933 55165 37967 55199
rect 32413 55097 32447 55131
rect 33517 55097 33551 55131
rect 32689 55029 32723 55063
rect 33885 55029 33919 55063
rect 37289 55029 37323 55063
rect 1409 54689 1443 54723
rect 33149 54689 33183 54723
rect 33297 54689 33331 54723
rect 33425 54689 33459 54723
rect 33517 54689 33551 54723
rect 33655 54689 33689 54723
rect 37197 54689 37231 54723
rect 33793 54485 33827 54519
rect 21557 54281 21591 54315
rect 32137 54281 32171 54315
rect 33241 54281 33275 54315
rect 37565 54281 37599 54315
rect 34253 54213 34287 54247
rect 33149 54077 33183 54111
rect 21465 54009 21499 54043
rect 32045 54009 32079 54043
rect 34069 54009 34103 54043
rect 37289 54009 37323 54043
rect 19349 53737 19383 53771
rect 22937 53737 22971 53771
rect 25053 53737 25087 53771
rect 27997 53737 28031 53771
rect 24961 53669 24995 53703
rect 29377 53669 29411 53703
rect 1409 53601 1443 53635
rect 19073 53601 19107 53635
rect 22845 53601 22879 53635
rect 27905 53601 27939 53635
rect 29009 53601 29043 53635
rect 36737 53601 36771 53635
rect 37197 53601 37231 53635
rect 36553 53397 36587 53431
rect 1409 52989 1443 53023
rect 37289 52989 37323 53023
rect 37933 52989 37967 53023
rect 1409 52513 1443 52547
rect 33701 52037 33735 52071
rect 33057 51901 33091 51935
rect 33150 51901 33184 51935
rect 33563 51901 33597 51935
rect 37473 51901 37507 51935
rect 37933 51901 37967 51935
rect 33333 51833 33367 51867
rect 33425 51833 33459 51867
rect 32873 51765 32907 51799
rect 37289 51765 37323 51799
rect 33701 51493 33735 51527
rect 1409 51425 1443 51459
rect 33333 51425 33367 51459
rect 33426 51425 33460 51459
rect 33609 51425 33643 51459
rect 33839 51425 33873 51459
rect 37197 51425 37231 51459
rect 33149 51221 33183 51255
rect 33977 51221 34011 51255
rect 33333 50813 33367 50847
rect 33426 50813 33460 50847
rect 33563 50813 33597 50847
rect 33817 50813 33851 50847
rect 37473 50813 37507 50847
rect 37933 50813 37967 50847
rect 1869 50745 1903 50779
rect 33709 50745 33743 50779
rect 1961 50677 1995 50711
rect 33241 50677 33275 50711
rect 33977 50677 34011 50711
rect 37289 50677 37323 50711
rect 33609 50405 33643 50439
rect 28917 50337 28951 50371
rect 33333 50337 33367 50371
rect 33426 50337 33460 50371
rect 33714 50337 33748 50371
rect 33839 50337 33873 50371
rect 34621 50337 34655 50371
rect 28733 50201 28767 50235
rect 29101 50201 29135 50235
rect 34805 50201 34839 50235
rect 33977 50133 34011 50167
rect 2053 49861 2087 49895
rect 1869 49725 1903 49759
rect 32045 49725 32079 49759
rect 32229 49725 32263 49759
rect 32413 49725 32447 49759
rect 32689 49725 32723 49759
rect 37933 49725 37967 49759
rect 32045 49589 32079 49623
rect 1869 49249 1903 49283
rect 37381 49249 37415 49283
rect 1961 49045 1995 49079
rect 37197 49045 37231 49079
rect 16681 48637 16715 48671
rect 27629 48637 27663 48671
rect 28089 48637 28123 48671
rect 28365 48637 28399 48671
rect 28549 48637 28583 48671
rect 37289 48637 37323 48671
rect 37933 48637 37967 48671
rect 28825 48569 28859 48603
rect 16865 48501 16899 48535
rect 2053 48229 2087 48263
rect 1869 48161 1903 48195
rect 37381 48161 37415 48195
rect 37197 47957 37231 47991
rect 16773 47549 16807 47583
rect 37289 47549 37323 47583
rect 37933 47549 37967 47583
rect 1869 47481 1903 47515
rect 1961 47413 1995 47447
rect 16957 47413 16991 47447
rect 33977 47073 34011 47107
rect 34070 47073 34104 47107
rect 34253 47073 34287 47107
rect 34345 47073 34379 47107
rect 34483 47073 34517 47107
rect 34621 46937 34655 46971
rect 34621 46597 34655 46631
rect 1869 46461 1903 46495
rect 33977 46461 34011 46495
rect 34070 46461 34104 46495
rect 34483 46461 34517 46495
rect 37473 46461 37507 46495
rect 37933 46461 37967 46495
rect 34253 46393 34287 46427
rect 34345 46393 34379 46427
rect 1961 46325 1995 46359
rect 37289 46325 37323 46359
rect 1869 45985 1903 46019
rect 33977 45985 34011 46019
rect 34070 45985 34104 46019
rect 34253 45985 34287 46019
rect 34345 45985 34379 46019
rect 34483 45985 34517 46019
rect 37197 45985 37231 46019
rect 34621 45849 34655 45883
rect 1961 45781 1995 45815
rect 34621 45509 34655 45543
rect 33977 45373 34011 45407
rect 34070 45373 34104 45407
rect 34483 45373 34517 45407
rect 37473 45373 37507 45407
rect 37933 45373 37967 45407
rect 34253 45305 34287 45339
rect 34345 45305 34379 45339
rect 37289 45237 37323 45271
rect 1869 44965 1903 44999
rect 1961 44693 1995 44727
rect 33885 44285 33919 44319
rect 33978 44285 34012 44319
rect 34161 44285 34195 44319
rect 34391 44285 34425 44319
rect 37473 44285 37507 44319
rect 37933 44285 37967 44319
rect 1869 44217 1903 44251
rect 34253 44217 34287 44251
rect 1961 44149 1995 44183
rect 34529 44149 34563 44183
rect 37289 44149 37323 44183
rect 37197 43809 37231 43843
rect 15669 43401 15703 43435
rect 16589 43333 16623 43367
rect 15301 43265 15335 43299
rect 16221 43265 16255 43299
rect 1869 43197 1903 43231
rect 15485 43197 15519 43231
rect 16405 43197 16439 43231
rect 37933 43197 37967 43231
rect 1961 43061 1995 43095
rect 1869 42721 1903 42755
rect 16129 42721 16163 42755
rect 16313 42721 16347 42755
rect 17509 42721 17543 42755
rect 17693 42721 17727 42755
rect 37381 42721 37415 42755
rect 15945 42653 15979 42687
rect 17325 42653 17359 42687
rect 1961 42517 1995 42551
rect 37197 42517 37231 42551
rect 16589 42313 16623 42347
rect 16221 42177 16255 42211
rect 16405 42109 16439 42143
rect 33793 42109 33827 42143
rect 33886 42109 33920 42143
rect 34161 42109 34195 42143
rect 34299 42109 34333 42143
rect 37289 42109 37323 42143
rect 37933 42109 37967 42143
rect 34069 42041 34103 42075
rect 34437 41973 34471 42007
rect 1869 41701 1903 41735
rect 34069 41701 34103 41735
rect 33793 41633 33827 41667
rect 33886 41633 33920 41667
rect 34161 41633 34195 41667
rect 34299 41633 34333 41667
rect 37381 41633 37415 41667
rect 2053 41497 2087 41531
rect 37197 41497 37231 41531
rect 34437 41429 34471 41463
rect 33701 41021 33735 41055
rect 33794 41021 33828 41055
rect 33977 41021 34011 41055
rect 34207 41021 34241 41055
rect 37289 41021 37323 41055
rect 37933 41021 37967 41055
rect 1869 40953 1903 40987
rect 2053 40953 2087 40987
rect 34069 40953 34103 40987
rect 34345 40885 34379 40919
rect 1869 40545 1903 40579
rect 17509 40545 17543 40579
rect 17325 40477 17359 40511
rect 2053 40409 2087 40443
rect 17693 40341 17727 40375
rect 17693 40137 17727 40171
rect 16037 40001 16071 40035
rect 16497 40001 16531 40035
rect 16865 40001 16899 40035
rect 18153 40001 18187 40035
rect 18521 40001 18555 40035
rect 15761 39933 15795 39967
rect 15853 39933 15887 39967
rect 16681 39933 16715 39967
rect 17325 39933 17359 39967
rect 17509 39933 17543 39967
rect 18337 39933 18371 39967
rect 33701 39933 33735 39967
rect 33794 39933 33828 39967
rect 33977 39933 34011 39967
rect 34207 39933 34241 39967
rect 37473 39933 37507 39967
rect 37933 39933 37967 39967
rect 34069 39865 34103 39899
rect 34345 39797 34379 39831
rect 37289 39797 37323 39831
rect 33977 39525 34011 39559
rect 1869 39457 1903 39491
rect 33701 39457 33735 39491
rect 33794 39457 33828 39491
rect 34069 39457 34103 39491
rect 34207 39457 34241 39491
rect 2053 39321 2087 39355
rect 34345 39253 34379 39287
rect 37289 39049 37323 39083
rect 37473 38845 37507 38879
rect 37933 38845 37967 38879
rect 1869 38777 1903 38811
rect 2053 38777 2087 38811
rect 34069 38505 34103 38539
rect 29009 38437 29043 38471
rect 33425 38437 33459 38471
rect 33241 38369 33275 38403
rect 33977 38369 34011 38403
rect 34621 38369 34655 38403
rect 37197 38369 37231 38403
rect 29193 38233 29227 38267
rect 34805 38165 34839 38199
rect 1869 37757 1903 37791
rect 33333 37757 33367 37791
rect 33426 37757 33460 37791
rect 33609 37757 33643 37791
rect 33701 37757 33735 37791
rect 33839 37757 33873 37791
rect 37933 37757 37967 37791
rect 2053 37689 2087 37723
rect 33149 37621 33183 37655
rect 33977 37621 34011 37655
rect 37197 37417 37231 37451
rect 1869 37281 1903 37315
rect 2053 37281 2087 37315
rect 37381 37281 37415 37315
rect 34529 36873 34563 36907
rect 33241 36669 33275 36703
rect 33334 36669 33368 36703
rect 33517 36669 33551 36703
rect 33747 36669 33781 36703
rect 37289 36669 37323 36703
rect 37933 36669 37967 36703
rect 33609 36601 33643 36635
rect 34437 36601 34471 36635
rect 33149 36533 33183 36567
rect 33885 36533 33919 36567
rect 28825 36329 28859 36363
rect 34529 36329 34563 36363
rect 37197 36329 37231 36363
rect 28733 36261 28767 36295
rect 33517 36261 33551 36295
rect 1869 36193 1903 36227
rect 33149 36193 33183 36227
rect 33241 36193 33275 36227
rect 33334 36193 33368 36227
rect 33609 36193 33643 36227
rect 33747 36193 33781 36227
rect 34437 36193 34471 36227
rect 37381 36193 37415 36227
rect 2053 36057 2087 36091
rect 33885 35989 33919 36023
rect 33149 35581 33183 35615
rect 33241 35581 33275 35615
rect 33334 35581 33368 35615
rect 33517 35581 33551 35615
rect 33747 35581 33781 35615
rect 37289 35581 37323 35615
rect 37933 35581 37967 35615
rect 1869 35513 1903 35547
rect 2053 35513 2087 35547
rect 28825 35513 28859 35547
rect 29009 35513 29043 35547
rect 33609 35513 33643 35547
rect 34437 35513 34471 35547
rect 33885 35445 33919 35479
rect 34529 35445 34563 35479
rect 33425 35173 33459 35207
rect 34345 35173 34379 35207
rect 33149 35105 33183 35139
rect 33242 35105 33276 35139
rect 33517 35105 33551 35139
rect 33655 35105 33689 35139
rect 32965 34901 32999 34935
rect 33793 34901 33827 34935
rect 34437 34901 34471 34935
rect 37289 34697 37323 34731
rect 2053 34493 2087 34527
rect 37473 34493 37507 34527
rect 37933 34493 37967 34527
rect 1869 34425 1903 34459
rect 1869 34017 1903 34051
rect 2053 33881 2087 33915
rect 37289 33609 37323 33643
rect 28733 33405 28767 33439
rect 33701 33405 33735 33439
rect 37473 33405 37507 33439
rect 37933 33405 37967 33439
rect 28917 33337 28951 33371
rect 33793 33269 33827 33303
rect 1869 32997 1903 33031
rect 37197 32929 37231 32963
rect 1961 32725 1995 32759
rect 32873 32521 32907 32555
rect 33057 32317 33091 32351
rect 33150 32317 33184 32351
rect 33333 32317 33367 32351
rect 33425 32317 33459 32351
rect 33563 32317 33597 32351
rect 37933 32317 37967 32351
rect 1869 32249 1903 32283
rect 2053 32249 2087 32283
rect 33701 32181 33735 32215
rect 33701 31977 33735 32011
rect 37197 31977 37231 32011
rect 33333 31909 33367 31943
rect 33425 31909 33459 31943
rect 33057 31841 33091 31875
rect 33150 31841 33184 31875
rect 33563 31841 33597 31875
rect 37381 31841 37415 31875
rect 32873 31773 32907 31807
rect 1869 31229 1903 31263
rect 32781 31229 32815 31263
rect 32965 31229 32999 31263
rect 33058 31229 33092 31263
rect 33333 31229 33367 31263
rect 33471 31229 33505 31263
rect 37289 31229 37323 31263
rect 37933 31229 37967 31263
rect 2053 31161 2087 31195
rect 33241 31161 33275 31195
rect 33609 31093 33643 31127
rect 37197 30889 37231 30923
rect 33425 30821 33459 30855
rect 1869 30753 1903 30787
rect 33057 30753 33091 30787
rect 33150 30753 33184 30787
rect 33333 30753 33367 30787
rect 33563 30753 33597 30787
rect 37381 30753 37415 30787
rect 1961 30549 1995 30583
rect 32873 30549 32907 30583
rect 33701 30549 33735 30583
rect 32873 30141 32907 30175
rect 32966 30141 33000 30175
rect 33149 30141 33183 30175
rect 33241 30141 33275 30175
rect 33379 30141 33413 30175
rect 37289 30141 37323 30175
rect 37933 30141 37967 30175
rect 32689 30005 32723 30039
rect 33517 30005 33551 30039
rect 1869 29733 1903 29767
rect 2053 29529 2087 29563
rect 37289 29257 37323 29291
rect 1869 29053 1903 29087
rect 37473 29053 37507 29087
rect 37933 29053 37967 29087
rect 2053 28985 2087 29019
rect 37289 28169 37323 28203
rect 32597 28033 32631 28067
rect 1869 27965 1903 27999
rect 26801 27965 26835 27999
rect 26893 27965 26927 27999
rect 27077 27965 27111 27999
rect 27537 27965 27571 27999
rect 32781 27965 32815 27999
rect 32874 27965 32908 27999
rect 33149 27965 33183 27999
rect 33287 27965 33321 27999
rect 37473 27965 37507 27999
rect 37933 27965 37967 27999
rect 2053 27897 2087 27931
rect 33057 27897 33091 27931
rect 33425 27829 33459 27863
rect 33701 27625 33735 27659
rect 27813 27557 27847 27591
rect 28018 27557 28052 27591
rect 33333 27557 33367 27591
rect 33425 27557 33459 27591
rect 1869 27489 1903 27523
rect 33057 27489 33091 27523
rect 33150 27489 33184 27523
rect 33563 27489 33597 27523
rect 37197 27489 37231 27523
rect 32873 27421 32907 27455
rect 1961 27285 1995 27319
rect 27997 27285 28031 27319
rect 28181 27285 28215 27319
rect 26801 27081 26835 27115
rect 31861 27081 31895 27115
rect 32597 27013 32631 27047
rect 25329 26945 25363 26979
rect 26893 26945 26927 26979
rect 30757 26945 30791 26979
rect 25237 26877 25271 26911
rect 26617 26877 26651 26911
rect 26709 26877 26743 26911
rect 30481 26877 30515 26911
rect 32781 26877 32815 26911
rect 32874 26877 32908 26911
rect 33149 26877 33183 26911
rect 33287 26877 33321 26911
rect 37933 26877 37967 26911
rect 1869 26809 1903 26843
rect 2053 26809 2087 26843
rect 33057 26809 33091 26843
rect 33425 26741 33459 26775
rect 32873 26537 32907 26571
rect 37197 26537 37231 26571
rect 33425 26469 33459 26503
rect 25329 26401 25363 26435
rect 33057 26401 33091 26435
rect 33150 26401 33184 26435
rect 33333 26401 33367 26435
rect 33563 26401 33597 26435
rect 34161 26401 34195 26435
rect 34254 26401 34288 26435
rect 34437 26401 34471 26435
rect 34529 26401 34563 26435
rect 34667 26401 34701 26435
rect 37381 26401 37415 26435
rect 25053 26333 25087 26367
rect 26433 26333 26467 26367
rect 33701 26265 33735 26299
rect 34805 26197 34839 26231
rect 33425 25925 33459 25959
rect 1869 25789 1903 25823
rect 32781 25789 32815 25823
rect 32874 25789 32908 25823
rect 33149 25789 33183 25823
rect 33287 25789 33321 25823
rect 35909 25789 35943 25823
rect 36001 25789 36035 25823
rect 36185 25789 36219 25823
rect 36277 25789 36311 25823
rect 37289 25789 37323 25823
rect 37933 25789 37967 25823
rect 2053 25721 2087 25755
rect 33057 25721 33091 25755
rect 32597 25653 32631 25687
rect 35725 25653 35759 25687
rect 37381 25449 37415 25483
rect 33333 25381 33367 25415
rect 33425 25381 33459 25415
rect 1869 25313 1903 25347
rect 33057 25313 33091 25347
rect 33150 25313 33184 25347
rect 33563 25313 33597 25347
rect 34345 25313 34379 25347
rect 34437 25313 34471 25347
rect 34621 25313 34655 25347
rect 34713 25313 34747 25347
rect 35357 25313 35391 25347
rect 35449 25313 35483 25347
rect 35633 25313 35667 25347
rect 35725 25313 35759 25347
rect 36369 25313 36403 25347
rect 36461 25313 36495 25347
rect 36645 25313 36679 25347
rect 36737 25313 36771 25347
rect 37197 25313 37231 25347
rect 2145 25245 2179 25279
rect 34161 25177 34195 25211
rect 32873 25109 32907 25143
rect 33701 25109 33735 25143
rect 35173 25109 35207 25143
rect 36185 25109 36219 25143
rect 27169 24769 27203 24803
rect 27077 24701 27111 24735
rect 27721 24701 27755 24735
rect 32873 24701 32907 24735
rect 32966 24701 33000 24735
rect 33241 24701 33275 24735
rect 33379 24701 33413 24735
rect 35909 24701 35943 24735
rect 36001 24701 36035 24735
rect 36185 24701 36219 24735
rect 36277 24701 36311 24735
rect 37289 24701 37323 24735
rect 37933 24701 37967 24735
rect 32689 24633 32723 24667
rect 33149 24633 33183 24667
rect 27813 24565 27847 24599
rect 33517 24565 33551 24599
rect 35725 24565 35759 24599
rect 28917 24361 28951 24395
rect 37197 24361 37231 24395
rect 29469 24293 29503 24327
rect 1869 24225 1903 24259
rect 27997 24225 28031 24259
rect 28089 24225 28123 24259
rect 28365 24225 28399 24259
rect 29193 24225 29227 24259
rect 33241 24225 33275 24259
rect 33333 24225 33367 24259
rect 33609 24225 33643 24259
rect 35541 24225 35575 24259
rect 35633 24225 35667 24259
rect 35817 24225 35851 24259
rect 35909 24225 35943 24259
rect 37381 24225 37415 24259
rect 29101 24157 29135 24191
rect 29561 24157 29595 24191
rect 35357 24157 35391 24191
rect 28273 24089 28307 24123
rect 33517 24089 33551 24123
rect 2145 24021 2179 24055
rect 27813 24021 27847 24055
rect 33057 24021 33091 24055
rect 2145 23817 2179 23851
rect 33609 23681 33643 23715
rect 27261 23613 27295 23647
rect 27445 23613 27479 23647
rect 27905 23613 27939 23647
rect 28089 23613 28123 23647
rect 33333 23613 33367 23647
rect 33425 23613 33459 23647
rect 33701 23613 33735 23647
rect 35909 23613 35943 23647
rect 36001 23613 36035 23647
rect 36185 23613 36219 23647
rect 36277 23613 36311 23647
rect 37289 23613 37323 23647
rect 37933 23613 37967 23647
rect 1869 23545 1903 23579
rect 27353 23477 27387 23511
rect 27997 23477 28031 23511
rect 33149 23477 33183 23511
rect 35725 23477 35759 23511
rect 29193 23273 29227 23307
rect 28058 23205 28092 23239
rect 33241 23137 33275 23171
rect 33333 23137 33367 23171
rect 33609 23137 33643 23171
rect 34253 23137 34287 23171
rect 34345 23137 34379 23171
rect 34621 23137 34655 23171
rect 35449 23137 35483 23171
rect 35541 23137 35575 23171
rect 35725 23137 35759 23171
rect 35817 23137 35851 23171
rect 27813 23069 27847 23103
rect 33517 23001 33551 23035
rect 34529 23001 34563 23035
rect 33057 22933 33091 22967
rect 34069 22933 34103 22967
rect 35265 22933 35299 22967
rect 32321 22729 32355 22763
rect 37473 22729 37507 22763
rect 33333 22661 33367 22695
rect 26433 22593 26467 22627
rect 34345 22593 34379 22627
rect 1869 22525 1903 22559
rect 26700 22525 26734 22559
rect 32045 22525 32079 22559
rect 32137 22525 32171 22559
rect 32413 22525 32447 22559
rect 33057 22525 33091 22559
rect 33149 22525 33183 22559
rect 33379 22525 33413 22559
rect 34070 22525 34104 22559
rect 34161 22525 34195 22559
rect 34437 22525 34471 22559
rect 35909 22525 35943 22559
rect 36001 22525 36035 22559
rect 36185 22525 36219 22559
rect 36277 22525 36311 22559
rect 37289 22525 37323 22559
rect 37933 22525 37967 22559
rect 2145 22389 2179 22423
rect 27813 22389 27847 22423
rect 31861 22389 31895 22423
rect 32873 22389 32907 22423
rect 33885 22389 33919 22423
rect 35725 22389 35759 22423
rect 1869 22117 1903 22151
rect 33241 22049 33275 22083
rect 33333 22049 33367 22083
rect 33609 22049 33643 22083
rect 35081 22049 35115 22083
rect 35173 22049 35207 22083
rect 35357 22049 35391 22083
rect 35449 22049 35483 22083
rect 36093 22049 36127 22083
rect 36185 22049 36219 22083
rect 36369 22049 36403 22083
rect 36461 22049 36495 22083
rect 34897 21981 34931 22015
rect 1961 21845 1995 21879
rect 33057 21845 33091 21879
rect 33517 21845 33551 21879
rect 35909 21845 35943 21879
rect 32689 21641 32723 21675
rect 37473 21641 37507 21675
rect 32137 21505 32171 21539
rect 34345 21505 34379 21539
rect 31861 21437 31895 21471
rect 31953 21437 31987 21471
rect 32229 21437 32263 21471
rect 32873 21437 32907 21471
rect 37289 21437 37323 21471
rect 37933 21437 37967 21471
rect 34161 21369 34195 21403
rect 31677 21301 31711 21335
rect 33302 21029 33336 21063
rect 1869 20961 1903 20995
rect 30481 20961 30515 20995
rect 30573 20961 30607 20995
rect 30849 20961 30883 20995
rect 31493 20961 31527 20995
rect 31585 20961 31619 20995
rect 31861 20961 31895 20995
rect 33057 20961 33091 20995
rect 35081 20961 35115 20995
rect 35173 20961 35207 20995
rect 35357 20961 35391 20995
rect 35449 20961 35483 20995
rect 36093 20961 36127 20995
rect 36185 20961 36219 20995
rect 36369 20961 36403 20995
rect 36461 20961 36495 20995
rect 37197 20961 37231 20995
rect 31309 20825 31343 20859
rect 35909 20825 35943 20859
rect 1961 20757 1995 20791
rect 30297 20757 30331 20791
rect 30757 20757 30791 20791
rect 31769 20757 31803 20791
rect 34437 20757 34471 20791
rect 34897 20757 34931 20791
rect 27261 20553 27295 20587
rect 28089 20485 28123 20519
rect 31125 20485 31159 20519
rect 33701 20485 33735 20519
rect 36001 20485 36035 20519
rect 31677 20417 31711 20451
rect 27445 20349 27479 20383
rect 27905 20349 27939 20383
rect 30849 20349 30883 20383
rect 30941 20349 30975 20383
rect 31217 20349 31251 20383
rect 31944 20349 31978 20383
rect 33517 20349 33551 20383
rect 34437 20349 34471 20383
rect 34529 20349 34563 20383
rect 34672 20349 34706 20383
rect 34805 20349 34839 20383
rect 35817 20349 35851 20383
rect 37933 20349 37967 20383
rect 1869 20281 1903 20315
rect 28641 20281 28675 20315
rect 28825 20281 28859 20315
rect 1961 20213 1995 20247
rect 30665 20213 30699 20247
rect 33057 20213 33091 20247
rect 34253 20213 34287 20247
rect 34897 20009 34931 20043
rect 37381 20009 37415 20043
rect 36185 19941 36219 19975
rect 25697 19873 25731 19907
rect 25973 19873 26007 19907
rect 27905 19873 27939 19907
rect 28733 19873 28767 19907
rect 28825 19873 28859 19907
rect 29101 19873 29135 19907
rect 29745 19873 29779 19907
rect 29837 19873 29871 19907
rect 30113 19873 30147 19907
rect 30757 19873 30791 19907
rect 30849 19873 30883 19907
rect 31125 19873 31159 19907
rect 31585 19873 31619 19907
rect 33057 19873 33091 19907
rect 33324 19873 33358 19907
rect 35081 19873 35115 19907
rect 35173 19873 35207 19907
rect 35357 19873 35391 19907
rect 35449 19873 35483 19907
rect 36001 19873 36035 19907
rect 37197 19873 37231 19907
rect 26433 19805 26467 19839
rect 29561 19805 29595 19839
rect 25789 19737 25823 19771
rect 28089 19737 28123 19771
rect 30021 19737 30055 19771
rect 31769 19737 31803 19771
rect 34437 19737 34471 19771
rect 28549 19669 28583 19703
rect 29009 19669 29043 19703
rect 30573 19669 30607 19703
rect 31033 19669 31067 19703
rect 24133 19465 24167 19499
rect 27077 19465 27111 19499
rect 31861 19397 31895 19431
rect 26617 19329 26651 19363
rect 32321 19329 32355 19363
rect 1869 19261 1903 19295
rect 23949 19261 23983 19295
rect 24133 19261 24167 19295
rect 26157 19261 26191 19295
rect 26985 19261 27019 19295
rect 30481 19261 30515 19295
rect 30748 19261 30782 19295
rect 34161 19261 34195 19295
rect 34348 19261 34382 19295
rect 34483 19261 34517 19295
rect 34621 19261 34655 19295
rect 34713 19261 34747 19295
rect 35725 19261 35759 19295
rect 37289 19261 37323 19295
rect 37933 19261 37967 19295
rect 2053 19193 2087 19227
rect 25973 19193 26007 19227
rect 27813 19193 27847 19227
rect 32588 19193 32622 19227
rect 24317 19125 24351 19159
rect 29285 19125 29319 19159
rect 33701 19125 33735 19159
rect 35909 19125 35943 19159
rect 29285 18921 29319 18955
rect 30757 18921 30791 18955
rect 31953 18921 31987 18955
rect 34437 18921 34471 18955
rect 37381 18921 37415 18955
rect 24317 18853 24351 18887
rect 1869 18785 1903 18819
rect 26341 18785 26375 18819
rect 26433 18785 26467 18819
rect 26709 18785 26743 18819
rect 27813 18785 27847 18819
rect 28089 18785 28123 18819
rect 28273 18785 28307 18819
rect 28457 18785 28491 18819
rect 24685 18717 24719 18751
rect 25053 18717 25087 18751
rect 28641 18717 28675 18751
rect 24482 18649 24516 18683
rect 29644 18853 29678 18887
rect 31493 18853 31527 18887
rect 33302 18853 33336 18887
rect 36001 18853 36035 18887
rect 36185 18853 36219 18887
rect 31309 18785 31343 18819
rect 32137 18785 32171 18819
rect 33057 18785 33091 18819
rect 35081 18785 35115 18819
rect 35173 18785 35207 18819
rect 35357 18785 35391 18819
rect 35449 18785 35483 18819
rect 37197 18785 37231 18819
rect 29377 18717 29411 18751
rect 34897 18649 34931 18683
rect 1961 18581 1995 18615
rect 24593 18581 24627 18615
rect 26157 18581 26191 18615
rect 26617 18581 26651 18615
rect 29285 18581 29319 18615
rect 26617 18377 26651 18411
rect 28457 18377 28491 18411
rect 29469 18309 29503 18343
rect 35909 18309 35943 18343
rect 25237 18241 25271 18275
rect 32321 18241 32355 18275
rect 27077 18173 27111 18207
rect 29193 18173 29227 18207
rect 29285 18173 29319 18207
rect 29561 18173 29595 18207
rect 30481 18173 30515 18207
rect 32577 18173 32611 18207
rect 34345 18173 34379 18207
rect 34437 18173 34471 18207
rect 34621 18173 34655 18207
rect 34713 18173 34747 18207
rect 35725 18173 35759 18207
rect 37289 18173 37323 18207
rect 37933 18173 37967 18207
rect 25504 18105 25538 18139
rect 27322 18105 27356 18139
rect 30748 18105 30782 18139
rect 34161 18105 34195 18139
rect 29009 18037 29043 18071
rect 31861 18037 31895 18071
rect 33701 18037 33735 18071
rect 26801 17833 26835 17867
rect 29193 17833 29227 17867
rect 31493 17833 31527 17867
rect 34437 17833 34471 17867
rect 1869 17765 1903 17799
rect 23848 17765 23882 17799
rect 25688 17765 25722 17799
rect 28080 17765 28114 17799
rect 29920 17765 29954 17799
rect 33302 17765 33336 17799
rect 23581 17697 23615 17731
rect 31677 17697 31711 17731
rect 31769 17697 31803 17731
rect 32045 17697 32079 17731
rect 33057 17697 33091 17731
rect 35081 17697 35115 17731
rect 35173 17697 35207 17731
rect 35369 17697 35403 17731
rect 35459 17697 35493 17731
rect 25421 17629 25455 17663
rect 27813 17629 27847 17663
rect 29653 17629 29687 17663
rect 24961 17561 24995 17595
rect 34897 17561 34931 17595
rect 1961 17493 1995 17527
rect 31033 17493 31067 17527
rect 31953 17493 31987 17527
rect 26617 17289 26651 17323
rect 28457 17289 28491 17323
rect 31861 17289 31895 17323
rect 37473 17289 37507 17323
rect 25237 17153 25271 17187
rect 29469 17153 29503 17187
rect 33793 17153 33827 17187
rect 24317 17085 24351 17119
rect 27077 17085 27111 17119
rect 29193 17085 29227 17119
rect 29331 17085 29365 17119
rect 29561 17085 29595 17119
rect 30481 17085 30515 17119
rect 32321 17085 32355 17119
rect 33977 17085 34011 17119
rect 34069 17085 34103 17119
rect 34253 17085 34287 17119
rect 34345 17085 34379 17119
rect 37289 17085 37323 17119
rect 37933 17085 37967 17119
rect 1869 17017 1903 17051
rect 24133 17017 24167 17051
rect 25482 17017 25516 17051
rect 27322 17017 27356 17051
rect 30726 17017 30760 17051
rect 1961 16949 1995 16983
rect 29009 16949 29043 16983
rect 32505 16949 32539 16983
rect 26433 16745 26467 16779
rect 29193 16745 29227 16779
rect 31033 16745 31067 16779
rect 25298 16677 25332 16711
rect 28080 16677 28114 16711
rect 29920 16677 29954 16711
rect 31493 16677 31527 16711
rect 23581 16609 23615 16643
rect 24041 16609 24075 16643
rect 24225 16609 24259 16643
rect 24317 16609 24351 16643
rect 24593 16609 24627 16643
rect 27813 16609 27847 16643
rect 29653 16609 29687 16643
rect 31677 16609 31711 16643
rect 31769 16609 31803 16643
rect 32045 16609 32079 16643
rect 33701 16609 33735 16643
rect 33793 16609 33827 16643
rect 33977 16609 34011 16643
rect 34069 16609 34103 16643
rect 34713 16609 34747 16643
rect 34805 16609 34839 16643
rect 34989 16609 35023 16643
rect 35081 16609 35115 16643
rect 25053 16541 25087 16575
rect 34529 16541 34563 16575
rect 33517 16473 33551 16507
rect 23397 16405 23431 16439
rect 24501 16405 24535 16439
rect 31953 16405 31987 16439
rect 23949 16201 23983 16235
rect 29561 16201 29595 16235
rect 32229 16201 32263 16235
rect 33241 16201 33275 16235
rect 37473 16201 37507 16235
rect 34529 16133 34563 16167
rect 25605 16065 25639 16099
rect 27537 16065 27571 16099
rect 30941 16065 30975 16099
rect 1869 15997 1903 16031
rect 22569 15997 22603 16031
rect 25872 15997 25906 16031
rect 27804 15997 27838 16031
rect 29377 15997 29411 16031
rect 30665 15997 30699 16031
rect 30757 15997 30791 16031
rect 31033 15997 31067 16031
rect 32413 15997 32447 16031
rect 32505 15997 32539 16031
rect 32648 15997 32682 16031
rect 32781 15997 32815 16031
rect 33425 15997 33459 16031
rect 33517 15997 33551 16031
rect 33701 15997 33735 16031
rect 33793 15997 33827 16031
rect 37289 15997 37323 16031
rect 37933 15997 37967 16031
rect 22836 15929 22870 15963
rect 31585 15929 31619 15963
rect 31769 15929 31803 15963
rect 34345 15929 34379 15963
rect 1961 15861 1995 15895
rect 26985 15861 27019 15895
rect 28917 15861 28951 15895
rect 30481 15861 30515 15895
rect 22753 15657 22787 15691
rect 28080 15589 28114 15623
rect 1869 15521 1903 15555
rect 22937 15521 22971 15555
rect 23581 15521 23615 15555
rect 23673 15521 23707 15555
rect 23949 15521 23983 15555
rect 24593 15521 24627 15555
rect 24685 15521 24719 15555
rect 24961 15521 24995 15555
rect 25421 15521 25455 15555
rect 25688 15521 25722 15555
rect 29837 15521 29871 15555
rect 29929 15521 29963 15555
rect 30205 15521 30239 15555
rect 30849 15521 30883 15555
rect 30987 15521 31021 15555
rect 31217 15521 31251 15555
rect 33333 15521 33367 15555
rect 33425 15521 33459 15555
rect 33609 15521 33643 15555
rect 33701 15521 33735 15555
rect 34345 15521 34379 15555
rect 34437 15521 34471 15555
rect 34621 15521 34655 15555
rect 34713 15521 34747 15555
rect 37197 15521 37231 15555
rect 27813 15453 27847 15487
rect 30113 15453 30147 15487
rect 29653 15385 29687 15419
rect 31125 15385 31159 15419
rect 1961 15317 1995 15351
rect 23397 15317 23431 15351
rect 23857 15317 23891 15351
rect 24409 15317 24443 15351
rect 24869 15317 24903 15351
rect 26801 15317 26835 15351
rect 29193 15317 29227 15351
rect 30665 15317 30699 15351
rect 33149 15317 33183 15351
rect 34161 15317 34195 15351
rect 33977 15113 34011 15147
rect 35909 15113 35943 15147
rect 23213 15045 23247 15079
rect 24225 15045 24259 15079
rect 29469 15045 29503 15079
rect 25237 14977 25271 15011
rect 32965 14977 32999 15011
rect 22937 14909 22971 14943
rect 23029 14909 23063 14943
rect 23305 14909 23339 14943
rect 23949 14909 23983 14943
rect 24041 14909 24075 14943
rect 24317 14909 24351 14943
rect 27261 14909 27295 14943
rect 28089 14909 28123 14943
rect 28457 14909 28491 14943
rect 29193 14909 29227 14943
rect 29285 14909 29319 14943
rect 29561 14909 29595 14943
rect 32137 14909 32171 14943
rect 32229 14909 32263 14943
rect 32413 14909 32447 14943
rect 32505 14909 32539 14943
rect 33149 14909 33183 14943
rect 33241 14909 33275 14943
rect 33425 14909 33459 14943
rect 33517 14909 33551 14943
rect 34161 14909 34195 14943
rect 34253 14909 34287 14943
rect 34437 14909 34471 14943
rect 34529 14909 34563 14943
rect 37933 14909 37967 14943
rect 25504 14841 25538 14875
rect 35817 14841 35851 14875
rect 22753 14773 22787 14807
rect 23765 14773 23799 14807
rect 26617 14773 26651 14807
rect 29009 14773 29043 14807
rect 31953 14773 31987 14807
rect 23489 14569 23523 14603
rect 37381 14569 37415 14603
rect 1869 14501 1903 14535
rect 28080 14501 28114 14535
rect 29745 14501 29779 14535
rect 23397 14433 23431 14467
rect 24041 14433 24075 14467
rect 24308 14433 24342 14467
rect 26525 14433 26559 14467
rect 26617 14433 26651 14467
rect 26893 14433 26927 14467
rect 33057 14433 33091 14467
rect 33241 14433 33275 14467
rect 33333 14433 33367 14467
rect 33517 14433 33551 14467
rect 33609 14433 33643 14467
rect 34253 14433 34287 14467
rect 34345 14433 34379 14467
rect 34529 14433 34563 14467
rect 34621 14433 34655 14467
rect 37197 14433 37231 14467
rect 27813 14365 27847 14399
rect 25421 14297 25455 14331
rect 1961 14229 1995 14263
rect 26341 14229 26375 14263
rect 26801 14229 26835 14263
rect 29193 14229 29227 14263
rect 29837 14229 29871 14263
rect 34069 14229 34103 14263
rect 2145 14025 2179 14059
rect 24317 14025 24351 14059
rect 28457 14025 28491 14059
rect 29285 14025 29319 14059
rect 32873 14025 32907 14059
rect 34161 14025 34195 14059
rect 34805 14025 34839 14059
rect 38117 14025 38151 14059
rect 26617 13957 26651 13991
rect 37473 13957 37507 13991
rect 22937 13889 22971 13923
rect 28917 13889 28951 13923
rect 1869 13821 1903 13855
rect 23204 13821 23238 13855
rect 25237 13821 25271 13855
rect 25493 13821 25527 13855
rect 27077 13821 27111 13855
rect 27344 13821 27378 13855
rect 29101 13821 29135 13855
rect 33057 13821 33091 13855
rect 33149 13821 33183 13855
rect 33333 13821 33367 13855
rect 33425 13821 33459 13855
rect 33977 13821 34011 13855
rect 34621 13821 34655 13855
rect 37289 13821 37323 13855
rect 37933 13821 37967 13855
rect 25881 13481 25915 13515
rect 29193 13481 29227 13515
rect 37381 13481 37415 13515
rect 24746 13413 24780 13447
rect 1869 13345 1903 13379
rect 22569 13345 22603 13379
rect 22836 13345 22870 13379
rect 26525 13345 26559 13379
rect 26617 13345 26651 13379
rect 26893 13345 26927 13379
rect 28080 13345 28114 13379
rect 37197 13345 37231 13379
rect 24501 13277 24535 13311
rect 27813 13277 27847 13311
rect 26801 13209 26835 13243
rect 2145 13141 2179 13175
rect 23949 13141 23983 13175
rect 26341 13141 26375 13175
rect 20913 12937 20947 12971
rect 26617 12937 26651 12971
rect 28825 12937 28859 12971
rect 37473 12937 37507 12971
rect 38117 12937 38151 12971
rect 23397 12869 23431 12903
rect 21557 12801 21591 12835
rect 25237 12801 25271 12835
rect 27537 12801 27571 12835
rect 21097 12733 21131 12767
rect 21281 12733 21315 12767
rect 21419 12733 21453 12767
rect 22017 12733 22051 12767
rect 22284 12733 22318 12767
rect 25504 12733 25538 12767
rect 27261 12733 27295 12767
rect 27353 12733 27387 12767
rect 27629 12733 27663 12767
rect 28733 12733 28767 12767
rect 37289 12733 37323 12767
rect 37933 12733 37967 12767
rect 21189 12665 21223 12699
rect 27077 12597 27111 12631
rect 23949 12393 23983 12427
rect 26341 12393 26375 12427
rect 22814 12325 22848 12359
rect 24768 12325 24802 12359
rect 1869 12257 1903 12291
rect 22569 12257 22603 12291
rect 24501 12257 24535 12291
rect 26525 12257 26559 12291
rect 2145 12121 2179 12155
rect 25881 12053 25915 12087
rect 37473 11849 37507 11883
rect 38117 11781 38151 11815
rect 22293 11713 22327 11747
rect 22560 11645 22594 11679
rect 37289 11645 37323 11679
rect 37933 11645 37967 11679
rect 38945 11645 38979 11679
rect 1869 11577 1903 11611
rect 2145 11509 2179 11543
rect 23673 11509 23707 11543
rect 37381 11305 37415 11339
rect 22836 11237 22870 11271
rect 22569 11169 22603 11203
rect 30757 11169 30791 11203
rect 31242 11169 31276 11203
rect 37197 11169 37231 11203
rect 31033 11101 31067 11135
rect 31125 11101 31159 11135
rect 23949 11033 23983 11067
rect 31401 11033 31435 11067
rect 38945 11033 38979 11067
rect 2145 10761 2179 10795
rect 37473 10761 37507 10795
rect 38117 10693 38151 10727
rect 1869 10557 1903 10591
rect 37289 10557 37323 10591
rect 37933 10557 37967 10591
rect 1869 10081 1903 10115
rect 30389 10081 30423 10115
rect 2145 9877 2179 9911
rect 30573 9877 30607 9911
rect 38117 9605 38151 9639
rect 37289 9469 37323 9503
rect 37933 9469 37967 9503
rect 37473 9333 37507 9367
rect 37381 9129 37415 9163
rect 1869 8993 1903 9027
rect 37197 8993 37231 9027
rect 2145 8789 2179 8823
rect 37473 8585 37507 8619
rect 38117 8517 38151 8551
rect 37289 8381 37323 8415
rect 37933 8381 37967 8415
rect 1869 8313 1903 8347
rect 2237 8313 2271 8347
rect 29469 8041 29503 8075
rect 29469 7905 29503 7939
rect 29653 7905 29687 7939
rect 29837 7905 29871 7939
rect 30113 7905 30147 7939
rect 2145 7497 2179 7531
rect 37473 7497 37507 7531
rect 38117 7429 38151 7463
rect 1869 7293 1903 7327
rect 37289 7293 37323 7327
rect 37933 7293 37967 7327
rect 1869 6817 1903 6851
rect 23673 6817 23707 6851
rect 24593 6817 24627 6851
rect 37197 6817 37231 6851
rect 2145 6749 2179 6783
rect 37381 6681 37415 6715
rect 36829 6409 36863 6443
rect 37473 6409 37507 6443
rect 38117 6341 38151 6375
rect 36645 6205 36679 6239
rect 37289 6205 37323 6239
rect 37933 6205 37967 6239
rect 38945 6205 38979 6239
rect 35449 5865 35483 5899
rect 36093 5865 36127 5899
rect 36737 5865 36771 5899
rect 1869 5797 1903 5831
rect 3893 5729 3927 5763
rect 34713 5729 34747 5763
rect 35265 5729 35299 5763
rect 35909 5729 35943 5763
rect 36553 5729 36587 5763
rect 37197 5729 37231 5763
rect 2145 5593 2179 5627
rect 3709 5593 3743 5627
rect 37381 5593 37415 5627
rect 3249 5525 3283 5559
rect 34529 5525 34563 5559
rect 38945 5525 38979 5559
rect 2145 5321 2179 5355
rect 34805 5321 34839 5355
rect 36737 5321 36771 5355
rect 36093 5253 36127 5287
rect 2973 5185 3007 5219
rect 34621 5117 34655 5151
rect 35909 5117 35943 5151
rect 36553 5117 36587 5151
rect 37197 5117 37231 5151
rect 1869 5049 1903 5083
rect 2789 5049 2823 5083
rect 37933 5049 37967 5083
rect 38117 5049 38151 5083
rect 37381 4981 37415 5015
rect 34713 4777 34747 4811
rect 36645 4777 36679 4811
rect 2237 4709 2271 4743
rect 2789 4709 2823 4743
rect 3525 4709 3559 4743
rect 35265 4709 35299 4743
rect 37197 4709 37231 4743
rect 1869 4641 1903 4675
rect 4353 4641 4387 4675
rect 4997 4641 5031 4675
rect 32137 4641 32171 4675
rect 33793 4641 33827 4675
rect 34529 4641 34563 4675
rect 36461 4641 36495 4675
rect 2973 4505 3007 4539
rect 31953 4505 31987 4539
rect 37381 4505 37415 4539
rect 3617 4437 3651 4471
rect 4813 4437 4847 4471
rect 33609 4437 33643 4471
rect 35357 4437 35391 4471
rect 2881 4233 2915 4267
rect 23489 4233 23523 4267
rect 5181 4165 5215 4199
rect 26157 4165 26191 4199
rect 2145 4097 2179 4131
rect 4353 4029 4387 4063
rect 4997 4029 5031 4063
rect 5641 4029 5675 4063
rect 6561 4029 6595 4063
rect 11897 4029 11931 4063
rect 12817 4029 12851 4063
rect 14749 4029 14783 4063
rect 18705 4029 18739 4063
rect 20177 4029 20211 4063
rect 22017 4029 22051 4063
rect 23029 4029 23063 4063
rect 23673 4029 23707 4063
rect 24317 4029 24351 4063
rect 25421 4029 25455 4063
rect 25973 4029 26007 4063
rect 26801 4029 26835 4063
rect 27445 4029 27479 4063
rect 28917 4029 28951 4063
rect 29561 4029 29595 4063
rect 30665 4029 30699 4063
rect 31309 4029 31343 4063
rect 31953 4029 31987 4063
rect 32781 4029 32815 4063
rect 33425 4029 33459 4063
rect 34253 4029 34287 4063
rect 35909 4029 35943 4063
rect 37933 4029 37967 4063
rect 1869 3961 1903 3995
rect 2789 3961 2823 3995
rect 16773 3961 16807 3995
rect 17693 3961 17727 3995
rect 36461 3961 36495 3995
rect 37197 3961 37231 3995
rect 38117 3961 38151 3995
rect 4445 3893 4479 3927
rect 11989 3893 12023 3927
rect 12909 3893 12943 3927
rect 14933 3893 14967 3927
rect 16865 3893 16899 3927
rect 17785 3893 17819 3927
rect 18797 3893 18831 3927
rect 19993 3893 20027 3927
rect 21833 3893 21867 3927
rect 22845 3893 22879 3927
rect 24133 3893 24167 3927
rect 25237 3893 25271 3927
rect 26617 3893 26651 3927
rect 27261 3893 27295 3927
rect 28733 3893 28767 3927
rect 29377 3893 29411 3927
rect 30481 3893 30515 3927
rect 31125 3893 31159 3927
rect 31769 3893 31803 3927
rect 32597 3893 32631 3927
rect 33609 3893 33643 3927
rect 34069 3893 34103 3927
rect 35725 3893 35759 3927
rect 36553 3893 36587 3927
rect 37289 3893 37323 3927
rect 3525 3689 3559 3723
rect 8401 3689 8435 3723
rect 18153 3689 18187 3723
rect 19441 3689 19475 3723
rect 2237 3621 2271 3655
rect 4353 3621 4387 3655
rect 6929 3621 6963 3655
rect 8953 3621 8987 3655
rect 10885 3621 10919 3655
rect 12495 3621 12529 3655
rect 13369 3621 13403 3655
rect 14105 3621 14139 3655
rect 29469 3621 29503 3655
rect 30389 3621 30423 3655
rect 35541 3621 35575 3655
rect 36277 3621 36311 3655
rect 37197 3621 37231 3655
rect 1869 3553 1903 3587
rect 3433 3553 3467 3587
rect 5089 3553 5123 3587
rect 5733 3553 5767 3587
rect 7573 3553 7607 3587
rect 8217 3553 8251 3587
rect 9597 3553 9631 3587
rect 13093 3553 13127 3587
rect 14841 3553 14875 3587
rect 15761 3553 15795 3587
rect 17969 3553 18003 3587
rect 19257 3553 19291 3587
rect 20085 3553 20119 3587
rect 20729 3553 20763 3587
rect 21557 3553 21591 3587
rect 22569 3553 22603 3587
rect 23213 3553 23247 3587
rect 24041 3553 24075 3587
rect 24593 3553 24627 3587
rect 25513 3553 25547 3587
rect 26433 3553 26467 3587
rect 27905 3553 27939 3587
rect 28733 3553 28767 3587
rect 31033 3553 31067 3587
rect 31677 3553 31711 3587
rect 33609 3553 33643 3587
rect 34345 3553 34379 3587
rect 12081 3485 12115 3519
rect 4537 3417 4571 3451
rect 9781 3417 9815 3451
rect 30573 3417 30607 3451
rect 31217 3417 31251 3451
rect 31861 3417 31895 3451
rect 35725 3417 35759 3451
rect 37381 3417 37415 3451
rect 5181 3349 5215 3383
rect 7021 3349 7055 3383
rect 9045 3349 9079 3383
rect 10977 3349 11011 3383
rect 12449 3349 12483 3383
rect 12633 3349 12667 3383
rect 14197 3349 14231 3383
rect 14933 3349 14967 3383
rect 15853 3349 15887 3383
rect 20177 3349 20211 3383
rect 20913 3349 20947 3383
rect 21373 3349 21407 3383
rect 22753 3349 22787 3383
rect 23397 3349 23431 3383
rect 23857 3349 23891 3383
rect 24685 3349 24719 3383
rect 25605 3349 25639 3383
rect 26617 3349 26651 3383
rect 27997 3349 28031 3383
rect 28549 3349 28583 3383
rect 29561 3349 29595 3383
rect 33701 3349 33735 3383
rect 34437 3349 34471 3383
rect 36369 3349 36403 3383
rect 2145 3145 2179 3179
rect 3065 3145 3099 3179
rect 7389 3145 7423 3179
rect 9689 3145 9723 3179
rect 16497 3145 16531 3179
rect 20269 3145 20303 3179
rect 25513 3145 25547 3179
rect 25881 3145 25915 3179
rect 27813 3145 27847 3179
rect 30849 3145 30883 3179
rect 30941 3145 30975 3179
rect 35909 3145 35943 3179
rect 20158 3077 20192 3111
rect 25375 3077 25409 3111
rect 27702 3077 27736 3111
rect 34437 3077 34471 3111
rect 34805 3077 34839 3111
rect 4813 3009 4847 3043
rect 6193 3009 6227 3043
rect 11437 3009 11471 3043
rect 12357 3009 12391 3043
rect 13277 3009 13311 3043
rect 15577 3009 15611 3043
rect 17601 3009 17635 3043
rect 18613 3009 18647 3043
rect 20361 3009 20395 3043
rect 25602 3009 25636 3043
rect 27905 3009 27939 3043
rect 28273 3009 28307 3043
rect 30481 3009 30515 3043
rect 31033 3009 31067 3043
rect 2789 2941 2823 2975
rect 4629 2941 4663 2975
rect 5917 2941 5951 2975
rect 7205 2941 7239 2975
rect 8033 2941 8067 2975
rect 9505 2941 9539 2975
rect 10333 2941 10367 2975
rect 11161 2941 11195 2975
rect 12081 2941 12115 2975
rect 13093 2941 13127 2975
rect 14749 2941 14783 2975
rect 15393 2941 15427 2975
rect 16313 2941 16347 2975
rect 17325 2941 17359 2975
rect 18337 2941 18371 2975
rect 19993 2941 20027 2975
rect 21465 2941 21499 2975
rect 22753 2941 22787 2975
rect 23581 2941 23615 2975
rect 25237 2941 25271 2975
rect 26525 2941 26559 2975
rect 27537 2941 27571 2975
rect 28825 2941 28859 2975
rect 31401 2941 31435 2975
rect 31953 2941 31987 2975
rect 32689 2941 32723 2975
rect 33425 2941 33459 2975
rect 34437 2941 34471 2975
rect 35725 2941 35759 2975
rect 37933 2941 37967 2975
rect 1869 2873 1903 2907
rect 21281 2873 21315 2907
rect 22017 2873 22051 2907
rect 34621 2873 34655 2907
rect 36645 2873 36679 2907
rect 38117 2873 38151 2907
rect 8125 2805 8159 2839
rect 10425 2805 10459 2839
rect 14933 2805 14967 2839
rect 20637 2805 20671 2839
rect 22109 2805 22143 2839
rect 22845 2805 22879 2839
rect 23673 2805 23707 2839
rect 26617 2805 26651 2839
rect 28917 2805 28951 2839
rect 32045 2805 32079 2839
rect 32781 2805 32815 2839
rect 33517 2805 33551 2839
rect 36737 2805 36771 2839
rect 3065 2601 3099 2635
rect 11253 2601 11287 2635
rect 23121 2601 23155 2635
rect 24593 2601 24627 2635
rect 28457 2601 28491 2635
rect 35633 2601 35667 2635
rect 36461 2601 36495 2635
rect 1869 2533 1903 2567
rect 5825 2533 5859 2567
rect 8493 2533 8527 2567
rect 10425 2533 10459 2567
rect 13737 2533 13771 2567
rect 16405 2533 16439 2567
rect 26341 2533 26375 2567
rect 32505 2533 32539 2567
rect 34069 2533 34103 2567
rect 2789 2465 2823 2499
rect 4261 2465 4295 2499
rect 5549 2465 5583 2499
rect 6929 2465 6963 2499
rect 8217 2465 8251 2499
rect 10149 2465 10183 2499
rect 11069 2465 11103 2499
rect 12265 2465 12299 2499
rect 13369 2465 13403 2499
rect 14933 2465 14967 2499
rect 16037 2465 16071 2499
rect 17693 2465 17727 2499
rect 18245 2465 18279 2499
rect 18981 2465 19015 2499
rect 20269 2465 20303 2499
rect 21189 2465 21223 2499
rect 21465 2465 21499 2499
rect 23029 2465 23063 2499
rect 24409 2465 24443 2499
rect 26065 2465 26099 2499
rect 27077 2465 27111 2499
rect 28273 2465 28307 2499
rect 29561 2465 29595 2499
rect 31033 2465 31067 2499
rect 33701 2465 33735 2499
rect 34529 2465 34563 2499
rect 37749 2533 37783 2567
rect 36369 2465 36403 2499
rect 37473 2465 37507 2499
rect 4445 2397 4479 2431
rect 7113 2397 7147 2431
rect 12449 2397 12483 2431
rect 15117 2397 15151 2431
rect 20453 2397 20487 2431
rect 29745 2397 29779 2431
rect 35633 2397 35667 2431
rect 27261 2329 27295 2363
rect 32689 2329 32723 2363
rect 2145 2261 2179 2295
rect 19257 2261 19291 2295
rect 31125 2261 31159 2295
rect 34713 2261 34747 2295
<< metal1 >>
rect 4706 118192 4712 118244
rect 4764 118192 4770 118244
rect 34790 118192 34796 118244
rect 34848 118192 34854 118244
rect 4724 117972 4752 118192
rect 34808 118040 34836 118192
rect 34790 117988 34796 118040
rect 34848 117988 34854 118040
rect 4706 117920 4712 117972
rect 4764 117920 4770 117972
rect 25038 117648 25044 117700
rect 25096 117688 25102 117700
rect 29270 117688 29276 117700
rect 25096 117660 29276 117688
rect 25096 117648 25102 117660
rect 29270 117648 29276 117660
rect 29328 117648 29334 117700
rect 34698 117648 34704 117700
rect 34756 117688 34762 117700
rect 34974 117688 34980 117700
rect 34756 117660 34980 117688
rect 34756 117648 34762 117660
rect 34974 117648 34980 117660
rect 35032 117648 35038 117700
rect 24394 117580 24400 117632
rect 24452 117620 24458 117632
rect 28810 117620 28816 117632
rect 24452 117592 28816 117620
rect 24452 117580 24458 117592
rect 28810 117580 28816 117592
rect 28868 117580 28874 117632
rect 1104 117530 38824 117552
rect 1104 117478 4246 117530
rect 4298 117478 4310 117530
rect 4362 117478 4374 117530
rect 4426 117478 4438 117530
rect 4490 117478 34966 117530
rect 35018 117478 35030 117530
rect 35082 117478 35094 117530
rect 35146 117478 35158 117530
rect 35210 117478 38824 117530
rect 1104 117456 38824 117478
rect 290 117376 296 117428
rect 348 117416 354 117428
rect 2685 117419 2743 117425
rect 2685 117416 2697 117419
rect 348 117388 2697 117416
rect 348 117376 354 117388
rect 2685 117385 2697 117388
rect 2731 117385 2743 117419
rect 2685 117379 2743 117385
rect 2958 117376 2964 117428
rect 3016 117416 3022 117428
rect 3016 117388 7328 117416
rect 3016 117376 3022 117388
rect 1210 117308 1216 117360
rect 1268 117348 1274 117360
rect 7193 117351 7251 117357
rect 7193 117348 7205 117351
rect 1268 117320 4660 117348
rect 1268 117308 1274 117320
rect 106 117240 112 117292
rect 164 117280 170 117292
rect 2041 117283 2099 117289
rect 2041 117280 2053 117283
rect 164 117252 2053 117280
rect 164 117240 170 117252
rect 2041 117249 2053 117252
rect 2087 117249 2099 117283
rect 4525 117283 4583 117289
rect 4525 117280 4537 117283
rect 2041 117243 2099 117249
rect 2746 117252 4537 117280
rect 750 117172 756 117224
rect 808 117212 814 117224
rect 2746 117212 2774 117252
rect 4525 117249 4537 117252
rect 4571 117249 4583 117283
rect 4632 117280 4660 117320
rect 6840 117320 7205 117348
rect 5997 117283 6055 117289
rect 5997 117280 6009 117283
rect 4632 117252 6009 117280
rect 4525 117243 4583 117249
rect 5997 117249 6009 117252
rect 6043 117249 6055 117283
rect 5997 117243 6055 117249
rect 6178 117240 6184 117292
rect 6236 117280 6242 117292
rect 6840 117280 6868 117320
rect 7193 117317 7205 117320
rect 7239 117317 7251 117351
rect 7193 117311 7251 117317
rect 6236 117252 6868 117280
rect 7300 117280 7328 117388
rect 11146 117376 11152 117428
rect 11204 117416 11210 117428
rect 12437 117419 12495 117425
rect 12437 117416 12449 117419
rect 11204 117388 12449 117416
rect 11204 117376 11210 117388
rect 12437 117385 12449 117388
rect 12483 117385 12495 117419
rect 12437 117379 12495 117385
rect 17402 117376 17408 117428
rect 17460 117416 17466 117428
rect 17954 117416 17960 117428
rect 17460 117388 17960 117416
rect 17460 117376 17466 117388
rect 17954 117376 17960 117388
rect 18012 117376 18018 117428
rect 18138 117376 18144 117428
rect 18196 117416 18202 117428
rect 18196 117388 19380 117416
rect 18196 117376 18202 117388
rect 16298 117308 16304 117360
rect 16356 117348 16362 117360
rect 16482 117348 16488 117360
rect 16356 117320 16488 117348
rect 16356 117308 16362 117320
rect 16482 117308 16488 117320
rect 16540 117308 16546 117360
rect 16758 117308 16764 117360
rect 16816 117348 16822 117360
rect 19352 117348 19380 117388
rect 20898 117376 20904 117428
rect 20956 117416 20962 117428
rect 20956 117388 22094 117416
rect 20956 117376 20962 117388
rect 16816 117320 18736 117348
rect 19352 117320 19472 117348
rect 16816 117308 16822 117320
rect 7929 117283 7987 117289
rect 7929 117280 7941 117283
rect 7300 117252 7941 117280
rect 6236 117240 6242 117252
rect 7929 117249 7941 117252
rect 7975 117249 7987 117283
rect 7929 117243 7987 117249
rect 9122 117240 9128 117292
rect 9180 117280 9186 117292
rect 9861 117283 9919 117289
rect 9861 117280 9873 117283
rect 9180 117252 9873 117280
rect 9180 117240 9186 117252
rect 9861 117249 9873 117252
rect 9907 117249 9919 117283
rect 9861 117243 9919 117249
rect 10502 117240 10508 117292
rect 10560 117280 10566 117292
rect 11333 117283 11391 117289
rect 11333 117280 11345 117283
rect 10560 117252 11345 117280
rect 10560 117240 10566 117252
rect 11333 117249 11345 117252
rect 11379 117249 11391 117283
rect 11333 117243 11391 117249
rect 11882 117240 11888 117292
rect 11940 117280 11946 117292
rect 13265 117283 13323 117289
rect 13265 117280 13277 117283
rect 11940 117252 13277 117280
rect 11940 117240 11946 117252
rect 13265 117249 13277 117252
rect 13311 117249 13323 117283
rect 13265 117243 13323 117249
rect 13354 117240 13360 117292
rect 13412 117280 13418 117292
rect 15197 117283 15255 117289
rect 15197 117280 15209 117283
rect 13412 117252 15209 117280
rect 13412 117240 13418 117252
rect 15197 117249 15209 117252
rect 15243 117249 15255 117283
rect 15197 117243 15255 117249
rect 17586 117240 17592 117292
rect 17644 117280 17650 117292
rect 18601 117283 18659 117289
rect 18601 117280 18613 117283
rect 17644 117252 18613 117280
rect 17644 117240 17650 117252
rect 18601 117249 18613 117252
rect 18647 117249 18659 117283
rect 18708 117280 18736 117320
rect 19337 117283 19395 117289
rect 19337 117280 19349 117283
rect 18708 117252 19349 117280
rect 18601 117243 18659 117249
rect 19337 117249 19349 117252
rect 19383 117249 19395 117283
rect 19444 117280 19472 117320
rect 19518 117308 19524 117360
rect 19576 117348 19582 117360
rect 19576 117320 21404 117348
rect 19576 117308 19582 117320
rect 21269 117283 21327 117289
rect 21269 117280 21281 117283
rect 19444 117252 21281 117280
rect 19337 117243 19395 117249
rect 21269 117249 21281 117252
rect 21315 117249 21327 117283
rect 21376 117280 21404 117320
rect 22066 117280 22094 117388
rect 22922 117376 22928 117428
rect 22980 117416 22986 117428
rect 27249 117419 27307 117425
rect 27249 117416 27261 117419
rect 22980 117388 27261 117416
rect 22980 117376 22986 117388
rect 27249 117385 27261 117388
rect 27295 117385 27307 117419
rect 27249 117379 27307 117385
rect 27338 117376 27344 117428
rect 27396 117416 27402 117428
rect 27396 117388 33088 117416
rect 27396 117376 27402 117388
rect 22278 117308 22284 117360
rect 22336 117348 22342 117360
rect 22336 117320 26280 117348
rect 22336 117308 22342 117320
rect 24673 117283 24731 117289
rect 24673 117280 24685 117283
rect 21376 117252 21956 117280
rect 22066 117252 24685 117280
rect 21269 117243 21327 117249
rect 5261 117215 5319 117221
rect 5261 117212 5273 117215
rect 808 117184 2774 117212
rect 4172 117184 5273 117212
rect 808 117172 814 117184
rect 1854 117144 1860 117156
rect 1815 117116 1860 117144
rect 1854 117104 1860 117116
rect 1912 117104 1918 117156
rect 2593 117147 2651 117153
rect 2593 117113 2605 117147
rect 2639 117144 2651 117147
rect 4062 117144 4068 117156
rect 2639 117116 4068 117144
rect 2639 117113 2651 117116
rect 2593 117107 2651 117113
rect 4062 117104 4068 117116
rect 4120 117104 4126 117156
rect 1026 117036 1032 117088
rect 1084 117076 1090 117088
rect 4172 117076 4200 117184
rect 5261 117181 5273 117184
rect 5307 117181 5319 117215
rect 5261 117175 5319 117181
rect 5442 117172 5448 117224
rect 5500 117212 5506 117224
rect 8481 117215 8539 117221
rect 8481 117212 8493 117215
rect 5500 117184 8493 117212
rect 5500 117172 5506 117184
rect 8481 117181 8493 117184
rect 8527 117181 8539 117215
rect 8481 117175 8539 117181
rect 9766 117172 9772 117224
rect 9824 117212 9830 117224
rect 10597 117215 10655 117221
rect 10597 117212 10609 117215
rect 9824 117184 10609 117212
rect 9824 117172 9830 117184
rect 10597 117181 10609 117184
rect 10643 117181 10655 117215
rect 10597 117175 10655 117181
rect 13906 117172 13912 117224
rect 13964 117212 13970 117224
rect 15933 117215 15991 117221
rect 15933 117212 15945 117215
rect 13964 117184 15945 117212
rect 13964 117172 13970 117184
rect 15933 117181 15945 117184
rect 15979 117181 15991 117215
rect 15933 117175 15991 117181
rect 17310 117172 17316 117224
rect 17368 117212 17374 117224
rect 18417 117215 18475 117221
rect 18417 117212 18429 117215
rect 17368 117184 18429 117212
rect 17368 117172 17374 117184
rect 18417 117181 18429 117184
rect 18463 117181 18475 117215
rect 18417 117175 18475 117181
rect 4341 117147 4399 117153
rect 4341 117113 4353 117147
rect 4387 117144 4399 117147
rect 4522 117144 4528 117156
rect 4387 117116 4528 117144
rect 4387 117113 4399 117116
rect 4341 117107 4399 117113
rect 4522 117104 4528 117116
rect 4580 117104 4586 117156
rect 5077 117147 5135 117153
rect 5077 117113 5089 117147
rect 5123 117113 5135 117147
rect 5077 117107 5135 117113
rect 5813 117147 5871 117153
rect 5813 117113 5825 117147
rect 5859 117144 5871 117147
rect 6822 117144 6828 117156
rect 5859 117116 6828 117144
rect 5859 117113 5871 117116
rect 5813 117107 5871 117113
rect 1084 117048 4200 117076
rect 5092 117076 5120 117107
rect 6822 117104 6828 117116
rect 6880 117104 6886 117156
rect 7009 117147 7067 117153
rect 7009 117113 7021 117147
rect 7055 117144 7067 117147
rect 7558 117144 7564 117156
rect 7055 117116 7564 117144
rect 7055 117113 7067 117116
rect 7009 117107 7067 117113
rect 7558 117104 7564 117116
rect 7616 117104 7622 117156
rect 7742 117144 7748 117156
rect 7703 117116 7748 117144
rect 7742 117104 7748 117116
rect 7800 117104 7806 117156
rect 9674 117144 9680 117156
rect 9635 117116 9680 117144
rect 9674 117104 9680 117116
rect 9732 117104 9738 117156
rect 10410 117144 10416 117156
rect 10371 117116 10416 117144
rect 10410 117104 10416 117116
rect 10468 117104 10474 117156
rect 11146 117144 11152 117156
rect 11107 117116 11152 117144
rect 11146 117104 11152 117116
rect 11204 117104 11210 117156
rect 11606 117104 11612 117156
rect 11664 117144 11670 117156
rect 12345 117147 12403 117153
rect 12345 117144 12357 117147
rect 11664 117116 12357 117144
rect 11664 117104 11670 117116
rect 12345 117113 12357 117116
rect 12391 117113 12403 117147
rect 13078 117144 13084 117156
rect 13039 117116 13084 117144
rect 12345 117107 12403 117113
rect 13078 117104 13084 117116
rect 13136 117104 13142 117156
rect 13814 117144 13820 117156
rect 13775 117116 13820 117144
rect 13814 117104 13820 117116
rect 13872 117104 13878 117156
rect 13998 117104 14004 117156
rect 14056 117144 14062 117156
rect 15013 117147 15071 117153
rect 15013 117144 15025 117147
rect 14056 117116 15025 117144
rect 14056 117104 14062 117116
rect 15013 117113 15025 117116
rect 15059 117113 15071 117147
rect 15013 117107 15071 117113
rect 15194 117104 15200 117156
rect 15252 117144 15258 117156
rect 15749 117147 15807 117153
rect 15749 117144 15761 117147
rect 15252 117116 15761 117144
rect 15252 117104 15258 117116
rect 15749 117113 15761 117116
rect 15795 117113 15807 117147
rect 15749 117107 15807 117113
rect 16206 117104 16212 117156
rect 16264 117144 16270 117156
rect 16485 117147 16543 117153
rect 16485 117144 16497 117147
rect 16264 117116 16497 117144
rect 16264 117104 16270 117116
rect 16485 117113 16497 117116
rect 16531 117113 16543 117147
rect 17678 117144 17684 117156
rect 17639 117116 17684 117144
rect 16485 117107 16543 117113
rect 17678 117104 17684 117116
rect 17736 117104 17742 117156
rect 19150 117144 19156 117156
rect 19111 117116 19156 117144
rect 19150 117104 19156 117116
rect 19208 117104 19214 117156
rect 19334 117104 19340 117156
rect 19392 117144 19398 117156
rect 20349 117147 20407 117153
rect 20349 117144 20361 117147
rect 19392 117116 20361 117144
rect 19392 117104 19398 117116
rect 20349 117113 20361 117116
rect 20395 117113 20407 117147
rect 20349 117107 20407 117113
rect 20530 117104 20536 117156
rect 20588 117144 20594 117156
rect 21085 117147 21143 117153
rect 21085 117144 21097 117147
rect 20588 117116 21097 117144
rect 20588 117104 20594 117116
rect 21085 117113 21097 117116
rect 21131 117113 21143 117147
rect 21085 117107 21143 117113
rect 21266 117104 21272 117156
rect 21324 117144 21330 117156
rect 21821 117147 21879 117153
rect 21821 117144 21833 117147
rect 21324 117116 21833 117144
rect 21324 117104 21330 117116
rect 21821 117113 21833 117116
rect 21867 117113 21879 117147
rect 21928 117144 21956 117252
rect 24673 117249 24685 117252
rect 24719 117249 24731 117283
rect 26252 117280 26280 117320
rect 26418 117308 26424 117360
rect 26476 117348 26482 117360
rect 28902 117348 28908 117360
rect 26476 117320 28908 117348
rect 26476 117308 26482 117320
rect 28902 117308 28908 117320
rect 28960 117308 28966 117360
rect 26605 117283 26663 117289
rect 26605 117280 26617 117283
rect 26252 117252 26617 117280
rect 24673 117243 24731 117249
rect 26605 117249 26617 117252
rect 26651 117249 26663 117283
rect 26605 117243 26663 117249
rect 27154 117240 27160 117292
rect 27212 117280 27218 117292
rect 32677 117283 32735 117289
rect 32677 117280 32689 117283
rect 27212 117252 32689 117280
rect 27212 117240 27218 117252
rect 32677 117249 32689 117252
rect 32723 117249 32735 117283
rect 33060 117280 33088 117388
rect 34790 117376 34796 117428
rect 34848 117416 34854 117428
rect 34977 117419 35035 117425
rect 34977 117416 34989 117419
rect 34848 117388 34989 117416
rect 34848 117376 34854 117388
rect 34977 117385 34989 117388
rect 35023 117385 35035 117419
rect 34977 117379 35035 117385
rect 33873 117283 33931 117289
rect 33873 117280 33885 117283
rect 33060 117252 33885 117280
rect 32677 117243 32735 117249
rect 33873 117249 33885 117252
rect 33919 117249 33931 117283
rect 33873 117243 33931 117249
rect 22922 117172 22928 117224
rect 22980 117212 22986 117224
rect 25869 117215 25927 117221
rect 25869 117212 25881 117215
rect 22980 117184 25881 117212
rect 22980 117172 22986 117184
rect 25869 117181 25881 117184
rect 25915 117181 25927 117215
rect 25869 117175 25927 117181
rect 27706 117172 27712 117224
rect 27764 117212 27770 117224
rect 32493 117215 32551 117221
rect 32493 117212 32505 117215
rect 27764 117184 32505 117212
rect 27764 117172 27770 117184
rect 32493 117181 32505 117184
rect 32539 117181 32551 117215
rect 32493 117175 32551 117181
rect 35434 117172 35440 117224
rect 35492 117212 35498 117224
rect 36357 117215 36415 117221
rect 36357 117212 36369 117215
rect 35492 117184 36369 117212
rect 35492 117172 35498 117184
rect 36357 117181 36369 117184
rect 36403 117181 36415 117215
rect 36357 117175 36415 117181
rect 37090 117172 37096 117224
rect 37148 117212 37154 117224
rect 37185 117215 37243 117221
rect 37185 117212 37197 117215
rect 37148 117184 37197 117212
rect 37148 117172 37154 117184
rect 37185 117181 37197 117184
rect 37231 117181 37243 117215
rect 37185 117175 37243 117181
rect 23014 117144 23020 117156
rect 21928 117116 22094 117144
rect 22975 117116 23020 117144
rect 21821 117107 21879 117113
rect 7374 117076 7380 117088
rect 5092 117048 7380 117076
rect 1084 117036 1090 117048
rect 7374 117036 7380 117048
rect 7432 117036 7438 117088
rect 7834 117036 7840 117088
rect 7892 117076 7898 117088
rect 8573 117079 8631 117085
rect 8573 117076 8585 117079
rect 7892 117048 8585 117076
rect 7892 117036 7898 117048
rect 8573 117045 8585 117048
rect 8619 117045 8631 117079
rect 8573 117039 8631 117045
rect 12526 117036 12532 117088
rect 12584 117076 12590 117088
rect 13909 117079 13967 117085
rect 13909 117076 13921 117079
rect 12584 117048 13921 117076
rect 12584 117036 12590 117048
rect 13909 117045 13921 117048
rect 13955 117045 13967 117079
rect 13909 117039 13967 117045
rect 14642 117036 14648 117088
rect 14700 117076 14706 117088
rect 16577 117079 16635 117085
rect 16577 117076 16589 117079
rect 14700 117048 16589 117076
rect 14700 117036 14706 117048
rect 16577 117045 16589 117048
rect 16623 117045 16635 117079
rect 16577 117039 16635 117045
rect 17034 117036 17040 117088
rect 17092 117076 17098 117088
rect 17773 117079 17831 117085
rect 17773 117076 17785 117079
rect 17092 117048 17785 117076
rect 17092 117036 17098 117048
rect 17773 117045 17785 117048
rect 17819 117045 17831 117079
rect 17773 117039 17831 117045
rect 17954 117036 17960 117088
rect 18012 117076 18018 117088
rect 20441 117079 20499 117085
rect 20441 117076 20453 117079
rect 18012 117048 20453 117076
rect 18012 117036 18018 117048
rect 20441 117045 20453 117048
rect 20487 117045 20499 117079
rect 21910 117076 21916 117088
rect 21871 117048 21916 117076
rect 20441 117039 20499 117045
rect 21910 117036 21916 117048
rect 21968 117036 21974 117088
rect 22066 117076 22094 117116
rect 23014 117104 23020 117116
rect 23072 117104 23078 117156
rect 23290 117104 23296 117156
rect 23348 117144 23354 117156
rect 23753 117147 23811 117153
rect 23753 117144 23765 117147
rect 23348 117116 23765 117144
rect 23348 117104 23354 117116
rect 23753 117113 23765 117116
rect 23799 117113 23811 117147
rect 24486 117144 24492 117156
rect 24447 117116 24492 117144
rect 23753 117107 23811 117113
rect 24486 117104 24492 117116
rect 24544 117104 24550 117156
rect 24670 117104 24676 117156
rect 24728 117144 24734 117156
rect 25685 117147 25743 117153
rect 25685 117144 25697 117147
rect 24728 117116 25697 117144
rect 24728 117104 24734 117116
rect 25685 117113 25697 117116
rect 25731 117113 25743 117147
rect 26418 117144 26424 117156
rect 26379 117116 26424 117144
rect 25685 117107 25743 117113
rect 26418 117104 26424 117116
rect 26476 117104 26482 117156
rect 27154 117144 27160 117156
rect 27115 117116 27160 117144
rect 27154 117104 27160 117116
rect 27212 117104 27218 117156
rect 28350 117144 28356 117156
rect 28311 117116 28356 117144
rect 28350 117104 28356 117116
rect 28408 117104 28414 117156
rect 28626 117104 28632 117156
rect 28684 117144 28690 117156
rect 29089 117147 29147 117153
rect 29089 117144 29101 117147
rect 28684 117116 29101 117144
rect 28684 117104 28690 117116
rect 29089 117113 29101 117116
rect 29135 117113 29147 117147
rect 29822 117144 29828 117156
rect 29783 117116 29828 117144
rect 29089 117107 29147 117113
rect 29822 117104 29828 117116
rect 29880 117104 29886 117156
rect 30006 117104 30012 117156
rect 30064 117144 30070 117156
rect 31021 117147 31079 117153
rect 31021 117144 31033 117147
rect 30064 117116 31033 117144
rect 30064 117104 30070 117116
rect 31021 117113 31033 117116
rect 31067 117113 31079 117147
rect 31021 117107 31079 117113
rect 31386 117104 31392 117156
rect 31444 117144 31450 117156
rect 31757 117147 31815 117153
rect 31757 117144 31769 117147
rect 31444 117116 31769 117144
rect 31444 117104 31450 117116
rect 31757 117113 31769 117116
rect 31803 117113 31815 117147
rect 31757 117107 31815 117113
rect 33318 117104 33324 117156
rect 33376 117144 33382 117156
rect 33689 117147 33747 117153
rect 33689 117144 33701 117147
rect 33376 117116 33701 117144
rect 33376 117104 33382 117116
rect 33689 117113 33701 117116
rect 33735 117113 33747 117147
rect 33689 117107 33747 117113
rect 34146 117104 34152 117156
rect 34204 117144 34210 117156
rect 34606 117144 34612 117156
rect 34204 117116 34612 117144
rect 34204 117104 34210 117116
rect 34606 117104 34612 117116
rect 34664 117104 34670 117156
rect 34885 117147 34943 117153
rect 34885 117113 34897 117147
rect 34931 117113 34943 117147
rect 34885 117107 34943 117113
rect 37461 117147 37519 117153
rect 37461 117113 37473 117147
rect 37507 117144 37519 117147
rect 38562 117144 38568 117156
rect 37507 117116 38568 117144
rect 37507 117113 37519 117116
rect 37461 117107 37519 117113
rect 23109 117079 23167 117085
rect 23109 117076 23121 117079
rect 22066 117048 23121 117076
rect 23109 117045 23121 117048
rect 23155 117045 23167 117079
rect 23109 117039 23167 117045
rect 23198 117036 23204 117088
rect 23256 117076 23262 117088
rect 23845 117079 23903 117085
rect 23845 117076 23857 117079
rect 23256 117048 23857 117076
rect 23256 117036 23262 117048
rect 23845 117045 23857 117048
rect 23891 117045 23903 117079
rect 23845 117039 23903 117045
rect 28166 117036 28172 117088
rect 28224 117076 28230 117088
rect 28445 117079 28503 117085
rect 28445 117076 28457 117079
rect 28224 117048 28457 117076
rect 28224 117036 28230 117048
rect 28445 117045 28457 117048
rect 28491 117045 28503 117079
rect 28445 117039 28503 117045
rect 28810 117036 28816 117088
rect 28868 117076 28874 117088
rect 29181 117079 29239 117085
rect 29181 117076 29193 117079
rect 28868 117048 29193 117076
rect 28868 117036 28874 117048
rect 29181 117045 29193 117048
rect 29227 117045 29239 117079
rect 29181 117039 29239 117045
rect 29270 117036 29276 117088
rect 29328 117076 29334 117088
rect 29917 117079 29975 117085
rect 29917 117076 29929 117079
rect 29328 117048 29929 117076
rect 29328 117036 29334 117048
rect 29917 117045 29929 117048
rect 29963 117045 29975 117079
rect 29917 117039 29975 117045
rect 30926 117036 30932 117088
rect 30984 117076 30990 117088
rect 31113 117079 31171 117085
rect 31113 117076 31125 117079
rect 30984 117048 31125 117076
rect 30984 117036 30990 117048
rect 31113 117045 31125 117048
rect 31159 117045 31171 117079
rect 31113 117039 31171 117045
rect 31202 117036 31208 117088
rect 31260 117076 31266 117088
rect 31849 117079 31907 117085
rect 31849 117076 31861 117079
rect 31260 117048 31861 117076
rect 31260 117036 31266 117048
rect 31849 117045 31861 117048
rect 31895 117045 31907 117079
rect 31849 117039 31907 117045
rect 33042 117036 33048 117088
rect 33100 117076 33106 117088
rect 34900 117076 34928 117107
rect 38562 117104 38568 117116
rect 38620 117104 38626 117156
rect 36446 117076 36452 117088
rect 33100 117048 34928 117076
rect 36407 117048 36452 117076
rect 33100 117036 33106 117048
rect 36446 117036 36452 117048
rect 36504 117036 36510 117088
rect 36538 117036 36544 117088
rect 36596 117076 36602 117088
rect 37734 117076 37740 117088
rect 36596 117048 37740 117076
rect 36596 117036 36602 117048
rect 37734 117036 37740 117048
rect 37792 117036 37798 117088
rect 1104 116986 38824 117008
rect 1104 116934 19606 116986
rect 19658 116934 19670 116986
rect 19722 116934 19734 116986
rect 19786 116934 19798 116986
rect 19850 116934 38824 116986
rect 1104 116912 38824 116934
rect 1670 116832 1676 116884
rect 1728 116872 1734 116884
rect 1949 116875 2007 116881
rect 1949 116872 1961 116875
rect 1728 116844 1961 116872
rect 1728 116832 1734 116844
rect 1949 116841 1961 116844
rect 1995 116841 2007 116875
rect 1949 116835 2007 116841
rect 4062 116832 4068 116884
rect 4120 116872 4126 116884
rect 4120 116844 4844 116872
rect 4120 116832 4126 116844
rect 2130 116764 2136 116816
rect 2188 116804 2194 116816
rect 2777 116807 2835 116813
rect 2777 116804 2789 116807
rect 2188 116776 2789 116804
rect 2188 116764 2194 116776
rect 2777 116773 2789 116776
rect 2823 116773 2835 116807
rect 2777 116767 2835 116773
rect 4525 116807 4583 116813
rect 4525 116773 4537 116807
rect 4571 116804 4583 116807
rect 4614 116804 4620 116816
rect 4571 116776 4620 116804
rect 4571 116773 4583 116776
rect 4525 116767 4583 116773
rect 4614 116764 4620 116776
rect 4672 116764 4678 116816
rect 4816 116804 4844 116844
rect 4890 116832 4896 116884
rect 4948 116872 4954 116884
rect 5169 116875 5227 116881
rect 5169 116872 5181 116875
rect 4948 116844 5181 116872
rect 4948 116832 4954 116844
rect 5169 116841 5181 116844
rect 5215 116841 5227 116875
rect 5169 116835 5227 116841
rect 6270 116832 6276 116884
rect 6328 116872 6334 116884
rect 7009 116875 7067 116881
rect 7009 116872 7021 116875
rect 6328 116844 7021 116872
rect 6328 116832 6334 116844
rect 7009 116841 7021 116844
rect 7055 116841 7067 116875
rect 7009 116835 7067 116841
rect 7098 116832 7104 116884
rect 7156 116872 7162 116884
rect 7745 116875 7803 116881
rect 7745 116872 7757 116875
rect 7156 116844 7757 116872
rect 7156 116832 7162 116844
rect 7745 116841 7757 116844
rect 7791 116841 7803 116875
rect 7745 116835 7803 116841
rect 8386 116832 8392 116884
rect 8444 116872 8450 116884
rect 9217 116875 9275 116881
rect 9217 116872 9229 116875
rect 8444 116844 9229 116872
rect 8444 116832 8450 116844
rect 9217 116841 9229 116844
rect 9263 116841 9275 116875
rect 9217 116835 9275 116841
rect 9306 116832 9312 116884
rect 9364 116872 9370 116884
rect 9953 116875 10011 116881
rect 9953 116872 9965 116875
rect 9364 116844 9965 116872
rect 9364 116832 9370 116844
rect 9953 116841 9965 116844
rect 9999 116841 10011 116875
rect 9953 116835 10011 116841
rect 10042 116832 10048 116884
rect 10100 116872 10106 116884
rect 10689 116875 10747 116881
rect 10689 116872 10701 116875
rect 10100 116844 10701 116872
rect 10100 116832 10106 116844
rect 10689 116841 10701 116844
rect 10735 116841 10747 116875
rect 10689 116835 10747 116841
rect 11422 116832 11428 116884
rect 11480 116872 11486 116884
rect 12253 116875 12311 116881
rect 12253 116872 12265 116875
rect 11480 116844 12265 116872
rect 11480 116832 11486 116844
rect 12253 116841 12265 116844
rect 12299 116841 12311 116875
rect 12253 116835 12311 116841
rect 12802 116832 12808 116884
rect 12860 116872 12866 116884
rect 13725 116875 13783 116881
rect 13725 116872 13737 116875
rect 12860 116844 13737 116872
rect 12860 116832 12866 116844
rect 13725 116841 13737 116844
rect 13771 116841 13783 116875
rect 13725 116835 13783 116841
rect 14182 116832 14188 116884
rect 14240 116872 14246 116884
rect 15197 116875 15255 116881
rect 15197 116872 15209 116875
rect 14240 116844 15209 116872
rect 14240 116832 14246 116844
rect 15197 116841 15209 116844
rect 15243 116841 15255 116875
rect 15197 116835 15255 116841
rect 15562 116832 15568 116884
rect 15620 116872 15626 116884
rect 15933 116875 15991 116881
rect 15933 116872 15945 116875
rect 15620 116844 15945 116872
rect 15620 116832 15626 116844
rect 15933 116841 15945 116844
rect 15979 116841 15991 116875
rect 15933 116835 15991 116841
rect 16942 116832 16948 116884
rect 17000 116872 17006 116884
rect 17497 116875 17555 116881
rect 17497 116872 17509 116875
rect 17000 116844 17509 116872
rect 17000 116832 17006 116844
rect 17497 116841 17509 116844
rect 17543 116841 17555 116875
rect 17497 116835 17555 116841
rect 17770 116832 17776 116884
rect 17828 116872 17834 116884
rect 18233 116875 18291 116881
rect 18233 116872 18245 116875
rect 17828 116844 18245 116872
rect 17828 116832 17834 116844
rect 18233 116841 18245 116844
rect 18279 116841 18291 116875
rect 18233 116835 18291 116841
rect 18322 116832 18328 116884
rect 18380 116872 18386 116884
rect 18969 116875 19027 116881
rect 18969 116872 18981 116875
rect 18380 116844 18981 116872
rect 18380 116832 18386 116844
rect 18969 116841 18981 116844
rect 19015 116841 19027 116875
rect 18969 116835 19027 116841
rect 19058 116832 19064 116884
rect 19116 116872 19122 116884
rect 19705 116875 19763 116881
rect 19705 116872 19717 116875
rect 19116 116844 19717 116872
rect 19116 116832 19122 116844
rect 19705 116841 19717 116844
rect 19751 116841 19763 116875
rect 19705 116835 19763 116841
rect 20438 116832 20444 116884
rect 20496 116872 20502 116884
rect 21177 116875 21235 116881
rect 21177 116872 21189 116875
rect 20496 116844 21189 116872
rect 20496 116832 20502 116844
rect 21177 116841 21189 116844
rect 21223 116841 21235 116875
rect 21177 116835 21235 116841
rect 21818 116832 21824 116884
rect 21876 116872 21882 116884
rect 22741 116875 22799 116881
rect 22741 116872 22753 116875
rect 21876 116844 22753 116872
rect 21876 116832 21882 116844
rect 22741 116841 22753 116844
rect 22787 116841 22799 116875
rect 22741 116835 22799 116841
rect 23106 116832 23112 116884
rect 23164 116872 23170 116884
rect 24213 116875 24271 116881
rect 24213 116872 24225 116875
rect 23164 116844 24225 116872
rect 23164 116832 23170 116844
rect 24213 116841 24225 116844
rect 24259 116841 24271 116875
rect 24213 116835 24271 116841
rect 24578 116832 24584 116884
rect 24636 116872 24642 116884
rect 24949 116875 25007 116881
rect 24949 116872 24961 116875
rect 24636 116844 24961 116872
rect 24636 116832 24642 116844
rect 24949 116841 24961 116844
rect 24995 116841 25007 116875
rect 24949 116835 25007 116841
rect 25314 116832 25320 116884
rect 25372 116872 25378 116884
rect 25685 116875 25743 116881
rect 25685 116872 25697 116875
rect 25372 116844 25697 116872
rect 25372 116832 25378 116844
rect 25685 116841 25697 116844
rect 25731 116841 25743 116875
rect 25685 116835 25743 116841
rect 25958 116832 25964 116884
rect 26016 116872 26022 116884
rect 26421 116875 26479 116881
rect 26421 116872 26433 116875
rect 26016 116844 26433 116872
rect 26016 116832 26022 116844
rect 26421 116841 26433 116844
rect 26467 116841 26479 116875
rect 26421 116835 26479 116841
rect 27798 116832 27804 116884
rect 27856 116872 27862 116884
rect 27985 116875 28043 116881
rect 27985 116872 27997 116875
rect 27856 116844 27997 116872
rect 27856 116832 27862 116844
rect 27985 116841 27997 116844
rect 28031 116841 28043 116875
rect 27985 116835 28043 116841
rect 28074 116832 28080 116884
rect 28132 116872 28138 116884
rect 28721 116875 28779 116881
rect 28721 116872 28733 116875
rect 28132 116844 28733 116872
rect 28132 116832 28138 116844
rect 28721 116841 28733 116844
rect 28767 116841 28779 116875
rect 28721 116835 28779 116841
rect 28902 116832 28908 116884
rect 28960 116872 28966 116884
rect 31202 116872 31208 116884
rect 28960 116844 31208 116872
rect 28960 116832 28966 116844
rect 31202 116832 31208 116844
rect 31260 116832 31266 116884
rect 31754 116832 31760 116884
rect 31812 116872 31818 116884
rect 32306 116872 32312 116884
rect 31812 116844 32312 116872
rect 31812 116832 31818 116844
rect 32306 116832 32312 116844
rect 32364 116832 32370 116884
rect 33597 116875 33655 116881
rect 33597 116841 33609 116875
rect 33643 116872 33655 116875
rect 36538 116872 36544 116884
rect 33643 116844 36544 116872
rect 33643 116841 33655 116844
rect 33597 116835 33655 116841
rect 36538 116832 36544 116844
rect 36596 116832 36602 116884
rect 36630 116832 36636 116884
rect 36688 116872 36694 116884
rect 37277 116875 37335 116881
rect 37277 116872 37289 116875
rect 36688 116844 37289 116872
rect 36688 116832 36694 116844
rect 37277 116841 37289 116844
rect 37323 116841 37335 116875
rect 37277 116835 37335 116841
rect 5994 116804 6000 116816
rect 4816 116776 6000 116804
rect 5994 116764 6000 116776
rect 6052 116764 6058 116816
rect 12066 116764 12072 116816
rect 12124 116804 12130 116816
rect 13081 116807 13139 116813
rect 13081 116804 13093 116807
rect 12124 116776 13093 116804
rect 12124 116764 12130 116776
rect 13081 116773 13093 116776
rect 13127 116773 13139 116807
rect 13081 116767 13139 116773
rect 13446 116764 13452 116816
rect 13504 116804 13510 116816
rect 14553 116807 14611 116813
rect 14553 116804 14565 116807
rect 13504 116776 14565 116804
rect 13504 116764 13510 116776
rect 14553 116773 14565 116776
rect 14599 116773 14611 116807
rect 14553 116767 14611 116773
rect 19886 116764 19892 116816
rect 19944 116804 19950 116816
rect 20533 116807 20591 116813
rect 20533 116804 20545 116807
rect 19944 116776 20545 116804
rect 19944 116764 19950 116776
rect 20533 116773 20545 116776
rect 20579 116773 20591 116807
rect 21266 116804 21272 116816
rect 20533 116767 20591 116773
rect 20640 116776 21272 116804
rect 1857 116739 1915 116745
rect 1857 116705 1869 116739
rect 1903 116705 1915 116739
rect 1857 116699 1915 116705
rect 2593 116739 2651 116745
rect 2593 116705 2605 116739
rect 2639 116736 2651 116739
rect 3234 116736 3240 116748
rect 2639 116708 3240 116736
rect 2639 116705 2651 116708
rect 2593 116699 2651 116705
rect 1872 116600 1900 116699
rect 3234 116696 3240 116708
rect 3292 116696 3298 116748
rect 3329 116739 3387 116745
rect 3329 116705 3341 116739
rect 3375 116736 3387 116739
rect 3878 116736 3884 116748
rect 3375 116708 3884 116736
rect 3375 116705 3387 116708
rect 3329 116699 3387 116705
rect 3878 116696 3884 116708
rect 3936 116696 3942 116748
rect 4341 116739 4399 116745
rect 4341 116705 4353 116739
rect 4387 116705 4399 116739
rect 5074 116736 5080 116748
rect 5035 116708 5080 116736
rect 4341 116699 4399 116705
rect 4356 116668 4384 116699
rect 5074 116696 5080 116708
rect 5132 116696 5138 116748
rect 6914 116736 6920 116748
rect 6875 116708 6920 116736
rect 6914 116696 6920 116708
rect 6972 116696 6978 116748
rect 7098 116696 7104 116748
rect 7156 116736 7162 116748
rect 7653 116739 7711 116745
rect 7653 116736 7665 116739
rect 7156 116708 7665 116736
rect 7156 116696 7162 116708
rect 7653 116705 7665 116708
rect 7699 116705 7711 116739
rect 8386 116736 8392 116748
rect 8347 116708 8392 116736
rect 7653 116699 7711 116705
rect 8386 116696 8392 116708
rect 8444 116696 8450 116748
rect 9122 116736 9128 116748
rect 9083 116708 9128 116736
rect 9122 116696 9128 116708
rect 9180 116696 9186 116748
rect 9858 116736 9864 116748
rect 9819 116708 9864 116736
rect 9858 116696 9864 116708
rect 9916 116696 9922 116748
rect 10594 116736 10600 116748
rect 10555 116708 10600 116736
rect 10594 116696 10600 116708
rect 10652 116696 10658 116748
rect 12158 116736 12164 116748
rect 12119 116708 12164 116736
rect 12158 116696 12164 116708
rect 12216 116696 12222 116748
rect 12894 116736 12900 116748
rect 12855 116708 12900 116736
rect 12894 116696 12900 116708
rect 12952 116696 12958 116748
rect 12986 116696 12992 116748
rect 13044 116736 13050 116748
rect 13633 116739 13691 116745
rect 13633 116736 13645 116739
rect 13044 116708 13645 116736
rect 13044 116696 13050 116708
rect 13633 116705 13645 116708
rect 13679 116705 13691 116739
rect 14366 116736 14372 116748
rect 14327 116708 14372 116736
rect 13633 116699 13691 116705
rect 14366 116696 14372 116708
rect 14424 116696 14430 116748
rect 15102 116736 15108 116748
rect 15063 116708 15108 116736
rect 15102 116696 15108 116708
rect 15160 116696 15166 116748
rect 15838 116736 15844 116748
rect 15799 116708 15844 116736
rect 15838 116696 15844 116708
rect 15896 116696 15902 116748
rect 17402 116736 17408 116748
rect 17363 116708 17408 116736
rect 17402 116696 17408 116708
rect 17460 116696 17466 116748
rect 18138 116736 18144 116748
rect 18099 116708 18144 116736
rect 18138 116696 18144 116708
rect 18196 116696 18202 116748
rect 18874 116736 18880 116748
rect 18835 116708 18880 116736
rect 18874 116696 18880 116708
rect 18932 116696 18938 116748
rect 19426 116696 19432 116748
rect 19484 116736 19490 116748
rect 19613 116739 19671 116745
rect 19613 116736 19625 116739
rect 19484 116708 19625 116736
rect 19484 116696 19490 116708
rect 19613 116705 19625 116708
rect 19659 116705 19671 116739
rect 20346 116736 20352 116748
rect 20307 116708 20352 116736
rect 19613 116699 19671 116705
rect 20346 116696 20352 116708
rect 20404 116696 20410 116748
rect 20438 116696 20444 116748
rect 20496 116736 20502 116748
rect 20640 116736 20668 116776
rect 21266 116764 21272 116776
rect 21324 116764 21330 116816
rect 22462 116764 22468 116816
rect 22520 116804 22526 116816
rect 23569 116807 23627 116813
rect 23569 116804 23581 116807
rect 22520 116776 23581 116804
rect 22520 116764 22526 116776
rect 23569 116773 23581 116776
rect 23615 116773 23627 116807
rect 28442 116804 28448 116816
rect 23569 116767 23627 116773
rect 25516 116776 28448 116804
rect 21082 116736 21088 116748
rect 20496 116708 20668 116736
rect 21043 116708 21088 116736
rect 20496 116696 20502 116708
rect 21082 116696 21088 116708
rect 21140 116696 21146 116748
rect 22646 116736 22652 116748
rect 22607 116708 22652 116736
rect 22646 116696 22652 116708
rect 22704 116696 22710 116748
rect 23385 116739 23443 116745
rect 23385 116705 23397 116739
rect 23431 116736 23443 116739
rect 24121 116739 24179 116745
rect 23431 116708 24072 116736
rect 23431 116705 23443 116708
rect 23385 116699 23443 116705
rect 4982 116668 4988 116680
rect 4356 116640 4988 116668
rect 4982 116628 4988 116640
rect 5040 116628 5046 116680
rect 5534 116628 5540 116680
rect 5592 116668 5598 116680
rect 7742 116668 7748 116680
rect 5592 116640 7748 116668
rect 5592 116628 5598 116640
rect 7742 116628 7748 116640
rect 7800 116628 7806 116680
rect 18782 116628 18788 116680
rect 18840 116668 18846 116680
rect 21910 116668 21916 116680
rect 18840 116640 21916 116668
rect 18840 116628 18846 116640
rect 21910 116628 21916 116640
rect 21968 116628 21974 116680
rect 22370 116628 22376 116680
rect 22428 116668 22434 116680
rect 24044 116668 24072 116708
rect 24121 116705 24133 116739
rect 24167 116736 24179 116739
rect 24762 116736 24768 116748
rect 24167 116708 24768 116736
rect 24167 116705 24179 116708
rect 24121 116699 24179 116705
rect 24762 116696 24768 116708
rect 24820 116696 24826 116748
rect 24857 116739 24915 116745
rect 24857 116705 24869 116739
rect 24903 116736 24915 116739
rect 25516 116736 25544 116776
rect 28442 116764 28448 116776
rect 28500 116764 28506 116816
rect 28534 116764 28540 116816
rect 28592 116804 28598 116816
rect 29549 116807 29607 116813
rect 29549 116804 29561 116807
rect 28592 116776 29561 116804
rect 28592 116764 28598 116776
rect 29549 116773 29561 116776
rect 29595 116773 29607 116807
rect 29549 116767 29607 116773
rect 31389 116807 31447 116813
rect 31389 116773 31401 116807
rect 31435 116804 31447 116807
rect 34146 116804 34152 116816
rect 31435 116776 34152 116804
rect 31435 116773 31447 116776
rect 31389 116767 31447 116773
rect 34146 116764 34152 116776
rect 34204 116764 34210 116816
rect 35161 116807 35219 116813
rect 35161 116773 35173 116807
rect 35207 116804 35219 116807
rect 35250 116804 35256 116816
rect 35207 116776 35256 116804
rect 35207 116773 35219 116776
rect 35161 116767 35219 116773
rect 35250 116764 35256 116776
rect 35308 116764 35314 116816
rect 35897 116807 35955 116813
rect 35897 116773 35909 116807
rect 35943 116804 35955 116807
rect 38194 116804 38200 116816
rect 35943 116776 38200 116804
rect 35943 116773 35955 116776
rect 35897 116767 35955 116773
rect 38194 116764 38200 116776
rect 38252 116764 38258 116816
rect 24903 116708 25544 116736
rect 25593 116739 25651 116745
rect 24903 116705 24915 116708
rect 24857 116699 24915 116705
rect 25593 116705 25605 116739
rect 25639 116736 25651 116739
rect 26329 116739 26387 116745
rect 25639 116708 26280 116736
rect 25639 116705 25651 116708
rect 25593 116699 25651 116705
rect 25682 116668 25688 116680
rect 22428 116640 23336 116668
rect 24044 116640 25688 116668
rect 22428 116628 22434 116640
rect 6270 116600 6276 116612
rect 1872 116572 6276 116600
rect 6270 116560 6276 116572
rect 6328 116560 6334 116612
rect 20254 116560 20260 116612
rect 20312 116600 20318 116612
rect 23198 116600 23204 116612
rect 20312 116572 23204 116600
rect 20312 116560 20318 116572
rect 23198 116560 23204 116572
rect 23256 116560 23262 116612
rect 23308 116600 23336 116640
rect 25682 116628 25688 116640
rect 25740 116628 25746 116680
rect 24486 116600 24492 116612
rect 23308 116572 24492 116600
rect 24486 116560 24492 116572
rect 24544 116560 24550 116612
rect 26252 116600 26280 116708
rect 26329 116705 26341 116739
rect 26375 116705 26387 116739
rect 27890 116736 27896 116748
rect 27851 116708 27896 116736
rect 26329 116699 26387 116705
rect 26344 116668 26372 116699
rect 27890 116696 27896 116708
rect 27948 116696 27954 116748
rect 28626 116736 28632 116748
rect 28587 116708 28632 116736
rect 28626 116696 28632 116708
rect 28684 116696 28690 116748
rect 28810 116696 28816 116748
rect 28868 116736 28874 116748
rect 29362 116736 29368 116748
rect 28868 116708 29224 116736
rect 29323 116708 29368 116736
rect 28868 116696 28874 116708
rect 28534 116668 28540 116680
rect 26344 116640 28540 116668
rect 28534 116628 28540 116640
rect 28592 116628 28598 116680
rect 29196 116668 29224 116708
rect 29362 116696 29368 116708
rect 29420 116696 29426 116748
rect 30466 116736 30472 116748
rect 30427 116708 30472 116736
rect 30466 116696 30472 116708
rect 30524 116696 30530 116748
rect 31018 116696 31024 116748
rect 31076 116736 31082 116748
rect 31205 116739 31263 116745
rect 31205 116736 31217 116739
rect 31076 116708 31217 116736
rect 31076 116696 31082 116708
rect 31205 116705 31217 116708
rect 31251 116705 31263 116739
rect 31205 116699 31263 116705
rect 31846 116696 31852 116748
rect 31904 116736 31910 116748
rect 31941 116739 31999 116745
rect 31941 116736 31953 116739
rect 31904 116708 31953 116736
rect 31904 116696 31910 116708
rect 31941 116705 31953 116708
rect 31987 116705 31999 116739
rect 31941 116699 31999 116705
rect 33505 116739 33563 116745
rect 33505 116705 33517 116739
rect 33551 116736 33563 116739
rect 33962 116736 33968 116748
rect 33551 116708 33968 116736
rect 33551 116705 33563 116708
rect 33505 116699 33563 116705
rect 33962 116696 33968 116708
rect 34020 116696 34026 116748
rect 34241 116739 34299 116745
rect 34241 116705 34253 116739
rect 34287 116705 34299 116739
rect 34241 116699 34299 116705
rect 31386 116668 31392 116680
rect 29196 116640 31392 116668
rect 31386 116628 31392 116640
rect 31444 116628 31450 116680
rect 34256 116668 34284 116699
rect 34698 116696 34704 116748
rect 34756 116736 34762 116748
rect 34977 116739 35035 116745
rect 34977 116736 34989 116739
rect 34756 116708 34989 116736
rect 34756 116696 34762 116708
rect 34977 116705 34989 116708
rect 35023 116705 35035 116739
rect 34977 116699 35035 116705
rect 35434 116696 35440 116748
rect 35492 116736 35498 116748
rect 35713 116739 35771 116745
rect 35713 116736 35725 116739
rect 35492 116708 35725 116736
rect 35492 116696 35498 116708
rect 35713 116705 35725 116708
rect 35759 116705 35771 116739
rect 36354 116736 36360 116748
rect 36315 116708 36360 116736
rect 35713 116699 35771 116705
rect 36354 116696 36360 116708
rect 36412 116696 36418 116748
rect 36538 116696 36544 116748
rect 36596 116736 36602 116748
rect 37185 116739 37243 116745
rect 37185 116736 37197 116739
rect 36596 116708 37197 116736
rect 36596 116696 36602 116708
rect 37185 116705 37197 116708
rect 37231 116705 37243 116739
rect 37185 116699 37243 116705
rect 36262 116668 36268 116680
rect 34256 116640 36268 116668
rect 36262 116628 36268 116640
rect 36320 116628 36326 116680
rect 28902 116600 28908 116612
rect 26252 116572 28908 116600
rect 28902 116560 28908 116572
rect 28960 116560 28966 116612
rect 30653 116603 30711 116609
rect 30653 116569 30665 116603
rect 30699 116600 30711 116603
rect 34238 116600 34244 116612
rect 30699 116572 34244 116600
rect 30699 116569 30711 116572
rect 30653 116563 30711 116569
rect 34238 116560 34244 116572
rect 34296 116560 34302 116612
rect 34425 116603 34483 116609
rect 34425 116569 34437 116603
rect 34471 116600 34483 116603
rect 36814 116600 36820 116612
rect 34471 116572 36820 116600
rect 34471 116569 34483 116572
rect 34425 116563 34483 116569
rect 36814 116560 36820 116572
rect 36872 116560 36878 116612
rect 2958 116492 2964 116544
rect 3016 116532 3022 116544
rect 3421 116535 3479 116541
rect 3421 116532 3433 116535
rect 3016 116504 3433 116532
rect 3016 116492 3022 116504
rect 3421 116501 3433 116504
rect 3467 116501 3479 116535
rect 3421 116495 3479 116501
rect 5718 116492 5724 116544
rect 5776 116532 5782 116544
rect 5905 116535 5963 116541
rect 5905 116532 5917 116535
rect 5776 116504 5917 116532
rect 5776 116492 5782 116504
rect 5905 116501 5917 116504
rect 5951 116501 5963 116535
rect 5905 116495 5963 116501
rect 7650 116492 7656 116544
rect 7708 116532 7714 116544
rect 8481 116535 8539 116541
rect 8481 116532 8493 116535
rect 7708 116504 8493 116532
rect 7708 116492 7714 116504
rect 8481 116501 8493 116504
rect 8527 116501 8539 116535
rect 8481 116495 8539 116501
rect 20714 116492 20720 116544
rect 20772 116532 20778 116544
rect 23290 116532 23296 116544
rect 20772 116504 23296 116532
rect 20772 116492 20778 116504
rect 23290 116492 23296 116504
rect 23348 116492 23354 116544
rect 25866 116492 25872 116544
rect 25924 116532 25930 116544
rect 30006 116532 30012 116544
rect 25924 116504 30012 116532
rect 25924 116492 25930 116504
rect 30006 116492 30012 116504
rect 30064 116492 30070 116544
rect 32033 116535 32091 116541
rect 32033 116501 32045 116535
rect 32079 116532 32091 116535
rect 32766 116532 32772 116544
rect 32079 116504 32772 116532
rect 32079 116501 32091 116504
rect 32033 116495 32091 116501
rect 32766 116492 32772 116504
rect 32824 116492 32830 116544
rect 33870 116492 33876 116544
rect 33928 116532 33934 116544
rect 34146 116532 34152 116544
rect 33928 116504 34152 116532
rect 33928 116492 33934 116504
rect 34146 116492 34152 116504
rect 34204 116492 34210 116544
rect 36541 116535 36599 116541
rect 36541 116501 36553 116535
rect 36587 116532 36599 116535
rect 36722 116532 36728 116544
rect 36587 116504 36728 116532
rect 36587 116501 36599 116504
rect 36541 116495 36599 116501
rect 36722 116492 36728 116504
rect 36780 116492 36786 116544
rect 1104 116442 38824 116464
rect 1104 116390 4246 116442
rect 4298 116390 4310 116442
rect 4362 116390 4374 116442
rect 4426 116390 4438 116442
rect 4490 116390 34966 116442
rect 35018 116390 35030 116442
rect 35082 116390 35094 116442
rect 35146 116390 35158 116442
rect 35210 116390 38824 116442
rect 1104 116368 38824 116390
rect 2406 116288 2412 116340
rect 2464 116328 2470 116340
rect 3237 116331 3295 116337
rect 3237 116328 3249 116331
rect 2464 116300 3249 116328
rect 2464 116288 2470 116300
rect 3237 116297 3249 116300
rect 3283 116297 3295 116331
rect 3237 116291 3295 116297
rect 3786 116288 3792 116340
rect 3844 116328 3850 116340
rect 4433 116331 4491 116337
rect 4433 116328 4445 116331
rect 3844 116300 4445 116328
rect 3844 116288 3850 116300
rect 4433 116297 4445 116300
rect 4479 116297 4491 116331
rect 4433 116291 4491 116297
rect 5169 116331 5227 116337
rect 5169 116297 5181 116331
rect 5215 116328 5227 116331
rect 5442 116328 5448 116340
rect 5215 116300 5448 116328
rect 5215 116297 5227 116300
rect 5169 116291 5227 116297
rect 5442 116288 5448 116300
rect 5500 116288 5506 116340
rect 5626 116288 5632 116340
rect 5684 116328 5690 116340
rect 5813 116331 5871 116337
rect 5813 116328 5825 116331
rect 5684 116300 5825 116328
rect 5684 116288 5690 116300
rect 5813 116297 5825 116300
rect 5859 116297 5871 116331
rect 5813 116291 5871 116297
rect 5902 116288 5908 116340
rect 5960 116328 5966 116340
rect 6549 116331 6607 116337
rect 6549 116328 6561 116331
rect 5960 116300 6561 116328
rect 5960 116288 5966 116300
rect 6549 116297 6561 116300
rect 6595 116297 6607 116331
rect 6549 116291 6607 116297
rect 6638 116288 6644 116340
rect 6696 116328 6702 116340
rect 7285 116331 7343 116337
rect 7285 116328 7297 116331
rect 6696 116300 7297 116328
rect 6696 116288 6702 116300
rect 7285 116297 7297 116300
rect 7331 116297 7343 116331
rect 7285 116291 7343 116297
rect 8662 116288 8668 116340
rect 8720 116328 8726 116340
rect 9677 116331 9735 116337
rect 9677 116328 9689 116331
rect 8720 116300 9689 116328
rect 8720 116288 8726 116300
rect 9677 116297 9689 116300
rect 9723 116297 9735 116331
rect 9677 116291 9735 116297
rect 10686 116288 10692 116340
rect 10744 116328 10750 116340
rect 10873 116331 10931 116337
rect 10873 116328 10885 116331
rect 10744 116300 10885 116328
rect 10744 116288 10750 116300
rect 10873 116297 10885 116300
rect 10919 116297 10931 116331
rect 11606 116328 11612 116340
rect 11567 116300 11612 116328
rect 10873 116291 10931 116297
rect 11606 116288 11612 116300
rect 11664 116288 11670 116340
rect 12253 116331 12311 116337
rect 12253 116297 12265 116331
rect 12299 116328 12311 116331
rect 13078 116328 13084 116340
rect 12299 116300 13084 116328
rect 12299 116297 12311 116300
rect 12253 116291 12311 116297
rect 13078 116288 13084 116300
rect 13136 116288 13142 116340
rect 13541 116331 13599 116337
rect 13541 116297 13553 116331
rect 13587 116328 13599 116331
rect 13998 116328 14004 116340
rect 13587 116300 14004 116328
rect 13587 116297 13599 116300
rect 13541 116291 13599 116297
rect 13998 116288 14004 116300
rect 14056 116288 14062 116340
rect 14826 116288 14832 116340
rect 14884 116328 14890 116340
rect 15013 116331 15071 116337
rect 15013 116328 15025 116331
rect 14884 116300 15025 116328
rect 14884 116288 14890 116300
rect 15013 116297 15025 116300
rect 15059 116297 15071 116331
rect 15013 116291 15071 116297
rect 15749 116331 15807 116337
rect 15749 116297 15761 116331
rect 15795 116328 15807 116331
rect 17678 116328 17684 116340
rect 15795 116300 17684 116328
rect 15795 116297 15807 116300
rect 15749 116291 15807 116297
rect 17678 116288 17684 116300
rect 17736 116288 17742 116340
rect 17865 116331 17923 116337
rect 17865 116297 17877 116331
rect 17911 116328 17923 116331
rect 19334 116328 19340 116340
rect 17911 116300 19340 116328
rect 17911 116297 17923 116300
rect 17865 116291 17923 116297
rect 19334 116288 19340 116300
rect 19392 116288 19398 116340
rect 21174 116288 21180 116340
rect 21232 116328 21238 116340
rect 21269 116331 21327 116337
rect 21269 116328 21281 116331
rect 21232 116300 21281 116328
rect 21232 116288 21238 116300
rect 21269 116297 21281 116300
rect 21315 116297 21327 116331
rect 23014 116328 23020 116340
rect 21269 116291 21327 116297
rect 21468 116300 23020 116328
rect 1854 116220 1860 116272
rect 1912 116260 1918 116272
rect 1912 116232 5488 116260
rect 1912 116220 1918 116232
rect 5460 116204 5488 116232
rect 7190 116220 7196 116272
rect 7248 116260 7254 116272
rect 8113 116263 8171 116269
rect 8113 116260 8125 116263
rect 7248 116232 8125 116260
rect 7248 116220 7254 116232
rect 8113 116229 8125 116232
rect 8159 116229 8171 116263
rect 8113 116223 8171 116229
rect 12897 116263 12955 116269
rect 12897 116229 12909 116263
rect 12943 116260 12955 116263
rect 13814 116260 13820 116272
rect 12943 116232 13820 116260
rect 12943 116229 12955 116232
rect 12897 116223 12955 116229
rect 13814 116220 13820 116232
rect 13872 116220 13878 116272
rect 16574 116220 16580 116272
rect 16632 116260 16638 116272
rect 17221 116263 17279 116269
rect 16632 116232 16677 116260
rect 16632 116220 16638 116232
rect 17221 116229 17233 116263
rect 17267 116260 17279 116263
rect 19150 116260 19156 116272
rect 17267 116232 19156 116260
rect 17267 116229 17279 116232
rect 17221 116223 17279 116229
rect 19150 116220 19156 116232
rect 19208 116220 19214 116272
rect 20165 116263 20223 116269
rect 20165 116229 20177 116263
rect 20211 116260 20223 116263
rect 21468 116260 21496 116300
rect 23014 116288 23020 116300
rect 23072 116288 23078 116340
rect 23842 116288 23848 116340
rect 23900 116328 23906 116340
rect 24029 116331 24087 116337
rect 24029 116328 24041 116331
rect 23900 116300 24041 116328
rect 23900 116288 23906 116300
rect 24029 116297 24041 116300
rect 24075 116297 24087 116331
rect 24029 116291 24087 116297
rect 24762 116288 24768 116340
rect 24820 116328 24826 116340
rect 26602 116328 26608 116340
rect 24820 116300 26608 116328
rect 24820 116288 24826 116300
rect 26602 116288 26608 116300
rect 26660 116288 26666 116340
rect 26694 116288 26700 116340
rect 26752 116328 26758 116340
rect 26881 116331 26939 116337
rect 26881 116328 26893 116331
rect 26752 116300 26893 116328
rect 26752 116288 26758 116300
rect 26881 116297 26893 116300
rect 26927 116297 26939 116331
rect 26881 116291 26939 116297
rect 26970 116288 26976 116340
rect 27028 116328 27034 116340
rect 27617 116331 27675 116337
rect 27028 116300 27568 116328
rect 27028 116288 27034 116300
rect 20211 116232 21496 116260
rect 20211 116229 20223 116232
rect 20165 116223 20223 116229
rect 21542 116220 21548 116272
rect 21600 116260 21606 116272
rect 22922 116260 22928 116272
rect 21600 116232 22928 116260
rect 21600 116220 21606 116232
rect 22922 116220 22928 116232
rect 22980 116220 22986 116272
rect 27154 116260 27160 116272
rect 23124 116232 27160 116260
rect 2038 116192 2044 116204
rect 1999 116164 2044 116192
rect 2038 116152 2044 116164
rect 2096 116152 2102 116204
rect 5442 116152 5448 116204
rect 5500 116152 5506 116204
rect 18509 116195 18567 116201
rect 18509 116161 18521 116195
rect 18555 116192 18567 116195
rect 20530 116192 20536 116204
rect 18555 116164 20536 116192
rect 18555 116161 18567 116164
rect 18509 116155 18567 116161
rect 20530 116152 20536 116164
rect 20588 116152 20594 116204
rect 21821 116195 21879 116201
rect 21821 116161 21833 116195
rect 21867 116192 21879 116195
rect 22462 116192 22468 116204
rect 21867 116164 22094 116192
rect 22423 116164 22468 116192
rect 21867 116161 21879 116164
rect 21821 116155 21879 116161
rect 5718 116124 5724 116136
rect 5679 116096 5724 116124
rect 5718 116084 5724 116096
rect 5776 116084 5782 116136
rect 15286 116084 15292 116136
rect 15344 116124 15350 116136
rect 17034 116124 17040 116136
rect 15344 116096 17040 116124
rect 15344 116084 15350 116096
rect 17034 116084 17040 116096
rect 17092 116084 17098 116136
rect 1762 116016 1768 116068
rect 1820 116056 1826 116068
rect 1857 116059 1915 116065
rect 1857 116056 1869 116059
rect 1820 116028 1869 116056
rect 1820 116016 1826 116028
rect 1857 116025 1869 116028
rect 1903 116025 1915 116059
rect 3142 116056 3148 116068
rect 3103 116028 3148 116056
rect 1857 116019 1915 116025
rect 3142 116016 3148 116028
rect 3200 116016 3206 116068
rect 4341 116059 4399 116065
rect 4341 116025 4353 116059
rect 4387 116056 4399 116059
rect 4890 116056 4896 116068
rect 4387 116028 4896 116056
rect 4387 116025 4399 116028
rect 4341 116019 4399 116025
rect 4890 116016 4896 116028
rect 4948 116016 4954 116068
rect 6454 116056 6460 116068
rect 6415 116028 6460 116056
rect 6454 116016 6460 116028
rect 6512 116016 6518 116068
rect 7006 116016 7012 116068
rect 7064 116056 7070 116068
rect 7193 116059 7251 116065
rect 7193 116056 7205 116059
rect 7064 116028 7205 116056
rect 7064 116016 7070 116028
rect 7193 116025 7205 116028
rect 7239 116025 7251 116059
rect 7926 116056 7932 116068
rect 7887 116028 7932 116056
rect 7193 116019 7251 116025
rect 7926 116016 7932 116028
rect 7984 116016 7990 116068
rect 9582 116056 9588 116068
rect 9543 116028 9588 116056
rect 9582 116016 9588 116028
rect 9640 116016 9646 116068
rect 10778 116056 10784 116068
rect 10739 116028 10784 116056
rect 10778 116016 10784 116028
rect 10836 116016 10842 116068
rect 14918 116056 14924 116068
rect 14879 116028 14924 116056
rect 14918 116016 14924 116028
rect 14976 116016 14982 116068
rect 16390 116056 16396 116068
rect 16351 116028 16396 116056
rect 16390 116016 16396 116028
rect 16448 116016 16454 116068
rect 21174 116056 21180 116068
rect 21135 116028 21180 116056
rect 21174 116016 21180 116028
rect 21232 116016 21238 116068
rect 22066 115988 22094 116164
rect 22462 116152 22468 116164
rect 22520 116152 22526 116204
rect 23124 116133 23152 116232
rect 27154 116220 27160 116232
rect 27212 116220 27218 116272
rect 27540 116260 27568 116300
rect 27617 116297 27629 116331
rect 27663 116328 27675 116331
rect 27706 116328 27712 116340
rect 27663 116300 27712 116328
rect 27663 116297 27675 116300
rect 27617 116291 27675 116297
rect 27706 116288 27712 116300
rect 27764 116288 27770 116340
rect 28258 116288 28264 116340
rect 28316 116328 28322 116340
rect 28445 116331 28503 116337
rect 28445 116328 28457 116331
rect 28316 116300 28457 116328
rect 28316 116288 28322 116300
rect 28445 116297 28457 116300
rect 28491 116297 28503 116331
rect 28445 116291 28503 116297
rect 28718 116288 28724 116340
rect 28776 116328 28782 116340
rect 29181 116331 29239 116337
rect 29181 116328 29193 116331
rect 28776 116300 29193 116328
rect 28776 116288 28782 116300
rect 29181 116297 29193 116300
rect 29227 116297 29239 116331
rect 29181 116291 29239 116297
rect 29270 116288 29276 116340
rect 29328 116328 29334 116340
rect 29328 116300 31616 116328
rect 29328 116288 29334 116300
rect 30926 116260 30932 116272
rect 27540 116232 30932 116260
rect 30926 116220 30932 116232
rect 30984 116220 30990 116272
rect 31297 116263 31355 116269
rect 31297 116229 31309 116263
rect 31343 116260 31355 116263
rect 31478 116260 31484 116272
rect 31343 116232 31484 116260
rect 31343 116229 31355 116232
rect 31297 116223 31355 116229
rect 31478 116220 31484 116232
rect 31536 116220 31542 116272
rect 31588 116260 31616 116300
rect 32398 116288 32404 116340
rect 32456 116328 32462 116340
rect 32677 116331 32735 116337
rect 32677 116328 32689 116331
rect 32456 116300 32689 116328
rect 32456 116288 32462 116300
rect 32677 116297 32689 116300
rect 32723 116297 32735 116331
rect 32677 116291 32735 116297
rect 32766 116288 32772 116340
rect 32824 116328 32830 116340
rect 35710 116328 35716 116340
rect 32824 116300 35716 116328
rect 32824 116288 32830 116300
rect 35710 116288 35716 116300
rect 35768 116288 35774 116340
rect 35894 116328 35900 116340
rect 35855 116300 35900 116328
rect 35894 116288 35900 116300
rect 35952 116288 35958 116340
rect 31665 116263 31723 116269
rect 31665 116260 31677 116263
rect 31588 116232 31677 116260
rect 31665 116229 31677 116232
rect 31711 116229 31723 116263
rect 32214 116260 32220 116272
rect 31665 116223 31723 116229
rect 31864 116232 32220 116260
rect 25225 116195 25283 116201
rect 25225 116161 25237 116195
rect 25271 116192 25283 116195
rect 29822 116192 29828 116204
rect 25271 116164 29828 116192
rect 25271 116161 25283 116164
rect 25225 116155 25283 116161
rect 29822 116152 29828 116164
rect 29880 116152 29886 116204
rect 31386 116192 31392 116204
rect 31347 116164 31392 116192
rect 31386 116152 31392 116164
rect 31444 116152 31450 116204
rect 31570 116152 31576 116204
rect 31628 116192 31634 116204
rect 31864 116192 31892 116232
rect 32214 116220 32220 116232
rect 32272 116220 32278 116272
rect 32493 116263 32551 116269
rect 32493 116229 32505 116263
rect 32539 116260 32551 116263
rect 32858 116260 32864 116272
rect 32539 116232 32864 116260
rect 32539 116229 32551 116232
rect 32493 116223 32551 116229
rect 32858 116220 32864 116232
rect 32916 116220 32922 116272
rect 33686 116260 33692 116272
rect 33647 116232 33692 116260
rect 33686 116220 33692 116232
rect 33744 116220 33750 116272
rect 34238 116220 34244 116272
rect 34296 116260 34302 116272
rect 36354 116260 36360 116272
rect 34296 116232 36360 116260
rect 34296 116220 34302 116232
rect 36354 116220 36360 116232
rect 36412 116220 36418 116272
rect 37093 116263 37151 116269
rect 37093 116229 37105 116263
rect 37139 116260 37151 116263
rect 38010 116260 38016 116272
rect 37139 116232 38016 116260
rect 37139 116229 37151 116232
rect 37093 116223 37151 116229
rect 38010 116220 38016 116232
rect 38068 116220 38074 116272
rect 31628 116164 31892 116192
rect 31628 116152 31634 116164
rect 32030 116152 32036 116204
rect 32088 116192 32094 116204
rect 32364 116195 32422 116201
rect 32364 116192 32376 116195
rect 32088 116164 32376 116192
rect 32088 116152 32094 116164
rect 32364 116161 32376 116164
rect 32410 116161 32422 116195
rect 32582 116192 32588 116204
rect 32543 116164 32588 116192
rect 32364 116155 32422 116161
rect 32582 116152 32588 116164
rect 32640 116152 32646 116204
rect 33502 116152 33508 116204
rect 33560 116201 33566 116204
rect 33560 116195 33618 116201
rect 33560 116161 33572 116195
rect 33606 116161 33618 116195
rect 33778 116192 33784 116204
rect 33739 116164 33784 116192
rect 33560 116155 33618 116161
rect 33560 116152 33566 116155
rect 33778 116152 33784 116164
rect 33836 116152 33842 116204
rect 37737 116195 37795 116201
rect 37737 116192 37749 116195
rect 33888 116164 37749 116192
rect 23109 116127 23167 116133
rect 23109 116093 23121 116127
rect 23155 116093 23167 116127
rect 23109 116087 23167 116093
rect 23474 116084 23480 116136
rect 23532 116124 23538 116136
rect 23532 116096 26924 116124
rect 23532 116084 23538 116096
rect 23937 116059 23995 116065
rect 23937 116025 23949 116059
rect 23983 116056 23995 116059
rect 26694 116056 26700 116068
rect 23983 116028 26700 116056
rect 23983 116025 23995 116028
rect 23937 116019 23995 116025
rect 26694 116016 26700 116028
rect 26752 116016 26758 116068
rect 26789 116059 26847 116065
rect 26789 116025 26801 116059
rect 26835 116025 26847 116059
rect 26896 116056 26924 116096
rect 26970 116084 26976 116136
rect 27028 116124 27034 116136
rect 29089 116127 29147 116133
rect 29089 116124 29101 116127
rect 27028 116096 29101 116124
rect 27028 116084 27034 116096
rect 29089 116093 29101 116096
rect 29135 116093 29147 116127
rect 29089 116087 29147 116093
rect 31168 116127 31226 116133
rect 31168 116093 31180 116127
rect 31214 116124 31226 116127
rect 31662 116124 31668 116136
rect 31214 116096 31668 116124
rect 31214 116093 31226 116096
rect 31168 116087 31226 116093
rect 31662 116084 31668 116096
rect 31720 116084 31726 116136
rect 31754 116084 31760 116136
rect 31812 116124 31818 116136
rect 33888 116124 33916 116164
rect 37737 116161 37749 116164
rect 37783 116161 37795 116195
rect 37737 116155 37795 116161
rect 31812 116096 33916 116124
rect 31812 116084 31818 116096
rect 34514 116084 34520 116136
rect 34572 116124 34578 116136
rect 34793 116127 34851 116133
rect 34793 116124 34805 116127
rect 34572 116096 34805 116124
rect 34572 116084 34578 116096
rect 34793 116093 34805 116096
rect 34839 116093 34851 116127
rect 34793 116087 34851 116093
rect 34882 116084 34888 116136
rect 34940 116124 34946 116136
rect 36078 116124 36084 116136
rect 34940 116096 36084 116124
rect 34940 116084 34946 116096
rect 36078 116084 36084 116096
rect 36136 116084 36142 116136
rect 37550 116124 37556 116136
rect 37511 116096 37556 116124
rect 37550 116084 37556 116096
rect 37608 116084 37614 116136
rect 28353 116059 28411 116065
rect 28353 116056 28365 116059
rect 26896 116028 28365 116056
rect 26789 116019 26847 116025
rect 28353 116025 28365 116028
rect 28399 116025 28411 116059
rect 28353 116019 28411 116025
rect 24670 115988 24676 116000
rect 22066 115960 24676 115988
rect 24670 115948 24676 115960
rect 24728 115948 24734 116000
rect 25866 115988 25872 116000
rect 25827 115960 25872 115988
rect 25866 115948 25872 115960
rect 25924 115948 25930 116000
rect 26804 115988 26832 116019
rect 28718 116016 28724 116068
rect 28776 116056 28782 116068
rect 30926 116056 30932 116068
rect 28776 116028 30932 116056
rect 28776 116016 28782 116028
rect 30926 116016 30932 116028
rect 30984 116016 30990 116068
rect 31021 116059 31079 116065
rect 31021 116025 31033 116059
rect 31067 116025 31079 116059
rect 31021 116019 31079 116025
rect 32217 116059 32275 116065
rect 32217 116025 32229 116059
rect 32263 116056 32275 116059
rect 33226 116056 33232 116068
rect 32263 116028 33232 116056
rect 32263 116025 32275 116028
rect 32217 116019 32275 116025
rect 30282 115988 30288 116000
rect 26804 115960 30288 115988
rect 30282 115948 30288 115960
rect 30340 115948 30346 116000
rect 31036 115988 31064 116019
rect 33226 116016 33232 116028
rect 33284 116016 33290 116068
rect 33413 116059 33471 116065
rect 33413 116025 33425 116059
rect 33459 116056 33471 116059
rect 35802 116056 35808 116068
rect 33459 116028 34652 116056
rect 35763 116028 35808 116056
rect 33459 116025 33471 116028
rect 33413 116019 33471 116025
rect 31202 115988 31208 116000
rect 31036 115960 31208 115988
rect 31202 115948 31208 115960
rect 31260 115948 31266 116000
rect 32766 115948 32772 116000
rect 32824 115988 32830 116000
rect 33042 115988 33048 116000
rect 32824 115960 33048 115988
rect 32824 115948 32830 115960
rect 33042 115948 33048 115960
rect 33100 115948 33106 116000
rect 34057 115991 34115 115997
rect 34057 115957 34069 115991
rect 34103 115988 34115 115991
rect 34330 115988 34336 116000
rect 34103 115960 34336 115988
rect 34103 115957 34115 115960
rect 34057 115951 34115 115957
rect 34330 115948 34336 115960
rect 34388 115948 34394 116000
rect 34624 115997 34652 116028
rect 35802 116016 35808 116028
rect 35860 116016 35866 116068
rect 36909 116059 36967 116065
rect 36909 116025 36921 116059
rect 36955 116056 36967 116059
rect 36998 116056 37004 116068
rect 36955 116028 37004 116056
rect 36955 116025 36967 116028
rect 36909 116019 36967 116025
rect 36998 116016 37004 116028
rect 37056 116016 37062 116068
rect 34609 115991 34667 115997
rect 34609 115957 34621 115991
rect 34655 115957 34667 115991
rect 34609 115951 34667 115957
rect 1104 115898 38824 115920
rect 1104 115846 19606 115898
rect 19658 115846 19670 115898
rect 19722 115846 19734 115898
rect 19786 115846 19798 115898
rect 19850 115846 38824 115898
rect 1104 115824 38824 115846
rect 566 115744 572 115796
rect 624 115784 630 115796
rect 2958 115784 2964 115796
rect 624 115756 2964 115784
rect 624 115744 630 115756
rect 2958 115744 2964 115756
rect 3016 115744 3022 115796
rect 3050 115744 3056 115796
rect 3108 115784 3114 115796
rect 3237 115787 3295 115793
rect 3237 115784 3249 115787
rect 3108 115756 3249 115784
rect 3108 115744 3114 115756
rect 3237 115753 3249 115756
rect 3283 115753 3295 115787
rect 3237 115747 3295 115753
rect 3510 115744 3516 115796
rect 3568 115784 3574 115796
rect 3568 115756 5120 115784
rect 3568 115744 3574 115756
rect 4709 115719 4767 115725
rect 4709 115685 4721 115719
rect 4755 115716 4767 115719
rect 4798 115716 4804 115728
rect 4755 115688 4804 115716
rect 4755 115685 4767 115688
rect 4709 115679 4767 115685
rect 4798 115676 4804 115688
rect 4856 115676 4862 115728
rect 5092 115716 5120 115756
rect 5166 115744 5172 115796
rect 5224 115784 5230 115796
rect 5353 115787 5411 115793
rect 5353 115784 5365 115787
rect 5224 115756 5365 115784
rect 5224 115744 5230 115756
rect 5353 115753 5365 115756
rect 5399 115753 5411 115787
rect 7834 115784 7840 115796
rect 5353 115747 5411 115753
rect 7208 115756 7840 115784
rect 7208 115716 7236 115756
rect 7834 115744 7840 115756
rect 7892 115744 7898 115796
rect 8018 115744 8024 115796
rect 8076 115784 8082 115796
rect 8113 115787 8171 115793
rect 8113 115784 8125 115787
rect 8076 115756 8125 115784
rect 8076 115744 8082 115756
rect 8113 115753 8125 115756
rect 8159 115753 8171 115787
rect 8113 115747 8171 115753
rect 8665 115787 8723 115793
rect 8665 115753 8677 115787
rect 8711 115784 8723 115787
rect 9122 115784 9128 115796
rect 8711 115756 9128 115784
rect 8711 115753 8723 115756
rect 8665 115747 8723 115753
rect 9122 115744 9128 115756
rect 9180 115744 9186 115796
rect 22557 115787 22615 115793
rect 22557 115753 22569 115787
rect 22603 115784 22615 115787
rect 23474 115784 23480 115796
rect 22603 115756 23480 115784
rect 22603 115753 22615 115756
rect 22557 115747 22615 115753
rect 23474 115744 23480 115756
rect 23532 115744 23538 115796
rect 23569 115787 23627 115793
rect 23569 115753 23581 115787
rect 23615 115784 23627 115787
rect 24762 115784 24768 115796
rect 23615 115756 24768 115784
rect 23615 115753 23627 115756
rect 23569 115747 23627 115753
rect 24762 115744 24768 115756
rect 24820 115744 24826 115796
rect 24949 115787 25007 115793
rect 24949 115753 24961 115787
rect 24995 115784 25007 115787
rect 24995 115756 29132 115784
rect 24995 115753 25007 115756
rect 24949 115747 25007 115753
rect 5092 115688 7236 115716
rect 7285 115719 7343 115725
rect 7285 115685 7297 115719
rect 7331 115716 7343 115719
rect 8386 115716 8392 115728
rect 7331 115688 8392 115716
rect 7331 115685 7343 115688
rect 7285 115679 7343 115685
rect 8386 115676 8392 115688
rect 8444 115676 8450 115728
rect 21358 115676 21364 115728
rect 21416 115716 21422 115728
rect 21910 115716 21916 115728
rect 21416 115688 21916 115716
rect 21416 115676 21422 115688
rect 21910 115676 21916 115688
rect 21968 115676 21974 115728
rect 23400 115688 25176 115716
rect 1857 115651 1915 115657
rect 1857 115617 1869 115651
rect 1903 115617 1915 115651
rect 1857 115611 1915 115617
rect 3145 115651 3203 115657
rect 3145 115617 3157 115651
rect 3191 115648 3203 115651
rect 4062 115648 4068 115660
rect 3191 115620 4068 115648
rect 3191 115617 3203 115620
rect 3145 115611 3203 115617
rect 1872 115580 1900 115611
rect 4062 115608 4068 115620
rect 4120 115608 4126 115660
rect 4525 115651 4583 115657
rect 4525 115617 4537 115651
rect 4571 115648 4583 115651
rect 4614 115648 4620 115660
rect 4571 115620 4620 115648
rect 4571 115617 4583 115620
rect 4525 115611 4583 115617
rect 4614 115608 4620 115620
rect 4672 115608 4678 115660
rect 5258 115648 5264 115660
rect 5219 115620 5264 115648
rect 5258 115608 5264 115620
rect 5316 115608 5322 115660
rect 8021 115651 8079 115657
rect 8021 115617 8033 115651
rect 8067 115648 8079 115651
rect 8294 115648 8300 115660
rect 8067 115620 8300 115648
rect 8067 115617 8079 115620
rect 8021 115611 8079 115617
rect 8294 115608 8300 115620
rect 8352 115608 8358 115660
rect 9493 115651 9551 115657
rect 9493 115617 9505 115651
rect 9539 115648 9551 115651
rect 9674 115648 9680 115660
rect 9539 115620 9680 115648
rect 9539 115617 9551 115620
rect 9493 115611 9551 115617
rect 9674 115608 9680 115620
rect 9732 115608 9738 115660
rect 10137 115651 10195 115657
rect 10137 115617 10149 115651
rect 10183 115648 10195 115651
rect 10410 115648 10416 115660
rect 10183 115620 10416 115648
rect 10183 115617 10195 115620
rect 10137 115611 10195 115617
rect 10410 115608 10416 115620
rect 10468 115608 10474 115660
rect 10781 115651 10839 115657
rect 10781 115617 10793 115651
rect 10827 115648 10839 115651
rect 11146 115648 11152 115660
rect 10827 115620 11152 115648
rect 10827 115617 10839 115620
rect 10781 115611 10839 115617
rect 11146 115608 11152 115620
rect 11204 115608 11210 115660
rect 12158 115608 12164 115660
rect 12216 115648 12222 115660
rect 12253 115651 12311 115657
rect 12253 115648 12265 115651
rect 12216 115620 12265 115648
rect 12216 115608 12222 115620
rect 12253 115617 12265 115620
rect 12299 115617 12311 115651
rect 12894 115648 12900 115660
rect 12855 115620 12900 115648
rect 12253 115611 12311 115617
rect 12894 115608 12900 115620
rect 12952 115608 12958 115660
rect 15102 115608 15108 115660
rect 15160 115648 15166 115660
rect 15289 115651 15347 115657
rect 15289 115648 15301 115651
rect 15160 115620 15301 115648
rect 15160 115608 15166 115620
rect 15289 115617 15301 115620
rect 15335 115617 15347 115651
rect 15289 115611 15347 115617
rect 16025 115651 16083 115657
rect 16025 115617 16037 115651
rect 16071 115648 16083 115651
rect 17310 115648 17316 115660
rect 16071 115620 17316 115648
rect 16071 115617 16083 115620
rect 16025 115611 16083 115617
rect 17310 115608 17316 115620
rect 17368 115608 17374 115660
rect 17402 115608 17408 115660
rect 17460 115648 17466 115660
rect 17497 115651 17555 115657
rect 17497 115648 17509 115651
rect 17460 115620 17509 115648
rect 17460 115608 17466 115620
rect 17497 115617 17509 115620
rect 17543 115617 17555 115651
rect 18138 115648 18144 115660
rect 18099 115620 18144 115648
rect 17497 115611 17555 115617
rect 18138 115608 18144 115620
rect 18196 115608 18202 115660
rect 19426 115648 19432 115660
rect 19387 115620 19432 115648
rect 19426 115608 19432 115620
rect 19484 115608 19490 115660
rect 20165 115651 20223 115657
rect 20165 115617 20177 115651
rect 20211 115648 20223 115651
rect 20714 115648 20720 115660
rect 20211 115620 20720 115648
rect 20211 115617 20223 115620
rect 20165 115611 20223 115617
rect 20714 115608 20720 115620
rect 20772 115608 20778 115660
rect 21174 115608 21180 115660
rect 21232 115648 21238 115660
rect 21545 115651 21603 115657
rect 21545 115648 21557 115651
rect 21232 115620 21557 115648
rect 21232 115608 21238 115620
rect 21545 115617 21557 115620
rect 21591 115617 21603 115651
rect 21545 115611 21603 115617
rect 22741 115651 22799 115657
rect 22741 115617 22753 115651
rect 22787 115617 22799 115651
rect 22741 115611 22799 115617
rect 2961 115583 3019 115589
rect 2961 115580 2973 115583
rect 1872 115552 2973 115580
rect 2961 115549 2973 115552
rect 3007 115549 3019 115583
rect 2961 115543 3019 115549
rect 3234 115540 3240 115592
rect 3292 115580 3298 115592
rect 3973 115583 4031 115589
rect 3973 115580 3985 115583
rect 3292 115552 3985 115580
rect 3292 115540 3298 115552
rect 3973 115549 3985 115552
rect 4019 115549 4031 115583
rect 3973 115543 4031 115549
rect 4430 115540 4436 115592
rect 4488 115580 4494 115592
rect 4798 115580 4804 115592
rect 4488 115552 4804 115580
rect 4488 115540 4494 115552
rect 4798 115540 4804 115552
rect 4856 115540 4862 115592
rect 5166 115540 5172 115592
rect 5224 115580 5230 115592
rect 8478 115580 8484 115592
rect 5224 115552 8484 115580
rect 5224 115540 5230 115552
rect 8478 115540 8484 115552
rect 8536 115540 8542 115592
rect 13909 115583 13967 115589
rect 13909 115549 13921 115583
rect 13955 115580 13967 115583
rect 15194 115580 15200 115592
rect 13955 115552 15200 115580
rect 13955 115549 13967 115552
rect 13909 115543 13967 115549
rect 15194 115540 15200 115552
rect 15252 115540 15258 115592
rect 16114 115540 16120 115592
rect 16172 115580 16178 115592
rect 17586 115580 17592 115592
rect 16172 115552 17592 115580
rect 16172 115540 16178 115552
rect 17586 115540 17592 115552
rect 17644 115540 17650 115592
rect 18785 115583 18843 115589
rect 18785 115549 18797 115583
rect 18831 115580 18843 115583
rect 20438 115580 20444 115592
rect 18831 115552 20444 115580
rect 18831 115549 18843 115552
rect 18785 115543 18843 115549
rect 20438 115540 20444 115552
rect 20496 115540 20502 115592
rect 20901 115583 20959 115589
rect 20901 115549 20913 115583
rect 20947 115580 20959 115583
rect 22370 115580 22376 115592
rect 20947 115552 22376 115580
rect 20947 115549 20959 115552
rect 20901 115543 20959 115549
rect 22370 115540 22376 115552
rect 22428 115540 22434 115592
rect 1486 115472 1492 115524
rect 1544 115512 1550 115524
rect 6178 115512 6184 115524
rect 1544 115484 6184 115512
rect 1544 115472 1550 115484
rect 6178 115472 6184 115484
rect 6236 115472 6242 115524
rect 14645 115515 14703 115521
rect 14645 115481 14657 115515
rect 14691 115512 14703 115515
rect 16206 115512 16212 115524
rect 14691 115484 16212 115512
rect 14691 115481 14703 115484
rect 14645 115475 14703 115481
rect 16206 115472 16212 115484
rect 16264 115472 16270 115524
rect 17770 115472 17776 115524
rect 17828 115512 17834 115524
rect 22756 115512 22784 115611
rect 17828 115484 22784 115512
rect 17828 115472 17834 115484
rect 1946 115444 1952 115456
rect 1907 115416 1952 115444
rect 1946 115404 1952 115416
rect 2004 115404 2010 115456
rect 2961 115447 3019 115453
rect 2961 115413 2973 115447
rect 3007 115444 3019 115447
rect 7742 115444 7748 115456
rect 3007 115416 7748 115444
rect 3007 115413 3019 115416
rect 2961 115407 3019 115413
rect 7742 115404 7748 115416
rect 7800 115404 7806 115456
rect 20990 115404 20996 115456
rect 21048 115444 21054 115456
rect 23400 115444 23428 115688
rect 23658 115608 23664 115660
rect 23716 115648 23722 115660
rect 25148 115657 25176 115688
rect 25222 115676 25228 115728
rect 25280 115716 25286 115728
rect 26970 115716 26976 115728
rect 25280 115688 26976 115716
rect 25280 115676 25286 115688
rect 26970 115676 26976 115688
rect 27028 115676 27034 115728
rect 27062 115676 27068 115728
rect 27120 115716 27126 115728
rect 29104 115725 29132 115756
rect 29546 115744 29552 115796
rect 29604 115784 29610 115796
rect 29917 115787 29975 115793
rect 29917 115784 29929 115787
rect 29604 115756 29929 115784
rect 29604 115744 29610 115756
rect 29917 115753 29929 115756
rect 29963 115753 29975 115787
rect 29917 115747 29975 115753
rect 30282 115744 30288 115796
rect 30340 115784 30346 115796
rect 31205 115787 31263 115793
rect 31205 115784 31217 115787
rect 30340 115756 31217 115784
rect 30340 115744 30346 115756
rect 31205 115753 31217 115756
rect 31251 115753 31263 115787
rect 31205 115747 31263 115753
rect 34333 115787 34391 115793
rect 34333 115753 34345 115787
rect 34379 115784 34391 115787
rect 35342 115784 35348 115796
rect 34379 115756 35348 115784
rect 34379 115753 34391 115756
rect 34333 115747 34391 115753
rect 35342 115744 35348 115756
rect 35400 115744 35406 115796
rect 35710 115744 35716 115796
rect 35768 115784 35774 115796
rect 38654 115784 38660 115796
rect 35768 115756 38660 115784
rect 35768 115744 35774 115756
rect 38654 115744 38660 115756
rect 38712 115744 38718 115796
rect 29089 115719 29147 115725
rect 27120 115688 28948 115716
rect 27120 115676 27126 115688
rect 25133 115651 25191 115657
rect 23716 115620 25084 115648
rect 23716 115608 23722 115620
rect 24305 115583 24363 115589
rect 24305 115549 24317 115583
rect 24351 115580 24363 115583
rect 24946 115580 24952 115592
rect 24351 115552 24952 115580
rect 24351 115549 24363 115552
rect 24305 115543 24363 115549
rect 24946 115540 24952 115552
rect 25004 115540 25010 115592
rect 25056 115580 25084 115620
rect 25133 115617 25145 115651
rect 25179 115617 25191 115651
rect 25133 115611 25191 115617
rect 25869 115651 25927 115657
rect 25869 115617 25881 115651
rect 25915 115648 25927 115651
rect 25915 115620 27844 115648
rect 25915 115617 25927 115620
rect 25869 115611 25927 115617
rect 26329 115583 26387 115589
rect 25056 115552 26280 115580
rect 23474 115472 23480 115524
rect 23532 115512 23538 115524
rect 25222 115512 25228 115524
rect 23532 115484 25228 115512
rect 23532 115472 23538 115484
rect 25222 115472 25228 115484
rect 25280 115472 25286 115524
rect 25682 115512 25688 115524
rect 25643 115484 25688 115512
rect 25682 115472 25688 115484
rect 25740 115472 25746 115524
rect 26252 115512 26280 115552
rect 26329 115549 26341 115583
rect 26375 115580 26387 115583
rect 27706 115580 27712 115592
rect 26375 115552 27712 115580
rect 26375 115549 26387 115552
rect 26329 115543 26387 115549
rect 27706 115540 27712 115552
rect 27764 115540 27770 115592
rect 27816 115580 27844 115620
rect 27890 115608 27896 115660
rect 27948 115648 27954 115660
rect 27985 115651 28043 115657
rect 27985 115648 27997 115651
rect 27948 115620 27997 115648
rect 27948 115608 27954 115620
rect 27985 115617 27997 115620
rect 28031 115617 28043 115651
rect 27985 115611 28043 115617
rect 28074 115608 28080 115660
rect 28132 115648 28138 115660
rect 28810 115648 28816 115660
rect 28132 115620 28816 115648
rect 28132 115608 28138 115620
rect 28810 115608 28816 115620
rect 28868 115608 28874 115660
rect 28920 115648 28948 115688
rect 29089 115685 29101 115719
rect 29135 115685 29147 115719
rect 29089 115679 29147 115685
rect 29454 115676 29460 115728
rect 29512 115716 29518 115728
rect 30745 115719 30803 115725
rect 30745 115716 30757 115719
rect 29512 115688 30757 115716
rect 29512 115676 29518 115688
rect 30745 115685 30757 115688
rect 30791 115685 30803 115719
rect 30745 115679 30803 115685
rect 32125 115719 32183 115725
rect 32125 115685 32137 115719
rect 32171 115716 32183 115719
rect 34514 115716 34520 115728
rect 32171 115688 34520 115716
rect 32171 115685 32183 115688
rect 32125 115679 32183 115685
rect 34514 115676 34520 115688
rect 34572 115676 34578 115728
rect 35897 115719 35955 115725
rect 34900 115688 35112 115716
rect 29825 115651 29883 115657
rect 29825 115648 29837 115651
rect 28920 115620 29837 115648
rect 29825 115617 29837 115620
rect 29871 115617 29883 115651
rect 29825 115611 29883 115617
rect 30561 115651 30619 115657
rect 30561 115617 30573 115651
rect 30607 115617 30619 115651
rect 30561 115611 30619 115617
rect 29273 115583 29331 115589
rect 27816 115552 29132 115580
rect 28166 115512 28172 115524
rect 26252 115484 28172 115512
rect 28166 115472 28172 115484
rect 28224 115472 28230 115524
rect 29104 115512 29132 115552
rect 29273 115549 29285 115583
rect 29319 115580 29331 115583
rect 29546 115580 29552 115592
rect 29319 115552 29552 115580
rect 29319 115549 29331 115552
rect 29273 115543 29331 115549
rect 29546 115540 29552 115552
rect 29604 115540 29610 115592
rect 29178 115512 29184 115524
rect 29104 115484 29184 115512
rect 29178 115472 29184 115484
rect 29236 115472 29242 115524
rect 21048 115416 23428 115444
rect 21048 115404 21054 115416
rect 24210 115404 24216 115456
rect 24268 115444 24274 115456
rect 30576 115444 30604 115611
rect 30926 115608 30932 115660
rect 30984 115648 30990 115660
rect 31389 115651 31447 115657
rect 31389 115648 31401 115651
rect 30984 115620 31401 115648
rect 30984 115608 30990 115620
rect 31389 115617 31401 115620
rect 31435 115617 31447 115651
rect 31389 115611 31447 115617
rect 31754 115608 31760 115660
rect 31812 115648 31818 115660
rect 31941 115651 31999 115657
rect 31941 115648 31953 115651
rect 31812 115620 31953 115648
rect 31812 115608 31818 115620
rect 31941 115617 31953 115620
rect 31987 115617 31999 115651
rect 31941 115611 31999 115617
rect 33505 115651 33563 115657
rect 33505 115617 33517 115651
rect 33551 115648 33563 115651
rect 33594 115648 33600 115660
rect 33551 115620 33600 115648
rect 33551 115617 33563 115620
rect 33505 115611 33563 115617
rect 33594 115608 33600 115620
rect 33652 115608 33658 115660
rect 34241 115651 34299 115657
rect 34241 115617 34253 115651
rect 34287 115648 34299 115651
rect 34900 115648 34928 115688
rect 34287 115620 34928 115648
rect 34977 115651 35035 115657
rect 34287 115617 34299 115620
rect 34241 115611 34299 115617
rect 34977 115617 34989 115651
rect 35023 115617 35035 115651
rect 34977 115611 35035 115617
rect 33689 115583 33747 115589
rect 33689 115549 33701 115583
rect 33735 115580 33747 115583
rect 34790 115580 34796 115592
rect 33735 115552 34796 115580
rect 33735 115549 33747 115552
rect 33689 115543 33747 115549
rect 34790 115540 34796 115552
rect 34848 115540 34854 115592
rect 24268 115416 30604 115444
rect 24268 115404 24274 115416
rect 31570 115404 31576 115456
rect 31628 115444 31634 115456
rect 33318 115444 33324 115456
rect 31628 115416 33324 115444
rect 31628 115404 31634 115416
rect 33318 115404 33324 115416
rect 33376 115404 33382 115456
rect 34992 115444 35020 115611
rect 35084 115512 35112 115688
rect 35897 115685 35909 115719
rect 35943 115716 35955 115719
rect 36170 115716 36176 115728
rect 35943 115688 36176 115716
rect 35943 115685 35955 115688
rect 35897 115679 35955 115685
rect 36170 115676 36176 115688
rect 36228 115676 36234 115728
rect 36354 115676 36360 115728
rect 36412 115716 36418 115728
rect 39574 115716 39580 115728
rect 36412 115688 39580 115716
rect 36412 115676 36418 115688
rect 39574 115676 39580 115688
rect 39632 115676 39638 115728
rect 35710 115648 35716 115660
rect 35671 115620 35716 115648
rect 35710 115608 35716 115620
rect 35768 115608 35774 115660
rect 35986 115608 35992 115660
rect 36044 115648 36050 115660
rect 36449 115651 36507 115657
rect 36449 115648 36461 115651
rect 36044 115620 36461 115648
rect 36044 115608 36050 115620
rect 36449 115617 36461 115620
rect 36495 115617 36507 115651
rect 36449 115611 36507 115617
rect 36814 115608 36820 115660
rect 36872 115648 36878 115660
rect 37185 115651 37243 115657
rect 37185 115648 37197 115651
rect 36872 115620 37197 115648
rect 36872 115608 36878 115620
rect 37185 115617 37197 115620
rect 37231 115617 37243 115651
rect 37185 115611 37243 115617
rect 35161 115583 35219 115589
rect 35161 115549 35173 115583
rect 35207 115580 35219 115583
rect 37274 115580 37280 115592
rect 35207 115552 37280 115580
rect 35207 115549 35219 115552
rect 35161 115543 35219 115549
rect 37274 115540 37280 115552
rect 37332 115540 37338 115592
rect 36354 115512 36360 115524
rect 35084 115484 36360 115512
rect 36354 115472 36360 115484
rect 36412 115472 36418 115524
rect 37366 115512 37372 115524
rect 37327 115484 37372 115512
rect 37366 115472 37372 115484
rect 37424 115472 37430 115524
rect 35250 115444 35256 115456
rect 34992 115416 35256 115444
rect 35250 115404 35256 115416
rect 35308 115404 35314 115456
rect 36538 115444 36544 115456
rect 36499 115416 36544 115444
rect 36538 115404 36544 115416
rect 36596 115404 36602 115456
rect 1104 115354 38824 115376
rect 1104 115302 4246 115354
rect 4298 115302 4310 115354
rect 4362 115302 4374 115354
rect 4426 115302 4438 115354
rect 4490 115302 34966 115354
rect 35018 115302 35030 115354
rect 35082 115302 35094 115354
rect 35146 115302 35158 115354
rect 35210 115302 38824 115354
rect 1104 115280 38824 115302
rect 1394 115200 1400 115252
rect 1452 115240 1458 115252
rect 1949 115243 2007 115249
rect 1949 115240 1961 115243
rect 1452 115212 1961 115240
rect 1452 115200 1458 115212
rect 1949 115209 1961 115212
rect 1995 115209 2007 115243
rect 1949 115203 2007 115209
rect 5074 115200 5080 115252
rect 5132 115240 5138 115252
rect 5721 115243 5779 115249
rect 5721 115240 5733 115243
rect 5132 115212 5733 115240
rect 5132 115200 5138 115212
rect 5721 115209 5733 115212
rect 5767 115209 5779 115243
rect 5721 115203 5779 115209
rect 6365 115243 6423 115249
rect 6365 115209 6377 115243
rect 6411 115240 6423 115243
rect 6914 115240 6920 115252
rect 6411 115212 6920 115240
rect 6411 115209 6423 115212
rect 6365 115203 6423 115209
rect 6914 115200 6920 115212
rect 6972 115200 6978 115252
rect 7009 115243 7067 115249
rect 7009 115209 7021 115243
rect 7055 115240 7067 115243
rect 7098 115240 7104 115252
rect 7055 115212 7104 115240
rect 7055 115209 7067 115212
rect 7009 115203 7067 115209
rect 7098 115200 7104 115212
rect 7156 115200 7162 115252
rect 7653 115243 7711 115249
rect 7653 115209 7665 115243
rect 7699 115240 7711 115243
rect 7926 115240 7932 115252
rect 7699 115212 7932 115240
rect 7699 115209 7711 115212
rect 7653 115203 7711 115209
rect 7926 115200 7932 115212
rect 7984 115200 7990 115252
rect 8294 115240 8300 115252
rect 8255 115212 8300 115240
rect 8294 115200 8300 115212
rect 8352 115200 8358 115252
rect 9677 115243 9735 115249
rect 9677 115209 9689 115243
rect 9723 115240 9735 115243
rect 9858 115240 9864 115252
rect 9723 115212 9864 115240
rect 9723 115209 9735 115212
rect 9677 115203 9735 115209
rect 9858 115200 9864 115212
rect 9916 115200 9922 115252
rect 10321 115243 10379 115249
rect 10321 115209 10333 115243
rect 10367 115240 10379 115243
rect 10594 115240 10600 115252
rect 10367 115212 10600 115240
rect 10367 115209 10379 115212
rect 10321 115203 10379 115209
rect 10594 115200 10600 115212
rect 10652 115200 10658 115252
rect 10778 115200 10784 115252
rect 10836 115240 10842 115252
rect 10965 115243 11023 115249
rect 10965 115240 10977 115243
rect 10836 115212 10977 115240
rect 10836 115200 10842 115212
rect 10965 115209 10977 115212
rect 11011 115209 11023 115243
rect 10965 115203 11023 115209
rect 12805 115243 12863 115249
rect 12805 115209 12817 115243
rect 12851 115240 12863 115243
rect 12986 115240 12992 115252
rect 12851 115212 12992 115240
rect 12851 115209 12863 115212
rect 12805 115203 12863 115209
rect 12986 115200 12992 115212
rect 13044 115200 13050 115252
rect 13449 115243 13507 115249
rect 13449 115209 13461 115243
rect 13495 115240 13507 115243
rect 14366 115240 14372 115252
rect 13495 115212 14372 115240
rect 13495 115209 13507 115212
rect 13449 115203 13507 115209
rect 14366 115200 14372 115212
rect 14424 115200 14430 115252
rect 14918 115240 14924 115252
rect 14879 115212 14924 115240
rect 14918 115200 14924 115212
rect 14976 115200 14982 115252
rect 15565 115243 15623 115249
rect 15565 115209 15577 115243
rect 15611 115240 15623 115243
rect 15838 115240 15844 115252
rect 15611 115212 15844 115240
rect 15611 115209 15623 115212
rect 15565 115203 15623 115209
rect 15838 115200 15844 115212
rect 15896 115200 15902 115252
rect 16301 115243 16359 115249
rect 16301 115209 16313 115243
rect 16347 115240 16359 115243
rect 16390 115240 16396 115252
rect 16347 115212 16396 115240
rect 16347 115209 16359 115212
rect 16301 115203 16359 115209
rect 16390 115200 16396 115212
rect 16448 115200 16454 115252
rect 18325 115243 18383 115249
rect 18325 115209 18337 115243
rect 18371 115240 18383 115243
rect 18874 115240 18880 115252
rect 18371 115212 18880 115240
rect 18371 115209 18383 115212
rect 18325 115203 18383 115209
rect 18874 115200 18880 115212
rect 18932 115200 18938 115252
rect 20165 115243 20223 115249
rect 20165 115209 20177 115243
rect 20211 115240 20223 115243
rect 20346 115240 20352 115252
rect 20211 115212 20352 115240
rect 20211 115209 20223 115212
rect 20165 115203 20223 115209
rect 20346 115200 20352 115212
rect 20404 115200 20410 115252
rect 20809 115243 20867 115249
rect 20809 115209 20821 115243
rect 20855 115240 20867 115243
rect 21082 115240 21088 115252
rect 20855 115212 21088 115240
rect 20855 115209 20867 115212
rect 20809 115203 20867 115209
rect 21082 115200 21088 115212
rect 21140 115200 21146 115252
rect 25406 115200 25412 115252
rect 25464 115240 25470 115252
rect 26237 115243 26295 115249
rect 26237 115240 26249 115243
rect 25464 115212 26249 115240
rect 25464 115200 25470 115212
rect 26237 115209 26249 115212
rect 26283 115209 26295 115243
rect 26237 115203 26295 115209
rect 28077 115243 28135 115249
rect 28077 115209 28089 115243
rect 28123 115240 28135 115243
rect 28626 115240 28632 115252
rect 28123 115212 28632 115240
rect 28123 115209 28135 115212
rect 28077 115203 28135 115209
rect 28626 115200 28632 115212
rect 28684 115200 28690 115252
rect 28902 115200 28908 115252
rect 28960 115240 28966 115252
rect 29181 115243 29239 115249
rect 29181 115240 29193 115243
rect 28960 115212 29193 115240
rect 28960 115200 28966 115212
rect 29181 115209 29193 115212
rect 29227 115209 29239 115243
rect 29181 115203 29239 115209
rect 29638 115200 29644 115252
rect 29696 115240 29702 115252
rect 30653 115243 30711 115249
rect 30653 115240 30665 115243
rect 29696 115212 30665 115240
rect 29696 115200 29702 115212
rect 30653 115209 30665 115212
rect 30699 115209 30711 115243
rect 30653 115203 30711 115209
rect 31297 115243 31355 115249
rect 31297 115209 31309 115243
rect 31343 115240 31355 115243
rect 31386 115240 31392 115252
rect 31343 115212 31392 115240
rect 31343 115209 31355 115212
rect 31297 115203 31355 115209
rect 31386 115200 31392 115212
rect 31444 115200 31450 115252
rect 31478 115200 31484 115252
rect 31536 115240 31542 115252
rect 31941 115243 31999 115249
rect 31941 115240 31953 115243
rect 31536 115212 31953 115240
rect 31536 115200 31542 115212
rect 31941 115209 31953 115212
rect 31987 115209 31999 115243
rect 31941 115203 31999 115209
rect 33965 115243 34023 115249
rect 33965 115209 33977 115243
rect 34011 115240 34023 115243
rect 35342 115240 35348 115252
rect 34011 115212 35348 115240
rect 34011 115209 34023 115212
rect 33965 115203 34023 115209
rect 35342 115200 35348 115212
rect 35400 115200 35406 115252
rect 2774 115132 2780 115184
rect 2832 115172 2838 115184
rect 4433 115175 4491 115181
rect 2832 115144 2877 115172
rect 2832 115132 2838 115144
rect 4433 115141 4445 115175
rect 4479 115172 4491 115175
rect 5534 115172 5540 115184
rect 4479 115144 5540 115172
rect 4479 115141 4491 115144
rect 4433 115135 4491 115141
rect 5534 115132 5540 115144
rect 5592 115132 5598 115184
rect 11425 115175 11483 115181
rect 11425 115172 11437 115175
rect 6932 115144 11437 115172
rect 6932 115116 6960 115144
rect 11425 115141 11437 115144
rect 11471 115141 11483 115175
rect 11425 115135 11483 115141
rect 18785 115175 18843 115181
rect 18785 115141 18797 115175
rect 18831 115172 18843 115175
rect 21450 115172 21456 115184
rect 18831 115144 21456 115172
rect 18831 115141 18843 115144
rect 18785 115135 18843 115141
rect 21450 115132 21456 115144
rect 21508 115132 21514 115184
rect 22741 115175 22799 115181
rect 22741 115141 22753 115175
rect 22787 115172 22799 115175
rect 24026 115172 24032 115184
rect 22787 115144 24032 115172
rect 22787 115141 22799 115144
rect 22741 115135 22799 115141
rect 24026 115132 24032 115144
rect 24084 115132 24090 115184
rect 24121 115175 24179 115181
rect 24121 115141 24133 115175
rect 24167 115172 24179 115175
rect 24210 115172 24216 115184
rect 24167 115144 24216 115172
rect 24167 115141 24179 115144
rect 24121 115135 24179 115141
rect 24210 115132 24216 115144
rect 24268 115132 24274 115184
rect 25225 115175 25283 115181
rect 25225 115141 25237 115175
rect 25271 115172 25283 115175
rect 30006 115172 30012 115184
rect 25271 115144 30012 115172
rect 25271 115141 25283 115144
rect 25225 115135 25283 115141
rect 30006 115132 30012 115144
rect 30064 115132 30070 115184
rect 32122 115172 32128 115184
rect 31726 115144 32128 115172
rect 2608 115076 4936 115104
rect 2608 115045 2636 115076
rect 2593 115039 2651 115045
rect 2593 115005 2605 115039
rect 2639 115005 2651 115039
rect 2593 114999 2651 115005
rect 1857 114971 1915 114977
rect 1857 114937 1869 114971
rect 1903 114968 1915 114971
rect 4908 114968 4936 115076
rect 4982 115064 4988 115116
rect 5040 115104 5046 115116
rect 5077 115107 5135 115113
rect 5077 115104 5089 115107
rect 5040 115076 5089 115104
rect 5040 115064 5046 115076
rect 5077 115073 5089 115076
rect 5123 115073 5135 115107
rect 5077 115067 5135 115073
rect 6914 115064 6920 115116
rect 6972 115064 6978 115116
rect 8754 115064 8760 115116
rect 8812 115104 8818 115116
rect 15286 115104 15292 115116
rect 8812 115076 15292 115104
rect 8812 115064 8818 115076
rect 15286 115064 15292 115076
rect 15344 115064 15350 115116
rect 21818 115064 21824 115116
rect 21876 115104 21882 115116
rect 21876 115076 24348 115104
rect 21876 115064 21882 115076
rect 8662 115036 8668 115048
rect 7208 115008 8668 115036
rect 7208 114968 7236 115008
rect 8662 114996 8668 115008
rect 8720 114996 8726 115048
rect 10962 114996 10968 115048
rect 11020 115036 11026 115048
rect 11609 115039 11667 115045
rect 11609 115036 11621 115039
rect 11020 115008 11621 115036
rect 11020 114996 11026 115008
rect 11609 115005 11621 115008
rect 11655 115005 11667 115039
rect 11609 114999 11667 115005
rect 16482 114996 16488 115048
rect 16540 115036 16546 115048
rect 16945 115039 17003 115045
rect 16945 115036 16957 115039
rect 16540 115008 16957 115036
rect 16540 114996 16546 115008
rect 16945 115005 16957 115008
rect 16991 115005 17003 115039
rect 16945 114999 17003 115005
rect 17218 114996 17224 115048
rect 17276 115036 17282 115048
rect 17589 115039 17647 115045
rect 17589 115036 17601 115039
rect 17276 115008 17601 115036
rect 17276 114996 17282 115008
rect 17589 115005 17601 115008
rect 17635 115005 17647 115039
rect 17589 114999 17647 115005
rect 18598 114996 18604 115048
rect 18656 115036 18662 115048
rect 18969 115039 19027 115045
rect 18969 115036 18981 115039
rect 18656 115008 18981 115036
rect 18656 114996 18662 115008
rect 18969 115005 18981 115008
rect 19015 115005 19027 115039
rect 18969 114999 19027 115005
rect 20622 114996 20628 115048
rect 20680 115036 20686 115048
rect 21453 115039 21511 115045
rect 21453 115036 21465 115039
rect 20680 115008 21465 115036
rect 20680 114996 20686 115008
rect 21453 115005 21465 115008
rect 21499 115005 21511 115039
rect 21453 114999 21511 115005
rect 21910 114996 21916 115048
rect 21968 115036 21974 115048
rect 21968 115008 22013 115036
rect 21968 114996 21974 115008
rect 22462 114996 22468 115048
rect 22520 115036 22526 115048
rect 22925 115039 22983 115045
rect 22925 115036 22937 115039
rect 22520 115008 22937 115036
rect 22520 114996 22526 115008
rect 22925 115005 22937 115008
rect 22971 115005 22983 115039
rect 22925 114999 22983 115005
rect 23014 114996 23020 115048
rect 23072 115036 23078 115048
rect 24320 115045 24348 115076
rect 24394 115064 24400 115116
rect 24452 115104 24458 115116
rect 27062 115104 27068 115116
rect 24452 115076 27068 115104
rect 24452 115064 24458 115076
rect 27062 115064 27068 115076
rect 27120 115064 27126 115116
rect 27341 115107 27399 115113
rect 27341 115073 27353 115107
rect 27387 115104 27399 115107
rect 31570 115104 31576 115116
rect 27387 115076 31576 115104
rect 27387 115073 27399 115076
rect 27341 115067 27399 115073
rect 31570 115064 31576 115076
rect 31628 115064 31634 115116
rect 23661 115039 23719 115045
rect 23661 115036 23673 115039
rect 23072 115008 23673 115036
rect 23072 114996 23078 115008
rect 23661 115005 23673 115008
rect 23707 115005 23719 115039
rect 23661 114999 23719 115005
rect 24305 115039 24363 115045
rect 24305 115005 24317 115039
rect 24351 115005 24363 115039
rect 24305 114999 24363 115005
rect 25417 115039 25475 115045
rect 25417 115005 25429 115039
rect 25463 115005 25475 115039
rect 26418 115036 26424 115048
rect 26379 115008 26424 115036
rect 25417 114999 25475 115005
rect 1903 114940 2774 114968
rect 4908 114940 7236 114968
rect 1903 114937 1915 114940
rect 1857 114931 1915 114937
rect 2746 114900 2774 114940
rect 7650 114928 7656 114980
rect 7708 114968 7714 114980
rect 13354 114968 13360 114980
rect 7708 114940 13360 114968
rect 7708 114928 7714 114940
rect 13354 114928 13360 114940
rect 13412 114928 13418 114980
rect 22830 114968 22836 114980
rect 16776 114940 22836 114968
rect 5166 114900 5172 114912
rect 2746 114872 5172 114900
rect 5166 114860 5172 114872
rect 5224 114860 5230 114912
rect 5534 114860 5540 114912
rect 5592 114900 5598 114912
rect 10686 114900 10692 114912
rect 5592 114872 10692 114900
rect 5592 114860 5598 114872
rect 10686 114860 10692 114872
rect 10744 114860 10750 114912
rect 16776 114909 16804 114940
rect 22830 114928 22836 114940
rect 22888 114928 22894 114980
rect 25424 114968 25452 114999
rect 26418 114996 26424 115008
rect 26476 114996 26482 115048
rect 28721 115039 28779 115045
rect 28721 115005 28733 115039
rect 28767 115005 28779 115039
rect 28721 114999 28779 115005
rect 28728 114968 28756 114999
rect 28810 114996 28816 115048
rect 28868 115036 28874 115048
rect 29178 115036 29184 115048
rect 28868 115008 29184 115036
rect 28868 114996 28874 115008
rect 29178 114996 29184 115008
rect 29236 114996 29242 115048
rect 29362 115036 29368 115048
rect 29323 115008 29368 115036
rect 29362 114996 29368 115008
rect 29420 114996 29426 115048
rect 31481 115039 31539 115045
rect 31481 115005 31493 115039
rect 31527 115036 31539 115039
rect 31726 115036 31754 115144
rect 32122 115132 32128 115144
rect 32180 115132 32186 115184
rect 33321 115175 33379 115181
rect 33321 115141 33333 115175
rect 33367 115172 33379 115175
rect 34793 115175 34851 115181
rect 33367 115144 34744 115172
rect 33367 115141 33379 115144
rect 33321 115135 33379 115141
rect 34146 115104 34152 115116
rect 32324 115076 34152 115104
rect 31527 115008 31754 115036
rect 31527 115005 31539 115008
rect 31481 114999 31539 115005
rect 31938 114996 31944 115048
rect 31996 115036 32002 115048
rect 32125 115039 32183 115045
rect 32125 115036 32137 115039
rect 31996 115008 32137 115036
rect 31996 114996 32002 115008
rect 32125 115005 32137 115008
rect 32171 115005 32183 115039
rect 32125 114999 32183 115005
rect 30374 114968 30380 114980
rect 23308 114940 25452 114968
rect 25516 114940 28672 114968
rect 28728 114940 30380 114968
rect 16761 114903 16819 114909
rect 16761 114869 16773 114903
rect 16807 114869 16819 114903
rect 16761 114863 16819 114869
rect 17405 114903 17463 114909
rect 17405 114869 17417 114903
rect 17451 114900 17463 114903
rect 21082 114900 21088 114912
rect 17451 114872 21088 114900
rect 17451 114869 17463 114872
rect 17405 114863 17463 114869
rect 21082 114860 21088 114872
rect 21140 114860 21146 114912
rect 21269 114903 21327 114909
rect 21269 114869 21281 114903
rect 21315 114900 21327 114903
rect 23308 114900 23336 114940
rect 23474 114900 23480 114912
rect 21315 114872 23336 114900
rect 23435 114872 23480 114900
rect 21315 114869 21327 114872
rect 21269 114863 21327 114869
rect 23474 114860 23480 114872
rect 23532 114860 23538 114912
rect 23566 114860 23572 114912
rect 23624 114900 23630 114912
rect 24302 114900 24308 114912
rect 23624 114872 24308 114900
rect 23624 114860 23630 114872
rect 24302 114860 24308 114872
rect 24360 114860 24366 114912
rect 24394 114860 24400 114912
rect 24452 114900 24458 114912
rect 25516 114900 25544 114940
rect 24452 114872 25544 114900
rect 24452 114860 24458 114872
rect 26694 114860 26700 114912
rect 26752 114900 26758 114912
rect 28537 114903 28595 114909
rect 28537 114900 28549 114903
rect 26752 114872 28549 114900
rect 26752 114860 26758 114872
rect 28537 114869 28549 114872
rect 28583 114869 28595 114903
rect 28644 114900 28672 114940
rect 30374 114928 30380 114940
rect 30432 114928 30438 114980
rect 30561 114971 30619 114977
rect 30561 114937 30573 114971
rect 30607 114937 30619 114971
rect 30561 114931 30619 114937
rect 30576 114900 30604 114931
rect 28644 114872 30604 114900
rect 28537 114863 28595 114869
rect 30650 114860 30656 114912
rect 30708 114900 30714 114912
rect 31386 114900 31392 114912
rect 30708 114872 31392 114900
rect 30708 114860 30714 114872
rect 31386 114860 31392 114872
rect 31444 114860 31450 114912
rect 31478 114860 31484 114912
rect 31536 114900 31542 114912
rect 32324 114900 32352 115076
rect 34146 115064 34152 115076
rect 34204 115064 34210 115116
rect 34716 115104 34744 115144
rect 34793 115141 34805 115175
rect 34839 115172 34851 115175
rect 35526 115172 35532 115184
rect 34839 115144 35532 115172
rect 34839 115141 34851 115144
rect 34793 115135 34851 115141
rect 35526 115132 35532 115144
rect 35584 115132 35590 115184
rect 39850 115104 39856 115116
rect 34716 115076 39856 115104
rect 39850 115064 39856 115076
rect 39908 115064 39914 115116
rect 32398 114996 32404 115048
rect 32456 115036 32462 115048
rect 33873 115039 33931 115045
rect 33873 115036 33885 115039
rect 32456 115008 33885 115036
rect 32456 114996 32462 115008
rect 33873 115005 33885 115008
rect 33919 115005 33931 115039
rect 33873 114999 33931 115005
rect 34790 114996 34796 115048
rect 34848 115036 34854 115048
rect 35713 115039 35771 115045
rect 35713 115036 35725 115039
rect 34848 115008 35725 115036
rect 34848 114996 34854 115008
rect 35713 115005 35725 115008
rect 35759 115005 35771 115039
rect 35713 114999 35771 115005
rect 36078 114996 36084 115048
rect 36136 115036 36142 115048
rect 36173 115039 36231 115045
rect 36173 115036 36185 115039
rect 36136 115008 36185 115036
rect 36136 114996 36142 115008
rect 36173 115005 36185 115008
rect 36219 115005 36231 115039
rect 36173 114999 36231 115005
rect 36541 115039 36599 115045
rect 36541 115005 36553 115039
rect 36587 115005 36599 115039
rect 36541 114999 36599 115005
rect 33137 114971 33195 114977
rect 33137 114937 33149 114971
rect 33183 114968 33195 114971
rect 34238 114968 34244 114980
rect 33183 114940 34244 114968
rect 33183 114937 33195 114940
rect 33137 114931 33195 114937
rect 34238 114928 34244 114940
rect 34296 114928 34302 114980
rect 34514 114928 34520 114980
rect 34572 114968 34578 114980
rect 34609 114971 34667 114977
rect 34609 114968 34621 114971
rect 34572 114940 34621 114968
rect 34572 114928 34578 114940
rect 34609 114937 34621 114940
rect 34655 114937 34667 114971
rect 34609 114931 34667 114937
rect 35526 114928 35532 114980
rect 35584 114968 35590 114980
rect 36556 114968 36584 114999
rect 37918 114968 37924 114980
rect 35584 114940 36584 114968
rect 37879 114940 37924 114968
rect 35584 114928 35590 114940
rect 37918 114928 37924 114940
rect 37976 114928 37982 114980
rect 31536 114872 32352 114900
rect 31536 114860 31542 114872
rect 35250 114860 35256 114912
rect 35308 114900 35314 114912
rect 35805 114903 35863 114909
rect 35805 114900 35817 114903
rect 35308 114872 35817 114900
rect 35308 114860 35314 114872
rect 35805 114869 35817 114872
rect 35851 114869 35863 114903
rect 35805 114863 35863 114869
rect 37734 114860 37740 114912
rect 37792 114900 37798 114912
rect 38013 114903 38071 114909
rect 38013 114900 38025 114903
rect 37792 114872 38025 114900
rect 37792 114860 37798 114872
rect 38013 114869 38025 114872
rect 38059 114869 38071 114903
rect 38013 114863 38071 114869
rect 1104 114810 38824 114832
rect 1104 114758 19606 114810
rect 19658 114758 19670 114810
rect 19722 114758 19734 114810
rect 19786 114758 19798 114810
rect 19850 114758 38824 114810
rect 1104 114736 38824 114758
rect 3418 114696 3424 114708
rect 3379 114668 3424 114696
rect 3418 114656 3424 114668
rect 3476 114656 3482 114708
rect 6822 114656 6828 114708
rect 6880 114696 6886 114708
rect 8113 114699 8171 114705
rect 8113 114696 8125 114699
rect 6880 114668 8125 114696
rect 6880 114656 6886 114668
rect 8113 114665 8125 114668
rect 8159 114665 8171 114699
rect 8113 114659 8171 114665
rect 8294 114656 8300 114708
rect 8352 114696 8358 114708
rect 12069 114699 12127 114705
rect 12069 114696 12081 114699
rect 8352 114668 12081 114696
rect 8352 114656 8358 114668
rect 12069 114665 12081 114668
rect 12115 114665 12127 114699
rect 13354 114696 13360 114708
rect 13315 114668 13360 114696
rect 12069 114659 12127 114665
rect 13354 114656 13360 114668
rect 13412 114656 13418 114708
rect 14001 114699 14059 114705
rect 14001 114665 14013 114699
rect 14047 114665 14059 114699
rect 15286 114696 15292 114708
rect 15247 114668 15292 114696
rect 14001 114659 14059 114665
rect 1857 114631 1915 114637
rect 1857 114597 1869 114631
rect 1903 114628 1915 114631
rect 7190 114628 7196 114640
rect 1903 114600 7196 114628
rect 1903 114597 1915 114600
rect 1857 114591 1915 114597
rect 7190 114588 7196 114600
rect 7248 114588 7254 114640
rect 14016 114628 14044 114659
rect 15286 114656 15292 114668
rect 15344 114656 15350 114708
rect 15933 114699 15991 114705
rect 15933 114665 15945 114699
rect 15979 114696 15991 114699
rect 17770 114696 17776 114708
rect 15979 114668 17776 114696
rect 15979 114665 15991 114668
rect 15933 114659 15991 114665
rect 17770 114656 17776 114668
rect 17828 114656 17834 114708
rect 17865 114699 17923 114705
rect 17865 114665 17877 114699
rect 17911 114696 17923 114699
rect 21818 114696 21824 114708
rect 17911 114668 21824 114696
rect 17911 114665 17923 114668
rect 17865 114659 17923 114665
rect 21818 114656 21824 114668
rect 21876 114656 21882 114708
rect 22649 114699 22707 114705
rect 22649 114665 22661 114699
rect 22695 114696 22707 114699
rect 23566 114696 23572 114708
rect 22695 114668 23572 114696
rect 22695 114665 22707 114668
rect 22649 114659 22707 114665
rect 23566 114656 23572 114668
rect 23624 114656 23630 114708
rect 24118 114656 24124 114708
rect 24176 114696 24182 114708
rect 24176 114668 24624 114696
rect 24176 114656 24182 114668
rect 7300 114600 8248 114628
rect 2590 114560 2596 114572
rect 2551 114532 2596 114560
rect 2590 114520 2596 114532
rect 2648 114520 2654 114572
rect 3329 114563 3387 114569
rect 3329 114529 3341 114563
rect 3375 114560 3387 114563
rect 3694 114560 3700 114572
rect 3375 114532 3700 114560
rect 3375 114529 3387 114532
rect 3329 114523 3387 114529
rect 3694 114520 3700 114532
rect 3752 114520 3758 114572
rect 5258 114520 5264 114572
rect 5316 114560 5322 114572
rect 5445 114563 5503 114569
rect 5445 114560 5457 114563
rect 5316 114532 5457 114560
rect 5316 114520 5322 114532
rect 5445 114529 5457 114532
rect 5491 114529 5503 114563
rect 5445 114523 5503 114529
rect 6270 114520 6276 114572
rect 6328 114560 6334 114572
rect 7300 114560 7328 114600
rect 6328 114532 7328 114560
rect 6328 114520 6334 114532
rect 7374 114520 7380 114572
rect 7432 114560 7438 114572
rect 7650 114560 7656 114572
rect 7432 114532 7512 114560
rect 7611 114532 7656 114560
rect 7432 114520 7438 114532
rect 2038 114492 2044 114504
rect 1999 114464 2044 114492
rect 2038 114452 2044 114464
rect 2096 114452 2102 114504
rect 2777 114495 2835 114501
rect 2777 114461 2789 114495
rect 2823 114492 2835 114495
rect 2866 114492 2872 114504
rect 2823 114464 2872 114492
rect 2823 114461 2835 114464
rect 2777 114455 2835 114461
rect 2866 114452 2872 114464
rect 2924 114452 2930 114504
rect 4062 114452 4068 114504
rect 4120 114492 4126 114504
rect 4157 114495 4215 114501
rect 4157 114492 4169 114495
rect 4120 114464 4169 114492
rect 4120 114452 4126 114464
rect 4157 114461 4169 114464
rect 4203 114461 4215 114495
rect 4157 114455 4215 114461
rect 4801 114495 4859 114501
rect 4801 114461 4813 114495
rect 4847 114492 4859 114495
rect 4890 114492 4896 114504
rect 4847 114464 4896 114492
rect 4847 114461 4859 114464
rect 4801 114455 4859 114461
rect 4890 114452 4896 114464
rect 4948 114452 4954 114504
rect 7006 114492 7012 114504
rect 6967 114464 7012 114492
rect 7006 114452 7012 114464
rect 7064 114452 7070 114504
rect 7484 114433 7512 114532
rect 7650 114520 7656 114532
rect 7708 114520 7714 114572
rect 7469 114427 7527 114433
rect 7469 114393 7481 114427
rect 7515 114393 7527 114427
rect 8220 114424 8248 114600
rect 8312 114600 14044 114628
rect 19536 114600 24532 114628
rect 8312 114569 8340 114600
rect 8297 114563 8355 114569
rect 8297 114529 8309 114563
rect 8343 114529 8355 114563
rect 8754 114560 8760 114572
rect 8715 114532 8760 114560
rect 8297 114523 8355 114529
rect 8754 114520 8760 114532
rect 8812 114520 8818 114572
rect 8846 114520 8852 114572
rect 8904 114560 8910 114572
rect 9401 114563 9459 114569
rect 9401 114560 9413 114563
rect 8904 114532 9413 114560
rect 8904 114520 8910 114532
rect 9401 114529 9413 114532
rect 9447 114529 9459 114563
rect 9401 114523 9459 114529
rect 9490 114520 9496 114572
rect 9548 114560 9554 114572
rect 10045 114563 10103 114569
rect 10045 114560 10057 114563
rect 9548 114532 10057 114560
rect 9548 114520 9554 114532
rect 10045 114529 10057 114532
rect 10091 114529 10103 114563
rect 10045 114523 10103 114529
rect 10226 114520 10232 114572
rect 10284 114560 10290 114572
rect 10873 114563 10931 114569
rect 10873 114560 10885 114563
rect 10284 114532 10885 114560
rect 10284 114520 10290 114532
rect 10873 114529 10885 114532
rect 10919 114529 10931 114563
rect 10873 114523 10931 114529
rect 11698 114520 11704 114572
rect 11756 114560 11762 114572
rect 12253 114563 12311 114569
rect 12253 114560 12265 114563
rect 11756 114532 12265 114560
rect 11756 114520 11762 114532
rect 12253 114529 12265 114532
rect 12299 114529 12311 114563
rect 12253 114523 12311 114529
rect 12342 114520 12348 114572
rect 12400 114560 12406 114572
rect 12897 114563 12955 114569
rect 12897 114560 12909 114563
rect 12400 114532 12909 114560
rect 12400 114520 12406 114532
rect 12897 114529 12909 114532
rect 12943 114529 12955 114563
rect 12897 114523 12955 114529
rect 13170 114520 13176 114572
rect 13228 114560 13234 114572
rect 13541 114563 13599 114569
rect 13541 114560 13553 114563
rect 13228 114532 13553 114560
rect 13228 114520 13234 114532
rect 13541 114529 13553 114532
rect 13587 114529 13599 114563
rect 13541 114523 13599 114529
rect 13722 114520 13728 114572
rect 13780 114560 13786 114572
rect 14185 114563 14243 114569
rect 14185 114560 14197 114563
rect 13780 114532 14197 114560
rect 13780 114520 13786 114532
rect 14185 114529 14197 114532
rect 14231 114529 14243 114563
rect 14185 114523 14243 114529
rect 14458 114520 14464 114572
rect 14516 114560 14522 114572
rect 14829 114563 14887 114569
rect 14829 114560 14841 114563
rect 14516 114532 14841 114560
rect 14516 114520 14522 114532
rect 14829 114529 14841 114532
rect 14875 114529 14887 114563
rect 14829 114523 14887 114529
rect 15010 114520 15016 114572
rect 15068 114560 15074 114572
rect 15473 114563 15531 114569
rect 15473 114560 15485 114563
rect 15068 114532 15485 114560
rect 15068 114520 15074 114532
rect 15473 114529 15485 114532
rect 15519 114529 15531 114563
rect 15473 114523 15531 114529
rect 15746 114520 15752 114572
rect 15804 114560 15810 114572
rect 16117 114563 16175 114569
rect 16117 114560 16129 114563
rect 15804 114532 16129 114560
rect 15804 114520 15810 114532
rect 16117 114529 16129 114532
rect 16163 114529 16175 114563
rect 16117 114523 16175 114529
rect 17862 114520 17868 114572
rect 17920 114560 17926 114572
rect 18049 114563 18107 114569
rect 18049 114560 18061 114563
rect 17920 114532 18061 114560
rect 17920 114520 17926 114532
rect 18049 114529 18061 114532
rect 18095 114529 18107 114563
rect 18049 114523 18107 114529
rect 19242 114520 19248 114572
rect 19300 114560 19306 114572
rect 19429 114563 19487 114569
rect 19429 114560 19441 114563
rect 19300 114532 19441 114560
rect 19300 114520 19306 114532
rect 19429 114529 19441 114532
rect 19475 114529 19487 114563
rect 19429 114523 19487 114529
rect 19536 114492 19564 114600
rect 19978 114520 19984 114572
rect 20036 114560 20042 114572
rect 20165 114563 20223 114569
rect 20165 114560 20177 114563
rect 20036 114532 20177 114560
rect 20036 114520 20042 114532
rect 20165 114529 20177 114532
rect 20211 114529 20223 114563
rect 20990 114560 20996 114572
rect 20165 114523 20223 114529
rect 20272 114532 20996 114560
rect 19260 114464 19564 114492
rect 8941 114427 8999 114433
rect 8941 114424 8953 114427
rect 8220 114396 8953 114424
rect 7469 114387 7527 114393
rect 8941 114393 8953 114396
rect 8987 114393 8999 114427
rect 10686 114424 10692 114436
rect 10647 114396 10692 114424
rect 8941 114387 8999 114393
rect 10686 114384 10692 114396
rect 10744 114384 10750 114436
rect 19260 114433 19288 114464
rect 19245 114427 19303 114433
rect 19245 114393 19257 114427
rect 19291 114393 19303 114427
rect 19245 114387 19303 114393
rect 19981 114427 20039 114433
rect 19981 114393 19993 114427
rect 20027 114424 20039 114427
rect 20272 114424 20300 114532
rect 20990 114520 20996 114532
rect 21048 114520 21054 114572
rect 21082 114520 21088 114572
rect 21140 114560 21146 114572
rect 22462 114560 22468 114572
rect 21140 114532 22468 114560
rect 21140 114520 21146 114532
rect 22462 114520 22468 114532
rect 22520 114520 22526 114572
rect 22830 114560 22836 114572
rect 22791 114532 22836 114560
rect 22830 114520 22836 114532
rect 22888 114520 22894 114572
rect 22922 114520 22928 114572
rect 22980 114560 22986 114572
rect 23293 114563 23351 114569
rect 23293 114560 23305 114563
rect 22980 114532 23305 114560
rect 22980 114520 22986 114532
rect 23293 114529 23305 114532
rect 23339 114529 23351 114563
rect 24394 114560 24400 114572
rect 23293 114523 23351 114529
rect 24320 114532 24400 114560
rect 24320 114433 24348 114532
rect 24394 114520 24400 114532
rect 24452 114520 24458 114572
rect 24504 114569 24532 114600
rect 24489 114563 24547 114569
rect 24489 114529 24501 114563
rect 24535 114529 24547 114563
rect 24596 114560 24624 114668
rect 25498 114656 25504 114708
rect 25556 114696 25562 114708
rect 25556 114668 25912 114696
rect 25556 114656 25562 114668
rect 24854 114588 24860 114640
rect 24912 114628 24918 114640
rect 24912 114600 25636 114628
rect 24912 114588 24918 114600
rect 25608 114569 25636 114600
rect 24949 114563 25007 114569
rect 24949 114560 24961 114563
rect 24596 114532 24961 114560
rect 24489 114523 24547 114529
rect 24949 114529 24961 114532
rect 24995 114529 25007 114563
rect 24949 114523 25007 114529
rect 25593 114563 25651 114569
rect 25593 114529 25605 114563
rect 25639 114529 25651 114563
rect 25884 114560 25912 114668
rect 26602 114656 26608 114708
rect 26660 114696 26666 114708
rect 27801 114699 27859 114705
rect 27801 114696 27813 114699
rect 26660 114668 27813 114696
rect 26660 114656 26666 114668
rect 27801 114665 27813 114668
rect 27847 114665 27859 114699
rect 28442 114696 28448 114708
rect 28403 114668 28448 114696
rect 27801 114659 27859 114665
rect 28442 114656 28448 114668
rect 28500 114656 28506 114708
rect 28534 114656 28540 114708
rect 28592 114696 28598 114708
rect 29089 114699 29147 114705
rect 29089 114696 29101 114699
rect 28592 114668 29101 114696
rect 28592 114656 28598 114668
rect 29089 114665 29101 114668
rect 29135 114665 29147 114699
rect 29089 114659 29147 114665
rect 29914 114656 29920 114708
rect 29972 114696 29978 114708
rect 30101 114699 30159 114705
rect 30101 114696 30113 114699
rect 29972 114668 30113 114696
rect 29972 114656 29978 114668
rect 30101 114665 30113 114668
rect 30147 114665 30159 114699
rect 30101 114659 30159 114665
rect 30282 114656 30288 114708
rect 30340 114696 30346 114708
rect 30653 114699 30711 114705
rect 30653 114696 30665 114699
rect 30340 114668 30665 114696
rect 30340 114656 30346 114668
rect 30653 114665 30665 114668
rect 30699 114665 30711 114699
rect 30653 114659 30711 114665
rect 31297 114699 31355 114705
rect 31297 114665 31309 114699
rect 31343 114665 31355 114699
rect 31297 114659 31355 114665
rect 31312 114628 31340 114659
rect 31662 114656 31668 114708
rect 31720 114696 31726 114708
rect 31941 114699 31999 114705
rect 31941 114696 31953 114699
rect 31720 114668 31953 114696
rect 31720 114656 31726 114668
rect 31941 114665 31953 114668
rect 31987 114665 31999 114699
rect 35894 114696 35900 114708
rect 31941 114659 31999 114665
rect 34624 114668 35900 114696
rect 33686 114628 33692 114640
rect 28000 114600 29224 114628
rect 28000 114569 28028 114600
rect 26237 114563 26295 114569
rect 26237 114560 26249 114563
rect 25884 114532 26249 114560
rect 25593 114523 25651 114529
rect 26237 114529 26249 114532
rect 26283 114529 26295 114563
rect 26237 114523 26295 114529
rect 27985 114563 28043 114569
rect 27985 114529 27997 114563
rect 28031 114529 28043 114563
rect 27985 114523 28043 114529
rect 28629 114563 28687 114569
rect 28629 114529 28641 114563
rect 28675 114560 28687 114563
rect 28675 114532 29132 114560
rect 28675 114529 28687 114532
rect 28629 114523 28687 114529
rect 20027 114396 20300 114424
rect 24305 114427 24363 114433
rect 20027 114393 20039 114396
rect 19981 114387 20039 114393
rect 24305 114393 24317 114427
rect 24351 114393 24363 114427
rect 29104 114424 29132 114532
rect 29196 114492 29224 114600
rect 29288 114600 31248 114628
rect 31312 114600 33692 114628
rect 29288 114569 29316 114600
rect 29273 114563 29331 114569
rect 29273 114529 29285 114563
rect 29319 114529 29331 114563
rect 30006 114560 30012 114572
rect 29967 114532 30012 114560
rect 29273 114523 29331 114529
rect 30006 114520 30012 114532
rect 30064 114520 30070 114572
rect 30098 114520 30104 114572
rect 30156 114560 30162 114572
rect 30837 114563 30895 114569
rect 30837 114560 30849 114563
rect 30156 114532 30849 114560
rect 30156 114520 30162 114532
rect 30837 114529 30849 114532
rect 30883 114529 30895 114563
rect 31220 114560 31248 114600
rect 33686 114588 33692 114600
rect 33744 114588 33750 114640
rect 31478 114560 31484 114572
rect 31220 114532 31340 114560
rect 31439 114532 31484 114560
rect 30837 114523 30895 114529
rect 30650 114492 30656 114504
rect 29196 114464 30656 114492
rect 30650 114452 30656 114464
rect 30708 114452 30714 114504
rect 30742 114424 30748 114436
rect 29104 114396 30748 114424
rect 24305 114387 24363 114393
rect 30742 114384 30748 114396
rect 30800 114384 30806 114436
rect 31312 114424 31340 114532
rect 31478 114520 31484 114532
rect 31536 114520 31542 114572
rect 32125 114563 32183 114569
rect 32125 114529 32137 114563
rect 32171 114560 32183 114563
rect 32674 114560 32680 114572
rect 32171 114532 32680 114560
rect 32171 114529 32183 114532
rect 32125 114523 32183 114529
rect 32674 114520 32680 114532
rect 32732 114520 32738 114572
rect 33042 114520 33048 114572
rect 33100 114560 33106 114572
rect 33229 114563 33287 114569
rect 33229 114560 33241 114563
rect 33100 114532 33241 114560
rect 33100 114520 33106 114532
rect 33229 114529 33241 114532
rect 33275 114529 33287 114563
rect 33229 114523 33287 114529
rect 33318 114520 33324 114572
rect 33376 114560 33382 114572
rect 33965 114563 34023 114569
rect 33965 114560 33977 114563
rect 33376 114532 33977 114560
rect 33376 114520 33382 114532
rect 33965 114529 33977 114532
rect 34011 114529 34023 114563
rect 33965 114523 34023 114529
rect 33413 114495 33471 114501
rect 33413 114461 33425 114495
rect 33459 114492 33471 114495
rect 34624 114492 34652 114668
rect 35894 114656 35900 114668
rect 35952 114656 35958 114708
rect 36262 114696 36268 114708
rect 36223 114668 36268 114696
rect 36262 114656 36268 114668
rect 36320 114656 36326 114708
rect 35544 114600 37044 114628
rect 35544 114572 35572 114600
rect 34790 114560 34796 114572
rect 34751 114532 34796 114560
rect 34790 114520 34796 114532
rect 34848 114520 34854 114572
rect 35437 114563 35495 114569
rect 34900 114532 35296 114560
rect 33459 114464 34652 114492
rect 33459 114461 33471 114464
rect 33413 114455 33471 114461
rect 32122 114424 32128 114436
rect 31312 114396 32128 114424
rect 32122 114384 32128 114396
rect 32180 114384 32186 114436
rect 34146 114384 34152 114436
rect 34204 114424 34210 114436
rect 34900 114424 34928 114532
rect 35268 114492 35296 114532
rect 35437 114529 35449 114563
rect 35483 114560 35495 114563
rect 35526 114560 35532 114572
rect 35483 114532 35532 114560
rect 35483 114529 35495 114532
rect 35437 114523 35495 114529
rect 35526 114520 35532 114532
rect 35584 114520 35590 114572
rect 35710 114560 35716 114572
rect 35671 114532 35716 114560
rect 35710 114520 35716 114532
rect 35768 114520 35774 114572
rect 36170 114560 36176 114572
rect 36131 114532 36176 114560
rect 36170 114520 36176 114532
rect 36228 114520 36234 114572
rect 37016 114569 37044 114600
rect 37001 114563 37059 114569
rect 37001 114529 37013 114563
rect 37047 114529 37059 114563
rect 37001 114523 37059 114529
rect 35345 114495 35403 114501
rect 35345 114492 35357 114495
rect 35268 114464 35357 114492
rect 35345 114461 35357 114464
rect 35391 114492 35403 114495
rect 36909 114495 36967 114501
rect 36909 114492 36921 114495
rect 35391 114464 36921 114492
rect 35391 114461 35403 114464
rect 35345 114455 35403 114461
rect 36909 114461 36921 114464
rect 36955 114461 36967 114495
rect 36909 114455 36967 114461
rect 34204 114396 34928 114424
rect 34204 114384 34210 114396
rect 36078 114384 36084 114436
rect 36136 114424 36142 114436
rect 36262 114424 36268 114436
rect 36136 114396 36268 114424
rect 36136 114384 36142 114396
rect 36262 114384 36268 114396
rect 36320 114384 36326 114436
rect 12710 114356 12716 114368
rect 12671 114328 12716 114356
rect 12710 114316 12716 114328
rect 12768 114316 12774 114368
rect 14642 114356 14648 114368
rect 14603 114328 14648 114356
rect 14642 114316 14648 114328
rect 14700 114316 14706 114368
rect 34057 114359 34115 114365
rect 34057 114325 34069 114359
rect 34103 114356 34115 114359
rect 34422 114356 34428 114368
rect 34103 114328 34428 114356
rect 34103 114325 34115 114328
rect 34057 114319 34115 114325
rect 34422 114316 34428 114328
rect 34480 114316 34486 114368
rect 1104 114266 38824 114288
rect 1104 114214 4246 114266
rect 4298 114214 4310 114266
rect 4362 114214 4374 114266
rect 4426 114214 4438 114266
rect 4490 114214 34966 114266
rect 35018 114214 35030 114266
rect 35082 114214 35094 114266
rect 35146 114214 35158 114266
rect 35210 114214 38824 114266
rect 1104 114192 38824 114214
rect 3053 114155 3111 114161
rect 3053 114121 3065 114155
rect 3099 114152 3111 114155
rect 3142 114152 3148 114164
rect 3099 114124 3148 114152
rect 3099 114121 3111 114124
rect 3053 114115 3111 114121
rect 3142 114112 3148 114124
rect 3200 114112 3206 114164
rect 4433 114155 4491 114161
rect 4433 114121 4445 114155
rect 4479 114152 4491 114155
rect 4614 114152 4620 114164
rect 4479 114124 4620 114152
rect 4479 114121 4491 114124
rect 4433 114115 4491 114121
rect 4614 114112 4620 114124
rect 4672 114112 4678 114164
rect 4985 114155 5043 114161
rect 4985 114121 4997 114155
rect 5031 114152 5043 114155
rect 5442 114152 5448 114164
rect 5031 114124 5448 114152
rect 5031 114121 5043 114124
rect 4985 114115 5043 114121
rect 5442 114112 5448 114124
rect 5500 114112 5506 114164
rect 5813 114155 5871 114161
rect 5813 114121 5825 114155
rect 5859 114152 5871 114155
rect 6454 114152 6460 114164
rect 5859 114124 6460 114152
rect 5859 114121 5871 114124
rect 5813 114115 5871 114121
rect 6454 114112 6460 114124
rect 6512 114112 6518 114164
rect 7558 114112 7564 114164
rect 7616 114152 7622 114164
rect 8205 114155 8263 114161
rect 8205 114152 8217 114155
rect 7616 114124 8217 114152
rect 7616 114112 7622 114124
rect 8205 114121 8217 114124
rect 8251 114121 8263 114155
rect 8205 114115 8263 114121
rect 30374 114112 30380 114164
rect 30432 114152 30438 114164
rect 30469 114155 30527 114161
rect 30469 114152 30481 114155
rect 30432 114124 30481 114152
rect 30432 114112 30438 114124
rect 30469 114121 30481 114124
rect 30515 114121 30527 114155
rect 30469 114115 30527 114121
rect 31849 114155 31907 114161
rect 31849 114121 31861 114155
rect 31895 114152 31907 114155
rect 32030 114152 32036 114164
rect 31895 114124 32036 114152
rect 31895 114121 31907 114124
rect 31849 114115 31907 114121
rect 32030 114112 32036 114124
rect 32088 114112 32094 114164
rect 32858 114112 32864 114164
rect 32916 114152 32922 114164
rect 33137 114155 33195 114161
rect 33137 114152 33149 114155
rect 32916 114124 33149 114152
rect 32916 114112 32922 114124
rect 33137 114121 33149 114124
rect 33183 114121 33195 114155
rect 33137 114115 33195 114121
rect 33502 114112 33508 114164
rect 33560 114152 33566 114164
rect 33873 114155 33931 114161
rect 33873 114152 33885 114155
rect 33560 114124 33885 114152
rect 33560 114112 33566 114124
rect 33873 114121 33885 114124
rect 33919 114121 33931 114155
rect 33873 114115 33931 114121
rect 35526 114112 35532 114164
rect 35584 114152 35590 114164
rect 35584 114124 36124 114152
rect 35584 114112 35590 114124
rect 3878 114044 3884 114096
rect 3936 114084 3942 114096
rect 6917 114087 6975 114093
rect 6917 114084 6929 114087
rect 3936 114056 6929 114084
rect 3936 114044 3942 114056
rect 6917 114053 6929 114056
rect 6963 114053 6975 114087
rect 6917 114047 6975 114053
rect 29362 114044 29368 114096
rect 29420 114084 29426 114096
rect 31113 114087 31171 114093
rect 31113 114084 31125 114087
rect 29420 114056 31125 114084
rect 29420 114044 29426 114056
rect 31113 114053 31125 114056
rect 31159 114053 31171 114087
rect 31113 114047 31171 114053
rect 31202 114044 31208 114096
rect 31260 114084 31266 114096
rect 32493 114087 32551 114093
rect 32493 114084 32505 114087
rect 31260 114056 32505 114084
rect 31260 114044 31266 114056
rect 32493 114053 32505 114056
rect 32539 114053 32551 114087
rect 32493 114047 32551 114053
rect 34422 114044 34428 114096
rect 34480 114084 34486 114096
rect 34793 114087 34851 114093
rect 34480 114056 34744 114084
rect 34480 114044 34486 114056
rect 12710 114016 12716 114028
rect 7760 113988 12716 114016
rect 5169 113951 5227 113957
rect 5169 113917 5181 113951
rect 5215 113948 5227 113951
rect 5534 113948 5540 113960
rect 5215 113920 5540 113948
rect 5215 113917 5227 113920
rect 5169 113911 5227 113917
rect 5534 113908 5540 113920
rect 5592 113908 5598 113960
rect 6457 113951 6515 113957
rect 6457 113917 6469 113951
rect 6503 113948 6515 113951
rect 6914 113948 6920 113960
rect 6503 113920 6920 113948
rect 6503 113917 6515 113920
rect 6457 113911 6515 113917
rect 6914 113908 6920 113920
rect 6972 113908 6978 113960
rect 7760 113957 7788 113988
rect 12710 113976 12716 113988
rect 12768 113976 12774 114028
rect 33870 114016 33876 114028
rect 32048 113988 33876 114016
rect 7101 113951 7159 113957
rect 7101 113917 7113 113951
rect 7147 113917 7159 113951
rect 7101 113911 7159 113917
rect 7745 113951 7803 113957
rect 7745 113917 7757 113951
rect 7791 113917 7803 113951
rect 7745 113911 7803 113917
rect 8389 113951 8447 113957
rect 8389 113917 8401 113951
rect 8435 113948 8447 113951
rect 14642 113948 14648 113960
rect 8435 113920 14648 113948
rect 8435 113917 8447 113920
rect 8389 113911 8447 113917
rect 1854 113880 1860 113892
rect 1815 113852 1860 113880
rect 1854 113840 1860 113852
rect 1912 113840 1918 113892
rect 2041 113883 2099 113889
rect 2041 113849 2053 113883
rect 2087 113880 2099 113883
rect 2682 113880 2688 113892
rect 2087 113852 2688 113880
rect 2087 113849 2099 113852
rect 2041 113843 2099 113849
rect 2682 113840 2688 113852
rect 2740 113840 2746 113892
rect 4798 113840 4804 113892
rect 4856 113880 4862 113892
rect 7116 113880 7144 113911
rect 14642 113908 14648 113920
rect 14700 113908 14706 113960
rect 22002 113948 22008 113960
rect 21963 113920 22008 113948
rect 22002 113908 22008 113920
rect 22060 113908 22066 113960
rect 23382 113948 23388 113960
rect 23343 113920 23388 113948
rect 23382 113908 23388 113920
rect 23440 113908 23446 113960
rect 26234 113948 26240 113960
rect 26195 113920 26240 113948
rect 26234 113908 26240 113920
rect 26292 113908 26298 113960
rect 26878 113948 26884 113960
rect 26839 113920 26884 113948
rect 26878 113908 26884 113920
rect 26936 113908 26942 113960
rect 27614 113948 27620 113960
rect 27575 113920 27620 113948
rect 27614 113908 27620 113920
rect 27672 113908 27678 113960
rect 30558 113908 30564 113960
rect 30616 113948 30622 113960
rect 30653 113951 30711 113957
rect 30653 113948 30665 113951
rect 30616 113920 30665 113948
rect 30616 113908 30622 113920
rect 30653 113917 30665 113920
rect 30699 113917 30711 113951
rect 30653 113911 30711 113917
rect 31297 113951 31355 113957
rect 31297 113917 31309 113951
rect 31343 113948 31355 113951
rect 31386 113948 31392 113960
rect 31343 113920 31392 113948
rect 31343 113917 31355 113920
rect 31297 113911 31355 113917
rect 31386 113908 31392 113920
rect 31444 113908 31450 113960
rect 32048 113957 32076 113988
rect 33870 113976 33876 113988
rect 33928 113976 33934 114028
rect 34606 113976 34612 114028
rect 34664 113976 34670 114028
rect 32033 113951 32091 113957
rect 32033 113917 32045 113951
rect 32079 113917 32091 113951
rect 32033 113911 32091 113917
rect 32490 113908 32496 113960
rect 32548 113948 32554 113960
rect 32677 113951 32735 113957
rect 32677 113948 32689 113951
rect 32548 113920 32689 113948
rect 32548 113908 32554 113920
rect 32677 113917 32689 113920
rect 32723 113917 32735 113951
rect 32677 113911 32735 113917
rect 32950 113908 32956 113960
rect 33008 113948 33014 113960
rect 33321 113951 33379 113957
rect 33321 113948 33333 113951
rect 33008 113920 33333 113948
rect 33008 113908 33014 113920
rect 33321 113917 33333 113920
rect 33367 113917 33379 113951
rect 33321 113911 33379 113917
rect 34057 113951 34115 113957
rect 34057 113917 34069 113951
rect 34103 113948 34115 113951
rect 34624 113948 34652 113976
rect 34103 113920 34652 113948
rect 34103 113917 34115 113920
rect 34057 113911 34115 113917
rect 8294 113880 8300 113892
rect 4856 113852 6408 113880
rect 7116 113852 8300 113880
rect 4856 113840 4862 113852
rect 5994 113772 6000 113824
rect 6052 113812 6058 113824
rect 6273 113815 6331 113821
rect 6273 113812 6285 113815
rect 6052 113784 6285 113812
rect 6052 113772 6058 113784
rect 6273 113781 6285 113784
rect 6319 113781 6331 113815
rect 6380 113812 6408 113852
rect 8294 113840 8300 113852
rect 8352 113840 8358 113892
rect 25774 113840 25780 113892
rect 25832 113880 25838 113892
rect 31754 113880 31760 113892
rect 25832 113852 31760 113880
rect 25832 113840 25838 113852
rect 31754 113840 31760 113852
rect 31812 113840 31818 113892
rect 34606 113880 34612 113892
rect 34567 113852 34612 113880
rect 34606 113840 34612 113852
rect 34664 113840 34670 113892
rect 34716 113880 34744 114056
rect 34793 114053 34805 114087
rect 34839 114084 34851 114087
rect 35250 114084 35256 114096
rect 34839 114056 35256 114084
rect 34839 114053 34851 114056
rect 34793 114047 34851 114053
rect 35250 114044 35256 114056
rect 35308 114044 35314 114096
rect 36096 114016 36124 114124
rect 36096 113988 36584 114016
rect 35989 113951 36047 113957
rect 35989 113917 36001 113951
rect 36035 113948 36047 113951
rect 36078 113948 36084 113960
rect 36035 113920 36084 113948
rect 36035 113917 36047 113920
rect 35989 113911 36047 113917
rect 36078 113908 36084 113920
rect 36136 113908 36142 113960
rect 36262 113948 36268 113960
rect 36223 113920 36268 113948
rect 36262 113908 36268 113920
rect 36320 113908 36326 113960
rect 36556 113957 36584 113988
rect 36541 113951 36599 113957
rect 36541 113917 36553 113951
rect 36587 113917 36599 113951
rect 39390 113948 39396 113960
rect 36541 113911 36599 113917
rect 36648 113920 39396 113948
rect 36648 113880 36676 113920
rect 39390 113908 39396 113920
rect 39448 113908 39454 113960
rect 37918 113880 37924 113892
rect 34716 113852 36676 113880
rect 37879 113852 37924 113880
rect 37918 113840 37924 113852
rect 37976 113840 37982 113892
rect 7561 113815 7619 113821
rect 7561 113812 7573 113815
rect 6380 113784 7573 113812
rect 6273 113775 6331 113781
rect 7561 113781 7573 113784
rect 7607 113781 7619 113815
rect 7561 113775 7619 113781
rect 33962 113772 33968 113824
rect 34020 113812 34026 113824
rect 35805 113815 35863 113821
rect 35805 113812 35817 113815
rect 34020 113784 35817 113812
rect 34020 113772 34026 113784
rect 35805 113781 35817 113784
rect 35851 113781 35863 113815
rect 35805 113775 35863 113781
rect 37366 113772 37372 113824
rect 37424 113812 37430 113824
rect 38013 113815 38071 113821
rect 38013 113812 38025 113815
rect 37424 113784 38025 113812
rect 37424 113772 37430 113784
rect 38013 113781 38025 113784
rect 38059 113781 38071 113815
rect 38013 113775 38071 113781
rect 1104 113722 38824 113744
rect 1104 113670 19606 113722
rect 19658 113670 19670 113722
rect 19722 113670 19734 113722
rect 19786 113670 19798 113722
rect 19850 113670 38824 113722
rect 1104 113648 38824 113670
rect 30837 113611 30895 113617
rect 30837 113577 30849 113611
rect 30883 113608 30895 113611
rect 30926 113608 30932 113620
rect 30883 113580 30932 113608
rect 30883 113577 30895 113580
rect 30837 113571 30895 113577
rect 30926 113568 30932 113580
rect 30984 113568 30990 113620
rect 31726 113580 32536 113608
rect 6730 113500 6736 113552
rect 6788 113540 6794 113552
rect 6788 113512 7512 113540
rect 6788 113500 6794 113512
rect 2130 113472 2136 113484
rect 2091 113444 2136 113472
rect 2130 113432 2136 113444
rect 2188 113432 2194 113484
rect 2774 113432 2780 113484
rect 2832 113472 2838 113484
rect 2832 113444 2877 113472
rect 2832 113432 2838 113444
rect 3326 113432 3332 113484
rect 3384 113472 3390 113484
rect 3421 113475 3479 113481
rect 3421 113472 3433 113475
rect 3384 113444 3433 113472
rect 3384 113432 3390 113444
rect 3421 113441 3433 113444
rect 3467 113441 3479 113475
rect 3421 113435 3479 113441
rect 3970 113432 3976 113484
rect 4028 113472 4034 113484
rect 4249 113475 4307 113481
rect 4249 113472 4261 113475
rect 4028 113444 4261 113472
rect 4028 113432 4034 113444
rect 4249 113441 4261 113444
rect 4295 113441 4307 113475
rect 4249 113435 4307 113441
rect 4706 113432 4712 113484
rect 4764 113472 4770 113484
rect 4893 113475 4951 113481
rect 4893 113472 4905 113475
rect 4764 113444 4905 113472
rect 4764 113432 4770 113444
rect 4893 113441 4905 113444
rect 4939 113441 4951 113475
rect 4893 113435 4951 113441
rect 5350 113432 5356 113484
rect 5408 113472 5414 113484
rect 5537 113475 5595 113481
rect 5537 113472 5549 113475
rect 5408 113444 5549 113472
rect 5408 113432 5414 113444
rect 5537 113441 5549 113444
rect 5583 113441 5595 113475
rect 5537 113435 5595 113441
rect 6086 113432 6092 113484
rect 6144 113472 6150 113484
rect 7484 113481 7512 113512
rect 8202 113500 8208 113552
rect 8260 113540 8266 113552
rect 8260 113512 9076 113540
rect 8260 113500 8266 113512
rect 6825 113475 6883 113481
rect 6825 113472 6837 113475
rect 6144 113444 6837 113472
rect 6144 113432 6150 113444
rect 6825 113441 6837 113444
rect 6871 113441 6883 113475
rect 6825 113435 6883 113441
rect 7469 113475 7527 113481
rect 7469 113441 7481 113475
rect 7515 113441 7527 113475
rect 7469 113435 7527 113441
rect 7558 113432 7564 113484
rect 7616 113472 7622 113484
rect 9048 113481 9076 113512
rect 25038 113500 25044 113552
rect 25096 113540 25102 113552
rect 31726 113540 31754 113580
rect 25096 113512 31754 113540
rect 25096 113500 25102 113512
rect 8389 113475 8447 113481
rect 8389 113472 8401 113475
rect 7616 113444 8401 113472
rect 7616 113432 7622 113444
rect 8389 113441 8401 113444
rect 8435 113441 8447 113475
rect 8389 113435 8447 113441
rect 9033 113475 9091 113481
rect 9033 113441 9045 113475
rect 9079 113441 9091 113475
rect 9033 113435 9091 113441
rect 30834 113432 30840 113484
rect 30892 113472 30898 113484
rect 31021 113475 31079 113481
rect 31021 113472 31033 113475
rect 30892 113444 31033 113472
rect 30892 113432 30898 113444
rect 31021 113441 31033 113444
rect 31067 113441 31079 113475
rect 31021 113435 31079 113441
rect 31110 113432 31116 113484
rect 31168 113472 31174 113484
rect 31665 113475 31723 113481
rect 31665 113472 31677 113475
rect 31168 113444 31677 113472
rect 31168 113432 31174 113444
rect 31665 113441 31677 113444
rect 31711 113441 31723 113475
rect 31665 113435 31723 113441
rect 29178 113296 29184 113348
rect 29236 113336 29242 113348
rect 31481 113339 31539 113345
rect 31481 113336 31493 113339
rect 29236 113308 31493 113336
rect 29236 113296 29242 113308
rect 31481 113305 31493 113308
rect 31527 113305 31539 113339
rect 32508 113336 32536 113580
rect 32582 113568 32588 113620
rect 32640 113608 32646 113620
rect 33137 113611 33195 113617
rect 33137 113608 33149 113611
rect 32640 113580 33149 113608
rect 32640 113568 32646 113580
rect 33137 113577 33149 113580
rect 33183 113577 33195 113611
rect 33137 113571 33195 113577
rect 34146 113568 34152 113620
rect 34204 113608 34210 113620
rect 34241 113611 34299 113617
rect 34241 113608 34253 113611
rect 34204 113580 34253 113608
rect 34204 113568 34210 113580
rect 34241 113577 34253 113580
rect 34287 113577 34299 113611
rect 34241 113571 34299 113577
rect 34609 113611 34667 113617
rect 34609 113577 34621 113611
rect 34655 113608 34667 113611
rect 35802 113608 35808 113620
rect 34655 113580 35808 113608
rect 34655 113577 34667 113580
rect 34609 113571 34667 113577
rect 33134 113432 33140 113484
rect 33192 113472 33198 113484
rect 33321 113475 33379 113481
rect 33321 113472 33333 113475
rect 33192 113444 33333 113472
rect 33192 113432 33198 113444
rect 33321 113441 33333 113444
rect 33367 113441 33379 113475
rect 33321 113435 33379 113441
rect 33965 113407 34023 113413
rect 33965 113373 33977 113407
rect 34011 113404 34023 113407
rect 34146 113404 34152 113416
rect 34011 113376 34152 113404
rect 34011 113373 34023 113376
rect 33965 113367 34023 113373
rect 34146 113364 34152 113376
rect 34204 113364 34210 113416
rect 34256 113404 34284 113571
rect 35802 113568 35808 113580
rect 35860 113568 35866 113620
rect 37182 113608 37188 113620
rect 35912 113580 37188 113608
rect 34450 113543 34508 113549
rect 34450 113509 34462 113543
rect 34496 113540 34508 113543
rect 34882 113540 34888 113552
rect 34496 113512 34888 113540
rect 34496 113509 34508 113512
rect 34450 113503 34508 113509
rect 34882 113500 34888 113512
rect 34940 113540 34946 113552
rect 35250 113540 35256 113552
rect 34940 113512 35256 113540
rect 34940 113500 34946 113512
rect 35250 113500 35256 113512
rect 35308 113500 35314 113552
rect 35912 113549 35940 113580
rect 37182 113568 37188 113580
rect 37240 113568 37246 113620
rect 35897 113543 35955 113549
rect 35897 113509 35909 113543
rect 35943 113509 35955 113543
rect 35897 113503 35955 113509
rect 36633 113543 36691 113549
rect 36633 113509 36645 113543
rect 36679 113540 36691 113543
rect 36906 113540 36912 113552
rect 36679 113512 36912 113540
rect 36679 113509 36691 113512
rect 36633 113503 36691 113509
rect 36906 113500 36912 113512
rect 36964 113500 36970 113552
rect 34333 113475 34391 113481
rect 34333 113441 34345 113475
rect 34379 113472 34391 113475
rect 34790 113472 34796 113484
rect 34379 113444 34796 113472
rect 34379 113441 34391 113444
rect 34333 113435 34391 113441
rect 34790 113432 34796 113444
rect 34848 113432 34854 113484
rect 35710 113472 35716 113484
rect 35671 113444 35716 113472
rect 35710 113432 35716 113444
rect 35768 113432 35774 113484
rect 36449 113475 36507 113481
rect 36449 113441 36461 113475
rect 36495 113472 36507 113475
rect 36538 113472 36544 113484
rect 36495 113444 36544 113472
rect 36495 113441 36507 113444
rect 36449 113435 36507 113441
rect 36538 113432 36544 113444
rect 36596 113432 36602 113484
rect 37182 113472 37188 113484
rect 37143 113444 37188 113472
rect 37182 113432 37188 113444
rect 37240 113432 37246 113484
rect 34422 113404 34428 113416
rect 34256 113376 34428 113404
rect 34422 113364 34428 113376
rect 34480 113364 34486 113416
rect 35526 113364 35532 113416
rect 35584 113404 35590 113416
rect 35802 113404 35808 113416
rect 35584 113376 35808 113404
rect 35584 113364 35590 113376
rect 35802 113364 35808 113376
rect 35860 113364 35866 113416
rect 36998 113336 37004 113348
rect 32508 113308 37004 113336
rect 31481 113299 31539 113305
rect 36998 113296 37004 113308
rect 37056 113296 37062 113348
rect 37274 113268 37280 113280
rect 37235 113240 37280 113268
rect 37274 113228 37280 113240
rect 37332 113228 37338 113280
rect 1104 113178 38824 113200
rect 1104 113126 4246 113178
rect 4298 113126 4310 113178
rect 4362 113126 4374 113178
rect 4426 113126 4438 113178
rect 4490 113126 34966 113178
rect 35018 113126 35030 113178
rect 35082 113126 35094 113178
rect 35146 113126 35158 113178
rect 35210 113126 38824 113178
rect 1104 113104 38824 113126
rect 1946 113064 1952 113076
rect 1907 113036 1952 113064
rect 1946 113024 1952 113036
rect 2004 113024 2010 113076
rect 30650 113024 30656 113076
rect 30708 113064 30714 113076
rect 31297 113067 31355 113073
rect 31297 113064 31309 113067
rect 30708 113036 31309 113064
rect 30708 113024 30714 113036
rect 31297 113033 31309 113036
rect 31343 113033 31355 113067
rect 31297 113027 31355 113033
rect 32122 113024 32128 113076
rect 32180 113064 32186 113076
rect 32585 113067 32643 113073
rect 32585 113064 32597 113067
rect 32180 113036 32597 113064
rect 32180 113024 32186 113036
rect 32585 113033 32597 113036
rect 32631 113033 32643 113067
rect 32585 113027 32643 113033
rect 33226 113024 33232 113076
rect 33284 113064 33290 113076
rect 33413 113067 33471 113073
rect 33413 113064 33425 113067
rect 33284 113036 33425 113064
rect 33284 113024 33290 113036
rect 33413 113033 33425 113036
rect 33459 113033 33471 113067
rect 34698 113064 34704 113076
rect 34659 113036 34704 113064
rect 33413 113027 33471 113033
rect 34698 113024 34704 113036
rect 34756 113024 34762 113076
rect 35161 113067 35219 113073
rect 35161 113033 35173 113067
rect 35207 113064 35219 113067
rect 36262 113064 36268 113076
rect 35207 113036 36268 113064
rect 35207 113033 35219 113036
rect 35161 113027 35219 113033
rect 36262 113024 36268 113036
rect 36320 113024 36326 113076
rect 36541 113067 36599 113073
rect 36541 113033 36553 113067
rect 36587 113064 36599 113067
rect 39114 113064 39120 113076
rect 36587 113036 39120 113064
rect 36587 113033 36599 113036
rect 36541 113027 36599 113033
rect 39114 113024 39120 113036
rect 39172 113024 39178 113076
rect 28905 112999 28963 113005
rect 28905 112965 28917 112999
rect 28951 112996 28963 112999
rect 29270 112996 29276 113008
rect 28951 112968 29276 112996
rect 28951 112965 28963 112968
rect 28905 112959 28963 112965
rect 29270 112956 29276 112968
rect 29328 112956 29334 113008
rect 30742 112956 30748 113008
rect 30800 112996 30806 113008
rect 31941 112999 31999 113005
rect 31941 112996 31953 112999
rect 30800 112968 31953 112996
rect 30800 112956 30806 112968
rect 31941 112965 31953 112968
rect 31987 112965 31999 112999
rect 31941 112959 31999 112965
rect 37369 112999 37427 113005
rect 37369 112965 37381 112999
rect 37415 112996 37427 112999
rect 38930 112996 38936 113008
rect 37415 112968 38936 112996
rect 37415 112965 37427 112968
rect 37369 112959 37427 112965
rect 38930 112956 38936 112968
rect 38988 112956 38994 113008
rect 34542 112931 34600 112937
rect 34542 112897 34554 112931
rect 34588 112928 34600 112931
rect 35250 112928 35256 112940
rect 34588 112900 35256 112928
rect 34588 112897 34600 112900
rect 34542 112891 34600 112897
rect 35250 112888 35256 112900
rect 35308 112888 35314 112940
rect 38470 112928 38476 112940
rect 35728 112900 38476 112928
rect 28813 112863 28871 112869
rect 28813 112829 28825 112863
rect 28859 112829 28871 112863
rect 28813 112823 28871 112829
rect 29089 112863 29147 112869
rect 29089 112829 29101 112863
rect 29135 112860 29147 112863
rect 30374 112860 30380 112872
rect 29135 112832 30380 112860
rect 29135 112829 29147 112832
rect 29089 112823 29147 112829
rect 1857 112795 1915 112801
rect 1857 112761 1869 112795
rect 1903 112792 1915 112795
rect 2222 112792 2228 112804
rect 1903 112764 2228 112792
rect 1903 112761 1915 112764
rect 1857 112755 1915 112761
rect 2222 112752 2228 112764
rect 2280 112752 2286 112804
rect 28828 112792 28856 112823
rect 30374 112820 30380 112832
rect 30432 112820 30438 112872
rect 31294 112820 31300 112872
rect 31352 112860 31358 112872
rect 31481 112863 31539 112869
rect 31481 112860 31493 112863
rect 31352 112832 31493 112860
rect 31352 112820 31358 112832
rect 31481 112829 31493 112832
rect 31527 112829 31539 112863
rect 31481 112823 31539 112829
rect 32125 112863 32183 112869
rect 32125 112829 32137 112863
rect 32171 112860 32183 112863
rect 32214 112860 32220 112872
rect 32171 112832 32220 112860
rect 32171 112829 32183 112832
rect 32125 112823 32183 112829
rect 32214 112820 32220 112832
rect 32272 112820 32278 112872
rect 32306 112820 32312 112872
rect 32364 112860 32370 112872
rect 32769 112863 32827 112869
rect 32769 112860 32781 112863
rect 32364 112832 32781 112860
rect 32364 112820 32370 112832
rect 32769 112829 32781 112832
rect 32815 112829 32827 112863
rect 32769 112823 32827 112829
rect 33410 112820 33416 112872
rect 33468 112860 33474 112872
rect 33597 112863 33655 112869
rect 33597 112860 33609 112863
rect 33468 112832 33609 112860
rect 33468 112820 33474 112832
rect 33597 112829 33609 112832
rect 33643 112829 33655 112863
rect 33597 112823 33655 112829
rect 34057 112863 34115 112869
rect 34057 112829 34069 112863
rect 34103 112860 34115 112863
rect 34146 112860 34152 112872
rect 34103 112832 34152 112860
rect 34103 112829 34115 112832
rect 34057 112823 34115 112829
rect 34146 112820 34152 112832
rect 34204 112820 34210 112872
rect 34330 112820 34336 112872
rect 34388 112820 34394 112872
rect 34425 112863 34483 112869
rect 34425 112829 34437 112863
rect 34471 112860 34483 112863
rect 34790 112860 34796 112872
rect 34471 112832 34796 112860
rect 34471 112829 34483 112832
rect 34425 112823 34483 112829
rect 34790 112820 34796 112832
rect 34848 112860 34854 112872
rect 35618 112860 35624 112872
rect 34848 112832 35624 112860
rect 34848 112820 34854 112832
rect 35618 112820 35624 112832
rect 35676 112820 35682 112872
rect 35728 112869 35756 112900
rect 38470 112888 38476 112900
rect 38528 112888 38534 112940
rect 35713 112863 35771 112869
rect 35713 112829 35725 112863
rect 35759 112829 35771 112863
rect 37918 112860 37924 112872
rect 37879 112832 37924 112860
rect 35713 112823 35771 112829
rect 37918 112820 37924 112832
rect 37976 112820 37982 112872
rect 34348 112792 34376 112820
rect 35161 112795 35219 112801
rect 35161 112792 35173 112795
rect 28828 112764 34376 112792
rect 34624 112764 35173 112792
rect 28994 112684 29000 112736
rect 29052 112724 29058 112736
rect 29273 112727 29331 112733
rect 29273 112724 29285 112727
rect 29052 112696 29285 112724
rect 29052 112684 29058 112696
rect 29273 112693 29285 112696
rect 29319 112693 29331 112727
rect 29273 112687 29331 112693
rect 31846 112684 31852 112736
rect 31904 112724 31910 112736
rect 32766 112724 32772 112736
rect 31904 112696 32772 112724
rect 31904 112684 31910 112696
rect 32766 112684 32772 112696
rect 32824 112684 32830 112736
rect 34330 112724 34336 112736
rect 34291 112696 34336 112724
rect 34330 112684 34336 112696
rect 34388 112724 34394 112736
rect 34624 112724 34652 112764
rect 35161 112761 35173 112764
rect 35207 112761 35219 112795
rect 35161 112755 35219 112761
rect 36262 112752 36268 112804
rect 36320 112792 36326 112804
rect 36449 112795 36507 112801
rect 36449 112792 36461 112795
rect 36320 112764 36461 112792
rect 36320 112752 36326 112764
rect 36449 112761 36461 112764
rect 36495 112761 36507 112795
rect 37182 112792 37188 112804
rect 37143 112764 37188 112792
rect 36449 112755 36507 112761
rect 37182 112752 37188 112764
rect 37240 112752 37246 112804
rect 34388 112696 34652 112724
rect 34388 112684 34394 112696
rect 34698 112684 34704 112736
rect 34756 112724 34762 112736
rect 35897 112727 35955 112733
rect 35897 112724 35909 112727
rect 34756 112696 35909 112724
rect 34756 112684 34762 112696
rect 35897 112693 35909 112696
rect 35943 112693 35955 112727
rect 35897 112687 35955 112693
rect 37642 112684 37648 112736
rect 37700 112724 37706 112736
rect 38013 112727 38071 112733
rect 38013 112724 38025 112727
rect 37700 112696 38025 112724
rect 37700 112684 37706 112696
rect 38013 112693 38025 112696
rect 38059 112693 38071 112727
rect 38013 112687 38071 112693
rect 1104 112634 38824 112656
rect 1104 112582 19606 112634
rect 19658 112582 19670 112634
rect 19722 112582 19734 112634
rect 19786 112582 19798 112634
rect 19850 112582 38824 112634
rect 1104 112560 38824 112582
rect 33778 112480 33784 112532
rect 33836 112520 33842 112532
rect 34057 112523 34115 112529
rect 34057 112520 34069 112523
rect 33836 112492 34069 112520
rect 33836 112480 33842 112492
rect 34057 112489 34069 112492
rect 34103 112489 34115 112523
rect 34057 112483 34115 112489
rect 35526 112480 35532 112532
rect 35584 112520 35590 112532
rect 36541 112523 36599 112529
rect 36541 112520 36553 112523
rect 35584 112492 36553 112520
rect 35584 112480 35590 112492
rect 36541 112489 36553 112492
rect 36587 112489 36599 112523
rect 36541 112483 36599 112489
rect 29454 112412 29460 112464
rect 29512 112452 29518 112464
rect 37182 112452 37188 112464
rect 29512 112424 37188 112452
rect 29512 112412 29518 112424
rect 37182 112412 37188 112424
rect 37240 112412 37246 112464
rect 1857 112387 1915 112393
rect 1857 112353 1869 112387
rect 1903 112384 1915 112387
rect 6270 112384 6276 112396
rect 1903 112356 6276 112384
rect 1903 112353 1915 112356
rect 1857 112347 1915 112353
rect 6270 112344 6276 112356
rect 6328 112344 6334 112396
rect 34054 112344 34060 112396
rect 34112 112384 34118 112396
rect 34241 112387 34299 112393
rect 34241 112384 34253 112387
rect 34112 112356 34253 112384
rect 34112 112344 34118 112356
rect 34241 112353 34253 112356
rect 34287 112353 34299 112387
rect 34241 112347 34299 112353
rect 35342 112344 35348 112396
rect 35400 112384 35406 112396
rect 35713 112387 35771 112393
rect 35713 112384 35725 112387
rect 35400 112356 35725 112384
rect 35400 112344 35406 112356
rect 35713 112353 35725 112356
rect 35759 112353 35771 112387
rect 35713 112347 35771 112353
rect 36078 112344 36084 112396
rect 36136 112384 36142 112396
rect 36449 112387 36507 112393
rect 36449 112384 36461 112387
rect 36136 112356 36461 112384
rect 36136 112344 36142 112356
rect 36449 112353 36461 112356
rect 36495 112353 36507 112387
rect 37090 112384 37096 112396
rect 37051 112356 37096 112384
rect 36449 112347 36507 112353
rect 37090 112344 37096 112356
rect 37148 112344 37154 112396
rect 2038 112316 2044 112328
rect 1999 112288 2044 112316
rect 2038 112276 2044 112288
rect 2096 112276 2102 112328
rect 35342 112208 35348 112260
rect 35400 112248 35406 112260
rect 37277 112251 37335 112257
rect 37277 112248 37289 112251
rect 35400 112220 37289 112248
rect 35400 112208 35406 112220
rect 37277 112217 37289 112220
rect 37323 112217 37335 112251
rect 37277 112211 37335 112217
rect 35894 112180 35900 112192
rect 35855 112152 35900 112180
rect 35894 112140 35900 112152
rect 35952 112140 35958 112192
rect 1104 112090 38824 112112
rect 1104 112038 4246 112090
rect 4298 112038 4310 112090
rect 4362 112038 4374 112090
rect 4426 112038 4438 112090
rect 4490 112038 34966 112090
rect 35018 112038 35030 112090
rect 35082 112038 35094 112090
rect 35146 112038 35158 112090
rect 35210 112038 38824 112090
rect 1104 112016 38824 112038
rect 34790 111800 34796 111852
rect 34848 111840 34854 111852
rect 35713 111843 35771 111849
rect 35713 111840 35725 111843
rect 34848 111812 35725 111840
rect 34848 111800 34854 111812
rect 35713 111809 35725 111812
rect 35759 111809 35771 111843
rect 35713 111803 35771 111809
rect 35618 111732 35624 111784
rect 35676 111772 35682 111784
rect 36081 111775 36139 111781
rect 36081 111772 36093 111775
rect 35676 111744 36093 111772
rect 35676 111732 35682 111744
rect 36081 111741 36093 111744
rect 36127 111741 36139 111775
rect 37090 111772 37096 111784
rect 37051 111744 37096 111772
rect 36081 111735 36139 111741
rect 37090 111732 37096 111744
rect 37148 111732 37154 111784
rect 37826 111772 37832 111784
rect 37787 111744 37832 111772
rect 37826 111732 37832 111744
rect 37884 111732 37890 111784
rect 35526 111664 35532 111716
rect 35584 111704 35590 111716
rect 36170 111704 36176 111716
rect 36228 111713 36234 111716
rect 36228 111707 36256 111713
rect 35584 111676 36176 111704
rect 35584 111664 35590 111676
rect 36170 111664 36176 111676
rect 36244 111673 36256 111707
rect 38470 111704 38476 111716
rect 36228 111667 36256 111673
rect 37292 111676 38476 111704
rect 36228 111664 36234 111667
rect 33778 111596 33784 111648
rect 33836 111636 33842 111648
rect 34330 111636 34336 111648
rect 33836 111608 34336 111636
rect 33836 111596 33842 111608
rect 34330 111596 34336 111608
rect 34388 111636 34394 111648
rect 35989 111639 36047 111645
rect 35989 111636 36001 111639
rect 34388 111608 36001 111636
rect 34388 111596 34394 111608
rect 35989 111605 36001 111608
rect 36035 111605 36047 111639
rect 36354 111636 36360 111648
rect 36315 111608 36360 111636
rect 35989 111599 36047 111605
rect 36354 111596 36360 111608
rect 36412 111596 36418 111648
rect 37292 111645 37320 111676
rect 38470 111664 38476 111676
rect 38528 111664 38534 111716
rect 37277 111639 37335 111645
rect 37277 111605 37289 111639
rect 37323 111605 37335 111639
rect 37277 111599 37335 111605
rect 38013 111639 38071 111645
rect 38013 111605 38025 111639
rect 38059 111636 38071 111639
rect 39114 111636 39120 111648
rect 38059 111608 39120 111636
rect 38059 111605 38071 111608
rect 38013 111599 38071 111605
rect 39114 111596 39120 111608
rect 39172 111596 39178 111648
rect 1104 111546 38824 111568
rect 1104 111494 19606 111546
rect 19658 111494 19670 111546
rect 19722 111494 19734 111546
rect 19786 111494 19798 111546
rect 19850 111494 38824 111546
rect 1104 111472 38824 111494
rect 1946 111432 1952 111444
rect 1907 111404 1952 111432
rect 1946 111392 1952 111404
rect 2004 111392 2010 111444
rect 35986 111432 35992 111444
rect 35947 111404 35992 111432
rect 35986 111392 35992 111404
rect 36044 111392 36050 111444
rect 35618 111324 35624 111376
rect 35676 111364 35682 111376
rect 35713 111367 35771 111373
rect 35713 111364 35725 111367
rect 35676 111336 35725 111364
rect 35676 111324 35682 111336
rect 35713 111333 35725 111336
rect 35759 111333 35771 111367
rect 35713 111327 35771 111333
rect 1857 111299 1915 111305
rect 1857 111265 1869 111299
rect 1903 111296 1915 111299
rect 2498 111296 2504 111308
rect 1903 111268 2504 111296
rect 1903 111265 1915 111268
rect 1857 111259 1915 111265
rect 2498 111256 2504 111268
rect 2556 111256 2562 111308
rect 34054 111256 34060 111308
rect 34112 111296 34118 111308
rect 34422 111296 34428 111308
rect 34112 111268 34428 111296
rect 34112 111256 34118 111268
rect 34422 111256 34428 111268
rect 34480 111296 34486 111308
rect 34480 111268 35480 111296
rect 34480 111256 34486 111268
rect 33502 111188 33508 111240
rect 33560 111228 33566 111240
rect 34146 111228 34152 111240
rect 33560 111200 34152 111228
rect 33560 111188 33566 111200
rect 34146 111188 34152 111200
rect 34204 111228 34210 111240
rect 35345 111231 35403 111237
rect 35345 111228 35357 111231
rect 34204 111200 35357 111228
rect 34204 111188 34210 111200
rect 35345 111197 35357 111200
rect 35391 111197 35403 111231
rect 35452 111228 35480 111268
rect 35526 111256 35532 111308
rect 35584 111296 35590 111308
rect 35830 111299 35888 111305
rect 35830 111296 35842 111299
rect 35584 111268 35842 111296
rect 35584 111256 35590 111268
rect 35830 111265 35842 111268
rect 35876 111265 35888 111299
rect 37090 111296 37096 111308
rect 37051 111268 37096 111296
rect 35830 111259 35888 111265
rect 37090 111256 37096 111268
rect 37148 111256 37154 111308
rect 35621 111231 35679 111237
rect 35621 111228 35633 111231
rect 35452 111200 35633 111228
rect 35345 111191 35403 111197
rect 35621 111197 35633 111200
rect 35667 111197 35679 111231
rect 35621 111191 35679 111197
rect 34422 111052 34428 111104
rect 34480 111092 34486 111104
rect 37277 111095 37335 111101
rect 37277 111092 37289 111095
rect 34480 111064 37289 111092
rect 34480 111052 34486 111064
rect 37277 111061 37289 111064
rect 37323 111061 37335 111095
rect 37277 111055 37335 111061
rect 1104 111002 38824 111024
rect 1104 110950 4246 111002
rect 4298 110950 4310 111002
rect 4362 110950 4374 111002
rect 4426 110950 4438 111002
rect 4490 110950 34966 111002
rect 35018 110950 35030 111002
rect 35082 110950 35094 111002
rect 35146 110950 35158 111002
rect 35210 110950 38824 111002
rect 1104 110928 38824 110950
rect 1857 110687 1915 110693
rect 1857 110653 1869 110687
rect 1903 110684 1915 110687
rect 2130 110684 2136 110696
rect 1903 110656 2136 110684
rect 1903 110653 1915 110656
rect 1857 110647 1915 110653
rect 2130 110644 2136 110656
rect 2188 110644 2194 110696
rect 13722 110644 13728 110696
rect 13780 110684 13786 110696
rect 26605 110687 26663 110693
rect 26605 110684 26617 110687
rect 13780 110656 26617 110684
rect 13780 110644 13786 110656
rect 26605 110653 26617 110656
rect 26651 110653 26663 110687
rect 37826 110684 37832 110696
rect 37787 110656 37832 110684
rect 26605 110647 26663 110653
rect 37826 110644 37832 110656
rect 37884 110644 37890 110696
rect 2038 110616 2044 110628
rect 1999 110588 2044 110616
rect 2038 110576 2044 110588
rect 2096 110576 2102 110628
rect 36078 110616 36084 110628
rect 31726 110588 36084 110616
rect 26789 110551 26847 110557
rect 26789 110517 26801 110551
rect 26835 110548 26847 110551
rect 31726 110548 31754 110588
rect 36078 110576 36084 110588
rect 36136 110576 36142 110628
rect 26835 110520 31754 110548
rect 26835 110517 26847 110520
rect 26789 110511 26847 110517
rect 32582 110508 32588 110560
rect 32640 110548 32646 110560
rect 38013 110551 38071 110557
rect 38013 110548 38025 110551
rect 32640 110520 38025 110548
rect 32640 110508 32646 110520
rect 38013 110517 38025 110520
rect 38059 110517 38071 110551
rect 38013 110511 38071 110517
rect 1104 110458 38824 110480
rect 1104 110406 19606 110458
rect 19658 110406 19670 110458
rect 19722 110406 19734 110458
rect 19786 110406 19798 110458
rect 19850 110406 38824 110458
rect 1104 110384 38824 110406
rect 37090 110208 37096 110220
rect 37051 110180 37096 110208
rect 37090 110168 37096 110180
rect 37148 110168 37154 110220
rect 33226 110032 33232 110084
rect 33284 110072 33290 110084
rect 34698 110072 34704 110084
rect 33284 110044 34704 110072
rect 33284 110032 33290 110044
rect 34698 110032 34704 110044
rect 34756 110032 34762 110084
rect 31938 109964 31944 110016
rect 31996 110004 32002 110016
rect 35802 110004 35808 110016
rect 31996 109976 35808 110004
rect 31996 109964 32002 109976
rect 35802 109964 35808 109976
rect 35860 109964 35866 110016
rect 37277 110007 37335 110013
rect 37277 109973 37289 110007
rect 37323 110004 37335 110007
rect 38654 110004 38660 110016
rect 37323 109976 38660 110004
rect 37323 109973 37335 109976
rect 37277 109967 37335 109973
rect 38654 109964 38660 109976
rect 38712 109964 38718 110016
rect 1104 109914 38824 109936
rect 1104 109862 4246 109914
rect 4298 109862 4310 109914
rect 4362 109862 4374 109914
rect 4426 109862 4438 109914
rect 4490 109862 34966 109914
rect 35018 109862 35030 109914
rect 35082 109862 35094 109914
rect 35146 109862 35158 109914
rect 35210 109862 38824 109914
rect 1104 109840 38824 109862
rect 1946 109800 1952 109812
rect 1907 109772 1952 109800
rect 1946 109760 1952 109772
rect 2004 109760 2010 109812
rect 34609 109803 34667 109809
rect 33060 109772 33364 109800
rect 2682 109556 2688 109608
rect 2740 109596 2746 109608
rect 32674 109596 32680 109608
rect 2740 109568 22094 109596
rect 32635 109568 32680 109596
rect 2740 109556 2746 109568
rect 1857 109531 1915 109537
rect 1857 109497 1869 109531
rect 1903 109528 1915 109531
rect 1946 109528 1952 109540
rect 1903 109500 1952 109528
rect 1903 109497 1915 109500
rect 1857 109491 1915 109497
rect 1946 109488 1952 109500
rect 2004 109488 2010 109540
rect 22066 109528 22094 109568
rect 32674 109556 32680 109568
rect 32732 109556 32738 109608
rect 32953 109599 33011 109605
rect 32953 109565 32965 109599
rect 32999 109596 33011 109599
rect 33060 109596 33088 109772
rect 33336 109664 33364 109772
rect 34609 109769 34621 109803
rect 34655 109800 34667 109803
rect 35434 109800 35440 109812
rect 34655 109772 35440 109800
rect 34655 109769 34667 109772
rect 34609 109763 34667 109769
rect 35434 109760 35440 109772
rect 35492 109760 35498 109812
rect 35802 109760 35808 109812
rect 35860 109800 35866 109812
rect 37277 109803 37335 109809
rect 37277 109800 37289 109803
rect 35860 109772 37289 109800
rect 35860 109760 35866 109772
rect 37277 109769 37289 109772
rect 37323 109769 37335 109803
rect 37277 109763 37335 109769
rect 35894 109664 35900 109676
rect 33336 109636 35900 109664
rect 35894 109624 35900 109636
rect 35952 109624 35958 109676
rect 33226 109596 33232 109608
rect 32999 109568 33088 109596
rect 33187 109568 33232 109596
rect 32999 109565 33011 109568
rect 32953 109559 33011 109565
rect 33226 109556 33232 109568
rect 33284 109556 33290 109608
rect 33321 109599 33379 109605
rect 33321 109565 33333 109599
rect 33367 109565 33379 109599
rect 33321 109559 33379 109565
rect 33965 109599 34023 109605
rect 33965 109565 33977 109599
rect 34011 109596 34023 109599
rect 34790 109596 34796 109608
rect 34011 109568 34796 109596
rect 34011 109565 34023 109568
rect 33965 109559 34023 109565
rect 33336 109528 33364 109559
rect 34790 109556 34796 109568
rect 34848 109556 34854 109608
rect 37090 109596 37096 109608
rect 37051 109568 37096 109596
rect 37090 109556 37096 109568
rect 37148 109556 37154 109608
rect 37826 109596 37832 109608
rect 37787 109568 37832 109596
rect 37826 109556 37832 109568
rect 37884 109556 37890 109608
rect 22066 109500 33364 109528
rect 34146 109488 34152 109540
rect 34204 109528 34210 109540
rect 34450 109531 34508 109537
rect 34450 109528 34462 109531
rect 34204 109500 34462 109528
rect 34204 109488 34210 109500
rect 34450 109497 34462 109500
rect 34496 109497 34508 109531
rect 34450 109491 34508 109497
rect 33134 109420 33140 109472
rect 33192 109460 33198 109472
rect 33229 109463 33287 109469
rect 33229 109460 33241 109463
rect 33192 109432 33241 109460
rect 33192 109420 33198 109432
rect 33229 109429 33241 109432
rect 33275 109429 33287 109463
rect 33229 109423 33287 109429
rect 34054 109420 34060 109472
rect 34112 109460 34118 109472
rect 34241 109463 34299 109469
rect 34241 109460 34253 109463
rect 34112 109432 34253 109460
rect 34112 109420 34118 109432
rect 34241 109429 34253 109432
rect 34287 109429 34299 109463
rect 34241 109423 34299 109429
rect 34330 109420 34336 109472
rect 34388 109460 34394 109472
rect 38013 109463 38071 109469
rect 34388 109432 34433 109460
rect 34388 109420 34394 109432
rect 38013 109429 38025 109463
rect 38059 109460 38071 109463
rect 38838 109460 38844 109472
rect 38059 109432 38844 109460
rect 38059 109429 38071 109432
rect 38013 109423 38071 109429
rect 38838 109420 38844 109432
rect 38896 109420 38902 109472
rect 1104 109370 38824 109392
rect 1104 109318 19606 109370
rect 19658 109318 19670 109370
rect 19722 109318 19734 109370
rect 19786 109318 19798 109370
rect 19850 109318 38824 109370
rect 1104 109296 38824 109318
rect 34425 109259 34483 109265
rect 34425 109225 34437 109259
rect 34471 109256 34483 109259
rect 34514 109256 34520 109268
rect 34471 109228 34520 109256
rect 34471 109225 34483 109228
rect 34425 109219 34483 109225
rect 34514 109216 34520 109228
rect 34572 109216 34578 109268
rect 36906 109216 36912 109268
rect 36964 109256 36970 109268
rect 37277 109259 37335 109265
rect 37277 109256 37289 109259
rect 36964 109228 37289 109256
rect 36964 109216 36970 109228
rect 37277 109225 37289 109228
rect 37323 109225 37335 109259
rect 37277 109219 37335 109225
rect 33410 109148 33416 109200
rect 33468 109188 33474 109200
rect 34149 109191 34207 109197
rect 34149 109188 34161 109191
rect 33468 109160 34161 109188
rect 33468 109148 33474 109160
rect 34149 109157 34161 109160
rect 34195 109188 34207 109191
rect 34330 109188 34336 109200
rect 34195 109160 34336 109188
rect 34195 109157 34207 109160
rect 34149 109151 34207 109157
rect 34330 109148 34336 109160
rect 34388 109148 34394 109200
rect 1854 109120 1860 109132
rect 1815 109092 1860 109120
rect 1854 109080 1860 109092
rect 1912 109080 1918 109132
rect 33226 109080 33232 109132
rect 33284 109120 33290 109132
rect 34057 109123 34115 109129
rect 34057 109120 34069 109123
rect 33284 109092 34069 109120
rect 33284 109080 33290 109092
rect 34057 109089 34069 109092
rect 34103 109089 34115 109123
rect 34790 109120 34796 109132
rect 34057 109083 34115 109089
rect 34164 109092 34796 109120
rect 2133 109055 2191 109061
rect 2133 109021 2145 109055
rect 2179 109052 2191 109055
rect 27154 109052 27160 109064
rect 2179 109024 27160 109052
rect 2179 109021 2191 109024
rect 2133 109015 2191 109021
rect 27154 109012 27160 109024
rect 27212 109012 27218 109064
rect 30558 109012 30564 109064
rect 30616 109052 30622 109064
rect 33781 109055 33839 109061
rect 33781 109052 33793 109055
rect 30616 109024 33793 109052
rect 30616 109012 30622 109024
rect 33781 109021 33793 109024
rect 33827 109052 33839 109055
rect 34164 109052 34192 109092
rect 34790 109080 34796 109092
rect 34848 109080 34854 109132
rect 37090 109120 37096 109132
rect 37051 109092 37096 109120
rect 37090 109080 37096 109092
rect 37148 109080 37154 109132
rect 33827 109024 34192 109052
rect 34266 109055 34324 109061
rect 33827 109021 33839 109024
rect 33781 109015 33839 109021
rect 34266 109021 34278 109055
rect 34312 109052 34324 109055
rect 34882 109052 34888 109064
rect 34312 109024 34888 109052
rect 34312 109021 34324 109024
rect 34266 109015 34324 109021
rect 34882 109012 34888 109024
rect 34940 109012 34946 109064
rect 1104 108826 38824 108848
rect 1104 108774 4246 108826
rect 4298 108774 4310 108826
rect 4362 108774 4374 108826
rect 4426 108774 4438 108826
rect 4490 108774 34966 108826
rect 35018 108774 35030 108826
rect 35082 108774 35094 108826
rect 35146 108774 35158 108826
rect 35210 108774 38824 108826
rect 1104 108752 38824 108774
rect 8478 108672 8484 108724
rect 8536 108712 8542 108724
rect 13081 108715 13139 108721
rect 13081 108712 13093 108715
rect 8536 108684 13093 108712
rect 8536 108672 8542 108684
rect 13081 108681 13093 108684
rect 13127 108681 13139 108715
rect 13081 108675 13139 108681
rect 28721 108715 28779 108721
rect 28721 108681 28733 108715
rect 28767 108712 28779 108715
rect 36538 108712 36544 108724
rect 28767 108684 36544 108712
rect 28767 108681 28779 108684
rect 28721 108675 28779 108681
rect 36538 108672 36544 108684
rect 36596 108672 36602 108724
rect 32858 108604 32864 108656
rect 32916 108644 32922 108656
rect 38013 108647 38071 108653
rect 38013 108644 38025 108647
rect 32916 108616 38025 108644
rect 32916 108604 32922 108616
rect 38013 108613 38025 108616
rect 38059 108613 38071 108647
rect 38013 108607 38071 108613
rect 33689 108579 33747 108585
rect 33689 108545 33701 108579
rect 33735 108576 33747 108579
rect 35434 108576 35440 108588
rect 33735 108548 35440 108576
rect 33735 108545 33747 108548
rect 33689 108539 33747 108545
rect 35434 108536 35440 108548
rect 35492 108536 35498 108588
rect 12894 108508 12900 108520
rect 12855 108480 12900 108508
rect 12894 108468 12900 108480
rect 12952 108468 12958 108520
rect 17586 108468 17592 108520
rect 17644 108508 17650 108520
rect 28537 108511 28595 108517
rect 28537 108508 28549 108511
rect 17644 108480 28549 108508
rect 17644 108468 17650 108480
rect 28537 108477 28549 108480
rect 28583 108477 28595 108511
rect 28537 108471 28595 108477
rect 33321 108511 33379 108517
rect 33321 108477 33333 108511
rect 33367 108508 33379 108511
rect 33410 108508 33416 108520
rect 33367 108480 33416 108508
rect 33367 108477 33379 108480
rect 33321 108471 33379 108477
rect 33410 108468 33416 108480
rect 33468 108468 33474 108520
rect 34146 108508 34152 108520
rect 34107 108480 34152 108508
rect 34146 108468 34152 108480
rect 34204 108468 34210 108520
rect 37826 108508 37832 108520
rect 37787 108480 37832 108508
rect 37826 108468 37832 108480
rect 37884 108468 37890 108520
rect 33137 108443 33195 108449
rect 33137 108409 33149 108443
rect 33183 108440 33195 108443
rect 33502 108440 33508 108452
rect 33183 108412 33508 108440
rect 33183 108409 33195 108412
rect 33137 108403 33195 108409
rect 33502 108400 33508 108412
rect 33560 108400 33566 108452
rect 34333 108375 34391 108381
rect 34333 108341 34345 108375
rect 34379 108372 34391 108375
rect 34514 108372 34520 108384
rect 34379 108344 34520 108372
rect 34379 108341 34391 108344
rect 34333 108335 34391 108341
rect 34514 108332 34520 108344
rect 34572 108372 34578 108384
rect 35526 108372 35532 108384
rect 34572 108344 35532 108372
rect 34572 108332 34578 108344
rect 35526 108332 35532 108344
rect 35584 108332 35590 108384
rect 1104 108282 38824 108304
rect 1104 108230 19606 108282
rect 19658 108230 19670 108282
rect 19722 108230 19734 108282
rect 19786 108230 19798 108282
rect 19850 108230 38824 108282
rect 1104 108208 38824 108230
rect 1946 108168 1952 108180
rect 1907 108140 1952 108168
rect 1946 108128 1952 108140
rect 2004 108128 2010 108180
rect 34238 108060 34244 108112
rect 34296 108100 34302 108112
rect 34422 108100 34428 108112
rect 34296 108072 34428 108100
rect 34296 108060 34302 108072
rect 34422 108060 34428 108072
rect 34480 108060 34486 108112
rect 1857 108035 1915 108041
rect 1857 108001 1869 108035
rect 1903 108032 1915 108035
rect 3510 108032 3516 108044
rect 1903 108004 3516 108032
rect 1903 108001 1915 108004
rect 1857 107995 1915 108001
rect 3510 107992 3516 108004
rect 3568 107992 3574 108044
rect 33226 107992 33232 108044
rect 33284 108032 33290 108044
rect 33321 108035 33379 108041
rect 33321 108032 33333 108035
rect 33284 108004 33333 108032
rect 33284 107992 33290 108004
rect 33321 108001 33333 108004
rect 33367 108001 33379 108035
rect 37182 108032 37188 108044
rect 37143 108004 37188 108032
rect 33321 107995 33379 108001
rect 37182 107992 37188 108004
rect 37240 107992 37246 108044
rect 32490 107856 32496 107908
rect 32548 107896 32554 107908
rect 37369 107899 37427 107905
rect 37369 107896 37381 107899
rect 32548 107868 37381 107896
rect 32548 107856 32554 107868
rect 37369 107865 37381 107868
rect 37415 107865 37427 107899
rect 37369 107859 37427 107865
rect 33505 107831 33563 107837
rect 33505 107797 33517 107831
rect 33551 107828 33563 107831
rect 33778 107828 33784 107840
rect 33551 107800 33784 107828
rect 33551 107797 33563 107800
rect 33505 107791 33563 107797
rect 33778 107788 33784 107800
rect 33836 107828 33842 107840
rect 35250 107828 35256 107840
rect 33836 107800 35256 107828
rect 33836 107788 33842 107800
rect 35250 107788 35256 107800
rect 35308 107788 35314 107840
rect 1104 107738 38824 107760
rect 1104 107686 4246 107738
rect 4298 107686 4310 107738
rect 4362 107686 4374 107738
rect 4426 107686 4438 107738
rect 4490 107686 34966 107738
rect 35018 107686 35030 107738
rect 35082 107686 35094 107738
rect 35146 107686 35158 107738
rect 35210 107686 38824 107738
rect 1104 107664 38824 107686
rect 33137 107559 33195 107565
rect 33137 107525 33149 107559
rect 33183 107556 33195 107559
rect 35434 107556 35440 107568
rect 33183 107528 35440 107556
rect 33183 107525 33195 107528
rect 33137 107519 33195 107525
rect 35434 107516 35440 107528
rect 35492 107516 35498 107568
rect 1857 107423 1915 107429
rect 1857 107389 1869 107423
rect 1903 107420 1915 107423
rect 2406 107420 2412 107432
rect 1903 107392 2412 107420
rect 1903 107389 1915 107392
rect 1857 107383 1915 107389
rect 2406 107380 2412 107392
rect 2464 107380 2470 107432
rect 31110 107380 31116 107432
rect 31168 107420 31174 107432
rect 32953 107423 33011 107429
rect 32953 107420 32965 107423
rect 31168 107392 32965 107420
rect 31168 107380 31174 107392
rect 32953 107389 32965 107392
rect 32999 107420 33011 107423
rect 33410 107420 33416 107432
rect 32999 107392 33416 107420
rect 32999 107389 33011 107392
rect 32953 107383 33011 107389
rect 33410 107380 33416 107392
rect 33468 107380 33474 107432
rect 37182 107420 37188 107432
rect 37143 107392 37188 107420
rect 37182 107380 37188 107392
rect 37240 107380 37246 107432
rect 2038 107352 2044 107364
rect 1999 107324 2044 107352
rect 2038 107312 2044 107324
rect 2096 107312 2102 107364
rect 35618 107312 35624 107364
rect 35676 107352 35682 107364
rect 37918 107352 37924 107364
rect 35676 107324 37412 107352
rect 37879 107324 37924 107352
rect 35676 107312 35682 107324
rect 34330 107244 34336 107296
rect 34388 107284 34394 107296
rect 37277 107287 37335 107293
rect 37277 107284 37289 107287
rect 34388 107256 37289 107284
rect 34388 107244 34394 107256
rect 37277 107253 37289 107256
rect 37323 107253 37335 107287
rect 37384 107284 37412 107324
rect 37918 107312 37924 107324
rect 37976 107312 37982 107364
rect 38013 107287 38071 107293
rect 38013 107284 38025 107287
rect 37384 107256 38025 107284
rect 37277 107247 37335 107253
rect 38013 107253 38025 107256
rect 38059 107253 38071 107287
rect 38013 107247 38071 107253
rect 1104 107194 38824 107216
rect 1104 107142 19606 107194
rect 19658 107142 19670 107194
rect 19722 107142 19734 107194
rect 19786 107142 19798 107194
rect 19850 107142 38824 107194
rect 1104 107120 38824 107142
rect 1857 106947 1915 106953
rect 1857 106913 1869 106947
rect 1903 106944 1915 106947
rect 2866 106944 2872 106956
rect 1903 106916 2872 106944
rect 1903 106913 1915 106916
rect 1857 106907 1915 106913
rect 2866 106904 2872 106916
rect 2924 106904 2930 106956
rect 37182 106944 37188 106956
rect 37143 106916 37188 106944
rect 37182 106904 37188 106916
rect 37240 106904 37246 106956
rect 1946 106740 1952 106752
rect 1907 106712 1952 106740
rect 1946 106700 1952 106712
rect 2004 106700 2010 106752
rect 35526 106700 35532 106752
rect 35584 106740 35590 106752
rect 37277 106743 37335 106749
rect 37277 106740 37289 106743
rect 35584 106712 37289 106740
rect 35584 106700 35590 106712
rect 37277 106709 37289 106712
rect 37323 106709 37335 106743
rect 37277 106703 37335 106709
rect 1104 106650 38824 106672
rect 1104 106598 4246 106650
rect 4298 106598 4310 106650
rect 4362 106598 4374 106650
rect 4426 106598 4438 106650
rect 4490 106598 34966 106650
rect 35018 106598 35030 106650
rect 35082 106598 35094 106650
rect 35146 106598 35158 106650
rect 35210 106598 38824 106650
rect 1104 106576 38824 106598
rect 34054 106360 34060 106412
rect 34112 106400 34118 106412
rect 38105 106403 38163 106409
rect 38105 106400 38117 106403
rect 34112 106372 38117 106400
rect 34112 106360 34118 106372
rect 38105 106369 38117 106372
rect 38151 106369 38163 106403
rect 38105 106363 38163 106369
rect 37918 106332 37924 106344
rect 37879 106304 37924 106332
rect 37918 106292 37924 106304
rect 37976 106292 37982 106344
rect 1104 106106 38824 106128
rect 1104 106054 19606 106106
rect 19658 106054 19670 106106
rect 19722 106054 19734 106106
rect 19786 106054 19798 106106
rect 19850 106054 38824 106106
rect 1104 106032 38824 106054
rect 8662 105952 8668 106004
rect 8720 105992 8726 106004
rect 10137 105995 10195 106001
rect 10137 105992 10149 105995
rect 8720 105964 10149 105992
rect 8720 105952 8726 105964
rect 10137 105961 10149 105964
rect 10183 105961 10195 105995
rect 10137 105955 10195 105961
rect 33134 105924 33140 105936
rect 33095 105896 33140 105924
rect 33134 105884 33140 105896
rect 33192 105884 33198 105936
rect 35250 105924 35256 105936
rect 35211 105896 35256 105924
rect 35250 105884 35256 105896
rect 35308 105884 35314 105936
rect 1394 105856 1400 105868
rect 1355 105828 1400 105856
rect 1394 105816 1400 105828
rect 1452 105816 1458 105868
rect 9950 105856 9956 105868
rect 9911 105828 9956 105856
rect 9950 105816 9956 105828
rect 10008 105816 10014 105868
rect 34514 105816 34520 105868
rect 34572 105856 34578 105868
rect 35069 105859 35127 105865
rect 35069 105856 35081 105859
rect 34572 105828 35081 105856
rect 34572 105816 34578 105828
rect 35069 105825 35081 105828
rect 35115 105825 35127 105859
rect 35069 105819 35127 105825
rect 35161 105859 35219 105865
rect 35161 105825 35173 105859
rect 35207 105856 35219 105859
rect 35434 105856 35440 105868
rect 35207 105828 35440 105856
rect 35207 105825 35219 105828
rect 35161 105819 35219 105825
rect 35434 105816 35440 105828
rect 35492 105816 35498 105868
rect 37182 105856 37188 105868
rect 37143 105828 37188 105856
rect 37182 105816 37188 105828
rect 37240 105816 37246 105868
rect 1578 105788 1584 105800
rect 1539 105760 1584 105788
rect 1578 105748 1584 105760
rect 1636 105748 1642 105800
rect 27062 105748 27068 105800
rect 27120 105788 27126 105800
rect 33502 105788 33508 105800
rect 27120 105760 33508 105788
rect 27120 105748 27126 105760
rect 33502 105748 33508 105760
rect 33560 105788 33566 105800
rect 34609 105791 34667 105797
rect 34609 105788 34621 105791
rect 33560 105760 34621 105788
rect 33560 105748 33566 105760
rect 34609 105757 34621 105760
rect 34655 105757 34667 105791
rect 34609 105751 34667 105757
rect 34698 105748 34704 105800
rect 34756 105788 34762 105800
rect 34756 105760 34801 105788
rect 34756 105748 34762 105760
rect 27614 105612 27620 105664
rect 27672 105652 27678 105664
rect 33229 105655 33287 105661
rect 33229 105652 33241 105655
rect 27672 105624 33241 105652
rect 27672 105612 27678 105624
rect 33229 105621 33241 105624
rect 33275 105621 33287 105655
rect 33229 105615 33287 105621
rect 35434 105612 35440 105664
rect 35492 105652 35498 105664
rect 37277 105655 37335 105661
rect 37277 105652 37289 105655
rect 35492 105624 37289 105652
rect 35492 105612 35498 105624
rect 37277 105621 37289 105624
rect 37323 105621 37335 105655
rect 37277 105615 37335 105621
rect 1104 105562 38824 105584
rect 1104 105510 4246 105562
rect 4298 105510 4310 105562
rect 4362 105510 4374 105562
rect 4426 105510 4438 105562
rect 4490 105510 34966 105562
rect 35018 105510 35030 105562
rect 35082 105510 35094 105562
rect 35146 105510 35158 105562
rect 35210 105510 38824 105562
rect 1104 105488 38824 105510
rect 37918 105244 37924 105256
rect 37879 105216 37924 105244
rect 37918 105204 37924 105216
rect 37976 105204 37982 105256
rect 1857 105179 1915 105185
rect 1857 105145 1869 105179
rect 1903 105176 1915 105179
rect 2314 105176 2320 105188
rect 1903 105148 2320 105176
rect 1903 105145 1915 105148
rect 1857 105139 1915 105145
rect 2314 105136 2320 105148
rect 2372 105136 2378 105188
rect 1946 105108 1952 105120
rect 1907 105080 1952 105108
rect 1946 105068 1952 105080
rect 2004 105068 2010 105120
rect 33962 105068 33968 105120
rect 34020 105108 34026 105120
rect 38013 105111 38071 105117
rect 38013 105108 38025 105111
rect 34020 105080 38025 105108
rect 34020 105068 34026 105080
rect 38013 105077 38025 105080
rect 38059 105077 38071 105111
rect 38013 105071 38071 105077
rect 1104 105018 38824 105040
rect 1104 104966 19606 105018
rect 19658 104966 19670 105018
rect 19722 104966 19734 105018
rect 19786 104966 19798 105018
rect 19850 104966 38824 105018
rect 1104 104944 38824 104966
rect 37182 104836 37188 104848
rect 37143 104808 37188 104836
rect 37182 104796 37188 104808
rect 37240 104796 37246 104848
rect 35986 104524 35992 104576
rect 36044 104564 36050 104576
rect 37277 104567 37335 104573
rect 37277 104564 37289 104567
rect 36044 104536 37289 104564
rect 36044 104524 36050 104536
rect 37277 104533 37289 104536
rect 37323 104533 37335 104567
rect 37277 104527 37335 104533
rect 1104 104474 38824 104496
rect 1104 104422 4246 104474
rect 4298 104422 4310 104474
rect 4362 104422 4374 104474
rect 4426 104422 4438 104474
rect 4490 104422 34966 104474
rect 35018 104422 35030 104474
rect 35082 104422 35094 104474
rect 35146 104422 35158 104474
rect 35210 104422 38824 104474
rect 1104 104400 38824 104422
rect 30653 104363 30711 104369
rect 30653 104329 30665 104363
rect 30699 104360 30711 104363
rect 34790 104360 34796 104372
rect 30699 104332 34796 104360
rect 30699 104329 30711 104332
rect 30653 104323 30711 104329
rect 34790 104320 34796 104332
rect 34848 104320 34854 104372
rect 1486 104156 1492 104168
rect 1447 104128 1492 104156
rect 1486 104116 1492 104128
rect 1544 104116 1550 104168
rect 30469 104159 30527 104165
rect 30469 104125 30481 104159
rect 30515 104156 30527 104159
rect 30650 104156 30656 104168
rect 30515 104128 30656 104156
rect 30515 104125 30527 104128
rect 30469 104119 30527 104125
rect 30650 104116 30656 104128
rect 30708 104116 30714 104168
rect 37182 104156 37188 104168
rect 37143 104128 37188 104156
rect 37182 104116 37188 104128
rect 37240 104116 37246 104168
rect 2041 104091 2099 104097
rect 2041 104057 2053 104091
rect 2087 104088 2099 104091
rect 3602 104088 3608 104100
rect 2087 104060 3608 104088
rect 2087 104057 2099 104060
rect 2041 104051 2099 104057
rect 3602 104048 3608 104060
rect 3660 104048 3666 104100
rect 31202 104048 31208 104100
rect 31260 104088 31266 104100
rect 37918 104088 37924 104100
rect 31260 104060 37412 104088
rect 37879 104060 37924 104088
rect 31260 104048 31266 104060
rect 36170 103980 36176 104032
rect 36228 104020 36234 104032
rect 37277 104023 37335 104029
rect 37277 104020 37289 104023
rect 36228 103992 37289 104020
rect 36228 103980 36234 103992
rect 37277 103989 37289 103992
rect 37323 103989 37335 104023
rect 37384 104020 37412 104060
rect 37918 104048 37924 104060
rect 37976 104048 37982 104100
rect 38013 104023 38071 104029
rect 38013 104020 38025 104023
rect 37384 103992 38025 104020
rect 37277 103983 37335 103989
rect 38013 103989 38025 103992
rect 38059 103989 38071 104023
rect 38013 103983 38071 103989
rect 1104 103930 38824 103952
rect 1104 103878 19606 103930
rect 19658 103878 19670 103930
rect 19722 103878 19734 103930
rect 19786 103878 19798 103930
rect 19850 103878 38824 103930
rect 1104 103856 38824 103878
rect 30929 103819 30987 103825
rect 30929 103785 30941 103819
rect 30975 103816 30987 103819
rect 33226 103816 33232 103828
rect 30975 103788 33232 103816
rect 30975 103785 30987 103788
rect 30929 103779 30987 103785
rect 33226 103776 33232 103788
rect 33284 103776 33290 103828
rect 30377 103751 30435 103757
rect 30377 103717 30389 103751
rect 30423 103748 30435 103751
rect 33870 103748 33876 103760
rect 30423 103720 33876 103748
rect 30423 103717 30435 103720
rect 30377 103711 30435 103717
rect 33870 103708 33876 103720
rect 33928 103708 33934 103760
rect 1670 103640 1676 103692
rect 1728 103680 1734 103692
rect 1857 103683 1915 103689
rect 1857 103680 1869 103683
rect 1728 103652 1869 103680
rect 1728 103640 1734 103652
rect 1857 103649 1869 103652
rect 1903 103649 1915 103683
rect 30006 103680 30012 103692
rect 29919 103652 30012 103680
rect 1857 103643 1915 103649
rect 30006 103640 30012 103652
rect 30064 103680 30070 103692
rect 30837 103683 30895 103689
rect 30837 103680 30849 103683
rect 30064 103652 30849 103680
rect 30064 103640 30070 103652
rect 30837 103649 30849 103652
rect 30883 103649 30895 103683
rect 37182 103680 37188 103692
rect 37143 103652 37188 103680
rect 30837 103643 30895 103649
rect 37182 103640 37188 103652
rect 37240 103640 37246 103692
rect 2038 103544 2044 103556
rect 1999 103516 2044 103544
rect 2038 103504 2044 103516
rect 2096 103504 2102 103556
rect 37369 103547 37427 103553
rect 37369 103513 37381 103547
rect 37415 103544 37427 103547
rect 38194 103544 38200 103556
rect 37415 103516 38200 103544
rect 37415 103513 37427 103516
rect 37369 103507 37427 103513
rect 38194 103504 38200 103516
rect 38252 103504 38258 103556
rect 1104 103386 38824 103408
rect 1104 103334 4246 103386
rect 4298 103334 4310 103386
rect 4362 103334 4374 103386
rect 4426 103334 4438 103386
rect 4490 103334 34966 103386
rect 35018 103334 35030 103386
rect 35082 103334 35094 103386
rect 35146 103334 35158 103386
rect 35210 103334 38824 103386
rect 1104 103312 38824 103334
rect 7098 103272 7104 103284
rect 7059 103244 7104 103272
rect 7098 103232 7104 103244
rect 7156 103232 7162 103284
rect 30561 103275 30619 103281
rect 30561 103241 30573 103275
rect 30607 103272 30619 103275
rect 34146 103272 34152 103284
rect 30607 103244 34152 103272
rect 30607 103241 30619 103244
rect 30561 103235 30619 103241
rect 34146 103232 34152 103244
rect 34204 103232 34210 103284
rect 25685 103139 25743 103145
rect 25685 103105 25697 103139
rect 25731 103136 25743 103139
rect 36814 103136 36820 103148
rect 25731 103108 36820 103136
rect 25731 103105 25743 103108
rect 25685 103099 25743 103105
rect 36814 103096 36820 103108
rect 36872 103096 36878 103148
rect 6917 103071 6975 103077
rect 6917 103037 6929 103071
rect 6963 103068 6975 103071
rect 7006 103068 7012 103080
rect 6963 103040 7012 103068
rect 6963 103037 6975 103040
rect 6917 103031 6975 103037
rect 7006 103028 7012 103040
rect 7064 103028 7070 103080
rect 30469 103071 30527 103077
rect 30469 103037 30481 103071
rect 30515 103068 30527 103071
rect 30650 103068 30656 103080
rect 30515 103040 30656 103068
rect 30515 103037 30527 103040
rect 30469 103031 30527 103037
rect 30650 103028 30656 103040
rect 30708 103028 30714 103080
rect 11422 102960 11428 103012
rect 11480 103000 11486 103012
rect 25501 103003 25559 103009
rect 25501 103000 25513 103003
rect 11480 102972 25513 103000
rect 11480 102960 11486 102972
rect 25501 102969 25513 102972
rect 25547 102969 25559 103003
rect 37918 103000 37924 103012
rect 37879 102972 37924 103000
rect 25501 102963 25559 102969
rect 37918 102960 37924 102972
rect 37976 102960 37982 103012
rect 31570 102892 31576 102944
rect 31628 102932 31634 102944
rect 38013 102935 38071 102941
rect 38013 102932 38025 102935
rect 31628 102904 38025 102932
rect 31628 102892 31634 102904
rect 38013 102901 38025 102904
rect 38059 102901 38071 102935
rect 38013 102895 38071 102901
rect 1104 102842 38824 102864
rect 1104 102790 19606 102842
rect 19658 102790 19670 102842
rect 19722 102790 19734 102842
rect 19786 102790 19798 102842
rect 19850 102790 38824 102842
rect 1104 102768 38824 102790
rect 7742 102728 7748 102740
rect 7703 102700 7748 102728
rect 7742 102688 7748 102700
rect 7800 102688 7806 102740
rect 1486 102552 1492 102604
rect 1544 102592 1550 102604
rect 1857 102595 1915 102601
rect 1857 102592 1869 102595
rect 1544 102564 1869 102592
rect 1544 102552 1550 102564
rect 1857 102561 1869 102564
rect 1903 102561 1915 102595
rect 2038 102592 2044 102604
rect 1999 102564 2044 102592
rect 1857 102555 1915 102561
rect 2038 102552 2044 102564
rect 2096 102552 2102 102604
rect 7558 102592 7564 102604
rect 7519 102564 7564 102592
rect 7558 102552 7564 102564
rect 7616 102552 7622 102604
rect 37182 102592 37188 102604
rect 37143 102564 37188 102592
rect 37182 102552 37188 102564
rect 37240 102552 37246 102604
rect 36998 102348 37004 102400
rect 37056 102388 37062 102400
rect 37277 102391 37335 102397
rect 37277 102388 37289 102391
rect 37056 102360 37289 102388
rect 37056 102348 37062 102360
rect 37277 102357 37289 102360
rect 37323 102357 37335 102391
rect 37277 102351 37335 102357
rect 1104 102298 38824 102320
rect 1104 102246 4246 102298
rect 4298 102246 4310 102298
rect 4362 102246 4374 102298
rect 4426 102246 4438 102298
rect 4490 102246 34966 102298
rect 35018 102246 35030 102298
rect 35082 102246 35094 102298
rect 35146 102246 35158 102298
rect 35210 102246 38824 102298
rect 1104 102224 38824 102246
rect 30650 102144 30656 102196
rect 30708 102184 30714 102196
rect 31294 102184 31300 102196
rect 30708 102156 31300 102184
rect 30708 102144 30714 102156
rect 31294 102144 31300 102156
rect 31352 102144 31358 102196
rect 32766 102144 32772 102196
rect 32824 102184 32830 102196
rect 36722 102184 36728 102196
rect 32824 102156 36728 102184
rect 32824 102144 32830 102156
rect 36722 102144 36728 102156
rect 36780 102144 36786 102196
rect 25774 102076 25780 102128
rect 25832 102116 25838 102128
rect 25869 102119 25927 102125
rect 25869 102116 25881 102119
rect 25832 102088 25881 102116
rect 25832 102076 25838 102088
rect 25869 102085 25881 102088
rect 25915 102085 25927 102119
rect 25869 102079 25927 102085
rect 1394 101980 1400 101992
rect 1355 101952 1400 101980
rect 1394 101940 1400 101952
rect 1452 101940 1458 101992
rect 9493 101983 9551 101989
rect 9493 101949 9505 101983
rect 9539 101980 9551 101983
rect 18598 101980 18604 101992
rect 9539 101952 18604 101980
rect 9539 101949 9551 101952
rect 9493 101943 9551 101949
rect 18598 101940 18604 101952
rect 18656 101940 18662 101992
rect 37182 101980 37188 101992
rect 37143 101952 37188 101980
rect 37182 101940 37188 101952
rect 37240 101940 37246 101992
rect 37369 101983 37427 101989
rect 37369 101949 37381 101983
rect 37415 101980 37427 101983
rect 38746 101980 38752 101992
rect 37415 101952 38752 101980
rect 37415 101949 37427 101952
rect 37369 101943 37427 101949
rect 38746 101940 38752 101952
rect 38804 101940 38810 101992
rect 12342 101872 12348 101924
rect 12400 101912 12406 101924
rect 25685 101915 25743 101921
rect 25685 101912 25697 101915
rect 12400 101884 25697 101912
rect 12400 101872 12406 101884
rect 25685 101881 25697 101884
rect 25731 101881 25743 101915
rect 37918 101912 37924 101924
rect 37879 101884 37924 101912
rect 25685 101875 25743 101881
rect 37918 101872 37924 101884
rect 37976 101872 37982 101924
rect 1854 101804 1860 101856
rect 1912 101844 1918 101856
rect 9677 101847 9735 101853
rect 9677 101844 9689 101847
rect 1912 101816 9689 101844
rect 1912 101804 1918 101816
rect 9677 101813 9689 101816
rect 9723 101813 9735 101847
rect 9677 101807 9735 101813
rect 36722 101804 36728 101856
rect 36780 101844 36786 101856
rect 38013 101847 38071 101853
rect 38013 101844 38025 101847
rect 36780 101816 38025 101844
rect 36780 101804 36786 101816
rect 38013 101813 38025 101816
rect 38059 101813 38071 101847
rect 38013 101807 38071 101813
rect 1104 101754 38824 101776
rect 1104 101702 19606 101754
rect 19658 101702 19670 101754
rect 19722 101702 19734 101754
rect 19786 101702 19798 101754
rect 19850 101702 38824 101754
rect 1104 101680 38824 101702
rect 37182 101504 37188 101516
rect 37143 101476 37188 101504
rect 37182 101464 37188 101476
rect 37240 101464 37246 101516
rect 35802 101396 35808 101448
rect 35860 101436 35866 101448
rect 37734 101436 37740 101448
rect 35860 101408 37740 101436
rect 35860 101396 35866 101408
rect 37734 101396 37740 101408
rect 37792 101396 37798 101448
rect 31386 101260 31392 101312
rect 31444 101300 31450 101312
rect 37277 101303 37335 101309
rect 37277 101300 37289 101303
rect 31444 101272 37289 101300
rect 31444 101260 31450 101272
rect 37277 101269 37289 101272
rect 37323 101269 37335 101303
rect 37277 101263 37335 101269
rect 1104 101210 38824 101232
rect 1104 101158 4246 101210
rect 4298 101158 4310 101210
rect 4362 101158 4374 101210
rect 4426 101158 4438 101210
rect 4490 101158 34966 101210
rect 35018 101158 35030 101210
rect 35082 101158 35094 101210
rect 35146 101158 35158 101210
rect 35210 101158 38824 101210
rect 1104 101136 38824 101158
rect 2222 101056 2228 101108
rect 2280 101096 2286 101108
rect 6549 101099 6607 101105
rect 6549 101096 6561 101099
rect 2280 101068 6561 101096
rect 2280 101056 2286 101068
rect 6549 101065 6561 101068
rect 6595 101065 6607 101099
rect 6549 101059 6607 101065
rect 1394 100892 1400 100904
rect 1355 100864 1400 100892
rect 1394 100852 1400 100864
rect 1452 100852 1458 100904
rect 6365 100895 6423 100901
rect 6365 100861 6377 100895
rect 6411 100892 6423 100895
rect 10502 100892 10508 100904
rect 6411 100864 10508 100892
rect 6411 100861 6423 100864
rect 6365 100855 6423 100861
rect 10502 100852 10508 100864
rect 10560 100852 10566 100904
rect 37918 100824 37924 100836
rect 37879 100796 37924 100824
rect 37918 100784 37924 100796
rect 37976 100784 37982 100836
rect 36262 100716 36268 100768
rect 36320 100756 36326 100768
rect 38013 100759 38071 100765
rect 38013 100756 38025 100759
rect 36320 100728 38025 100756
rect 36320 100716 36326 100728
rect 38013 100725 38025 100728
rect 38059 100725 38071 100759
rect 38013 100719 38071 100725
rect 1104 100666 38824 100688
rect 1104 100614 19606 100666
rect 19658 100614 19670 100666
rect 19722 100614 19734 100666
rect 19786 100614 19798 100666
rect 19850 100614 38824 100666
rect 1104 100592 38824 100614
rect 34146 100444 34152 100496
rect 34204 100484 34210 100496
rect 37642 100484 37648 100496
rect 34204 100456 37648 100484
rect 34204 100444 34210 100456
rect 37642 100444 37648 100456
rect 37700 100444 37706 100496
rect 1394 100416 1400 100428
rect 1355 100388 1400 100416
rect 1394 100376 1400 100388
rect 1452 100376 1458 100428
rect 37182 100416 37188 100428
rect 37143 100388 37188 100416
rect 37182 100376 37188 100388
rect 37240 100376 37246 100428
rect 33042 100172 33048 100224
rect 33100 100212 33106 100224
rect 37277 100215 37335 100221
rect 37277 100212 37289 100215
rect 33100 100184 37289 100212
rect 33100 100172 33106 100184
rect 37277 100181 37289 100184
rect 37323 100181 37335 100215
rect 37277 100175 37335 100181
rect 1104 100122 38824 100144
rect 1104 100070 4246 100122
rect 4298 100070 4310 100122
rect 4362 100070 4374 100122
rect 4426 100070 4438 100122
rect 4490 100070 34966 100122
rect 35018 100070 35030 100122
rect 35082 100070 35094 100122
rect 35146 100070 35158 100122
rect 35210 100070 38824 100122
rect 1104 100048 38824 100070
rect 6270 100008 6276 100020
rect 6231 99980 6276 100008
rect 6270 99968 6276 99980
rect 6328 99968 6334 100020
rect 36538 99968 36544 100020
rect 36596 100008 36602 100020
rect 37274 100008 37280 100020
rect 36596 99980 37280 100008
rect 36596 99968 36602 99980
rect 37274 99968 37280 99980
rect 37332 99968 37338 100020
rect 34514 99900 34520 99952
rect 34572 99940 34578 99952
rect 38105 99943 38163 99949
rect 38105 99940 38117 99943
rect 34572 99912 38117 99940
rect 34572 99900 34578 99912
rect 38105 99909 38117 99912
rect 38151 99909 38163 99943
rect 38105 99903 38163 99909
rect 6089 99807 6147 99813
rect 6089 99773 6101 99807
rect 6135 99804 6147 99807
rect 13262 99804 13268 99816
rect 6135 99776 13268 99804
rect 6135 99773 6147 99776
rect 6089 99767 6147 99773
rect 13262 99764 13268 99776
rect 13320 99764 13326 99816
rect 37274 99804 37280 99816
rect 37235 99776 37280 99804
rect 37274 99764 37280 99776
rect 37332 99764 37338 99816
rect 37918 99804 37924 99816
rect 37879 99776 37924 99804
rect 37918 99764 37924 99776
rect 37976 99764 37982 99816
rect 36814 99628 36820 99680
rect 36872 99668 36878 99680
rect 37461 99671 37519 99677
rect 37461 99668 37473 99671
rect 36872 99640 37473 99668
rect 36872 99628 36878 99640
rect 37461 99637 37473 99640
rect 37507 99637 37519 99671
rect 37461 99631 37519 99637
rect 1104 99578 38824 99600
rect 1104 99526 19606 99578
rect 19658 99526 19670 99578
rect 19722 99526 19734 99578
rect 19786 99526 19798 99578
rect 19850 99526 38824 99578
rect 1104 99504 38824 99526
rect 1394 99328 1400 99340
rect 1355 99300 1400 99328
rect 1394 99288 1400 99300
rect 1452 99288 1458 99340
rect 5074 99328 5080 99340
rect 5035 99300 5080 99328
rect 5074 99288 5080 99300
rect 5132 99288 5138 99340
rect 37182 99328 37188 99340
rect 37143 99300 37188 99328
rect 37182 99288 37188 99300
rect 37240 99288 37246 99340
rect 2498 99152 2504 99204
rect 2556 99192 2562 99204
rect 5261 99195 5319 99201
rect 5261 99192 5273 99195
rect 2556 99164 5273 99192
rect 2556 99152 2562 99164
rect 5261 99161 5273 99164
rect 5307 99161 5319 99195
rect 5261 99155 5319 99161
rect 34790 99084 34796 99136
rect 34848 99124 34854 99136
rect 37369 99127 37427 99133
rect 37369 99124 37381 99127
rect 34848 99096 37381 99124
rect 34848 99084 34854 99096
rect 37369 99093 37381 99096
rect 37415 99093 37427 99127
rect 37369 99087 37427 99093
rect 1104 99034 38824 99056
rect 1104 98982 4246 99034
rect 4298 98982 4310 99034
rect 4362 98982 4374 99034
rect 4426 98982 4438 99034
rect 4490 98982 34966 99034
rect 35018 98982 35030 99034
rect 35082 98982 35094 99034
rect 35146 98982 35158 99034
rect 35210 98982 38824 99034
rect 1104 98960 38824 98982
rect 35342 98880 35348 98932
rect 35400 98880 35406 98932
rect 1394 98716 1400 98728
rect 1355 98688 1400 98716
rect 1394 98676 1400 98688
rect 1452 98676 1458 98728
rect 35360 98660 35388 98880
rect 37918 98716 37924 98728
rect 37879 98688 37924 98716
rect 37918 98676 37924 98688
rect 37976 98676 37982 98728
rect 35342 98608 35348 98660
rect 35400 98608 35406 98660
rect 35434 98540 35440 98592
rect 35492 98580 35498 98592
rect 38105 98583 38163 98589
rect 38105 98580 38117 98583
rect 35492 98552 38117 98580
rect 35492 98540 35498 98552
rect 38105 98549 38117 98552
rect 38151 98549 38163 98583
rect 38105 98543 38163 98549
rect 1104 98490 38824 98512
rect 1104 98438 19606 98490
rect 19658 98438 19670 98490
rect 19722 98438 19734 98490
rect 19786 98438 19798 98490
rect 19850 98438 38824 98490
rect 1104 98416 38824 98438
rect 2130 98336 2136 98388
rect 2188 98376 2194 98388
rect 5077 98379 5135 98385
rect 5077 98376 5089 98379
rect 2188 98348 5089 98376
rect 2188 98336 2194 98348
rect 5077 98345 5089 98348
rect 5123 98345 5135 98379
rect 5077 98339 5135 98345
rect 4890 98240 4896 98252
rect 4851 98212 4896 98240
rect 4890 98200 4896 98212
rect 4948 98200 4954 98252
rect 37090 98240 37096 98252
rect 37051 98212 37096 98240
rect 37090 98200 37096 98212
rect 37148 98200 37154 98252
rect 33410 97996 33416 98048
rect 33468 98036 33474 98048
rect 37277 98039 37335 98045
rect 37277 98036 37289 98039
rect 33468 98008 37289 98036
rect 33468 97996 33474 98008
rect 37277 98005 37289 98008
rect 37323 98005 37335 98039
rect 37277 97999 37335 98005
rect 1104 97946 38824 97968
rect 1104 97894 4246 97946
rect 4298 97894 4310 97946
rect 4362 97894 4374 97946
rect 4426 97894 4438 97946
rect 4490 97894 34966 97946
rect 35018 97894 35030 97946
rect 35082 97894 35094 97946
rect 35146 97894 35158 97946
rect 35210 97894 38824 97946
rect 1104 97872 38824 97894
rect 1946 97792 1952 97844
rect 2004 97832 2010 97844
rect 4433 97835 4491 97841
rect 4433 97832 4445 97835
rect 2004 97804 4445 97832
rect 2004 97792 2010 97804
rect 4433 97801 4445 97804
rect 4479 97801 4491 97835
rect 4433 97795 4491 97801
rect 1394 97628 1400 97640
rect 1355 97600 1400 97628
rect 1394 97588 1400 97600
rect 1452 97588 1458 97640
rect 4249 97631 4307 97637
rect 4249 97597 4261 97631
rect 4295 97628 4307 97631
rect 8386 97628 8392 97640
rect 4295 97600 8392 97628
rect 4295 97597 4307 97600
rect 4249 97591 4307 97597
rect 8386 97588 8392 97600
rect 8444 97588 8450 97640
rect 37826 97628 37832 97640
rect 37787 97600 37832 97628
rect 37826 97588 37832 97600
rect 37884 97588 37890 97640
rect 33502 97452 33508 97504
rect 33560 97492 33566 97504
rect 38013 97495 38071 97501
rect 38013 97492 38025 97495
rect 33560 97464 38025 97492
rect 33560 97452 33566 97464
rect 38013 97461 38025 97464
rect 38059 97461 38071 97495
rect 38013 97455 38071 97461
rect 1104 97402 38824 97424
rect 1104 97350 19606 97402
rect 19658 97350 19670 97402
rect 19722 97350 19734 97402
rect 19786 97350 19798 97402
rect 19850 97350 38824 97402
rect 1104 97328 38824 97350
rect 1394 97152 1400 97164
rect 1355 97124 1400 97152
rect 1394 97112 1400 97124
rect 1452 97112 1458 97164
rect 37090 97152 37096 97164
rect 37051 97124 37096 97152
rect 37090 97112 37096 97124
rect 37148 97112 37154 97164
rect 33134 96908 33140 96960
rect 33192 96948 33198 96960
rect 37277 96951 37335 96957
rect 37277 96948 37289 96951
rect 33192 96920 37289 96948
rect 33192 96908 33198 96920
rect 37277 96917 37289 96920
rect 37323 96917 37335 96951
rect 37277 96911 37335 96917
rect 1104 96858 38824 96880
rect 1104 96806 4246 96858
rect 4298 96806 4310 96858
rect 4362 96806 4374 96858
rect 4426 96806 4438 96858
rect 4490 96806 34966 96858
rect 35018 96806 35030 96858
rect 35082 96806 35094 96858
rect 35146 96806 35158 96858
rect 35210 96806 38824 96858
rect 1104 96784 38824 96806
rect 37090 96540 37096 96552
rect 37051 96512 37096 96540
rect 37090 96500 37096 96512
rect 37148 96500 37154 96552
rect 32214 96432 32220 96484
rect 32272 96472 32278 96484
rect 37918 96472 37924 96484
rect 32272 96444 37412 96472
rect 37879 96444 37924 96472
rect 32272 96432 32278 96444
rect 33686 96364 33692 96416
rect 33744 96404 33750 96416
rect 37277 96407 37335 96413
rect 37277 96404 37289 96407
rect 33744 96376 37289 96404
rect 33744 96364 33750 96376
rect 37277 96373 37289 96376
rect 37323 96373 37335 96407
rect 37384 96404 37412 96444
rect 37918 96432 37924 96444
rect 37976 96432 37982 96484
rect 38013 96407 38071 96413
rect 38013 96404 38025 96407
rect 37384 96376 38025 96404
rect 37277 96367 37335 96373
rect 38013 96373 38025 96376
rect 38059 96373 38071 96407
rect 38013 96367 38071 96373
rect 1104 96314 38824 96336
rect 1104 96262 19606 96314
rect 19658 96262 19670 96314
rect 19722 96262 19734 96314
rect 19786 96262 19798 96314
rect 19850 96262 38824 96314
rect 1104 96240 38824 96262
rect 3510 96200 3516 96212
rect 3471 96172 3516 96200
rect 3510 96160 3516 96172
rect 3568 96160 3574 96212
rect 1394 96064 1400 96076
rect 1355 96036 1400 96064
rect 1394 96024 1400 96036
rect 1452 96024 1458 96076
rect 3329 96067 3387 96073
rect 3329 96033 3341 96067
rect 3375 96064 3387 96067
rect 5258 96064 5264 96076
rect 3375 96036 5264 96064
rect 3375 96033 3387 96036
rect 3329 96027 3387 96033
rect 5258 96024 5264 96036
rect 5316 96024 5322 96076
rect 37182 96064 37188 96076
rect 37143 96036 37188 96064
rect 37182 96024 37188 96036
rect 37240 96024 37246 96076
rect 38562 95996 38568 96008
rect 26206 95968 38568 95996
rect 23474 95888 23480 95940
rect 23532 95928 23538 95940
rect 26206 95928 26234 95968
rect 38562 95956 38568 95968
rect 38620 95956 38626 96008
rect 23532 95900 26234 95928
rect 37369 95931 37427 95937
rect 23532 95888 23538 95900
rect 37369 95897 37381 95931
rect 37415 95928 37427 95931
rect 38378 95928 38384 95940
rect 37415 95900 38384 95928
rect 37415 95897 37427 95900
rect 37369 95891 37427 95897
rect 38378 95888 38384 95900
rect 38436 95888 38442 95940
rect 1104 95770 38824 95792
rect 1104 95718 4246 95770
rect 4298 95718 4310 95770
rect 4362 95718 4374 95770
rect 4426 95718 4438 95770
rect 4490 95718 34966 95770
rect 35018 95718 35030 95770
rect 35082 95718 35094 95770
rect 35146 95718 35158 95770
rect 35210 95718 38824 95770
rect 1104 95696 38824 95718
rect 2406 95616 2412 95668
rect 2464 95656 2470 95668
rect 2961 95659 3019 95665
rect 2961 95656 2973 95659
rect 2464 95628 2973 95656
rect 2464 95616 2470 95628
rect 2961 95625 2973 95628
rect 3007 95625 3019 95659
rect 2961 95619 3019 95625
rect 30742 95616 30748 95668
rect 30800 95656 30806 95668
rect 32398 95656 32404 95668
rect 30800 95628 32404 95656
rect 30800 95616 30806 95628
rect 32398 95616 32404 95628
rect 32456 95616 32462 95668
rect 1394 95452 1400 95464
rect 1355 95424 1400 95452
rect 1394 95412 1400 95424
rect 1452 95412 1458 95464
rect 2777 95455 2835 95461
rect 2777 95421 2789 95455
rect 2823 95452 2835 95455
rect 6178 95452 6184 95464
rect 2823 95424 6184 95452
rect 2823 95421 2835 95424
rect 2777 95415 2835 95421
rect 6178 95412 6184 95424
rect 6236 95412 6242 95464
rect 31478 95412 31484 95464
rect 31536 95452 31542 95464
rect 38105 95455 38163 95461
rect 38105 95452 38117 95455
rect 31536 95424 38117 95452
rect 31536 95412 31542 95424
rect 38105 95421 38117 95424
rect 38151 95421 38163 95455
rect 38105 95415 38163 95421
rect 37918 95384 37924 95396
rect 37879 95356 37924 95384
rect 37918 95344 37924 95356
rect 37976 95344 37982 95396
rect 1104 95226 38824 95248
rect 1104 95174 19606 95226
rect 19658 95174 19670 95226
rect 19722 95174 19734 95226
rect 19786 95174 19798 95226
rect 19850 95174 38824 95226
rect 1104 95152 38824 95174
rect 37182 94976 37188 94988
rect 37143 94948 37188 94976
rect 37182 94936 37188 94948
rect 37240 94936 37246 94988
rect 32030 94800 32036 94852
rect 32088 94840 32094 94852
rect 35250 94840 35256 94852
rect 32088 94812 35256 94840
rect 32088 94800 32094 94812
rect 35250 94800 35256 94812
rect 35308 94800 35314 94852
rect 33870 94732 33876 94784
rect 33928 94772 33934 94784
rect 34054 94772 34060 94784
rect 33928 94744 34060 94772
rect 33928 94732 33934 94744
rect 34054 94732 34060 94744
rect 34112 94732 34118 94784
rect 35434 94732 35440 94784
rect 35492 94772 35498 94784
rect 35894 94772 35900 94784
rect 35492 94744 35900 94772
rect 35492 94732 35498 94744
rect 35894 94732 35900 94744
rect 35952 94732 35958 94784
rect 36998 94732 37004 94784
rect 37056 94772 37062 94784
rect 37277 94775 37335 94781
rect 37277 94772 37289 94775
rect 37056 94744 37289 94772
rect 37056 94732 37062 94744
rect 37277 94741 37289 94744
rect 37323 94741 37335 94775
rect 37277 94735 37335 94741
rect 1104 94682 38824 94704
rect 1104 94630 4246 94682
rect 4298 94630 4310 94682
rect 4362 94630 4374 94682
rect 4426 94630 4438 94682
rect 4490 94630 34966 94682
rect 35018 94630 35030 94682
rect 35082 94630 35094 94682
rect 35146 94630 35158 94682
rect 35210 94630 38824 94682
rect 1104 94608 38824 94630
rect 2866 94568 2872 94580
rect 2827 94540 2872 94568
rect 2866 94528 2872 94540
rect 2924 94528 2930 94580
rect 32398 94460 32404 94512
rect 32456 94500 32462 94512
rect 34330 94500 34336 94512
rect 32456 94472 34336 94500
rect 32456 94460 32462 94472
rect 34330 94460 34336 94472
rect 34388 94460 34394 94512
rect 35250 94460 35256 94512
rect 35308 94500 35314 94512
rect 35618 94500 35624 94512
rect 35308 94472 35624 94500
rect 35308 94460 35314 94472
rect 35618 94460 35624 94472
rect 35676 94460 35682 94512
rect 1394 94364 1400 94376
rect 1355 94336 1400 94364
rect 1394 94324 1400 94336
rect 1452 94324 1458 94376
rect 2685 94367 2743 94373
rect 2685 94333 2697 94367
rect 2731 94364 2743 94367
rect 5350 94364 5356 94376
rect 2731 94336 5356 94364
rect 2731 94333 2743 94336
rect 2685 94327 2743 94333
rect 5350 94324 5356 94336
rect 5408 94324 5414 94376
rect 35434 94324 35440 94376
rect 35492 94364 35498 94376
rect 35802 94364 35808 94376
rect 35492 94336 35808 94364
rect 35492 94324 35498 94336
rect 35802 94324 35808 94336
rect 35860 94324 35866 94376
rect 37182 94364 37188 94376
rect 37143 94336 37188 94364
rect 37182 94324 37188 94336
rect 37240 94324 37246 94376
rect 37918 94296 37924 94308
rect 37879 94268 37924 94296
rect 37918 94256 37924 94268
rect 37976 94256 37982 94308
rect 35802 94188 35808 94240
rect 35860 94228 35866 94240
rect 37277 94231 37335 94237
rect 37277 94228 37289 94231
rect 35860 94200 37289 94228
rect 35860 94188 35866 94200
rect 37277 94197 37289 94200
rect 37323 94197 37335 94231
rect 37277 94191 37335 94197
rect 37550 94188 37556 94240
rect 37608 94228 37614 94240
rect 38013 94231 38071 94237
rect 38013 94228 38025 94231
rect 37608 94200 38025 94228
rect 37608 94188 37614 94200
rect 38013 94197 38025 94200
rect 38059 94197 38071 94231
rect 38013 94191 38071 94197
rect 1104 94138 38824 94160
rect 1104 94086 19606 94138
rect 19658 94086 19670 94138
rect 19722 94086 19734 94138
rect 19786 94086 19798 94138
rect 19850 94086 38824 94138
rect 1104 94064 38824 94086
rect 33962 93984 33968 94036
rect 34020 94024 34026 94036
rect 37369 94027 37427 94033
rect 37369 94024 37381 94027
rect 34020 93996 37381 94024
rect 34020 93984 34026 93996
rect 37369 93993 37381 93996
rect 37415 93993 37427 94027
rect 37369 93987 37427 93993
rect 1394 93888 1400 93900
rect 1355 93860 1400 93888
rect 1394 93848 1400 93860
rect 1452 93848 1458 93900
rect 37182 93888 37188 93900
rect 37143 93860 37188 93888
rect 37182 93848 37188 93860
rect 37240 93848 37246 93900
rect 36630 93780 36636 93832
rect 36688 93820 36694 93832
rect 37366 93820 37372 93832
rect 36688 93792 37372 93820
rect 36688 93780 36694 93792
rect 37366 93780 37372 93792
rect 37424 93780 37430 93832
rect 1104 93594 38824 93616
rect 1104 93542 4246 93594
rect 4298 93542 4310 93594
rect 4362 93542 4374 93594
rect 4426 93542 4438 93594
rect 4490 93542 34966 93594
rect 35018 93542 35030 93594
rect 35082 93542 35094 93594
rect 35146 93542 35158 93594
rect 35210 93542 38824 93594
rect 1104 93520 38824 93542
rect 30834 93304 30840 93356
rect 30892 93344 30898 93356
rect 33870 93344 33876 93356
rect 30892 93316 33876 93344
rect 30892 93304 30898 93316
rect 33870 93304 33876 93316
rect 33928 93304 33934 93356
rect 1394 93276 1400 93288
rect 1355 93248 1400 93276
rect 1394 93236 1400 93248
rect 1452 93236 1458 93288
rect 37274 93276 37280 93288
rect 37235 93248 37280 93276
rect 37274 93236 37280 93248
rect 37332 93236 37338 93288
rect 37918 93276 37924 93288
rect 37879 93248 37924 93276
rect 37918 93236 37924 93248
rect 37976 93236 37982 93288
rect 35618 93100 35624 93152
rect 35676 93140 35682 93152
rect 37461 93143 37519 93149
rect 37461 93140 37473 93143
rect 35676 93112 37473 93140
rect 35676 93100 35682 93112
rect 37461 93109 37473 93112
rect 37507 93109 37519 93143
rect 38102 93140 38108 93152
rect 38063 93112 38108 93140
rect 37461 93103 37519 93109
rect 38102 93100 38108 93112
rect 38160 93100 38166 93152
rect 1104 93050 38824 93072
rect 1104 92998 19606 93050
rect 19658 92998 19670 93050
rect 19722 92998 19734 93050
rect 19786 92998 19798 93050
rect 19850 92998 38824 93050
rect 1104 92976 38824 92998
rect 2314 92936 2320 92948
rect 2275 92908 2320 92936
rect 2314 92896 2320 92908
rect 2372 92896 2378 92948
rect 30742 92868 30748 92880
rect 30703 92840 30748 92868
rect 30742 92828 30748 92840
rect 30800 92828 30806 92880
rect 2133 92803 2191 92809
rect 2133 92769 2145 92803
rect 2179 92800 2191 92803
rect 4798 92800 4804 92812
rect 2179 92772 4804 92800
rect 2179 92769 2191 92772
rect 2133 92763 2191 92769
rect 4798 92760 4804 92772
rect 4856 92760 4862 92812
rect 21358 92760 21364 92812
rect 21416 92800 21422 92812
rect 30561 92803 30619 92809
rect 30561 92800 30573 92803
rect 21416 92772 30573 92800
rect 21416 92760 21422 92772
rect 30561 92769 30573 92772
rect 30607 92769 30619 92803
rect 30561 92763 30619 92769
rect 1104 92506 38824 92528
rect 1104 92454 4246 92506
rect 4298 92454 4310 92506
rect 4362 92454 4374 92506
rect 4426 92454 4438 92506
rect 4490 92454 34966 92506
rect 35018 92454 35030 92506
rect 35082 92454 35094 92506
rect 35146 92454 35158 92506
rect 35210 92454 38824 92506
rect 1104 92432 38824 92454
rect 1394 92188 1400 92200
rect 1355 92160 1400 92188
rect 1394 92148 1400 92160
rect 1452 92148 1458 92200
rect 37274 92188 37280 92200
rect 37235 92160 37280 92188
rect 37274 92148 37280 92160
rect 37332 92148 37338 92200
rect 37918 92188 37924 92200
rect 37879 92160 37924 92188
rect 37918 92148 37924 92160
rect 37976 92148 37982 92200
rect 37366 92012 37372 92064
rect 37424 92052 37430 92064
rect 37461 92055 37519 92061
rect 37461 92052 37473 92055
rect 37424 92024 37473 92052
rect 37424 92012 37430 92024
rect 37461 92021 37473 92024
rect 37507 92021 37519 92055
rect 37461 92015 37519 92021
rect 37826 92012 37832 92064
rect 37884 92052 37890 92064
rect 38105 92055 38163 92061
rect 38105 92052 38117 92055
rect 37884 92024 38117 92052
rect 37884 92012 37890 92024
rect 38105 92021 38117 92024
rect 38151 92021 38163 92055
rect 38105 92015 38163 92021
rect 1104 91962 38824 91984
rect 1104 91910 19606 91962
rect 19658 91910 19670 91962
rect 19722 91910 19734 91962
rect 19786 91910 19798 91962
rect 19850 91910 38824 91962
rect 1104 91888 38824 91910
rect 21542 91808 21548 91860
rect 21600 91848 21606 91860
rect 32950 91848 32956 91860
rect 21600 91820 32956 91848
rect 21600 91808 21606 91820
rect 32950 91808 32956 91820
rect 33008 91808 33014 91860
rect 19334 91740 19340 91792
rect 19392 91780 19398 91792
rect 33594 91780 33600 91792
rect 19392 91752 33600 91780
rect 19392 91740 19398 91752
rect 33594 91740 33600 91752
rect 33652 91740 33658 91792
rect 1394 91712 1400 91724
rect 1355 91684 1400 91712
rect 1394 91672 1400 91684
rect 1452 91672 1458 91724
rect 37182 91712 37188 91724
rect 37143 91684 37188 91712
rect 37182 91672 37188 91684
rect 37240 91672 37246 91724
rect 33962 91536 33968 91588
rect 34020 91576 34026 91588
rect 35618 91576 35624 91588
rect 34020 91548 35624 91576
rect 34020 91536 34026 91548
rect 35618 91536 35624 91548
rect 35676 91536 35682 91588
rect 37274 91468 37280 91520
rect 37332 91508 37338 91520
rect 37369 91511 37427 91517
rect 37369 91508 37381 91511
rect 37332 91480 37381 91508
rect 37332 91468 37338 91480
rect 37369 91477 37381 91480
rect 37415 91477 37427 91511
rect 37369 91471 37427 91477
rect 1104 91418 38824 91440
rect 1104 91366 4246 91418
rect 4298 91366 4310 91418
rect 4362 91366 4374 91418
rect 4426 91366 4438 91418
rect 4490 91366 34966 91418
rect 35018 91366 35030 91418
rect 35082 91366 35094 91418
rect 35146 91366 35158 91418
rect 35210 91366 38824 91418
rect 1104 91344 38824 91366
rect 1581 91307 1639 91313
rect 1581 91273 1593 91307
rect 1627 91304 1639 91307
rect 1670 91304 1676 91316
rect 1627 91276 1676 91304
rect 1627 91273 1639 91276
rect 1581 91267 1639 91273
rect 1670 91264 1676 91276
rect 1728 91264 1734 91316
rect 37734 91196 37740 91248
rect 37792 91236 37798 91248
rect 38105 91239 38163 91245
rect 38105 91236 38117 91239
rect 37792 91208 38117 91236
rect 37792 91196 37798 91208
rect 38105 91205 38117 91208
rect 38151 91205 38163 91239
rect 38105 91199 38163 91205
rect 27982 91128 27988 91180
rect 28040 91168 28046 91180
rect 31754 91168 31760 91180
rect 28040 91140 31760 91168
rect 28040 91128 28046 91140
rect 31754 91128 31760 91140
rect 31812 91128 31818 91180
rect 1394 91100 1400 91112
rect 1355 91072 1400 91100
rect 1394 91060 1400 91072
rect 1452 91060 1458 91112
rect 31662 91060 31668 91112
rect 31720 91100 31726 91112
rect 33042 91100 33048 91112
rect 31720 91072 33048 91100
rect 31720 91060 31726 91072
rect 33042 91060 33048 91072
rect 33100 91060 33106 91112
rect 37182 91060 37188 91112
rect 37240 91100 37246 91112
rect 37277 91103 37335 91109
rect 37277 91100 37289 91103
rect 37240 91072 37289 91100
rect 37240 91060 37246 91072
rect 37277 91069 37289 91072
rect 37323 91069 37335 91103
rect 37918 91100 37924 91112
rect 37879 91072 37924 91100
rect 37277 91063 37335 91069
rect 37918 91060 37924 91072
rect 37976 91060 37982 91112
rect 37458 90964 37464 90976
rect 37419 90936 37464 90964
rect 37458 90924 37464 90936
rect 37516 90924 37522 90976
rect 1104 90874 38824 90896
rect 1104 90822 19606 90874
rect 19658 90822 19670 90874
rect 19722 90822 19734 90874
rect 19786 90822 19798 90874
rect 19850 90822 38824 90874
rect 1104 90800 38824 90822
rect 1486 90720 1492 90772
rect 1544 90760 1550 90772
rect 1581 90763 1639 90769
rect 1581 90760 1593 90763
rect 1544 90732 1593 90760
rect 1544 90720 1550 90732
rect 1581 90729 1593 90732
rect 1627 90729 1639 90763
rect 1581 90723 1639 90729
rect 1397 90627 1455 90633
rect 1397 90593 1409 90627
rect 1443 90593 1455 90627
rect 2038 90624 2044 90636
rect 1999 90596 2044 90624
rect 1397 90587 1455 90593
rect 1412 90556 1440 90587
rect 2038 90584 2044 90596
rect 2096 90584 2102 90636
rect 2866 90556 2872 90568
rect 1412 90528 2872 90556
rect 2866 90516 2872 90528
rect 2924 90516 2930 90568
rect 1104 90330 38824 90352
rect 1104 90278 4246 90330
rect 4298 90278 4310 90330
rect 4362 90278 4374 90330
rect 4426 90278 4438 90330
rect 4490 90278 34966 90330
rect 35018 90278 35030 90330
rect 35082 90278 35094 90330
rect 35146 90278 35158 90330
rect 35210 90278 38824 90330
rect 1104 90256 38824 90278
rect 35158 90108 35164 90160
rect 35216 90148 35222 90160
rect 35894 90148 35900 90160
rect 35216 90120 35900 90148
rect 35216 90108 35222 90120
rect 35894 90108 35900 90120
rect 35952 90108 35958 90160
rect 36078 90108 36084 90160
rect 36136 90148 36142 90160
rect 38105 90151 38163 90157
rect 38105 90148 38117 90151
rect 36136 90120 38117 90148
rect 36136 90108 36142 90120
rect 38105 90117 38117 90120
rect 38151 90117 38163 90151
rect 38105 90111 38163 90117
rect 34882 90040 34888 90092
rect 34940 90080 34946 90092
rect 35434 90080 35440 90092
rect 34940 90052 35440 90080
rect 34940 90040 34946 90052
rect 35434 90040 35440 90052
rect 35492 90040 35498 90092
rect 1394 90012 1400 90024
rect 1355 89984 1400 90012
rect 1394 89972 1400 89984
rect 1452 89972 1458 90024
rect 37274 90012 37280 90024
rect 37235 89984 37280 90012
rect 37274 89972 37280 89984
rect 37332 89972 37338 90024
rect 37458 89972 37464 90024
rect 37516 89972 37522 90024
rect 37918 90012 37924 90024
rect 37879 89984 37924 90012
rect 37918 89972 37924 89984
rect 37976 89972 37982 90024
rect 33594 89904 33600 89956
rect 33652 89944 33658 89956
rect 35250 89944 35256 89956
rect 33652 89916 35256 89944
rect 33652 89904 33658 89916
rect 35250 89904 35256 89916
rect 35308 89904 35314 89956
rect 35894 89904 35900 89956
rect 35952 89944 35958 89956
rect 37476 89944 37504 89972
rect 35952 89916 37504 89944
rect 35952 89904 35958 89916
rect 34790 89836 34796 89888
rect 34848 89876 34854 89888
rect 35434 89876 35440 89888
rect 34848 89848 35440 89876
rect 34848 89836 34854 89848
rect 35434 89836 35440 89848
rect 35492 89836 35498 89888
rect 37458 89876 37464 89888
rect 37419 89848 37464 89876
rect 37458 89836 37464 89848
rect 37516 89836 37522 89888
rect 1104 89786 38824 89808
rect 1104 89734 19606 89786
rect 19658 89734 19670 89786
rect 19722 89734 19734 89786
rect 19786 89734 19798 89786
rect 19850 89734 38824 89786
rect 1104 89712 38824 89734
rect 37182 89536 37188 89548
rect 37143 89508 37188 89536
rect 37182 89496 37188 89508
rect 37240 89496 37246 89548
rect 37369 89335 37427 89341
rect 37369 89301 37381 89335
rect 37415 89332 37427 89335
rect 37642 89332 37648 89344
rect 37415 89304 37648 89332
rect 37415 89301 37427 89304
rect 37369 89295 37427 89301
rect 37642 89292 37648 89304
rect 37700 89292 37706 89344
rect 1104 89242 38824 89264
rect 1104 89190 4246 89242
rect 4298 89190 4310 89242
rect 4362 89190 4374 89242
rect 4426 89190 4438 89242
rect 4490 89190 34966 89242
rect 35018 89190 35030 89242
rect 35082 89190 35094 89242
rect 35146 89190 35158 89242
rect 35210 89190 38824 89242
rect 1104 89168 38824 89190
rect 1394 88924 1400 88936
rect 1355 88896 1400 88924
rect 1394 88884 1400 88896
rect 1452 88884 1458 88936
rect 37274 88924 37280 88936
rect 37235 88896 37280 88924
rect 37274 88884 37280 88896
rect 37332 88884 37338 88936
rect 37918 88924 37924 88936
rect 37879 88896 37924 88924
rect 37918 88884 37924 88896
rect 37976 88884 37982 88936
rect 37461 88791 37519 88797
rect 37461 88757 37473 88791
rect 37507 88788 37519 88791
rect 37826 88788 37832 88800
rect 37507 88760 37832 88788
rect 37507 88757 37519 88760
rect 37461 88751 37519 88757
rect 37826 88748 37832 88760
rect 37884 88748 37890 88800
rect 38105 88791 38163 88797
rect 38105 88757 38117 88791
rect 38151 88788 38163 88791
rect 38286 88788 38292 88800
rect 38151 88760 38292 88788
rect 38151 88757 38163 88760
rect 38105 88751 38163 88757
rect 38286 88748 38292 88760
rect 38344 88748 38350 88800
rect 1104 88698 38824 88720
rect 1104 88646 19606 88698
rect 19658 88646 19670 88698
rect 19722 88646 19734 88698
rect 19786 88646 19798 88698
rect 19850 88646 38824 88698
rect 1104 88624 38824 88646
rect 1394 88448 1400 88460
rect 1355 88420 1400 88448
rect 1394 88408 1400 88420
rect 1452 88408 1458 88460
rect 35618 88340 35624 88392
rect 35676 88380 35682 88392
rect 37550 88380 37556 88392
rect 35676 88352 37556 88380
rect 35676 88340 35682 88352
rect 37550 88340 37556 88352
rect 37608 88340 37614 88392
rect 30742 88272 30748 88324
rect 30800 88312 30806 88324
rect 34054 88312 34060 88324
rect 30800 88284 34060 88312
rect 30800 88272 30806 88284
rect 34054 88272 34060 88284
rect 34112 88272 34118 88324
rect 1104 88154 38824 88176
rect 1104 88102 4246 88154
rect 4298 88102 4310 88154
rect 4362 88102 4374 88154
rect 4426 88102 4438 88154
rect 4490 88102 34966 88154
rect 35018 88102 35030 88154
rect 35082 88102 35094 88154
rect 35146 88102 35158 88154
rect 35210 88102 38824 88154
rect 1104 88080 38824 88102
rect 34146 87904 34152 87916
rect 33704 87876 34152 87904
rect 33704 87845 33732 87876
rect 34146 87864 34152 87876
rect 34204 87864 34210 87916
rect 33689 87839 33747 87845
rect 33689 87805 33701 87839
rect 33735 87805 33747 87839
rect 33689 87799 33747 87805
rect 33778 87796 33784 87848
rect 33836 87836 33842 87848
rect 34054 87836 34060 87848
rect 33836 87808 33881 87836
rect 34015 87808 34060 87836
rect 33836 87796 33842 87808
rect 34054 87796 34060 87808
rect 34112 87796 34118 87848
rect 34330 87836 34336 87848
rect 34291 87808 34336 87836
rect 34330 87796 34336 87808
rect 34388 87796 34394 87848
rect 34609 87839 34667 87845
rect 34609 87805 34621 87839
rect 34655 87836 34667 87839
rect 35250 87836 35256 87848
rect 34655 87808 35256 87836
rect 34655 87805 34667 87808
rect 34609 87799 34667 87805
rect 35250 87796 35256 87808
rect 35308 87796 35314 87848
rect 37274 87836 37280 87848
rect 37235 87808 37280 87836
rect 37274 87796 37280 87808
rect 37332 87796 37338 87848
rect 37918 87836 37924 87848
rect 37879 87808 37924 87836
rect 37918 87796 37924 87808
rect 37976 87796 37982 87848
rect 27890 87728 27896 87780
rect 27948 87768 27954 87780
rect 33229 87771 33287 87777
rect 33229 87768 33241 87771
rect 27948 87740 33241 87768
rect 27948 87728 27954 87740
rect 33229 87737 33241 87740
rect 33275 87737 33287 87771
rect 33229 87731 33287 87737
rect 35268 87740 38148 87768
rect 35268 87712 35296 87740
rect 35250 87660 35256 87712
rect 35308 87660 35314 87712
rect 37458 87700 37464 87712
rect 37419 87672 37464 87700
rect 37458 87660 37464 87672
rect 37516 87660 37522 87712
rect 38120 87709 38148 87740
rect 38105 87703 38163 87709
rect 38105 87669 38117 87703
rect 38151 87669 38163 87703
rect 38105 87663 38163 87669
rect 1104 87610 38824 87632
rect 1104 87558 19606 87610
rect 19658 87558 19670 87610
rect 19722 87558 19734 87610
rect 19786 87558 19798 87610
rect 19850 87558 38824 87610
rect 1104 87536 38824 87558
rect 36630 87496 36636 87508
rect 33520 87468 36636 87496
rect 1394 87360 1400 87372
rect 1355 87332 1400 87360
rect 1394 87320 1400 87332
rect 1452 87320 1458 87372
rect 21174 87320 21180 87372
rect 21232 87360 21238 87372
rect 33520 87360 33548 87468
rect 36630 87456 36636 87468
rect 36688 87456 36694 87508
rect 37093 87499 37151 87505
rect 37093 87465 37105 87499
rect 37139 87496 37151 87499
rect 37182 87496 37188 87508
rect 37139 87468 37188 87496
rect 37139 87465 37151 87468
rect 37093 87459 37151 87465
rect 37182 87456 37188 87468
rect 37240 87456 37246 87508
rect 34146 87388 34152 87440
rect 34204 87428 34210 87440
rect 35894 87428 35900 87440
rect 34204 87400 35900 87428
rect 34204 87388 34210 87400
rect 35894 87388 35900 87400
rect 35952 87388 35958 87440
rect 33689 87363 33747 87369
rect 33689 87360 33701 87363
rect 21232 87332 26234 87360
rect 33520 87332 33701 87360
rect 21232 87320 21238 87332
rect 26206 87292 26234 87332
rect 33689 87329 33701 87332
rect 33735 87329 33747 87363
rect 33689 87323 33747 87329
rect 33778 87320 33784 87372
rect 33836 87360 33842 87372
rect 34057 87363 34115 87369
rect 33836 87332 33881 87360
rect 33836 87320 33842 87332
rect 34057 87329 34069 87363
rect 34103 87329 34115 87363
rect 34330 87360 34336 87372
rect 34291 87332 34336 87360
rect 34057 87323 34115 87329
rect 34072 87292 34100 87323
rect 34330 87320 34336 87332
rect 34388 87320 34394 87372
rect 34609 87363 34667 87369
rect 34609 87329 34621 87363
rect 34655 87360 34667 87363
rect 35434 87360 35440 87372
rect 34655 87332 35440 87360
rect 34655 87329 34667 87332
rect 34609 87323 34667 87329
rect 35434 87320 35440 87332
rect 35492 87320 35498 87372
rect 37182 87360 37188 87372
rect 37143 87332 37188 87360
rect 37182 87320 37188 87332
rect 37240 87320 37246 87372
rect 26206 87264 34100 87292
rect 34698 87252 34704 87304
rect 34756 87252 34762 87304
rect 20346 87184 20352 87236
rect 20404 87224 20410 87236
rect 34054 87224 34060 87236
rect 20404 87196 34060 87224
rect 20404 87184 20410 87196
rect 34054 87184 34060 87196
rect 34112 87184 34118 87236
rect 34716 87168 34744 87252
rect 36630 87184 36636 87236
rect 36688 87224 36694 87236
rect 36906 87224 36912 87236
rect 36688 87196 36912 87224
rect 36688 87184 36694 87196
rect 36906 87184 36912 87196
rect 36964 87184 36970 87236
rect 37093 87227 37151 87233
rect 37093 87193 37105 87227
rect 37139 87224 37151 87227
rect 37182 87224 37188 87236
rect 37139 87196 37188 87224
rect 37139 87193 37151 87196
rect 37093 87187 37151 87193
rect 37182 87184 37188 87196
rect 37240 87184 37246 87236
rect 28626 87116 28632 87168
rect 28684 87156 28690 87168
rect 33321 87159 33379 87165
rect 33321 87156 33333 87159
rect 28684 87128 33333 87156
rect 28684 87116 28690 87128
rect 33321 87125 33333 87128
rect 33367 87125 33379 87159
rect 33321 87119 33379 87125
rect 34698 87116 34704 87168
rect 34756 87116 34762 87168
rect 35894 87116 35900 87168
rect 35952 87156 35958 87168
rect 37369 87159 37427 87165
rect 37369 87156 37381 87159
rect 35952 87128 37381 87156
rect 35952 87116 35958 87128
rect 37369 87125 37381 87128
rect 37415 87125 37427 87159
rect 37369 87119 37427 87125
rect 1104 87066 38824 87088
rect 1104 87014 4246 87066
rect 4298 87014 4310 87066
rect 4362 87014 4374 87066
rect 4426 87014 4438 87066
rect 4490 87014 34966 87066
rect 35018 87014 35030 87066
rect 35082 87014 35094 87066
rect 35146 87014 35158 87066
rect 35210 87014 38824 87066
rect 1104 86992 38824 87014
rect 27249 86887 27307 86893
rect 27249 86853 27261 86887
rect 27295 86853 27307 86887
rect 27249 86847 27307 86853
rect 27264 86816 27292 86847
rect 30926 86844 30932 86896
rect 30984 86884 30990 86896
rect 32677 86887 32735 86893
rect 32677 86884 32689 86887
rect 30984 86856 32689 86884
rect 30984 86844 30990 86856
rect 32677 86853 32689 86856
rect 32723 86884 32735 86887
rect 33778 86884 33784 86896
rect 32723 86856 33784 86884
rect 32723 86853 32735 86856
rect 32677 86847 32735 86853
rect 33778 86844 33784 86856
rect 33836 86844 33842 86896
rect 36722 86844 36728 86896
rect 36780 86884 36786 86896
rect 38105 86887 38163 86893
rect 38105 86884 38117 86887
rect 36780 86856 38117 86884
rect 36780 86844 36786 86856
rect 38105 86853 38117 86856
rect 38151 86853 38163 86887
rect 38105 86847 38163 86853
rect 33318 86816 33324 86828
rect 27264 86788 33324 86816
rect 33318 86776 33324 86788
rect 33376 86776 33382 86828
rect 34790 86816 34796 86828
rect 33704 86788 34796 86816
rect 1394 86748 1400 86760
rect 1355 86720 1400 86748
rect 1394 86708 1400 86720
rect 1452 86708 1458 86760
rect 27065 86751 27123 86757
rect 27065 86717 27077 86751
rect 27111 86748 27123 86751
rect 27154 86748 27160 86760
rect 27111 86720 27160 86748
rect 27111 86717 27123 86720
rect 27065 86711 27123 86717
rect 27154 86708 27160 86720
rect 27212 86748 27218 86760
rect 27801 86751 27859 86757
rect 27801 86748 27813 86751
rect 27212 86720 27813 86748
rect 27212 86708 27218 86720
rect 27801 86717 27813 86720
rect 27847 86717 27859 86751
rect 27801 86711 27859 86717
rect 31757 86751 31815 86757
rect 31757 86717 31769 86751
rect 31803 86748 31815 86751
rect 32122 86748 32128 86760
rect 31803 86720 32128 86748
rect 31803 86717 31815 86720
rect 31757 86711 31815 86717
rect 32122 86708 32128 86720
rect 32180 86748 32186 86760
rect 32493 86751 32551 86757
rect 32493 86748 32505 86751
rect 32180 86720 32505 86748
rect 32180 86708 32186 86720
rect 32493 86717 32505 86720
rect 32539 86748 32551 86751
rect 32766 86748 32772 86760
rect 32539 86720 32772 86748
rect 32539 86717 32551 86720
rect 32493 86711 32551 86717
rect 32766 86708 32772 86720
rect 32824 86708 32830 86760
rect 33704 86757 33732 86788
rect 34790 86776 34796 86788
rect 34848 86776 34854 86828
rect 35434 86776 35440 86828
rect 35492 86816 35498 86828
rect 35618 86816 35624 86828
rect 35492 86788 35624 86816
rect 35492 86776 35498 86788
rect 35618 86776 35624 86788
rect 35676 86776 35682 86828
rect 33689 86751 33747 86757
rect 33689 86717 33701 86751
rect 33735 86717 33747 86751
rect 33689 86711 33747 86717
rect 33778 86708 33784 86760
rect 33836 86748 33842 86760
rect 34057 86751 34115 86757
rect 33836 86720 33881 86748
rect 33836 86708 33842 86720
rect 34057 86717 34069 86751
rect 34103 86717 34115 86751
rect 34330 86748 34336 86760
rect 34291 86720 34336 86748
rect 34057 86711 34115 86717
rect 28350 86640 28356 86692
rect 28408 86680 28414 86692
rect 33229 86683 33287 86689
rect 33229 86680 33241 86683
rect 28408 86652 33241 86680
rect 28408 86640 28414 86652
rect 33229 86649 33241 86652
rect 33275 86649 33287 86683
rect 33229 86643 33287 86649
rect 27985 86615 28043 86621
rect 27985 86581 27997 86615
rect 28031 86612 28043 86615
rect 29638 86612 29644 86624
rect 28031 86584 29644 86612
rect 28031 86581 28043 86584
rect 27985 86575 28043 86581
rect 29638 86572 29644 86584
rect 29696 86572 29702 86624
rect 31941 86615 31999 86621
rect 31941 86581 31953 86615
rect 31987 86612 31999 86615
rect 32306 86612 32312 86624
rect 31987 86584 32312 86612
rect 31987 86581 31999 86584
rect 31941 86575 31999 86581
rect 32306 86572 32312 86584
rect 32364 86572 32370 86624
rect 32766 86572 32772 86624
rect 32824 86612 32830 86624
rect 34072 86612 34100 86711
rect 34330 86708 34336 86720
rect 34388 86708 34394 86760
rect 34609 86751 34667 86757
rect 34609 86717 34621 86751
rect 34655 86748 34667 86751
rect 36814 86748 36820 86760
rect 34655 86720 36820 86748
rect 34655 86717 34667 86720
rect 34609 86711 34667 86717
rect 36814 86708 36820 86720
rect 36872 86708 36878 86760
rect 37274 86748 37280 86760
rect 37235 86720 37280 86748
rect 37274 86708 37280 86720
rect 37332 86708 37338 86760
rect 37918 86748 37924 86760
rect 37879 86720 37924 86748
rect 37918 86708 37924 86720
rect 37976 86708 37982 86760
rect 34790 86640 34796 86692
rect 34848 86680 34854 86692
rect 37182 86680 37188 86692
rect 34848 86652 37188 86680
rect 34848 86640 34854 86652
rect 37182 86640 37188 86652
rect 37240 86640 37246 86692
rect 32824 86584 34100 86612
rect 32824 86572 32830 86584
rect 35618 86572 35624 86624
rect 35676 86612 35682 86624
rect 37461 86615 37519 86621
rect 37461 86612 37473 86615
rect 35676 86584 37473 86612
rect 35676 86572 35682 86584
rect 37461 86581 37473 86584
rect 37507 86581 37519 86615
rect 37461 86575 37519 86581
rect 1104 86522 38824 86544
rect 1104 86470 19606 86522
rect 19658 86470 19670 86522
rect 19722 86470 19734 86522
rect 19786 86470 19798 86522
rect 19850 86470 38824 86522
rect 1104 86448 38824 86470
rect 26206 86380 34100 86408
rect 20530 86232 20536 86284
rect 20588 86272 20594 86284
rect 26206 86272 26234 86380
rect 33689 86275 33747 86281
rect 33689 86272 33701 86275
rect 20588 86244 26234 86272
rect 33618 86244 33701 86272
rect 20588 86232 20594 86244
rect 20438 86096 20444 86148
rect 20496 86136 20502 86148
rect 32766 86136 32772 86148
rect 20496 86108 32772 86136
rect 20496 86096 20502 86108
rect 32766 86096 32772 86108
rect 32824 86096 32830 86148
rect 33618 86136 33646 86244
rect 33689 86241 33701 86244
rect 33735 86241 33747 86275
rect 33689 86235 33747 86241
rect 33778 86232 33784 86284
rect 33836 86272 33842 86284
rect 34072 86281 34100 86380
rect 34057 86275 34115 86281
rect 33836 86244 33881 86272
rect 33836 86232 33842 86244
rect 34057 86241 34069 86275
rect 34103 86241 34115 86275
rect 34330 86272 34336 86284
rect 34291 86244 34336 86272
rect 34057 86235 34115 86241
rect 34330 86232 34336 86244
rect 34388 86232 34394 86284
rect 34514 86272 34520 86284
rect 34475 86244 34520 86272
rect 34514 86232 34520 86244
rect 34572 86232 34578 86284
rect 36538 86204 36544 86216
rect 36096 86176 36544 86204
rect 36096 86136 36124 86176
rect 36538 86164 36544 86176
rect 36596 86164 36602 86216
rect 33618 86108 36124 86136
rect 36170 86096 36176 86148
rect 36228 86136 36234 86148
rect 37090 86136 37096 86148
rect 36228 86108 37096 86136
rect 36228 86096 36234 86108
rect 37090 86096 37096 86108
rect 37148 86096 37154 86148
rect 32950 86028 32956 86080
rect 33008 86068 33014 86080
rect 33321 86071 33379 86077
rect 33321 86068 33333 86071
rect 33008 86040 33333 86068
rect 33008 86028 33014 86040
rect 33321 86037 33333 86040
rect 33367 86037 33379 86071
rect 33321 86031 33379 86037
rect 34146 86028 34152 86080
rect 34204 86068 34210 86080
rect 34330 86068 34336 86080
rect 34204 86040 34336 86068
rect 34204 86028 34210 86040
rect 34330 86028 34336 86040
rect 34388 86028 34394 86080
rect 1104 85978 38824 86000
rect 1104 85926 4246 85978
rect 4298 85926 4310 85978
rect 4362 85926 4374 85978
rect 4426 85926 4438 85978
rect 4490 85926 34966 85978
rect 35018 85926 35030 85978
rect 35082 85926 35094 85978
rect 35146 85926 35158 85978
rect 35210 85926 38824 85978
rect 1104 85904 38824 85926
rect 27341 85867 27399 85873
rect 27341 85833 27353 85867
rect 27387 85864 27399 85867
rect 31754 85864 31760 85876
rect 27387 85836 31760 85864
rect 27387 85833 27399 85836
rect 27341 85827 27399 85833
rect 31754 85824 31760 85836
rect 31812 85824 31818 85876
rect 32306 85824 32312 85876
rect 32364 85864 32370 85876
rect 32766 85864 32772 85876
rect 32364 85836 32772 85864
rect 32364 85824 32370 85836
rect 32766 85824 32772 85836
rect 32824 85824 32830 85876
rect 36170 85824 36176 85876
rect 36228 85864 36234 85876
rect 38105 85867 38163 85873
rect 38105 85864 38117 85867
rect 36228 85836 38117 85864
rect 36228 85824 36234 85836
rect 38105 85833 38117 85836
rect 38151 85833 38163 85867
rect 38105 85827 38163 85833
rect 16942 85756 16948 85808
rect 17000 85796 17006 85808
rect 17000 85768 32812 85796
rect 17000 85756 17006 85768
rect 32306 85688 32312 85740
rect 32364 85728 32370 85740
rect 32364 85700 32536 85728
rect 32364 85688 32370 85700
rect 1394 85660 1400 85672
rect 1355 85632 1400 85660
rect 1394 85620 1400 85632
rect 1452 85620 1458 85672
rect 27154 85660 27160 85672
rect 27115 85632 27160 85660
rect 27154 85620 27160 85632
rect 27212 85620 27218 85672
rect 32398 85660 32404 85672
rect 32359 85632 32404 85660
rect 32398 85620 32404 85632
rect 32456 85620 32462 85672
rect 32508 85669 32536 85700
rect 32784 85669 32812 85768
rect 33318 85756 33324 85808
rect 33376 85756 33382 85808
rect 36630 85756 36636 85808
rect 36688 85796 36694 85808
rect 37461 85799 37519 85805
rect 37461 85796 37473 85799
rect 36688 85768 37473 85796
rect 36688 85756 36694 85768
rect 37461 85765 37473 85768
rect 37507 85765 37519 85799
rect 37461 85759 37519 85765
rect 33336 85728 33364 85756
rect 33060 85700 33364 85728
rect 33060 85669 33088 85700
rect 32493 85663 32551 85669
rect 32493 85629 32505 85663
rect 32539 85629 32551 85663
rect 32493 85623 32551 85629
rect 32769 85663 32827 85669
rect 32769 85629 32781 85663
rect 32815 85629 32827 85663
rect 32769 85623 32827 85629
rect 33045 85663 33103 85669
rect 33045 85629 33057 85663
rect 33091 85629 33103 85663
rect 33045 85623 33103 85629
rect 33321 85663 33379 85669
rect 33321 85629 33333 85663
rect 33367 85660 33379 85663
rect 33962 85660 33968 85672
rect 33367 85632 33968 85660
rect 33367 85629 33379 85632
rect 33321 85623 33379 85629
rect 33962 85620 33968 85632
rect 34020 85620 34026 85672
rect 37274 85660 37280 85672
rect 37235 85632 37280 85660
rect 37274 85620 37280 85632
rect 37332 85620 37338 85672
rect 37918 85660 37924 85672
rect 37879 85632 37924 85660
rect 37918 85620 37924 85632
rect 37976 85620 37982 85672
rect 28258 85552 28264 85604
rect 28316 85592 28322 85604
rect 31941 85595 31999 85601
rect 31941 85592 31953 85595
rect 28316 85564 31953 85592
rect 28316 85552 28322 85564
rect 31941 85561 31953 85564
rect 31987 85561 31999 85595
rect 31941 85555 31999 85561
rect 34514 85552 34520 85604
rect 34572 85592 34578 85604
rect 35618 85592 35624 85604
rect 34572 85564 35624 85592
rect 34572 85552 34578 85564
rect 35618 85552 35624 85564
rect 35676 85552 35682 85604
rect 32398 85484 32404 85536
rect 32456 85524 32462 85536
rect 33594 85524 33600 85536
rect 32456 85496 33600 85524
rect 32456 85484 32462 85496
rect 33594 85484 33600 85496
rect 33652 85484 33658 85536
rect 1104 85434 38824 85456
rect 1104 85382 19606 85434
rect 19658 85382 19670 85434
rect 19722 85382 19734 85434
rect 19786 85382 19798 85434
rect 19850 85382 38824 85434
rect 1104 85360 38824 85382
rect 1394 85184 1400 85196
rect 1355 85156 1400 85184
rect 1394 85144 1400 85156
rect 1452 85144 1458 85196
rect 32122 85144 32128 85196
rect 32180 85184 32186 85196
rect 33045 85187 33103 85193
rect 33045 85184 33057 85187
rect 32180 85156 33057 85184
rect 32180 85144 32186 85156
rect 33045 85153 33057 85156
rect 33091 85153 33103 85187
rect 33045 85147 33103 85153
rect 33229 84983 33287 84989
rect 33229 84949 33241 84983
rect 33275 84980 33287 84983
rect 33594 84980 33600 84992
rect 33275 84952 33600 84980
rect 33275 84949 33287 84952
rect 33229 84943 33287 84949
rect 33594 84940 33600 84952
rect 33652 84940 33658 84992
rect 1104 84890 38824 84912
rect 1104 84838 4246 84890
rect 4298 84838 4310 84890
rect 4362 84838 4374 84890
rect 4426 84838 4438 84890
rect 4490 84838 34966 84890
rect 35018 84838 35030 84890
rect 35082 84838 35094 84890
rect 35146 84838 35158 84890
rect 35210 84838 38824 84890
rect 1104 84816 38824 84838
rect 33042 84736 33048 84788
rect 33100 84776 33106 84788
rect 36538 84776 36544 84788
rect 33100 84748 36544 84776
rect 33100 84736 33106 84748
rect 36538 84736 36544 84748
rect 36596 84736 36602 84788
rect 27157 84711 27215 84717
rect 27157 84677 27169 84711
rect 27203 84708 27215 84711
rect 34146 84708 34152 84720
rect 27203 84680 34152 84708
rect 27203 84677 27215 84680
rect 27157 84671 27215 84677
rect 34146 84668 34152 84680
rect 34204 84668 34210 84720
rect 17678 84600 17684 84652
rect 17736 84640 17742 84652
rect 17736 84612 32904 84640
rect 17736 84600 17742 84612
rect 26970 84572 26976 84584
rect 26883 84544 26976 84572
rect 26970 84532 26976 84544
rect 27028 84572 27034 84584
rect 27154 84572 27160 84584
rect 27028 84544 27160 84572
rect 27028 84532 27034 84544
rect 27154 84532 27160 84544
rect 27212 84532 27218 84584
rect 31297 84575 31355 84581
rect 31297 84541 31309 84575
rect 31343 84572 31355 84575
rect 32122 84572 32128 84584
rect 31343 84544 32128 84572
rect 31343 84541 31355 84544
rect 31297 84535 31355 84541
rect 32122 84532 32128 84544
rect 32180 84532 32186 84584
rect 32490 84572 32496 84584
rect 32451 84544 32496 84572
rect 32490 84532 32496 84544
rect 32548 84532 32554 84584
rect 32766 84572 32772 84584
rect 32727 84544 32772 84572
rect 32766 84532 32772 84544
rect 32824 84532 32830 84584
rect 32876 84581 32904 84612
rect 32861 84575 32919 84581
rect 32861 84541 32873 84575
rect 32907 84541 32919 84575
rect 32861 84535 32919 84541
rect 33137 84575 33195 84581
rect 33137 84541 33149 84575
rect 33183 84572 33195 84575
rect 33318 84572 33324 84584
rect 33183 84544 33324 84572
rect 33183 84541 33195 84544
rect 33137 84535 33195 84541
rect 33318 84532 33324 84544
rect 33376 84532 33382 84584
rect 33413 84575 33471 84581
rect 33413 84541 33425 84575
rect 33459 84572 33471 84575
rect 33870 84572 33876 84584
rect 33459 84544 33876 84572
rect 33459 84541 33471 84544
rect 33413 84535 33471 84541
rect 33870 84532 33876 84544
rect 33928 84532 33934 84584
rect 37274 84572 37280 84584
rect 37235 84544 37280 84572
rect 37274 84532 37280 84544
rect 37332 84532 37338 84584
rect 37918 84572 37924 84584
rect 37879 84544 37924 84572
rect 37918 84532 37924 84544
rect 37976 84532 37982 84584
rect 29362 84464 29368 84516
rect 29420 84504 29426 84516
rect 32033 84507 32091 84513
rect 32033 84504 32045 84507
rect 29420 84476 32045 84504
rect 29420 84464 29426 84476
rect 32033 84473 32045 84476
rect 32079 84473 32091 84507
rect 32784 84504 32812 84532
rect 34054 84504 34060 84516
rect 32784 84476 34060 84504
rect 32033 84467 32091 84473
rect 34054 84464 34060 84476
rect 34112 84464 34118 84516
rect 31481 84439 31539 84445
rect 31481 84405 31493 84439
rect 31527 84436 31539 84439
rect 33778 84436 33784 84448
rect 31527 84408 33784 84436
rect 31527 84405 31539 84408
rect 31481 84399 31539 84405
rect 33778 84396 33784 84408
rect 33836 84396 33842 84448
rect 36814 84396 36820 84448
rect 36872 84436 36878 84448
rect 37461 84439 37519 84445
rect 37461 84436 37473 84439
rect 36872 84408 37473 84436
rect 36872 84396 36878 84408
rect 37461 84405 37473 84408
rect 37507 84405 37519 84439
rect 37461 84399 37519 84405
rect 38105 84439 38163 84445
rect 38105 84405 38117 84439
rect 38151 84436 38163 84439
rect 39390 84436 39396 84448
rect 38151 84408 39396 84436
rect 38151 84405 38163 84408
rect 38105 84399 38163 84405
rect 39390 84396 39396 84408
rect 39448 84396 39454 84448
rect 1104 84346 38824 84368
rect 1104 84294 19606 84346
rect 19658 84294 19670 84346
rect 19722 84294 19734 84346
rect 19786 84294 19798 84346
rect 19850 84294 38824 84346
rect 1104 84272 38824 84294
rect 32122 84192 32128 84244
rect 32180 84232 32186 84244
rect 32490 84232 32496 84244
rect 32180 84204 32496 84232
rect 32180 84192 32186 84204
rect 32490 84192 32496 84204
rect 32548 84192 32554 84244
rect 33318 84192 33324 84244
rect 33376 84232 33382 84244
rect 33376 84204 34192 84232
rect 33376 84192 33382 84204
rect 32398 84164 32404 84176
rect 31404 84136 32404 84164
rect 1394 84096 1400 84108
rect 1355 84068 1400 84096
rect 1394 84056 1400 84068
rect 1452 84056 1458 84108
rect 30834 84056 30840 84108
rect 30892 84096 30898 84108
rect 31404 84105 31432 84136
rect 32398 84124 32404 84136
rect 32456 84164 32462 84176
rect 32766 84164 32772 84176
rect 32456 84136 32772 84164
rect 32456 84124 32462 84136
rect 32766 84124 32772 84136
rect 32824 84124 32830 84176
rect 34054 84164 34060 84176
rect 33796 84136 34060 84164
rect 33796 84105 33824 84136
rect 34054 84124 34060 84136
rect 34112 84124 34118 84176
rect 33962 84105 33968 84108
rect 31113 84099 31171 84105
rect 31113 84096 31125 84099
rect 30892 84068 31125 84096
rect 30892 84056 30898 84068
rect 31113 84065 31125 84068
rect 31159 84065 31171 84099
rect 31113 84059 31171 84065
rect 31389 84099 31447 84105
rect 31389 84065 31401 84099
rect 31435 84065 31447 84099
rect 31389 84059 31447 84065
rect 31481 84099 31539 84105
rect 31481 84065 31493 84099
rect 31527 84065 31539 84099
rect 31481 84059 31539 84065
rect 31757 84099 31815 84105
rect 31757 84065 31769 84099
rect 31803 84065 31815 84099
rect 31757 84059 31815 84065
rect 32033 84099 32091 84105
rect 32033 84065 32045 84099
rect 32079 84096 32091 84099
rect 33505 84099 33563 84105
rect 32079 84068 33364 84096
rect 32079 84065 32091 84068
rect 32033 84059 32091 84065
rect 16482 83988 16488 84040
rect 16540 84028 16546 84040
rect 31496 84028 31524 84059
rect 16540 84000 31524 84028
rect 31772 84028 31800 84059
rect 31772 84000 33272 84028
rect 16540 83988 16546 84000
rect 30374 83920 30380 83972
rect 30432 83960 30438 83972
rect 30432 83932 30880 83960
rect 30432 83920 30438 83932
rect 29178 83852 29184 83904
rect 29236 83892 29242 83904
rect 30745 83895 30803 83901
rect 30745 83892 30757 83895
rect 29236 83864 30757 83892
rect 29236 83852 29242 83864
rect 30745 83861 30757 83864
rect 30791 83861 30803 83895
rect 30852 83892 30880 83932
rect 33137 83895 33195 83901
rect 33137 83892 33149 83895
rect 30852 83864 33149 83892
rect 30745 83855 30803 83861
rect 33137 83861 33149 83864
rect 33183 83861 33195 83895
rect 33244 83892 33272 84000
rect 33336 83960 33364 84068
rect 33505 84065 33517 84099
rect 33551 84096 33563 84099
rect 33781 84099 33839 84105
rect 33551 84068 33732 84096
rect 33551 84065 33563 84068
rect 33505 84059 33563 84065
rect 33704 83960 33732 84068
rect 33781 84065 33793 84099
rect 33827 84065 33839 84099
rect 33781 84059 33839 84065
rect 33919 84099 33968 84105
rect 33919 84065 33931 84099
rect 33965 84065 33968 84099
rect 33919 84059 33968 84065
rect 33962 84056 33968 84059
rect 34020 84056 34026 84108
rect 34164 84105 34192 84204
rect 37366 84164 37372 84176
rect 34440 84136 37372 84164
rect 34440 84105 34468 84136
rect 37366 84124 37372 84136
rect 37424 84124 37430 84176
rect 34149 84099 34207 84105
rect 34149 84065 34161 84099
rect 34195 84065 34207 84099
rect 34149 84059 34207 84065
rect 34425 84099 34483 84105
rect 34425 84065 34437 84099
rect 34471 84065 34483 84099
rect 37182 84096 37188 84108
rect 37143 84068 37188 84096
rect 34425 84059 34483 84065
rect 37182 84056 37188 84068
rect 37240 84056 37246 84108
rect 35526 83960 35532 83972
rect 33336 83932 33646 83960
rect 33704 83932 35532 83960
rect 33318 83892 33324 83904
rect 33244 83864 33324 83892
rect 33137 83855 33195 83861
rect 33318 83852 33324 83864
rect 33376 83852 33382 83904
rect 33618 83892 33646 83932
rect 35526 83920 35532 83932
rect 35584 83920 35590 83972
rect 34790 83892 34796 83904
rect 33618 83864 34796 83892
rect 34790 83852 34796 83864
rect 34848 83852 34854 83904
rect 37366 83892 37372 83904
rect 37327 83864 37372 83892
rect 37366 83852 37372 83864
rect 37424 83852 37430 83904
rect 1104 83802 38824 83824
rect 1104 83750 4246 83802
rect 4298 83750 4310 83802
rect 4362 83750 4374 83802
rect 4426 83750 4438 83802
rect 4490 83750 34966 83802
rect 35018 83750 35030 83802
rect 35082 83750 35094 83802
rect 35146 83750 35158 83802
rect 35210 83750 38824 83802
rect 1104 83728 38824 83750
rect 32766 83648 32772 83700
rect 32824 83688 32830 83700
rect 34330 83688 34336 83700
rect 32824 83660 34336 83688
rect 32824 83648 32830 83660
rect 34330 83648 34336 83660
rect 34388 83648 34394 83700
rect 17770 83512 17776 83564
rect 17828 83552 17834 83564
rect 29270 83552 29276 83564
rect 17828 83524 29276 83552
rect 17828 83512 17834 83524
rect 29270 83512 29276 83524
rect 29328 83512 29334 83564
rect 33318 83552 33324 83564
rect 29472 83524 32720 83552
rect 1394 83484 1400 83496
rect 1355 83456 1400 83484
rect 1394 83444 1400 83456
rect 1452 83444 1458 83496
rect 17862 83444 17868 83496
rect 17920 83484 17926 83496
rect 29472 83484 29500 83524
rect 32306 83484 32312 83496
rect 17920 83456 29500 83484
rect 32267 83456 32312 83484
rect 17920 83444 17926 83456
rect 32306 83444 32312 83456
rect 32364 83444 32370 83496
rect 32398 83444 32404 83496
rect 32456 83484 32462 83496
rect 32692 83493 32720 83524
rect 32968 83524 33324 83552
rect 32968 83493 32996 83524
rect 33318 83512 33324 83524
rect 33376 83512 33382 83564
rect 38102 83552 38108 83564
rect 36188 83524 38108 83552
rect 32677 83487 32735 83493
rect 32456 83456 32501 83484
rect 32456 83444 32462 83456
rect 32677 83453 32689 83487
rect 32723 83453 32735 83487
rect 32677 83447 32735 83453
rect 32953 83487 33011 83493
rect 32953 83453 32965 83487
rect 32999 83453 33011 83487
rect 32953 83447 33011 83453
rect 33229 83487 33287 83493
rect 33229 83453 33241 83487
rect 33275 83484 33287 83487
rect 36188 83484 36216 83524
rect 38102 83512 38108 83524
rect 38160 83512 38166 83564
rect 37274 83484 37280 83496
rect 33275 83456 36216 83484
rect 37235 83456 37280 83484
rect 33275 83453 33287 83456
rect 33229 83447 33287 83453
rect 37274 83444 37280 83456
rect 37332 83444 37338 83496
rect 37918 83484 37924 83496
rect 37879 83456 37924 83484
rect 37918 83444 37924 83456
rect 37976 83444 37982 83496
rect 29546 83376 29552 83428
rect 29604 83416 29610 83428
rect 31849 83419 31907 83425
rect 31849 83416 31861 83419
rect 29604 83388 31861 83416
rect 29604 83376 29610 83388
rect 31849 83385 31861 83388
rect 31895 83385 31907 83419
rect 33594 83416 33600 83428
rect 31849 83379 31907 83385
rect 32600 83388 33600 83416
rect 32122 83308 32128 83360
rect 32180 83348 32186 83360
rect 32600 83348 32628 83388
rect 33594 83376 33600 83388
rect 33652 83376 33658 83428
rect 32180 83320 32628 83348
rect 32180 83308 32186 83320
rect 36538 83308 36544 83360
rect 36596 83348 36602 83360
rect 37461 83351 37519 83357
rect 37461 83348 37473 83351
rect 36596 83320 37473 83348
rect 36596 83308 36602 83320
rect 37461 83317 37473 83320
rect 37507 83317 37519 83351
rect 37461 83311 37519 83317
rect 38105 83351 38163 83357
rect 38105 83317 38117 83351
rect 38151 83348 38163 83351
rect 39022 83348 39028 83360
rect 38151 83320 39028 83348
rect 38151 83317 38163 83320
rect 38105 83311 38163 83317
rect 39022 83308 39028 83320
rect 39080 83308 39086 83360
rect 1104 83258 38824 83280
rect 1104 83206 19606 83258
rect 19658 83206 19670 83258
rect 19722 83206 19734 83258
rect 19786 83206 19798 83258
rect 19850 83206 38824 83258
rect 1104 83184 38824 83206
rect 29270 83104 29276 83156
rect 29328 83144 29334 83156
rect 29328 83116 33916 83144
rect 29328 83104 29334 83116
rect 32122 83076 32128 83088
rect 31404 83048 32128 83076
rect 29270 82968 29276 83020
rect 29328 83008 29334 83020
rect 29546 83008 29552 83020
rect 29328 82980 29552 83008
rect 29328 82968 29334 82980
rect 29546 82968 29552 82980
rect 29604 82968 29610 83020
rect 30650 83008 30656 83020
rect 30611 82980 30656 83008
rect 30650 82968 30656 82980
rect 30708 82968 30714 83020
rect 30742 82968 30748 83020
rect 30800 83008 30806 83020
rect 31404 83017 31432 83048
rect 32122 83036 32128 83048
rect 32180 83036 32186 83088
rect 31113 83011 31171 83017
rect 31113 83008 31125 83011
rect 30800 82980 31125 83008
rect 30800 82968 30806 82980
rect 31113 82977 31125 82980
rect 31159 82977 31171 83011
rect 31113 82971 31171 82977
rect 31389 83011 31447 83017
rect 31389 82977 31401 83011
rect 31435 82977 31447 83011
rect 31389 82971 31447 82977
rect 31481 83011 31539 83017
rect 31481 82977 31493 83011
rect 31527 82977 31539 83011
rect 31481 82971 31539 82977
rect 16022 82900 16028 82952
rect 16080 82940 16086 82952
rect 31496 82940 31524 82971
rect 31754 82968 31760 83020
rect 31812 83008 31818 83020
rect 32033 83011 32091 83017
rect 31812 82980 31857 83008
rect 31812 82968 31818 82980
rect 32033 82977 32045 83011
rect 32079 83008 32091 83011
rect 32766 83008 32772 83020
rect 32079 82980 32772 83008
rect 32079 82977 32091 82980
rect 32033 82971 32091 82977
rect 32766 82968 32772 82980
rect 32824 82968 32830 83020
rect 33505 83011 33563 83017
rect 33505 82977 33517 83011
rect 33551 82977 33563 83011
rect 33505 82971 33563 82977
rect 16080 82912 31524 82940
rect 31772 82940 31800 82968
rect 33520 82940 33548 82971
rect 33594 82968 33600 83020
rect 33652 83008 33658 83020
rect 33888 83017 33916 83116
rect 35986 83076 35992 83088
rect 34072 83048 35992 83076
rect 33873 83011 33931 83017
rect 33652 82980 33697 83008
rect 33652 82968 33658 82980
rect 33873 82977 33885 83011
rect 33919 82977 33931 83011
rect 33873 82971 33931 82977
rect 34072 82940 34100 83048
rect 35986 83036 35992 83048
rect 36044 83036 36050 83088
rect 34149 83011 34207 83017
rect 34149 82977 34161 83011
rect 34195 82977 34207 83011
rect 34149 82971 34207 82977
rect 34425 83011 34483 83017
rect 34425 82977 34437 83011
rect 34471 83008 34483 83011
rect 37734 83008 37740 83020
rect 34471 82980 37740 83008
rect 34471 82977 34483 82980
rect 34425 82971 34483 82977
rect 31772 82912 33456 82940
rect 33520 82912 34100 82940
rect 16080 82900 16086 82912
rect 24210 82832 24216 82884
rect 24268 82872 24274 82884
rect 33137 82875 33195 82881
rect 33137 82872 33149 82875
rect 24268 82844 33149 82872
rect 24268 82832 24274 82844
rect 33137 82841 33149 82844
rect 33183 82841 33195 82875
rect 33428 82872 33456 82912
rect 34164 82872 34192 82971
rect 37734 82968 37740 82980
rect 37792 82968 37798 83020
rect 33428 82844 34192 82872
rect 33137 82835 33195 82841
rect 37550 82832 37556 82884
rect 37608 82872 37614 82884
rect 37734 82872 37740 82884
rect 37608 82844 37740 82872
rect 37608 82832 37614 82844
rect 37734 82832 37740 82844
rect 37792 82832 37798 82884
rect 32766 82764 32772 82816
rect 32824 82804 32830 82816
rect 37090 82804 37096 82816
rect 32824 82776 37096 82804
rect 32824 82764 32830 82776
rect 37090 82764 37096 82776
rect 37148 82764 37154 82816
rect 1104 82714 38824 82736
rect 1104 82662 4246 82714
rect 4298 82662 4310 82714
rect 4362 82662 4374 82714
rect 4426 82662 4438 82714
rect 4490 82662 34966 82714
rect 35018 82662 35030 82714
rect 35082 82662 35094 82714
rect 35146 82662 35158 82714
rect 35210 82662 38824 82714
rect 1104 82640 38824 82662
rect 32030 82532 32036 82544
rect 31956 82504 32036 82532
rect 1394 82396 1400 82408
rect 1355 82368 1400 82396
rect 1394 82356 1400 82368
rect 1452 82356 1458 82408
rect 31956 82405 31984 82504
rect 32030 82492 32036 82504
rect 32088 82492 32094 82544
rect 32122 82464 32128 82476
rect 32048 82436 32128 82464
rect 32048 82405 32076 82436
rect 32122 82424 32128 82436
rect 32180 82424 32186 82476
rect 38010 82464 38016 82476
rect 32876 82436 38016 82464
rect 31941 82399 31999 82405
rect 31941 82365 31953 82399
rect 31987 82365 31999 82399
rect 31941 82359 31999 82365
rect 32033 82399 32091 82405
rect 32033 82365 32045 82399
rect 32079 82365 32091 82399
rect 32306 82396 32312 82408
rect 32267 82368 32312 82396
rect 32033 82359 32091 82365
rect 32306 82356 32312 82368
rect 32364 82356 32370 82408
rect 32876 82405 32904 82436
rect 38010 82424 38016 82436
rect 38068 82424 38074 82476
rect 32585 82399 32643 82405
rect 32585 82365 32597 82399
rect 32631 82365 32643 82399
rect 32585 82359 32643 82365
rect 32861 82399 32919 82405
rect 32861 82365 32873 82399
rect 32907 82365 32919 82399
rect 37274 82396 37280 82408
rect 37235 82368 37280 82396
rect 32861 82359 32919 82365
rect 29822 82288 29828 82340
rect 29880 82328 29886 82340
rect 31481 82331 31539 82337
rect 31481 82328 31493 82331
rect 29880 82300 31493 82328
rect 29880 82288 29886 82300
rect 31481 82297 31493 82300
rect 31527 82297 31539 82331
rect 31481 82291 31539 82297
rect 31754 82220 31760 82272
rect 31812 82260 31818 82272
rect 32398 82260 32404 82272
rect 31812 82232 32404 82260
rect 31812 82220 31818 82232
rect 32398 82220 32404 82232
rect 32456 82260 32462 82272
rect 32600 82260 32628 82359
rect 37274 82356 37280 82368
rect 37332 82356 37338 82408
rect 37918 82396 37924 82408
rect 37879 82368 37924 82396
rect 37918 82356 37924 82368
rect 37976 82356 37982 82408
rect 32456 82232 32628 82260
rect 32456 82220 32462 82232
rect 35526 82220 35532 82272
rect 35584 82260 35590 82272
rect 35802 82260 35808 82272
rect 35584 82232 35808 82260
rect 35584 82220 35590 82232
rect 35802 82220 35808 82232
rect 35860 82220 35866 82272
rect 37461 82263 37519 82269
rect 37461 82229 37473 82263
rect 37507 82260 37519 82263
rect 37550 82260 37556 82272
rect 37507 82232 37556 82260
rect 37507 82229 37519 82232
rect 37461 82223 37519 82229
rect 37550 82220 37556 82232
rect 37608 82220 37614 82272
rect 38105 82263 38163 82269
rect 38105 82229 38117 82263
rect 38151 82260 38163 82263
rect 39942 82260 39948 82272
rect 38151 82232 39948 82260
rect 38151 82229 38163 82232
rect 38105 82223 38163 82229
rect 39942 82220 39948 82232
rect 40000 82220 40006 82272
rect 1104 82170 38824 82192
rect 1104 82118 19606 82170
rect 19658 82118 19670 82170
rect 19722 82118 19734 82170
rect 19786 82118 19798 82170
rect 19850 82118 38824 82170
rect 1104 82096 38824 82118
rect 31202 82056 31208 82068
rect 30944 82028 31208 82056
rect 1394 81920 1400 81932
rect 1355 81892 1400 81920
rect 1394 81880 1400 81892
rect 1452 81880 1458 81932
rect 30944 81920 30972 82028
rect 31202 82016 31208 82028
rect 31260 82016 31266 82068
rect 37642 82056 37648 82068
rect 32600 82028 37648 82056
rect 32122 81988 32128 82000
rect 31404 81960 32128 81988
rect 31404 81929 31432 81960
rect 32122 81948 32128 81960
rect 32180 81948 32186 82000
rect 31113 81923 31171 81929
rect 31113 81920 31125 81923
rect 30944 81892 31125 81920
rect 31113 81889 31125 81892
rect 31159 81889 31171 81923
rect 31113 81883 31171 81889
rect 31389 81923 31447 81929
rect 31389 81889 31401 81923
rect 31435 81889 31447 81923
rect 31389 81883 31447 81889
rect 31481 81923 31539 81929
rect 31481 81889 31493 81923
rect 31527 81889 31539 81923
rect 31481 81883 31539 81889
rect 16666 81812 16672 81864
rect 16724 81852 16730 81864
rect 31496 81852 31524 81883
rect 31754 81880 31760 81932
rect 31812 81920 31818 81932
rect 32033 81923 32091 81929
rect 31812 81892 31857 81920
rect 31812 81880 31818 81892
rect 32033 81889 32045 81923
rect 32079 81920 32091 81923
rect 32600 81920 32628 82028
rect 37642 82016 37648 82028
rect 37700 82016 37706 82068
rect 38194 81988 38200 82000
rect 33796 81960 38200 81988
rect 32079 81892 32628 81920
rect 33505 81923 33563 81929
rect 32079 81889 32091 81892
rect 32033 81883 32091 81889
rect 33505 81889 33517 81923
rect 33551 81889 33563 81923
rect 33505 81883 33563 81889
rect 16724 81824 31524 81852
rect 33520 81852 33548 81883
rect 33594 81880 33600 81932
rect 33652 81920 33658 81932
rect 33652 81892 33697 81920
rect 33652 81880 33658 81892
rect 33796 81852 33824 81960
rect 38194 81948 38200 81960
rect 38252 81948 38258 82000
rect 33873 81923 33931 81929
rect 33873 81889 33885 81923
rect 33919 81920 33931 81923
rect 34146 81920 34152 81932
rect 33919 81892 34008 81920
rect 34107 81892 34152 81920
rect 33919 81889 33931 81892
rect 33873 81883 33931 81889
rect 33520 81824 33824 81852
rect 16724 81812 16730 81824
rect 15838 81744 15844 81796
rect 15896 81784 15902 81796
rect 33980 81784 34008 81892
rect 34146 81880 34152 81892
rect 34204 81880 34210 81932
rect 34425 81923 34483 81929
rect 34425 81889 34437 81923
rect 34471 81920 34483 81923
rect 36078 81920 36084 81932
rect 34471 81892 36084 81920
rect 34471 81889 34483 81892
rect 34425 81883 34483 81889
rect 36078 81880 36084 81892
rect 36136 81880 36142 81932
rect 37182 81920 37188 81932
rect 37143 81892 37188 81920
rect 37182 81880 37188 81892
rect 37240 81880 37246 81932
rect 15896 81756 34008 81784
rect 15896 81744 15902 81756
rect 36262 81744 36268 81796
rect 36320 81784 36326 81796
rect 37182 81784 37188 81796
rect 36320 81756 37188 81784
rect 36320 81744 36326 81756
rect 37182 81744 37188 81756
rect 37240 81744 37246 81796
rect 26510 81676 26516 81728
rect 26568 81716 26574 81728
rect 30745 81719 30803 81725
rect 30745 81716 30757 81719
rect 26568 81688 30757 81716
rect 26568 81676 26574 81688
rect 30745 81685 30757 81688
rect 30791 81685 30803 81719
rect 30745 81679 30803 81685
rect 31754 81676 31760 81728
rect 31812 81716 31818 81728
rect 32766 81716 32772 81728
rect 31812 81688 32772 81716
rect 31812 81676 31818 81688
rect 32766 81676 32772 81688
rect 32824 81676 32830 81728
rect 33134 81716 33140 81728
rect 33095 81688 33140 81716
rect 33134 81676 33140 81688
rect 33192 81676 33198 81728
rect 33594 81676 33600 81728
rect 33652 81716 33658 81728
rect 33778 81716 33784 81728
rect 33652 81688 33784 81716
rect 33652 81676 33658 81688
rect 33778 81676 33784 81688
rect 33836 81676 33842 81728
rect 37369 81719 37427 81725
rect 37369 81685 37381 81719
rect 37415 81716 37427 81719
rect 39666 81716 39672 81728
rect 37415 81688 39672 81716
rect 37415 81685 37427 81688
rect 37369 81679 37427 81685
rect 39666 81676 39672 81688
rect 39724 81676 39730 81728
rect 1104 81626 38824 81648
rect 1104 81574 4246 81626
rect 4298 81574 4310 81626
rect 4362 81574 4374 81626
rect 4426 81574 4438 81626
rect 4490 81574 34966 81626
rect 35018 81574 35030 81626
rect 35082 81574 35094 81626
rect 35146 81574 35158 81626
rect 35210 81574 38824 81626
rect 1104 81552 38824 81574
rect 23566 81472 23572 81524
rect 23624 81512 23630 81524
rect 33134 81512 33140 81524
rect 23624 81484 33140 81512
rect 23624 81472 23630 81484
rect 33134 81472 33140 81484
rect 33192 81472 33198 81524
rect 36262 81472 36268 81524
rect 36320 81512 36326 81524
rect 36722 81512 36728 81524
rect 36320 81484 36728 81512
rect 36320 81472 36326 81484
rect 36722 81472 36728 81484
rect 36780 81472 36786 81524
rect 37461 81515 37519 81521
rect 37461 81481 37473 81515
rect 37507 81481 37519 81515
rect 37461 81475 37519 81481
rect 25590 81404 25596 81456
rect 25648 81444 25654 81456
rect 32306 81444 32312 81456
rect 25648 81416 32312 81444
rect 25648 81404 25654 81416
rect 32306 81404 32312 81416
rect 32364 81404 32370 81456
rect 37476 81444 37504 81475
rect 37476 81416 37596 81444
rect 15562 81336 15568 81388
rect 15620 81376 15626 81388
rect 33594 81376 33600 81388
rect 15620 81348 33600 81376
rect 15620 81336 15626 81348
rect 33594 81336 33600 81348
rect 33652 81336 33658 81388
rect 33962 81376 33968 81388
rect 33704 81348 33968 81376
rect 30834 81268 30840 81320
rect 30892 81308 30898 81320
rect 31570 81308 31576 81320
rect 30892 81280 31576 81308
rect 30892 81268 30898 81280
rect 31570 81268 31576 81280
rect 31628 81268 31634 81320
rect 31754 81268 31760 81320
rect 31812 81308 31818 81320
rect 32030 81308 32036 81320
rect 31812 81280 31857 81308
rect 31991 81280 32036 81308
rect 31812 81268 31818 81280
rect 32030 81268 32036 81280
rect 32088 81268 32094 81320
rect 32125 81311 32183 81317
rect 32125 81277 32137 81311
rect 32171 81277 32183 81311
rect 32398 81308 32404 81320
rect 32359 81280 32404 81308
rect 32125 81271 32183 81277
rect 31389 81175 31447 81181
rect 31389 81141 31401 81175
rect 31435 81172 31447 81175
rect 31570 81172 31576 81184
rect 31435 81144 31576 81172
rect 31435 81141 31447 81144
rect 31389 81135 31447 81141
rect 31570 81132 31576 81144
rect 31628 81132 31634 81184
rect 31754 81132 31760 81184
rect 31812 81172 31818 81184
rect 32140 81172 32168 81271
rect 32398 81268 32404 81280
rect 32456 81268 32462 81320
rect 33704 81317 33732 81348
rect 33962 81336 33968 81348
rect 34020 81336 34026 81388
rect 37458 81376 37464 81388
rect 34624 81348 37464 81376
rect 32677 81311 32735 81317
rect 32677 81277 32689 81311
rect 32723 81277 32735 81311
rect 32677 81271 32735 81277
rect 33689 81311 33747 81317
rect 33689 81277 33701 81311
rect 33735 81277 33747 81311
rect 33689 81271 33747 81277
rect 32692 81240 32720 81271
rect 33778 81268 33784 81320
rect 33836 81308 33842 81320
rect 34054 81308 34060 81320
rect 33836 81280 33881 81308
rect 34015 81280 34060 81308
rect 33836 81268 33842 81280
rect 34054 81268 34060 81280
rect 34112 81268 34118 81320
rect 34146 81268 34152 81320
rect 34204 81308 34210 81320
rect 34624 81317 34652 81348
rect 37458 81336 37464 81348
rect 37516 81336 37522 81388
rect 37568 81376 37596 81416
rect 37642 81376 37648 81388
rect 37568 81348 37648 81376
rect 37642 81336 37648 81348
rect 37700 81336 37706 81388
rect 34333 81311 34391 81317
rect 34333 81308 34345 81311
rect 34204 81280 34345 81308
rect 34204 81268 34210 81280
rect 34333 81277 34345 81280
rect 34379 81277 34391 81311
rect 34333 81271 34391 81277
rect 34609 81311 34667 81317
rect 34609 81277 34621 81311
rect 34655 81277 34667 81311
rect 37274 81308 37280 81320
rect 37235 81280 37280 81308
rect 34609 81271 34667 81277
rect 37274 81268 37280 81280
rect 37332 81268 37338 81320
rect 37734 81268 37740 81320
rect 37792 81268 37798 81320
rect 37918 81308 37924 81320
rect 37879 81280 37924 81308
rect 37918 81268 37924 81280
rect 37976 81268 37982 81320
rect 37752 81240 37780 81268
rect 32692 81212 33548 81240
rect 33318 81172 33324 81184
rect 31812 81144 32168 81172
rect 33279 81144 33324 81172
rect 31812 81132 31818 81144
rect 33318 81132 33324 81144
rect 33376 81132 33382 81184
rect 33520 81172 33548 81212
rect 37476 81212 37780 81240
rect 37476 81172 37504 81212
rect 33520 81144 37504 81172
rect 38105 81175 38163 81181
rect 38105 81141 38117 81175
rect 38151 81172 38163 81175
rect 38286 81172 38292 81184
rect 38151 81144 38292 81172
rect 38151 81141 38163 81144
rect 38105 81135 38163 81141
rect 38286 81132 38292 81144
rect 38344 81132 38350 81184
rect 1104 81082 38824 81104
rect 1104 81030 19606 81082
rect 19658 81030 19670 81082
rect 19722 81030 19734 81082
rect 19786 81030 19798 81082
rect 19850 81030 38824 81082
rect 1104 81008 38824 81030
rect 26418 80928 26424 80980
rect 26476 80968 26482 80980
rect 33137 80971 33195 80977
rect 33137 80968 33149 80971
rect 26476 80940 33149 80968
rect 26476 80928 26482 80940
rect 33137 80937 33149 80940
rect 33183 80937 33195 80971
rect 33137 80931 33195 80937
rect 33594 80928 33600 80980
rect 33652 80968 33658 80980
rect 33652 80940 33916 80968
rect 33652 80928 33658 80940
rect 1394 80832 1400 80844
rect 1355 80804 1400 80832
rect 1394 80792 1400 80804
rect 1452 80792 1458 80844
rect 30834 80792 30840 80844
rect 30892 80832 30898 80844
rect 31113 80835 31171 80841
rect 31113 80832 31125 80835
rect 30892 80804 31125 80832
rect 30892 80792 30898 80804
rect 31113 80801 31125 80804
rect 31159 80801 31171 80835
rect 31113 80795 31171 80801
rect 31202 80792 31208 80844
rect 31260 80832 31266 80844
rect 31481 80835 31539 80841
rect 31260 80804 31305 80832
rect 31260 80792 31266 80804
rect 31481 80801 31493 80835
rect 31527 80801 31539 80835
rect 31481 80795 31539 80801
rect 31757 80835 31815 80841
rect 31757 80801 31769 80835
rect 31803 80801 31815 80835
rect 31757 80795 31815 80801
rect 31941 80835 31999 80841
rect 31941 80801 31953 80835
rect 31987 80832 31999 80835
rect 32125 80835 32183 80841
rect 32125 80832 32137 80835
rect 31987 80804 32137 80832
rect 31987 80801 31999 80804
rect 31941 80795 31999 80801
rect 32125 80801 32137 80804
rect 32171 80801 32183 80835
rect 32125 80795 32183 80801
rect 33505 80835 33563 80841
rect 33505 80801 33517 80835
rect 33551 80801 33563 80835
rect 33778 80832 33784 80844
rect 33739 80804 33784 80832
rect 33505 80795 33563 80801
rect 17494 80724 17500 80776
rect 17552 80764 17558 80776
rect 31496 80764 31524 80795
rect 17552 80736 31524 80764
rect 31772 80764 31800 80795
rect 32030 80764 32036 80776
rect 31772 80736 32036 80764
rect 17552 80724 17558 80736
rect 32030 80724 32036 80736
rect 32088 80764 32094 80776
rect 33520 80764 33548 80795
rect 33778 80792 33784 80804
rect 33836 80792 33842 80844
rect 33888 80841 33916 80940
rect 33962 80928 33968 80980
rect 34020 80968 34026 80980
rect 38746 80968 38752 80980
rect 34020 80940 38752 80968
rect 34020 80928 34026 80940
rect 38746 80928 38752 80940
rect 38804 80928 38810 80980
rect 33873 80835 33931 80841
rect 33873 80801 33885 80835
rect 33919 80801 33931 80835
rect 34146 80832 34152 80844
rect 34107 80804 34152 80832
rect 33873 80795 33931 80801
rect 34146 80792 34152 80804
rect 34204 80792 34210 80844
rect 34425 80835 34483 80841
rect 34425 80801 34437 80835
rect 34471 80832 34483 80835
rect 35894 80832 35900 80844
rect 34471 80804 35900 80832
rect 34471 80801 34483 80804
rect 34425 80795 34483 80801
rect 35894 80792 35900 80804
rect 35952 80792 35958 80844
rect 36906 80764 36912 80776
rect 32088 80736 33456 80764
rect 33520 80736 36912 80764
rect 32088 80724 32094 80736
rect 23750 80656 23756 80708
rect 23808 80696 23814 80708
rect 33318 80696 33324 80708
rect 23808 80668 33324 80696
rect 23808 80656 23814 80668
rect 33318 80656 33324 80668
rect 33376 80656 33382 80708
rect 33428 80696 33456 80736
rect 36906 80724 36912 80736
rect 36964 80724 36970 80776
rect 34146 80696 34152 80708
rect 33428 80668 34152 80696
rect 34146 80656 34152 80668
rect 34204 80656 34210 80708
rect 25498 80588 25504 80640
rect 25556 80628 25562 80640
rect 30745 80631 30803 80637
rect 30745 80628 30757 80631
rect 25556 80600 30757 80628
rect 25556 80588 25562 80600
rect 30745 80597 30757 80600
rect 30791 80597 30803 80631
rect 30745 80591 30803 80597
rect 32125 80631 32183 80637
rect 32125 80597 32137 80631
rect 32171 80628 32183 80631
rect 37826 80628 37832 80640
rect 32171 80600 37832 80628
rect 32171 80597 32183 80600
rect 32125 80591 32183 80597
rect 37826 80588 37832 80600
rect 37884 80588 37890 80640
rect 1104 80538 38824 80560
rect 1104 80486 4246 80538
rect 4298 80486 4310 80538
rect 4362 80486 4374 80538
rect 4426 80486 4438 80538
rect 4490 80486 34966 80538
rect 35018 80486 35030 80538
rect 35082 80486 35094 80538
rect 35146 80486 35158 80538
rect 35210 80486 38824 80538
rect 1104 80464 38824 80486
rect 31202 80384 31208 80436
rect 31260 80424 31266 80436
rect 33778 80424 33784 80436
rect 31260 80396 33784 80424
rect 31260 80384 31266 80396
rect 26206 80260 31800 80288
rect 1394 80220 1400 80232
rect 1355 80192 1400 80220
rect 1394 80180 1400 80192
rect 1452 80180 1458 80232
rect 16206 80180 16212 80232
rect 16264 80220 16270 80232
rect 26206 80220 26234 80260
rect 31772 80229 31800 80260
rect 31389 80223 31447 80229
rect 31389 80220 31401 80223
rect 16264 80192 26234 80220
rect 31220 80192 31401 80220
rect 16264 80180 16270 80192
rect 26786 80112 26792 80164
rect 26844 80152 26850 80164
rect 30929 80155 30987 80161
rect 30929 80152 30941 80155
rect 26844 80124 30941 80152
rect 26844 80112 26850 80124
rect 30929 80121 30941 80124
rect 30975 80121 30987 80155
rect 30929 80115 30987 80121
rect 31220 80084 31248 80192
rect 31389 80189 31401 80192
rect 31435 80189 31447 80223
rect 31389 80183 31447 80189
rect 31665 80223 31723 80229
rect 31665 80189 31677 80223
rect 31711 80189 31723 80223
rect 31665 80183 31723 80189
rect 31757 80223 31815 80229
rect 31757 80189 31769 80223
rect 31803 80189 31815 80223
rect 31757 80183 31815 80189
rect 31680 80152 31708 80183
rect 31864 80152 31892 80396
rect 33778 80384 33784 80396
rect 33836 80384 33842 80436
rect 37461 80359 37519 80365
rect 37461 80325 37473 80359
rect 37507 80356 37519 80359
rect 39850 80356 39856 80368
rect 37507 80328 39856 80356
rect 37507 80325 37519 80328
rect 37461 80319 37519 80325
rect 39850 80316 39856 80328
rect 39908 80316 39914 80368
rect 38194 80288 38200 80300
rect 32324 80260 38200 80288
rect 32030 80220 32036 80232
rect 31991 80192 32036 80220
rect 32030 80180 32036 80192
rect 32088 80180 32094 80232
rect 32324 80229 32352 80260
rect 38194 80248 38200 80260
rect 38252 80248 38258 80300
rect 32309 80223 32367 80229
rect 32309 80189 32321 80223
rect 32355 80189 32367 80223
rect 37274 80220 37280 80232
rect 37235 80192 37280 80220
rect 32309 80183 32367 80189
rect 37274 80180 37280 80192
rect 37332 80180 37338 80232
rect 37918 80220 37924 80232
rect 37879 80192 37924 80220
rect 37918 80180 37924 80192
rect 37976 80180 37982 80232
rect 31680 80124 31892 80152
rect 37090 80084 37096 80096
rect 31220 80056 37096 80084
rect 37090 80044 37096 80056
rect 37148 80044 37154 80096
rect 38105 80087 38163 80093
rect 38105 80053 38117 80087
rect 38151 80084 38163 80087
rect 39482 80084 39488 80096
rect 38151 80056 39488 80084
rect 38151 80053 38163 80056
rect 38105 80047 38163 80053
rect 39482 80044 39488 80056
rect 39540 80044 39546 80096
rect 1104 79994 38824 80016
rect 1104 79942 19606 79994
rect 19658 79942 19670 79994
rect 19722 79942 19734 79994
rect 19786 79942 19798 79994
rect 19850 79942 38824 79994
rect 1104 79920 38824 79942
rect 30742 79840 30748 79892
rect 30800 79880 30806 79892
rect 37182 79880 37188 79892
rect 30800 79852 37188 79880
rect 30800 79840 30806 79852
rect 37182 79840 37188 79852
rect 37240 79840 37246 79892
rect 1394 79744 1400 79756
rect 1355 79716 1400 79744
rect 1394 79704 1400 79716
rect 1452 79704 1458 79756
rect 14826 79744 14832 79756
rect 14787 79716 14832 79744
rect 14826 79704 14832 79716
rect 14884 79704 14890 79756
rect 37182 79744 37188 79756
rect 37143 79716 37188 79744
rect 37182 79704 37188 79716
rect 37240 79704 37246 79756
rect 2590 79500 2596 79552
rect 2648 79540 2654 79552
rect 15013 79543 15071 79549
rect 15013 79540 15025 79543
rect 2648 79512 15025 79540
rect 2648 79500 2654 79512
rect 15013 79509 15025 79512
rect 15059 79509 15071 79543
rect 15013 79503 15071 79509
rect 17126 79500 17132 79552
rect 17184 79540 17190 79552
rect 33870 79540 33876 79552
rect 17184 79512 33876 79540
rect 17184 79500 17190 79512
rect 33870 79500 33876 79512
rect 33928 79500 33934 79552
rect 37369 79543 37427 79549
rect 37369 79509 37381 79543
rect 37415 79540 37427 79543
rect 38562 79540 38568 79552
rect 37415 79512 38568 79540
rect 37415 79509 37427 79512
rect 37369 79503 37427 79509
rect 38562 79500 38568 79512
rect 38620 79500 38626 79552
rect 1104 79450 38824 79472
rect 1104 79398 4246 79450
rect 4298 79398 4310 79450
rect 4362 79398 4374 79450
rect 4426 79398 4438 79450
rect 4490 79398 34966 79450
rect 35018 79398 35030 79450
rect 35082 79398 35094 79450
rect 35146 79398 35158 79450
rect 35210 79398 38824 79450
rect 1104 79376 38824 79398
rect 16298 79296 16304 79348
rect 16356 79336 16362 79348
rect 34054 79336 34060 79348
rect 16356 79308 34060 79336
rect 16356 79296 16362 79308
rect 34054 79296 34060 79308
rect 34112 79296 34118 79348
rect 37461 79271 37519 79277
rect 37461 79237 37473 79271
rect 37507 79268 37519 79271
rect 38746 79268 38752 79280
rect 37507 79240 38752 79268
rect 37507 79237 37519 79240
rect 37461 79231 37519 79237
rect 38746 79228 38752 79240
rect 38804 79228 38810 79280
rect 37274 79132 37280 79144
rect 37235 79104 37280 79132
rect 37274 79092 37280 79104
rect 37332 79092 37338 79144
rect 37918 79132 37924 79144
rect 37879 79104 37924 79132
rect 37918 79092 37924 79104
rect 37976 79092 37982 79144
rect 38105 78999 38163 79005
rect 38105 78965 38117 78999
rect 38151 78996 38163 78999
rect 39114 78996 39120 79008
rect 38151 78968 39120 78996
rect 38151 78965 38163 78968
rect 38105 78959 38163 78965
rect 39114 78956 39120 78968
rect 39172 78956 39178 79008
rect 1104 78906 38824 78928
rect 1104 78854 19606 78906
rect 19658 78854 19670 78906
rect 19722 78854 19734 78906
rect 19786 78854 19798 78906
rect 19850 78854 38824 78906
rect 1104 78832 38824 78854
rect 1394 78656 1400 78668
rect 1355 78628 1400 78656
rect 1394 78616 1400 78628
rect 1452 78616 1458 78668
rect 26970 78616 26976 78668
rect 27028 78656 27034 78668
rect 27801 78659 27859 78665
rect 27801 78656 27813 78659
rect 27028 78628 27813 78656
rect 27028 78616 27034 78628
rect 27801 78625 27813 78628
rect 27847 78625 27859 78659
rect 27801 78619 27859 78625
rect 27985 78455 28043 78461
rect 27985 78421 27997 78455
rect 28031 78452 28043 78455
rect 30834 78452 30840 78464
rect 28031 78424 30840 78452
rect 28031 78421 28043 78424
rect 27985 78415 28043 78421
rect 30834 78412 30840 78424
rect 30892 78412 30898 78464
rect 1104 78362 38824 78384
rect 1104 78310 4246 78362
rect 4298 78310 4310 78362
rect 4362 78310 4374 78362
rect 4426 78310 4438 78362
rect 4490 78310 34966 78362
rect 35018 78310 35030 78362
rect 35082 78310 35094 78362
rect 35146 78310 35158 78362
rect 35210 78310 38824 78362
rect 1104 78288 38824 78310
rect 37461 78183 37519 78189
rect 37461 78149 37473 78183
rect 37507 78180 37519 78183
rect 39298 78180 39304 78192
rect 37507 78152 39304 78180
rect 37507 78149 37519 78152
rect 37461 78143 37519 78149
rect 39298 78140 39304 78152
rect 39356 78140 39362 78192
rect 1394 78044 1400 78056
rect 1355 78016 1400 78044
rect 1394 78004 1400 78016
rect 1452 78004 1458 78056
rect 32401 78047 32459 78053
rect 32401 78013 32413 78047
rect 32447 78044 32459 78047
rect 32490 78044 32496 78056
rect 32447 78016 32496 78044
rect 32447 78013 32459 78016
rect 32401 78007 32459 78013
rect 32490 78004 32496 78016
rect 32548 78004 32554 78056
rect 37274 78044 37280 78056
rect 37235 78016 37280 78044
rect 37274 78004 37280 78016
rect 37332 78004 37338 78056
rect 37918 78044 37924 78056
rect 37879 78016 37924 78044
rect 37918 78004 37924 78016
rect 37976 78004 37982 78056
rect 16390 77936 16396 77988
rect 16448 77976 16454 77988
rect 31754 77976 31760 77988
rect 16448 77948 31760 77976
rect 16448 77936 16454 77948
rect 31754 77936 31760 77948
rect 31812 77936 31818 77988
rect 32490 77868 32496 77920
rect 32548 77908 32554 77920
rect 32585 77911 32643 77917
rect 32585 77908 32597 77911
rect 32548 77880 32597 77908
rect 32548 77868 32554 77880
rect 32585 77877 32597 77880
rect 32631 77877 32643 77911
rect 32585 77871 32643 77877
rect 38105 77911 38163 77917
rect 38105 77877 38117 77911
rect 38151 77908 38163 77911
rect 38194 77908 38200 77920
rect 38151 77880 38200 77908
rect 38151 77877 38163 77880
rect 38105 77871 38163 77877
rect 38194 77868 38200 77880
rect 38252 77868 38258 77920
rect 1104 77818 38824 77840
rect 1104 77766 19606 77818
rect 19658 77766 19670 77818
rect 19722 77766 19734 77818
rect 19786 77766 19798 77818
rect 19850 77766 38824 77818
rect 1104 77744 38824 77766
rect 33042 77324 33048 77376
rect 33100 77364 33106 77376
rect 36262 77364 36268 77376
rect 33100 77336 36268 77364
rect 33100 77324 33106 77336
rect 36262 77324 36268 77336
rect 36320 77324 36326 77376
rect 1104 77274 38824 77296
rect 1104 77222 4246 77274
rect 4298 77222 4310 77274
rect 4362 77222 4374 77274
rect 4426 77222 4438 77274
rect 4490 77222 34966 77274
rect 35018 77222 35030 77274
rect 35082 77222 35094 77274
rect 35146 77222 35158 77274
rect 35210 77222 38824 77274
rect 1104 77200 38824 77222
rect 1394 76956 1400 76968
rect 1355 76928 1400 76956
rect 1394 76916 1400 76928
rect 1452 76916 1458 76968
rect 37274 76956 37280 76968
rect 37235 76928 37280 76956
rect 37274 76916 37280 76928
rect 37332 76916 37338 76968
rect 37921 76959 37979 76965
rect 37921 76925 37933 76959
rect 37967 76956 37979 76959
rect 38010 76956 38016 76968
rect 37967 76928 38016 76956
rect 37967 76925 37979 76928
rect 37921 76919 37979 76925
rect 38010 76916 38016 76928
rect 38068 76916 38074 76968
rect 29914 76848 29920 76900
rect 29972 76888 29978 76900
rect 30926 76888 30932 76900
rect 29972 76860 30932 76888
rect 29972 76848 29978 76860
rect 30926 76848 30932 76860
rect 30984 76848 30990 76900
rect 37461 76823 37519 76829
rect 37461 76789 37473 76823
rect 37507 76820 37519 76823
rect 37642 76820 37648 76832
rect 37507 76792 37648 76820
rect 37507 76789 37519 76792
rect 37461 76783 37519 76789
rect 37642 76780 37648 76792
rect 37700 76780 37706 76832
rect 37826 76780 37832 76832
rect 37884 76820 37890 76832
rect 38105 76823 38163 76829
rect 38105 76820 38117 76823
rect 37884 76792 38117 76820
rect 37884 76780 37890 76792
rect 38105 76789 38117 76792
rect 38151 76789 38163 76823
rect 38105 76783 38163 76789
rect 1104 76730 38824 76752
rect 1104 76678 19606 76730
rect 19658 76678 19670 76730
rect 19722 76678 19734 76730
rect 19786 76678 19798 76730
rect 19850 76678 38824 76730
rect 1104 76656 38824 76678
rect 31018 76576 31024 76628
rect 31076 76616 31082 76628
rect 31113 76619 31171 76625
rect 31113 76616 31125 76619
rect 31076 76588 31125 76616
rect 31076 76576 31082 76588
rect 31113 76585 31125 76588
rect 31159 76585 31171 76619
rect 31113 76579 31171 76585
rect 23474 76548 23480 76560
rect 23435 76520 23480 76548
rect 23474 76508 23480 76520
rect 23532 76508 23538 76560
rect 1394 76480 1400 76492
rect 1355 76452 1400 76480
rect 1394 76440 1400 76452
rect 1452 76440 1458 76492
rect 23106 76440 23112 76492
rect 23164 76480 23170 76492
rect 30929 76483 30987 76489
rect 30929 76480 30941 76483
rect 23164 76452 30941 76480
rect 23164 76440 23170 76452
rect 30929 76449 30941 76452
rect 30975 76449 30987 76483
rect 30929 76443 30987 76449
rect 23661 76347 23719 76353
rect 23661 76313 23673 76347
rect 23707 76344 23719 76347
rect 23842 76344 23848 76356
rect 23707 76316 23848 76344
rect 23707 76313 23719 76316
rect 23661 76307 23719 76313
rect 23842 76304 23848 76316
rect 23900 76304 23906 76356
rect 1104 76186 38824 76208
rect 1104 76134 4246 76186
rect 4298 76134 4310 76186
rect 4362 76134 4374 76186
rect 4426 76134 4438 76186
rect 4490 76134 34966 76186
rect 35018 76134 35030 76186
rect 35082 76134 35094 76186
rect 35146 76134 35158 76186
rect 35210 76134 38824 76186
rect 1104 76112 38824 76134
rect 33778 75964 33784 76016
rect 33836 76004 33842 76016
rect 38378 76004 38384 76016
rect 33836 75976 38384 76004
rect 33836 75964 33842 75976
rect 38378 75964 38384 75976
rect 38436 75964 38442 76016
rect 35250 75896 35256 75948
rect 35308 75936 35314 75948
rect 39206 75936 39212 75948
rect 35308 75908 39212 75936
rect 35308 75896 35314 75908
rect 39206 75896 39212 75908
rect 39264 75896 39270 75948
rect 20070 75868 20076 75880
rect 20031 75840 20076 75868
rect 20070 75828 20076 75840
rect 20128 75828 20134 75880
rect 20165 75871 20223 75877
rect 20165 75837 20177 75871
rect 20211 75837 20223 75871
rect 20165 75831 20223 75837
rect 20349 75871 20407 75877
rect 20349 75837 20361 75871
rect 20395 75868 20407 75871
rect 20530 75868 20536 75880
rect 20395 75840 20536 75868
rect 20395 75837 20407 75840
rect 20349 75831 20407 75837
rect 9030 75760 9036 75812
rect 9088 75800 9094 75812
rect 20180 75800 20208 75831
rect 20530 75828 20536 75840
rect 20588 75828 20594 75880
rect 37274 75868 37280 75880
rect 37235 75840 37280 75868
rect 37274 75828 37280 75840
rect 37332 75828 37338 75880
rect 37918 75868 37924 75880
rect 37879 75840 37924 75868
rect 37918 75828 37924 75840
rect 37976 75828 37982 75880
rect 39758 75800 39764 75812
rect 9088 75772 20208 75800
rect 37476 75772 39764 75800
rect 9088 75760 9094 75772
rect 37476 75741 37504 75772
rect 39758 75760 39764 75772
rect 39816 75760 39822 75812
rect 37461 75735 37519 75741
rect 37461 75701 37473 75735
rect 37507 75701 37519 75735
rect 37461 75695 37519 75701
rect 38105 75735 38163 75741
rect 38105 75701 38117 75735
rect 38151 75732 38163 75735
rect 38654 75732 38660 75744
rect 38151 75704 38660 75732
rect 38151 75701 38163 75704
rect 38105 75695 38163 75701
rect 38654 75692 38660 75704
rect 38712 75692 38718 75744
rect 1104 75642 38824 75664
rect 1104 75590 19606 75642
rect 19658 75590 19670 75642
rect 19722 75590 19734 75642
rect 19786 75590 19798 75642
rect 19850 75590 38824 75642
rect 1104 75568 38824 75590
rect 20349 75531 20407 75537
rect 20349 75497 20361 75531
rect 20395 75528 20407 75531
rect 20438 75528 20444 75540
rect 20395 75500 20444 75528
rect 20395 75497 20407 75500
rect 20349 75491 20407 75497
rect 20438 75488 20444 75500
rect 20496 75488 20502 75540
rect 21174 75528 21180 75540
rect 21135 75500 21180 75528
rect 21174 75488 21180 75500
rect 21232 75488 21238 75540
rect 29546 75488 29552 75540
rect 29604 75528 29610 75540
rect 29641 75531 29699 75537
rect 29641 75528 29653 75531
rect 29604 75500 29653 75528
rect 29604 75488 29610 75500
rect 29641 75497 29653 75500
rect 29687 75497 29699 75531
rect 29641 75491 29699 75497
rect 29748 75500 30144 75528
rect 23842 75460 23848 75472
rect 20824 75432 23848 75460
rect 1394 75392 1400 75404
rect 1355 75364 1400 75392
rect 1394 75352 1400 75364
rect 1452 75352 1458 75404
rect 10318 75352 10324 75404
rect 10376 75392 10382 75404
rect 20824 75401 20852 75432
rect 23842 75420 23848 75432
rect 23900 75460 23906 75472
rect 29748 75460 29776 75500
rect 23900 75432 29776 75460
rect 23900 75420 23906 75432
rect 20165 75395 20223 75401
rect 20165 75392 20177 75395
rect 10376 75364 20177 75392
rect 10376 75352 10382 75364
rect 20165 75361 20177 75364
rect 20211 75361 20223 75395
rect 20165 75355 20223 75361
rect 20809 75395 20867 75401
rect 20809 75361 20821 75395
rect 20855 75361 20867 75395
rect 20990 75392 20996 75404
rect 20951 75364 20996 75392
rect 20809 75355 20867 75361
rect 19981 75327 20039 75333
rect 19981 75293 19993 75327
rect 20027 75324 20039 75327
rect 20070 75324 20076 75336
rect 20027 75296 20076 75324
rect 20027 75293 20039 75296
rect 19981 75287 20039 75293
rect 20070 75284 20076 75296
rect 20128 75324 20134 75336
rect 20824 75324 20852 75355
rect 20990 75352 20996 75364
rect 21048 75352 21054 75404
rect 29457 75395 29515 75401
rect 29457 75361 29469 75395
rect 29503 75361 29515 75395
rect 29638 75392 29644 75404
rect 29599 75364 29644 75392
rect 29457 75355 29515 75361
rect 20128 75296 20852 75324
rect 29472 75324 29500 75355
rect 29638 75352 29644 75364
rect 29696 75352 29702 75404
rect 29914 75392 29920 75404
rect 29875 75364 29920 75392
rect 29914 75352 29920 75364
rect 29972 75352 29978 75404
rect 30116 75401 30144 75500
rect 32030 75488 32036 75540
rect 32088 75528 32094 75540
rect 34514 75528 34520 75540
rect 32088 75500 34520 75528
rect 32088 75488 32094 75500
rect 34514 75488 34520 75500
rect 34572 75488 34578 75540
rect 30101 75395 30159 75401
rect 30101 75361 30113 75395
rect 30147 75361 30159 75395
rect 37182 75392 37188 75404
rect 37143 75364 37188 75392
rect 30101 75355 30159 75361
rect 37182 75352 37188 75364
rect 37240 75352 37246 75404
rect 35894 75324 35900 75336
rect 29472 75296 35900 75324
rect 20128 75284 20134 75296
rect 35894 75284 35900 75296
rect 35952 75284 35958 75336
rect 32306 75216 32312 75268
rect 32364 75256 32370 75268
rect 32950 75256 32956 75268
rect 32364 75228 32956 75256
rect 32364 75216 32370 75228
rect 32950 75216 32956 75228
rect 33008 75216 33014 75268
rect 33870 75216 33876 75268
rect 33928 75256 33934 75268
rect 38930 75256 38936 75268
rect 33928 75228 38936 75256
rect 33928 75216 33934 75228
rect 38930 75216 38936 75228
rect 38988 75216 38994 75268
rect 39390 75216 39396 75268
rect 39448 75256 39454 75268
rect 39574 75256 39580 75268
rect 39448 75228 39580 75256
rect 39448 75216 39454 75228
rect 39574 75216 39580 75228
rect 39632 75216 39638 75268
rect 36262 75148 36268 75200
rect 36320 75188 36326 75200
rect 37369 75191 37427 75197
rect 37369 75188 37381 75191
rect 36320 75160 37381 75188
rect 36320 75148 36326 75160
rect 37369 75157 37381 75160
rect 37415 75157 37427 75191
rect 37369 75151 37427 75157
rect 39209 75123 39267 75129
rect 1104 75098 38824 75120
rect 1104 75046 4246 75098
rect 4298 75046 4310 75098
rect 4362 75046 4374 75098
rect 4426 75046 4438 75098
rect 4490 75046 34966 75098
rect 35018 75046 35030 75098
rect 35082 75046 35094 75098
rect 35146 75046 35158 75098
rect 35210 75046 38824 75098
rect 39209 75089 39221 75123
rect 39255 75120 39267 75123
rect 39666 75120 39672 75132
rect 39255 75092 39672 75120
rect 39255 75089 39267 75092
rect 39209 75083 39267 75089
rect 39666 75080 39672 75092
rect 39724 75080 39730 75132
rect 1104 75024 38824 75046
rect 39298 75012 39304 75064
rect 39356 75052 39362 75064
rect 39393 75055 39451 75061
rect 39393 75052 39405 75055
rect 39356 75024 39405 75052
rect 39356 75012 39362 75024
rect 39393 75021 39405 75024
rect 39439 75021 39451 75055
rect 39393 75015 39451 75021
rect 20346 74984 20352 74996
rect 20307 74956 20352 74984
rect 20346 74944 20352 74956
rect 20404 74944 20410 74996
rect 32950 74944 32956 74996
rect 33008 74984 33014 74996
rect 36354 74984 36360 74996
rect 33008 74956 36360 74984
rect 33008 74944 33014 74956
rect 36354 74944 36360 74956
rect 36412 74944 36418 74996
rect 38286 74944 38292 74996
rect 38344 74984 38350 74996
rect 39666 74984 39672 74996
rect 38344 74956 39672 74984
rect 38344 74944 38350 74956
rect 39666 74944 39672 74956
rect 39724 74944 39730 74996
rect 37461 74919 37519 74925
rect 37461 74885 37473 74919
rect 37507 74916 37519 74919
rect 39301 74919 39359 74925
rect 39301 74916 39313 74919
rect 37507 74888 39313 74916
rect 37507 74885 37519 74888
rect 37461 74879 37519 74885
rect 39301 74885 39313 74888
rect 39347 74885 39359 74919
rect 39301 74879 39359 74885
rect 19981 74851 20039 74857
rect 19981 74817 19993 74851
rect 20027 74848 20039 74851
rect 20070 74848 20076 74860
rect 20027 74820 20076 74848
rect 20027 74817 20039 74820
rect 19981 74811 20039 74817
rect 20070 74808 20076 74820
rect 20128 74808 20134 74860
rect 1394 74780 1400 74792
rect 1355 74752 1400 74780
rect 1394 74740 1400 74752
rect 1452 74740 1458 74792
rect 20165 74783 20223 74789
rect 20165 74749 20177 74783
rect 20211 74749 20223 74783
rect 37274 74780 37280 74792
rect 37235 74752 37280 74780
rect 20165 74743 20223 74749
rect 14550 74672 14556 74724
rect 14608 74712 14614 74724
rect 20180 74712 20208 74743
rect 37274 74740 37280 74752
rect 37332 74740 37338 74792
rect 37918 74780 37924 74792
rect 37879 74752 37924 74780
rect 37918 74740 37924 74752
rect 37976 74740 37982 74792
rect 14608 74684 20208 74712
rect 14608 74672 14614 74684
rect 35618 74604 35624 74656
rect 35676 74644 35682 74656
rect 38105 74647 38163 74653
rect 38105 74644 38117 74647
rect 35676 74616 38117 74644
rect 35676 74604 35682 74616
rect 38105 74613 38117 74616
rect 38151 74613 38163 74647
rect 38105 74607 38163 74613
rect 1104 74554 38824 74576
rect 1104 74502 19606 74554
rect 19658 74502 19670 74554
rect 19722 74502 19734 74554
rect 19786 74502 19798 74554
rect 19850 74502 38824 74554
rect 1104 74480 38824 74502
rect 34054 74400 34060 74452
rect 34112 74440 34118 74452
rect 38838 74440 38844 74452
rect 34112 74412 38844 74440
rect 34112 74400 34118 74412
rect 38838 74400 38844 74412
rect 38896 74400 38902 74452
rect 37182 74304 37188 74316
rect 37143 74276 37188 74304
rect 37182 74264 37188 74276
rect 37240 74264 37246 74316
rect 37369 74103 37427 74109
rect 37369 74069 37381 74103
rect 37415 74100 37427 74103
rect 38838 74100 38844 74112
rect 37415 74072 38844 74100
rect 37415 74069 37427 74072
rect 37369 74063 37427 74069
rect 38838 74060 38844 74072
rect 38896 74060 38902 74112
rect 1104 74010 38824 74032
rect 1104 73958 4246 74010
rect 4298 73958 4310 74010
rect 4362 73958 4374 74010
rect 4426 73958 4438 74010
rect 4490 73958 34966 74010
rect 35018 73958 35030 74010
rect 35082 73958 35094 74010
rect 35146 73958 35158 74010
rect 35210 73958 38824 74010
rect 1104 73936 38824 73958
rect 16114 73788 16120 73840
rect 16172 73828 16178 73840
rect 25590 73828 25596 73840
rect 16172 73800 25596 73828
rect 16172 73788 16178 73800
rect 25590 73788 25596 73800
rect 25648 73788 25654 73840
rect 37090 73788 37096 73840
rect 37148 73828 37154 73840
rect 38105 73831 38163 73837
rect 38105 73828 38117 73831
rect 37148 73800 38117 73828
rect 37148 73788 37154 73800
rect 38105 73797 38117 73800
rect 38151 73797 38163 73831
rect 38105 73791 38163 73797
rect 1394 73692 1400 73704
rect 1355 73664 1400 73692
rect 1394 73652 1400 73664
rect 1452 73652 1458 73704
rect 20073 73695 20131 73701
rect 20073 73661 20085 73695
rect 20119 73692 20131 73695
rect 20162 73692 20168 73704
rect 20119 73664 20168 73692
rect 20119 73661 20131 73664
rect 20073 73655 20131 73661
rect 20162 73652 20168 73664
rect 20220 73692 20226 73704
rect 20717 73695 20775 73701
rect 20717 73692 20729 73695
rect 20220 73664 20729 73692
rect 20220 73652 20226 73664
rect 20717 73661 20729 73664
rect 20763 73692 20775 73695
rect 23474 73692 23480 73704
rect 20763 73664 23480 73692
rect 20763 73661 20775 73664
rect 20717 73655 20775 73661
rect 23474 73652 23480 73664
rect 23532 73652 23538 73704
rect 37274 73692 37280 73704
rect 37235 73664 37280 73692
rect 37274 73652 37280 73664
rect 37332 73652 37338 73704
rect 37918 73692 37924 73704
rect 37879 73664 37924 73692
rect 37918 73652 37924 73664
rect 37976 73652 37982 73704
rect 17310 73584 17316 73636
rect 17368 73624 17374 73636
rect 17368 73596 20944 73624
rect 17368 73584 17374 73596
rect 17402 73516 17408 73568
rect 17460 73556 17466 73568
rect 20916 73565 20944 73596
rect 20257 73559 20315 73565
rect 20257 73556 20269 73559
rect 17460 73528 20269 73556
rect 17460 73516 17466 73528
rect 20257 73525 20269 73528
rect 20303 73525 20315 73559
rect 20257 73519 20315 73525
rect 20901 73559 20959 73565
rect 20901 73525 20913 73559
rect 20947 73525 20959 73559
rect 20901 73519 20959 73525
rect 36170 73516 36176 73568
rect 36228 73556 36234 73568
rect 37461 73559 37519 73565
rect 37461 73556 37473 73559
rect 36228 73528 37473 73556
rect 36228 73516 36234 73528
rect 37461 73525 37473 73528
rect 37507 73525 37519 73559
rect 37461 73519 37519 73525
rect 1104 73466 38824 73488
rect 1104 73414 19606 73466
rect 19658 73414 19670 73466
rect 19722 73414 19734 73466
rect 19786 73414 19798 73466
rect 19850 73414 38824 73466
rect 1104 73392 38824 73414
rect 1394 73216 1400 73228
rect 1355 73188 1400 73216
rect 1394 73176 1400 73188
rect 1452 73176 1458 73228
rect 32398 73108 32404 73160
rect 32456 73148 32462 73160
rect 34790 73148 34796 73160
rect 32456 73120 34796 73148
rect 32456 73108 32462 73120
rect 34790 73108 34796 73120
rect 34848 73108 34854 73160
rect 34330 73040 34336 73092
rect 34388 73080 34394 73092
rect 36998 73080 37004 73092
rect 34388 73052 37004 73080
rect 34388 73040 34394 73052
rect 36998 73040 37004 73052
rect 37056 73040 37062 73092
rect 37734 72972 37740 73024
rect 37792 73012 37798 73024
rect 37918 73012 37924 73024
rect 37792 72984 37924 73012
rect 37792 72972 37798 72984
rect 37918 72972 37924 72984
rect 37976 72972 37982 73024
rect 1104 72922 38824 72944
rect 1104 72870 4246 72922
rect 4298 72870 4310 72922
rect 4362 72870 4374 72922
rect 4426 72870 4438 72922
rect 4490 72870 34966 72922
rect 35018 72870 35030 72922
rect 35082 72870 35094 72922
rect 35146 72870 35158 72922
rect 35210 72870 38824 72922
rect 1104 72848 38824 72870
rect 16114 72808 16120 72820
rect 16075 72780 16120 72808
rect 16114 72768 16120 72780
rect 16172 72768 16178 72820
rect 16942 72808 16948 72820
rect 16903 72780 16948 72808
rect 16942 72768 16948 72780
rect 17000 72768 17006 72820
rect 17773 72811 17831 72817
rect 17773 72777 17785 72811
rect 17819 72808 17831 72811
rect 17862 72808 17868 72820
rect 17819 72780 17868 72808
rect 17819 72777 17831 72780
rect 17773 72771 17831 72777
rect 17862 72768 17868 72780
rect 17920 72768 17926 72820
rect 17310 72740 17316 72752
rect 15764 72712 17316 72740
rect 15764 72681 15792 72712
rect 17310 72700 17316 72712
rect 17368 72700 17374 72752
rect 15749 72675 15807 72681
rect 15749 72641 15761 72675
rect 15795 72641 15807 72675
rect 15749 72635 15807 72641
rect 16577 72675 16635 72681
rect 16577 72641 16589 72675
rect 16623 72672 16635 72675
rect 17402 72672 17408 72684
rect 16623 72644 17408 72672
rect 16623 72641 16635 72644
rect 16577 72635 16635 72641
rect 17402 72632 17408 72644
rect 17460 72632 17466 72684
rect 15930 72604 15936 72616
rect 15891 72576 15936 72604
rect 15930 72564 15936 72576
rect 15988 72564 15994 72616
rect 16761 72607 16819 72613
rect 16761 72573 16773 72607
rect 16807 72604 16819 72607
rect 17034 72604 17040 72616
rect 16807 72576 17040 72604
rect 16807 72573 16819 72576
rect 16761 72567 16819 72573
rect 17034 72564 17040 72576
rect 17092 72564 17098 72616
rect 17589 72607 17647 72613
rect 17589 72573 17601 72607
rect 17635 72573 17647 72607
rect 17589 72567 17647 72573
rect 19981 72607 20039 72613
rect 19981 72573 19993 72607
rect 20027 72604 20039 72607
rect 20162 72604 20168 72616
rect 20027 72576 20168 72604
rect 20027 72573 20039 72576
rect 19981 72567 20039 72573
rect 16942 72496 16948 72548
rect 17000 72536 17006 72548
rect 17604 72536 17632 72567
rect 20162 72564 20168 72576
rect 20220 72564 20226 72616
rect 37274 72604 37280 72616
rect 37235 72576 37280 72604
rect 37274 72564 37280 72576
rect 37332 72564 37338 72616
rect 37921 72607 37979 72613
rect 37921 72573 37933 72607
rect 37967 72604 37979 72607
rect 38933 72607 38991 72613
rect 38933 72604 38945 72607
rect 37967 72576 38945 72604
rect 37967 72573 37979 72576
rect 37921 72567 37979 72573
rect 38933 72573 38945 72576
rect 38979 72573 38991 72607
rect 38933 72567 38991 72573
rect 17000 72508 17632 72536
rect 17000 72496 17006 72508
rect 17218 72428 17224 72480
rect 17276 72468 17282 72480
rect 20165 72471 20223 72477
rect 20165 72468 20177 72471
rect 17276 72440 20177 72468
rect 17276 72428 17282 72440
rect 20165 72437 20177 72440
rect 20211 72437 20223 72471
rect 20165 72431 20223 72437
rect 36354 72428 36360 72480
rect 36412 72468 36418 72480
rect 37461 72471 37519 72477
rect 37461 72468 37473 72471
rect 36412 72440 37473 72468
rect 36412 72428 36418 72440
rect 37461 72437 37473 72440
rect 37507 72437 37519 72471
rect 37461 72431 37519 72437
rect 38105 72471 38163 72477
rect 38105 72437 38117 72471
rect 38151 72468 38163 72471
rect 38378 72468 38384 72480
rect 38151 72440 38384 72468
rect 38151 72437 38163 72440
rect 38105 72431 38163 72437
rect 38378 72428 38384 72440
rect 38436 72428 38442 72480
rect 1104 72378 38824 72400
rect 1104 72326 19606 72378
rect 19658 72326 19670 72378
rect 19722 72326 19734 72378
rect 19786 72326 19798 72378
rect 19850 72326 38824 72378
rect 1104 72304 38824 72326
rect 16393 72267 16451 72273
rect 16393 72233 16405 72267
rect 16439 72264 16451 72267
rect 16482 72264 16488 72276
rect 16439 72236 16488 72264
rect 16439 72233 16451 72236
rect 16393 72227 16451 72233
rect 16482 72224 16488 72236
rect 16540 72224 16546 72276
rect 17678 72264 17684 72276
rect 17639 72236 17684 72264
rect 17678 72224 17684 72236
rect 17736 72224 17742 72276
rect 17129 72199 17187 72205
rect 17129 72196 17141 72199
rect 6886 72168 17141 72196
rect 1394 72128 1400 72140
rect 1355 72100 1400 72128
rect 1394 72088 1400 72100
rect 1452 72088 1458 72140
rect 2222 72088 2228 72140
rect 2280 72128 2286 72140
rect 6886 72128 6914 72168
rect 17129 72165 17141 72168
rect 17175 72196 17187 72199
rect 17175 72168 17540 72196
rect 17175 72165 17187 72168
rect 17129 72159 17187 72165
rect 2280 72100 6914 72128
rect 2280 72088 2286 72100
rect 8938 72088 8944 72140
rect 8996 72128 9002 72140
rect 16209 72131 16267 72137
rect 16209 72128 16221 72131
rect 8996 72100 16221 72128
rect 8996 72088 9002 72100
rect 16209 72097 16221 72100
rect 16255 72097 16267 72131
rect 17402 72128 17408 72140
rect 17363 72100 17408 72128
rect 16209 72091 16267 72097
rect 17402 72088 17408 72100
rect 17460 72088 17466 72140
rect 17512 72137 17540 72168
rect 17497 72131 17555 72137
rect 17497 72097 17509 72131
rect 17543 72097 17555 72131
rect 37182 72128 37188 72140
rect 37143 72100 37188 72128
rect 17497 72091 17555 72097
rect 37182 72088 37188 72100
rect 37240 72088 37246 72140
rect 16025 72063 16083 72069
rect 16025 72029 16037 72063
rect 16071 72060 16083 72063
rect 16574 72060 16580 72072
rect 16071 72032 16580 72060
rect 16071 72029 16083 72032
rect 16025 72023 16083 72029
rect 16574 72020 16580 72032
rect 16632 72060 16638 72072
rect 17420 72060 17448 72088
rect 16632 72032 17448 72060
rect 16632 72020 16638 72032
rect 36906 71884 36912 71936
rect 36964 71924 36970 71936
rect 37369 71927 37427 71933
rect 37369 71924 37381 71927
rect 36964 71896 37381 71924
rect 36964 71884 36970 71896
rect 37369 71893 37381 71896
rect 37415 71893 37427 71927
rect 37369 71887 37427 71893
rect 1104 71834 38824 71856
rect 1104 71782 4246 71834
rect 4298 71782 4310 71834
rect 4362 71782 4374 71834
rect 4426 71782 4438 71834
rect 4490 71782 34966 71834
rect 35018 71782 35030 71834
rect 35082 71782 35094 71834
rect 35146 71782 35158 71834
rect 35210 71782 38824 71834
rect 38930 71788 38936 71800
rect 1104 71760 38824 71782
rect 38891 71760 38936 71788
rect 38930 71748 38936 71760
rect 38988 71748 38994 71800
rect 16850 71720 16856 71732
rect 15764 71692 16856 71720
rect 15764 71593 15792 71692
rect 16850 71680 16856 71692
rect 16908 71680 16914 71732
rect 16945 71723 17003 71729
rect 16945 71689 16957 71723
rect 16991 71720 17003 71723
rect 17126 71720 17132 71732
rect 16991 71692 17132 71720
rect 16991 71689 17003 71692
rect 16945 71683 17003 71689
rect 17126 71680 17132 71692
rect 17184 71680 17190 71732
rect 17770 71720 17776 71732
rect 17731 71692 17776 71720
rect 17770 71680 17776 71692
rect 17828 71680 17834 71732
rect 35894 71720 35900 71732
rect 35855 71692 35900 71720
rect 35894 71680 35900 71692
rect 35952 71680 35958 71732
rect 16022 71612 16028 71664
rect 16080 71652 16086 71664
rect 16117 71655 16175 71661
rect 16117 71652 16129 71655
rect 16080 71624 16129 71652
rect 16080 71612 16086 71624
rect 16117 71621 16129 71624
rect 16163 71621 16175 71655
rect 17862 71652 17868 71664
rect 16117 71615 16175 71621
rect 16776 71624 17868 71652
rect 15749 71587 15807 71593
rect 15749 71553 15761 71587
rect 15795 71553 15807 71587
rect 15749 71547 15807 71553
rect 16574 71544 16580 71596
rect 16632 71584 16638 71596
rect 16632 71556 16677 71584
rect 16632 71544 16638 71556
rect 1394 71516 1400 71528
rect 1355 71488 1400 71516
rect 1394 71476 1400 71488
rect 1452 71476 1458 71528
rect 15286 71476 15292 71528
rect 15344 71516 15350 71528
rect 16776 71525 16804 71624
rect 17862 71612 17868 71624
rect 17920 71612 17926 71664
rect 30834 71612 30840 71664
rect 30892 71652 30898 71664
rect 31018 71652 31024 71664
rect 30892 71624 31024 71652
rect 30892 71612 30898 71624
rect 31018 71612 31024 71624
rect 31076 71652 31082 71664
rect 32122 71652 32128 71664
rect 31076 71624 32128 71652
rect 31076 71612 31082 71624
rect 32122 71612 32128 71624
rect 32180 71612 32186 71664
rect 16850 71544 16856 71596
rect 16908 71584 16914 71596
rect 17310 71584 17316 71596
rect 16908 71556 17316 71584
rect 16908 71544 16914 71556
rect 17310 71544 17316 71556
rect 17368 71584 17374 71596
rect 17405 71587 17463 71593
rect 17405 71584 17417 71587
rect 17368 71556 17417 71584
rect 17368 71544 17374 71556
rect 17405 71553 17417 71556
rect 17451 71553 17463 71587
rect 26602 71584 26608 71596
rect 17405 71547 17463 71553
rect 17512 71556 26608 71584
rect 15933 71519 15991 71525
rect 15933 71516 15945 71519
rect 15344 71488 15945 71516
rect 15344 71476 15350 71488
rect 15933 71485 15945 71488
rect 15979 71485 15991 71519
rect 15933 71479 15991 71485
rect 16761 71519 16819 71525
rect 16761 71485 16773 71519
rect 16807 71485 16819 71519
rect 16761 71479 16819 71485
rect 15746 71408 15752 71460
rect 15804 71448 15810 71460
rect 17512 71448 17540 71556
rect 26602 71544 26608 71556
rect 26660 71544 26666 71596
rect 31386 71544 31392 71596
rect 31444 71544 31450 71596
rect 31754 71584 31760 71596
rect 31588 71556 31760 71584
rect 17589 71519 17647 71525
rect 17589 71485 17601 71519
rect 17635 71485 17647 71519
rect 31404 71516 31432 71544
rect 31588 71525 31616 71556
rect 31754 71544 31760 71556
rect 31812 71584 31818 71596
rect 32490 71584 32496 71596
rect 31812 71556 32496 71584
rect 31812 71544 31818 71556
rect 32490 71544 32496 71556
rect 32548 71544 32554 71596
rect 37550 71544 37556 71596
rect 37608 71584 37614 71596
rect 37608 71556 38884 71584
rect 37608 71544 37614 71556
rect 38856 71528 38884 71556
rect 31481 71519 31539 71525
rect 31481 71516 31493 71519
rect 31404 71488 31493 71516
rect 17589 71479 17647 71485
rect 31481 71485 31493 71488
rect 31527 71485 31539 71519
rect 31481 71479 31539 71485
rect 31573 71519 31631 71525
rect 31573 71485 31585 71519
rect 31619 71485 31631 71519
rect 31573 71479 31631 71485
rect 31849 71519 31907 71525
rect 31849 71485 31861 71519
rect 31895 71485 31907 71519
rect 32122 71516 32128 71528
rect 32083 71488 32128 71516
rect 31849 71479 31907 71485
rect 15804 71420 17540 71448
rect 15804 71408 15810 71420
rect 17402 71340 17408 71392
rect 17460 71380 17466 71392
rect 17604 71380 17632 71479
rect 30834 71408 30840 71460
rect 30892 71448 30898 71460
rect 31021 71451 31079 71457
rect 31021 71448 31033 71451
rect 30892 71420 31033 71448
rect 30892 71408 30898 71420
rect 31021 71417 31033 71420
rect 31067 71417 31079 71451
rect 31021 71411 31079 71417
rect 17460 71352 17632 71380
rect 17460 71340 17466 71352
rect 31202 71340 31208 71392
rect 31260 71380 31266 71392
rect 31864 71380 31892 71479
rect 32122 71476 32128 71488
rect 32180 71476 32186 71528
rect 32398 71516 32404 71528
rect 32359 71488 32404 71516
rect 32398 71476 32404 71488
rect 32456 71476 32462 71528
rect 35805 71519 35863 71525
rect 35805 71485 35817 71519
rect 35851 71516 35863 71519
rect 35986 71516 35992 71528
rect 35851 71488 35992 71516
rect 35851 71485 35863 71488
rect 35805 71479 35863 71485
rect 35986 71476 35992 71488
rect 36044 71516 36050 71528
rect 36446 71516 36452 71528
rect 36044 71488 36452 71516
rect 36044 71476 36050 71488
rect 36446 71476 36452 71488
rect 36504 71476 36510 71528
rect 37458 71516 37464 71528
rect 37419 71488 37464 71516
rect 37458 71476 37464 71488
rect 37516 71476 37522 71528
rect 38102 71516 38108 71528
rect 38063 71488 38108 71516
rect 38102 71476 38108 71488
rect 38160 71476 38166 71528
rect 38838 71476 38844 71528
rect 38896 71476 38902 71528
rect 37274 71380 37280 71392
rect 31260 71352 31892 71380
rect 37235 71352 37280 71380
rect 31260 71340 31266 71352
rect 37274 71340 37280 71352
rect 37332 71340 37338 71392
rect 37550 71340 37556 71392
rect 37608 71380 37614 71392
rect 37921 71383 37979 71389
rect 37921 71380 37933 71383
rect 37608 71352 37933 71380
rect 37608 71340 37614 71352
rect 37921 71349 37933 71352
rect 37967 71349 37979 71383
rect 37921 71343 37979 71349
rect 1104 71290 38824 71312
rect 1104 71238 19606 71290
rect 19658 71238 19670 71290
rect 19722 71238 19734 71290
rect 19786 71238 19798 71290
rect 19850 71238 38824 71290
rect 1104 71216 38824 71238
rect 15562 71176 15568 71188
rect 15523 71148 15568 71176
rect 15562 71136 15568 71148
rect 15620 71136 15626 71188
rect 16390 71176 16396 71188
rect 16351 71148 16396 71176
rect 16390 71136 16396 71148
rect 16448 71136 16454 71188
rect 16758 71136 16764 71188
rect 16816 71176 16822 71188
rect 31202 71176 31208 71188
rect 16816 71148 31208 71176
rect 16816 71136 16822 71148
rect 31202 71136 31208 71148
rect 31260 71136 31266 71188
rect 3418 71068 3424 71120
rect 3476 71108 3482 71120
rect 32122 71108 32128 71120
rect 3476 71080 16252 71108
rect 3476 71068 3482 71080
rect 2498 71000 2504 71052
rect 2556 71040 2562 71052
rect 16224 71049 16252 71080
rect 31772 71080 32128 71108
rect 15381 71043 15439 71049
rect 15381 71040 15393 71043
rect 2556 71012 15393 71040
rect 2556 71000 2562 71012
rect 15381 71009 15393 71012
rect 15427 71009 15439 71043
rect 15381 71003 15439 71009
rect 16209 71043 16267 71049
rect 16209 71009 16221 71043
rect 16255 71009 16267 71043
rect 16209 71003 16267 71009
rect 30742 71000 30748 71052
rect 30800 71040 30806 71052
rect 31113 71043 31171 71049
rect 31113 71040 31125 71043
rect 30800 71012 31125 71040
rect 30800 71000 30806 71012
rect 31113 71009 31125 71012
rect 31159 71009 31171 71043
rect 31386 71040 31392 71052
rect 31347 71012 31392 71040
rect 31113 71003 31171 71009
rect 31386 71000 31392 71012
rect 31444 71000 31450 71052
rect 31772 71049 31800 71080
rect 32122 71068 32128 71080
rect 32180 71108 32186 71120
rect 32398 71108 32404 71120
rect 32180 71080 32404 71108
rect 32180 71068 32186 71080
rect 32398 71068 32404 71080
rect 32456 71068 32462 71120
rect 31481 71043 31539 71049
rect 31481 71009 31493 71043
rect 31527 71009 31539 71043
rect 31481 71003 31539 71009
rect 31757 71043 31815 71049
rect 31757 71009 31769 71043
rect 31803 71009 31815 71043
rect 32030 71040 32036 71052
rect 31991 71012 32036 71040
rect 31757 71003 31815 71009
rect 15197 70975 15255 70981
rect 15197 70941 15209 70975
rect 15243 70972 15255 70975
rect 15470 70972 15476 70984
rect 15243 70944 15476 70972
rect 15243 70941 15255 70944
rect 15197 70935 15255 70941
rect 15470 70932 15476 70944
rect 15528 70932 15534 70984
rect 16025 70975 16083 70981
rect 16025 70941 16037 70975
rect 16071 70972 16083 70975
rect 16574 70972 16580 70984
rect 16071 70944 16580 70972
rect 16071 70941 16083 70944
rect 16025 70935 16083 70941
rect 16574 70932 16580 70944
rect 16632 70972 16638 70984
rect 16850 70972 16856 70984
rect 16632 70944 16856 70972
rect 16632 70932 16638 70944
rect 16850 70932 16856 70944
rect 16908 70932 16914 70984
rect 17770 70932 17776 70984
rect 17828 70972 17834 70984
rect 31496 70972 31524 71003
rect 32030 71000 32036 71012
rect 32088 71000 32094 71052
rect 37366 71040 37372 71052
rect 37327 71012 37372 71040
rect 37366 71000 37372 71012
rect 37424 71000 37430 71052
rect 17828 70944 31524 70972
rect 17828 70932 17834 70944
rect 32122 70932 32128 70984
rect 32180 70972 32186 70984
rect 32950 70972 32956 70984
rect 32180 70944 32956 70972
rect 32180 70932 32186 70944
rect 32950 70932 32956 70944
rect 33008 70932 33014 70984
rect 32030 70864 32036 70916
rect 32088 70904 32094 70916
rect 33042 70904 33048 70916
rect 32088 70876 33048 70904
rect 32088 70864 32094 70876
rect 33042 70864 33048 70876
rect 33100 70864 33106 70916
rect 15470 70796 15476 70848
rect 15528 70836 15534 70848
rect 17218 70836 17224 70848
rect 15528 70808 17224 70836
rect 15528 70796 15534 70808
rect 17218 70796 17224 70808
rect 17276 70796 17282 70848
rect 22830 70796 22836 70848
rect 22888 70836 22894 70848
rect 30745 70839 30803 70845
rect 30745 70836 30757 70839
rect 22888 70808 30757 70836
rect 22888 70796 22894 70808
rect 30745 70805 30757 70808
rect 30791 70805 30803 70839
rect 30745 70799 30803 70805
rect 37090 70796 37096 70848
rect 37148 70836 37154 70848
rect 37185 70839 37243 70845
rect 37185 70836 37197 70839
rect 37148 70808 37197 70836
rect 37148 70796 37154 70808
rect 37185 70805 37197 70808
rect 37231 70805 37243 70839
rect 37185 70799 37243 70805
rect 1104 70746 38824 70768
rect 1104 70694 4246 70746
rect 4298 70694 4310 70746
rect 4362 70694 4374 70746
rect 4426 70694 4438 70746
rect 4490 70694 34966 70746
rect 35018 70694 35030 70746
rect 35082 70694 35094 70746
rect 35146 70694 35158 70746
rect 35210 70694 38824 70746
rect 1104 70672 38824 70694
rect 2130 70592 2136 70644
rect 2188 70632 2194 70644
rect 15838 70632 15844 70644
rect 2188 70604 6914 70632
rect 15799 70604 15844 70632
rect 2188 70592 2194 70604
rect 6886 70564 6914 70604
rect 15838 70592 15844 70604
rect 15896 70592 15902 70644
rect 16666 70632 16672 70644
rect 16627 70604 16672 70632
rect 16666 70592 16672 70604
rect 16724 70592 16730 70644
rect 17494 70632 17500 70644
rect 17455 70604 17500 70632
rect 17494 70592 17500 70604
rect 17552 70592 17558 70644
rect 6886 70536 16574 70564
rect 6270 70456 6276 70508
rect 6328 70496 6334 70508
rect 16301 70499 16359 70505
rect 6328 70468 15792 70496
rect 6328 70456 6334 70468
rect 1394 70428 1400 70440
rect 1355 70400 1400 70428
rect 1394 70388 1400 70400
rect 1452 70388 1458 70440
rect 14458 70388 14464 70440
rect 14516 70428 14522 70440
rect 15470 70428 15476 70440
rect 14516 70400 15332 70428
rect 15431 70400 15476 70428
rect 14516 70388 14522 70400
rect 15304 70360 15332 70400
rect 15470 70388 15476 70400
rect 15528 70388 15534 70440
rect 15657 70431 15715 70437
rect 15657 70428 15669 70431
rect 15580 70400 15669 70428
rect 15580 70360 15608 70400
rect 15657 70397 15669 70400
rect 15703 70397 15715 70431
rect 15764 70428 15792 70468
rect 16301 70465 16313 70499
rect 16347 70496 16359 70499
rect 16390 70496 16396 70508
rect 16347 70468 16396 70496
rect 16347 70465 16359 70468
rect 16301 70459 16359 70465
rect 16390 70456 16396 70468
rect 16448 70456 16454 70508
rect 16546 70496 16574 70536
rect 31386 70524 31392 70576
rect 31444 70564 31450 70576
rect 31754 70564 31760 70576
rect 31444 70536 31760 70564
rect 31444 70524 31450 70536
rect 31754 70524 31760 70536
rect 31812 70524 31818 70576
rect 37277 70567 37335 70573
rect 37277 70533 37289 70567
rect 37323 70564 37335 70567
rect 37826 70564 37832 70576
rect 37323 70536 37832 70564
rect 37323 70533 37335 70536
rect 37277 70527 37335 70533
rect 37826 70524 37832 70536
rect 37884 70524 37890 70576
rect 37921 70567 37979 70573
rect 37921 70533 37933 70567
rect 37967 70564 37979 70567
rect 38010 70564 38016 70576
rect 37967 70536 38016 70564
rect 37967 70533 37979 70536
rect 37921 70527 37979 70533
rect 38010 70524 38016 70536
rect 38068 70524 38074 70576
rect 16500 70468 16574 70496
rect 16960 70468 17356 70496
rect 16500 70437 16528 70468
rect 16960 70437 16988 70468
rect 16485 70431 16543 70437
rect 15764 70400 16436 70428
rect 15657 70391 15715 70397
rect 15304 70332 15608 70360
rect 16408 70360 16436 70400
rect 16485 70397 16497 70431
rect 16531 70397 16543 70431
rect 16945 70431 17003 70437
rect 16945 70428 16957 70431
rect 16485 70391 16543 70397
rect 16592 70400 16957 70428
rect 16592 70360 16620 70400
rect 16945 70397 16957 70400
rect 16991 70397 17003 70431
rect 17218 70428 17224 70440
rect 17179 70400 17224 70428
rect 16945 70391 17003 70397
rect 17218 70388 17224 70400
rect 17276 70388 17282 70440
rect 17328 70437 17356 70468
rect 17313 70431 17371 70437
rect 17313 70397 17325 70431
rect 17359 70397 17371 70431
rect 17313 70391 17371 70397
rect 26602 70388 26608 70440
rect 26660 70428 26666 70440
rect 31386 70428 31392 70440
rect 26660 70400 31248 70428
rect 31347 70400 31392 70428
rect 26660 70388 26666 70400
rect 16408 70332 16620 70360
rect 26326 70320 26332 70372
rect 26384 70360 26390 70372
rect 30929 70363 30987 70369
rect 30929 70360 30941 70363
rect 26384 70332 30941 70360
rect 26384 70320 26390 70332
rect 30929 70329 30941 70332
rect 30975 70329 30987 70363
rect 30929 70323 30987 70329
rect 31220 70292 31248 70400
rect 31386 70388 31392 70400
rect 31444 70388 31450 70440
rect 31662 70428 31668 70440
rect 31623 70400 31668 70428
rect 31662 70388 31668 70400
rect 31720 70388 31726 70440
rect 31757 70431 31815 70437
rect 31757 70397 31769 70431
rect 31803 70397 31815 70431
rect 32030 70428 32036 70440
rect 31991 70400 32036 70428
rect 31757 70391 31815 70397
rect 31772 70292 31800 70391
rect 32030 70388 32036 70400
rect 32088 70388 32094 70440
rect 32309 70431 32367 70437
rect 32309 70397 32321 70431
rect 32355 70428 32367 70431
rect 32398 70428 32404 70440
rect 32355 70400 32404 70428
rect 32355 70397 32367 70400
rect 32309 70391 32367 70397
rect 32398 70388 32404 70400
rect 32456 70388 32462 70440
rect 37458 70428 37464 70440
rect 37419 70400 37464 70428
rect 37458 70388 37464 70400
rect 37516 70388 37522 70440
rect 38105 70431 38163 70437
rect 38105 70397 38117 70431
rect 38151 70428 38163 70431
rect 38286 70428 38292 70440
rect 38151 70400 38292 70428
rect 38151 70397 38163 70400
rect 38105 70391 38163 70397
rect 38286 70388 38292 70400
rect 38344 70388 38350 70440
rect 37734 70320 37740 70372
rect 37792 70320 37798 70372
rect 38654 70320 38660 70372
rect 38712 70360 38718 70372
rect 38712 70332 39160 70360
rect 38712 70320 38718 70332
rect 31220 70264 31800 70292
rect 37752 70292 37780 70320
rect 37918 70292 37924 70304
rect 37752 70264 37924 70292
rect 37918 70252 37924 70264
rect 37976 70252 37982 70304
rect 1104 70202 38824 70224
rect 1104 70150 19606 70202
rect 19658 70150 19670 70202
rect 19722 70150 19734 70202
rect 19786 70150 19798 70202
rect 19850 70150 38824 70202
rect 39132 70168 39160 70332
rect 39298 70320 39304 70372
rect 39356 70360 39362 70372
rect 39356 70332 39401 70360
rect 39356 70320 39362 70332
rect 1104 70128 38824 70150
rect 39114 70116 39120 70168
rect 39172 70116 39178 70168
rect 16206 70048 16212 70100
rect 16264 70088 16270 70100
rect 16393 70091 16451 70097
rect 16393 70088 16405 70091
rect 16264 70060 16405 70088
rect 16264 70048 16270 70060
rect 16393 70057 16405 70060
rect 16439 70057 16451 70091
rect 16393 70051 16451 70057
rect 37366 70048 37372 70100
rect 37424 70088 37430 70100
rect 37642 70088 37648 70100
rect 37424 70060 37648 70088
rect 37424 70048 37430 70060
rect 37642 70048 37648 70060
rect 37700 70048 37706 70100
rect 1394 69952 1400 69964
rect 1355 69924 1400 69952
rect 1394 69912 1400 69924
rect 1452 69912 1458 69964
rect 6362 69912 6368 69964
rect 6420 69952 6426 69964
rect 16209 69955 16267 69961
rect 16209 69952 16221 69955
rect 6420 69924 16221 69952
rect 6420 69912 6426 69924
rect 16209 69921 16221 69924
rect 16255 69921 16267 69955
rect 36722 69952 36728 69964
rect 36683 69924 36728 69952
rect 16209 69915 16267 69921
rect 36722 69912 36728 69924
rect 36780 69912 36786 69964
rect 37366 69952 37372 69964
rect 37327 69924 37372 69952
rect 37366 69912 37372 69924
rect 37424 69912 37430 69964
rect 15470 69844 15476 69896
rect 15528 69884 15534 69896
rect 16025 69887 16083 69893
rect 16025 69884 16037 69887
rect 15528 69856 16037 69884
rect 15528 69844 15534 69856
rect 16025 69853 16037 69856
rect 16071 69884 16083 69887
rect 16114 69884 16120 69896
rect 16071 69856 16120 69884
rect 16071 69853 16083 69856
rect 16025 69847 16083 69853
rect 16114 69844 16120 69856
rect 16172 69844 16178 69896
rect 36541 69819 36599 69825
rect 36541 69785 36553 69819
rect 36587 69816 36599 69819
rect 36998 69816 37004 69828
rect 36587 69788 37004 69816
rect 36587 69785 36599 69788
rect 36541 69779 36599 69785
rect 36998 69776 37004 69788
rect 37056 69776 37062 69828
rect 36906 69708 36912 69760
rect 36964 69748 36970 69760
rect 37185 69751 37243 69757
rect 37185 69748 37197 69751
rect 36964 69720 37197 69748
rect 36964 69708 36970 69720
rect 37185 69717 37197 69720
rect 37231 69717 37243 69751
rect 37185 69711 37243 69717
rect 39758 69680 39764 69692
rect 1104 69658 38824 69680
rect 1104 69606 4246 69658
rect 4298 69606 4310 69658
rect 4362 69606 4374 69658
rect 4426 69606 4438 69658
rect 4490 69606 34966 69658
rect 35018 69606 35030 69658
rect 35082 69606 35094 69658
rect 35146 69606 35158 69658
rect 35210 69606 38824 69658
rect 39719 69652 39764 69680
rect 39758 69640 39764 69652
rect 39816 69640 39822 69692
rect 1104 69584 38824 69606
rect 16298 69504 16304 69556
rect 16356 69544 16362 69556
rect 16485 69547 16543 69553
rect 16485 69544 16497 69547
rect 16356 69516 16497 69544
rect 16356 69504 16362 69516
rect 16485 69513 16497 69516
rect 16531 69513 16543 69547
rect 16485 69507 16543 69513
rect 38194 69504 38200 69556
rect 38252 69544 38258 69556
rect 39758 69544 39764 69556
rect 38252 69516 39764 69544
rect 38252 69504 38258 69516
rect 39758 69504 39764 69516
rect 39816 69504 39822 69556
rect 32398 69436 32404 69488
rect 32456 69476 32462 69488
rect 37185 69479 37243 69485
rect 37185 69476 37197 69479
rect 32456 69448 37197 69476
rect 32456 69436 32462 69448
rect 37185 69445 37197 69448
rect 37231 69445 37243 69479
rect 38378 69476 38384 69488
rect 37185 69439 37243 69445
rect 38212 69448 38384 69476
rect 38212 69420 38240 69448
rect 38378 69436 38384 69448
rect 38436 69436 38442 69488
rect 16114 69408 16120 69420
rect 16075 69380 16120 69408
rect 16114 69368 16120 69380
rect 16172 69368 16178 69420
rect 38194 69368 38200 69420
rect 38252 69368 38258 69420
rect 2038 69300 2044 69352
rect 2096 69340 2102 69352
rect 16301 69343 16359 69349
rect 2096 69312 6914 69340
rect 2096 69300 2102 69312
rect 6886 69272 6914 69312
rect 16301 69309 16313 69343
rect 16347 69309 16359 69343
rect 36630 69340 36636 69352
rect 36591 69312 36636 69340
rect 16301 69303 16359 69309
rect 16316 69272 16344 69303
rect 36630 69300 36636 69312
rect 36688 69300 36694 69352
rect 37001 69343 37059 69349
rect 37001 69309 37013 69343
rect 37047 69340 37059 69343
rect 37274 69340 37280 69352
rect 37047 69312 37280 69340
rect 37047 69309 37059 69312
rect 37001 69303 37059 69309
rect 37274 69300 37280 69312
rect 37332 69300 37338 69352
rect 38105 69343 38163 69349
rect 38105 69309 38117 69343
rect 38151 69340 38163 69343
rect 38378 69340 38384 69352
rect 38151 69312 38384 69340
rect 38151 69309 38163 69312
rect 38105 69303 38163 69309
rect 38378 69300 38384 69312
rect 38436 69300 38442 69352
rect 6886 69244 16344 69272
rect 35894 69232 35900 69284
rect 35952 69272 35958 69284
rect 36722 69272 36728 69284
rect 35952 69244 36728 69272
rect 35952 69232 35958 69244
rect 36722 69232 36728 69244
rect 36780 69272 36786 69284
rect 36817 69275 36875 69281
rect 36817 69272 36829 69275
rect 36780 69244 36829 69272
rect 36780 69232 36786 69244
rect 36817 69241 36829 69244
rect 36863 69241 36875 69275
rect 36817 69235 36875 69241
rect 36909 69275 36967 69281
rect 36909 69241 36921 69275
rect 36955 69272 36967 69275
rect 36955 69244 37320 69272
rect 36955 69241 36967 69244
rect 36909 69235 36967 69241
rect 37292 69216 37320 69244
rect 33962 69164 33968 69216
rect 34020 69204 34026 69216
rect 35342 69204 35348 69216
rect 34020 69176 35348 69204
rect 34020 69164 34026 69176
rect 35342 69164 35348 69176
rect 35400 69164 35406 69216
rect 37274 69164 37280 69216
rect 37332 69164 37338 69216
rect 37921 69207 37979 69213
rect 37921 69173 37933 69207
rect 37967 69204 37979 69207
rect 38010 69204 38016 69216
rect 37967 69176 38016 69204
rect 37967 69173 37979 69176
rect 37921 69167 37979 69173
rect 38010 69164 38016 69176
rect 38068 69164 38074 69216
rect 39206 69204 39212 69216
rect 39167 69176 39212 69204
rect 39206 69164 39212 69176
rect 39264 69164 39270 69216
rect 1104 69114 38824 69136
rect 1104 69062 19606 69114
rect 19658 69062 19670 69114
rect 19722 69062 19734 69114
rect 19786 69062 19798 69114
rect 19850 69062 38824 69114
rect 1104 69040 38824 69062
rect 36722 68960 36728 69012
rect 36780 69000 36786 69012
rect 36780 68972 36952 69000
rect 36780 68960 36786 68972
rect 36078 68892 36084 68944
rect 36136 68932 36142 68944
rect 36924 68941 36952 68972
rect 36909 68935 36967 68941
rect 36136 68904 36768 68932
rect 36136 68892 36142 68904
rect 1394 68864 1400 68876
rect 1355 68836 1400 68864
rect 1394 68824 1400 68836
rect 1452 68824 1458 68876
rect 35802 68824 35808 68876
rect 35860 68864 35866 68876
rect 36740 68873 36768 68904
rect 36909 68901 36921 68935
rect 36955 68901 36967 68935
rect 36909 68895 36967 68901
rect 37001 68935 37059 68941
rect 37001 68901 37013 68935
rect 37047 68932 37059 68935
rect 37274 68932 37280 68944
rect 37047 68904 37280 68932
rect 37047 68901 37059 68904
rect 37001 68895 37059 68901
rect 37274 68892 37280 68904
rect 37332 68892 37338 68944
rect 36265 68867 36323 68873
rect 36265 68864 36277 68867
rect 35860 68836 36277 68864
rect 35860 68824 35866 68836
rect 36265 68833 36277 68836
rect 36311 68833 36323 68867
rect 36265 68827 36323 68833
rect 36725 68867 36783 68873
rect 36725 68833 36737 68867
rect 36771 68833 36783 68867
rect 36725 68827 36783 68833
rect 37090 68824 37096 68876
rect 37148 68864 37154 68876
rect 37148 68836 37193 68864
rect 37148 68824 37154 68836
rect 36081 68731 36139 68737
rect 36081 68697 36093 68731
rect 36127 68728 36139 68731
rect 37182 68728 37188 68740
rect 36127 68700 37188 68728
rect 36127 68697 36139 68700
rect 36081 68691 36139 68697
rect 37182 68688 37188 68700
rect 37240 68688 37246 68740
rect 34514 68620 34520 68672
rect 34572 68660 34578 68672
rect 37277 68663 37335 68669
rect 37277 68660 37289 68663
rect 34572 68632 37289 68660
rect 34572 68620 34578 68632
rect 37277 68629 37289 68632
rect 37323 68629 37335 68663
rect 37277 68623 37335 68629
rect 1104 68570 38824 68592
rect 1104 68518 4246 68570
rect 4298 68518 4310 68570
rect 4362 68518 4374 68570
rect 4426 68518 4438 68570
rect 4490 68518 34966 68570
rect 35018 68518 35030 68570
rect 35082 68518 35094 68570
rect 35146 68518 35158 68570
rect 35210 68518 38824 68570
rect 1104 68496 38824 68518
rect 36262 68416 36268 68468
rect 36320 68456 36326 68468
rect 36446 68456 36452 68468
rect 36320 68428 36452 68456
rect 36320 68416 36326 68428
rect 36446 68416 36452 68428
rect 36504 68416 36510 68468
rect 37277 68459 37335 68465
rect 37277 68425 37289 68459
rect 37323 68456 37335 68459
rect 37366 68456 37372 68468
rect 37323 68428 37372 68456
rect 37323 68425 37335 68428
rect 37277 68419 37335 68425
rect 37366 68416 37372 68428
rect 37424 68416 37430 68468
rect 30098 68348 30104 68400
rect 30156 68388 30162 68400
rect 34514 68388 34520 68400
rect 30156 68360 34520 68388
rect 30156 68348 30162 68360
rect 34514 68348 34520 68360
rect 34572 68348 34578 68400
rect 36722 68348 36728 68400
rect 36780 68348 36786 68400
rect 36170 68280 36176 68332
rect 36228 68320 36234 68332
rect 36630 68320 36636 68332
rect 36228 68292 36636 68320
rect 36228 68280 36234 68292
rect 36630 68280 36636 68292
rect 36688 68280 36694 68332
rect 36740 68320 36768 68348
rect 36740 68292 36952 68320
rect 1394 68252 1400 68264
rect 1355 68224 1400 68252
rect 1394 68212 1400 68224
rect 1452 68212 1458 68264
rect 31941 68255 31999 68261
rect 31941 68221 31953 68255
rect 31987 68252 31999 68255
rect 36262 68252 36268 68264
rect 31987 68224 32021 68252
rect 36223 68224 36268 68252
rect 31987 68221 31999 68224
rect 31941 68215 31999 68221
rect 1578 68144 1584 68196
rect 1636 68184 1642 68196
rect 31849 68187 31907 68193
rect 31849 68184 31861 68187
rect 1636 68156 31861 68184
rect 1636 68144 1642 68156
rect 31849 68153 31861 68156
rect 31895 68184 31907 68187
rect 31956 68184 31984 68215
rect 36262 68212 36268 68224
rect 36320 68212 36326 68264
rect 36725 68255 36783 68261
rect 36725 68221 36737 68255
rect 36771 68252 36783 68255
rect 36814 68252 36820 68264
rect 36771 68224 36820 68252
rect 36771 68221 36783 68224
rect 36725 68215 36783 68221
rect 36814 68212 36820 68224
rect 36872 68212 36878 68264
rect 36924 68261 36952 68292
rect 37366 68280 37372 68332
rect 37424 68320 37430 68332
rect 37918 68320 37924 68332
rect 37424 68292 37924 68320
rect 37424 68280 37430 68292
rect 37918 68280 37924 68292
rect 37976 68280 37982 68332
rect 36909 68255 36967 68261
rect 36909 68221 36921 68255
rect 36955 68221 36967 68255
rect 36909 68215 36967 68221
rect 37093 68255 37151 68261
rect 37093 68221 37105 68255
rect 37139 68252 37151 68255
rect 37550 68252 37556 68264
rect 37139 68224 37556 68252
rect 37139 68221 37151 68224
rect 37093 68215 37151 68221
rect 37550 68212 37556 68224
rect 37608 68212 37614 68264
rect 38105 68255 38163 68261
rect 38105 68221 38117 68255
rect 38151 68252 38163 68255
rect 38194 68252 38200 68264
rect 38151 68224 38200 68252
rect 38151 68221 38163 68224
rect 38105 68215 38163 68221
rect 38194 68212 38200 68224
rect 38252 68212 38258 68264
rect 33042 68184 33048 68196
rect 31895 68156 33048 68184
rect 31895 68153 31907 68156
rect 31849 68147 31907 68153
rect 33042 68144 33048 68156
rect 33100 68144 33106 68196
rect 37001 68187 37059 68193
rect 37001 68184 37013 68187
rect 36004 68156 37013 68184
rect 32125 68119 32183 68125
rect 32125 68085 32137 68119
rect 32171 68116 32183 68119
rect 32950 68116 32956 68128
rect 32171 68088 32956 68116
rect 32171 68085 32183 68088
rect 32125 68079 32183 68085
rect 32950 68076 32956 68088
rect 33008 68116 33014 68128
rect 36004 68116 36032 68156
rect 37001 68153 37013 68156
rect 37047 68184 37059 68187
rect 37274 68184 37280 68196
rect 37047 68156 37280 68184
rect 37047 68153 37059 68156
rect 37001 68147 37059 68153
rect 37274 68144 37280 68156
rect 37332 68144 37338 68196
rect 33008 68088 36032 68116
rect 36081 68119 36139 68125
rect 33008 68076 33014 68088
rect 36081 68085 36093 68119
rect 36127 68116 36139 68119
rect 36170 68116 36176 68128
rect 36127 68088 36176 68116
rect 36127 68085 36139 68088
rect 36081 68079 36139 68085
rect 36170 68076 36176 68088
rect 36228 68076 36234 68128
rect 37918 68116 37924 68128
rect 37879 68088 37924 68116
rect 37918 68076 37924 68088
rect 37976 68076 37982 68128
rect 1104 68026 38824 68048
rect 1104 67974 19606 68026
rect 19658 67974 19670 68026
rect 19722 67974 19734 68026
rect 19786 67974 19798 68026
rect 19850 67974 38824 68026
rect 1104 67952 38824 67974
rect 27522 67872 27528 67924
rect 27580 67912 27586 67924
rect 35342 67912 35348 67924
rect 27580 67884 35348 67912
rect 27580 67872 27586 67884
rect 35342 67872 35348 67884
rect 35400 67872 35406 67924
rect 36722 67872 36728 67924
rect 36780 67872 36786 67924
rect 36814 67872 36820 67924
rect 36872 67912 36878 67924
rect 37642 67912 37648 67924
rect 36872 67884 37648 67912
rect 36872 67872 36878 67884
rect 37642 67872 37648 67884
rect 37700 67872 37706 67924
rect 29914 67804 29920 67856
rect 29972 67844 29978 67856
rect 36740 67844 36768 67872
rect 36909 67847 36967 67853
rect 36909 67844 36921 67847
rect 29972 67816 36308 67844
rect 36740 67816 36921 67844
rect 29972 67804 29978 67816
rect 35894 67736 35900 67788
rect 35952 67776 35958 67788
rect 35989 67779 36047 67785
rect 35989 67776 36001 67779
rect 35952 67748 36001 67776
rect 35952 67736 35958 67748
rect 35989 67745 36001 67748
rect 36035 67745 36047 67779
rect 35989 67739 36047 67745
rect 36280 67708 36308 67816
rect 36909 67813 36921 67816
rect 36955 67813 36967 67847
rect 36909 67807 36967 67813
rect 37001 67847 37059 67853
rect 37001 67813 37013 67847
rect 37047 67844 37059 67847
rect 37274 67844 37280 67856
rect 37047 67816 37280 67844
rect 37047 67813 37059 67816
rect 37001 67807 37059 67813
rect 37274 67804 37280 67816
rect 37332 67804 37338 67856
rect 36722 67776 36728 67788
rect 36683 67748 36728 67776
rect 36722 67736 36728 67748
rect 36780 67736 36786 67788
rect 37090 67736 37096 67788
rect 37148 67776 37154 67788
rect 37148 67748 37193 67776
rect 37148 67736 37154 67748
rect 36280 67680 37320 67708
rect 35710 67600 35716 67652
rect 35768 67640 35774 67652
rect 37292 67649 37320 67680
rect 37277 67643 37335 67649
rect 35768 67612 36216 67640
rect 35768 67600 35774 67612
rect 30190 67532 30196 67584
rect 30248 67572 30254 67584
rect 36078 67572 36084 67584
rect 30248 67544 36084 67572
rect 30248 67532 30254 67544
rect 36078 67532 36084 67544
rect 36136 67532 36142 67584
rect 36188 67581 36216 67612
rect 37277 67609 37289 67643
rect 37323 67609 37335 67643
rect 37277 67603 37335 67609
rect 36173 67575 36231 67581
rect 36173 67541 36185 67575
rect 36219 67541 36231 67575
rect 36173 67535 36231 67541
rect 36630 67532 36636 67584
rect 36688 67572 36694 67584
rect 39206 67572 39212 67584
rect 36688 67544 39212 67572
rect 36688 67532 36694 67544
rect 39206 67532 39212 67544
rect 39264 67532 39270 67584
rect 1104 67482 38824 67504
rect 1104 67430 4246 67482
rect 4298 67430 4310 67482
rect 4362 67430 4374 67482
rect 4426 67430 4438 67482
rect 4490 67430 34966 67482
rect 35018 67430 35030 67482
rect 35082 67430 35094 67482
rect 35146 67430 35158 67482
rect 35210 67430 38824 67482
rect 1104 67408 38824 67430
rect 36078 67328 36084 67380
rect 36136 67368 36142 67380
rect 38105 67371 38163 67377
rect 38105 67368 38117 67371
rect 36136 67340 38117 67368
rect 36136 67328 36142 67340
rect 38105 67337 38117 67340
rect 38151 67337 38163 67371
rect 38105 67331 38163 67337
rect 31202 67260 31208 67312
rect 31260 67300 31266 67312
rect 37093 67303 37151 67309
rect 37093 67300 37105 67303
rect 31260 67272 37105 67300
rect 31260 67260 31266 67272
rect 37093 67269 37105 67272
rect 37139 67269 37151 67303
rect 39574 67300 39580 67312
rect 37093 67263 37151 67269
rect 37752 67272 39580 67300
rect 1394 67164 1400 67176
rect 1355 67136 1400 67164
rect 1394 67124 1400 67136
rect 1452 67124 1458 67176
rect 32953 67167 33011 67173
rect 32953 67133 32965 67167
rect 32999 67164 33011 67167
rect 33042 67164 33048 67176
rect 32999 67136 33048 67164
rect 32999 67133 33011 67136
rect 32953 67127 33011 67133
rect 33042 67124 33048 67136
rect 33100 67124 33106 67176
rect 35897 67167 35955 67173
rect 35897 67133 35909 67167
rect 35943 67164 35955 67167
rect 35986 67164 35992 67176
rect 35943 67136 35992 67164
rect 35943 67133 35955 67136
rect 35897 67127 35955 67133
rect 35986 67124 35992 67136
rect 36044 67124 36050 67176
rect 36538 67164 36544 67176
rect 36499 67136 36544 67164
rect 36538 67124 36544 67136
rect 36596 67124 36602 67176
rect 36906 67164 36912 67176
rect 36867 67136 36912 67164
rect 36906 67124 36912 67136
rect 36964 67124 36970 67176
rect 37553 67167 37611 67173
rect 37108 67136 37509 67164
rect 37108 67108 37136 67136
rect 33137 67099 33195 67105
rect 33137 67065 33149 67099
rect 33183 67096 33195 67099
rect 34146 67096 34152 67108
rect 33183 67068 34152 67096
rect 33183 67065 33195 67068
rect 33137 67059 33195 67065
rect 34146 67056 34152 67068
rect 34204 67056 34210 67108
rect 36722 67096 36728 67108
rect 36683 67068 36728 67096
rect 36722 67056 36728 67068
rect 36780 67056 36786 67108
rect 36817 67099 36875 67105
rect 36817 67065 36829 67099
rect 36863 67096 36875 67099
rect 37090 67096 37096 67108
rect 36863 67068 37096 67096
rect 36863 67065 36875 67068
rect 36817 67059 36875 67065
rect 37090 67056 37096 67068
rect 37148 67056 37154 67108
rect 36078 67028 36084 67040
rect 36039 67000 36084 67028
rect 36078 66988 36084 67000
rect 36136 66988 36142 67040
rect 37481 67028 37509 67136
rect 37553 67133 37565 67167
rect 37599 67164 37611 67167
rect 37752 67164 37780 67272
rect 39574 67260 39580 67272
rect 39632 67260 39638 67312
rect 37826 67192 37832 67244
rect 37884 67192 37890 67244
rect 37599 67136 37780 67164
rect 37844 67164 37872 67192
rect 37921 67167 37979 67173
rect 37921 67164 37933 67167
rect 37844 67136 37933 67164
rect 37599 67133 37611 67136
rect 37553 67127 37611 67133
rect 37921 67133 37933 67136
rect 37967 67133 37979 67167
rect 37921 67127 37979 67133
rect 38378 67124 38384 67176
rect 38436 67164 38442 67176
rect 39393 67167 39451 67173
rect 39393 67164 39405 67167
rect 38436 67136 39405 67164
rect 38436 67124 38442 67136
rect 39393 67133 39405 67136
rect 39439 67133 39451 67167
rect 39393 67127 39451 67133
rect 39574 67124 39580 67176
rect 39632 67164 39638 67176
rect 39761 67167 39819 67173
rect 39761 67164 39773 67167
rect 39632 67136 39773 67164
rect 39632 67124 39638 67136
rect 39761 67133 39773 67136
rect 39807 67133 39819 67167
rect 39761 67127 39819 67133
rect 37642 67056 37648 67108
rect 37700 67096 37706 67108
rect 37737 67099 37795 67105
rect 37737 67096 37749 67099
rect 37700 67068 37749 67096
rect 37700 67056 37706 67068
rect 37737 67065 37749 67068
rect 37783 67065 37795 67099
rect 37737 67059 37795 67065
rect 37829 67099 37887 67105
rect 37829 67065 37841 67099
rect 37875 67065 37887 67099
rect 37829 67059 37887 67065
rect 37844 67028 37872 67059
rect 37481 67000 37872 67028
rect 1104 66938 38824 66960
rect 1104 66886 19606 66938
rect 19658 66886 19670 66938
rect 19722 66886 19734 66938
rect 19786 66886 19798 66938
rect 19850 66886 38824 66938
rect 1104 66864 38824 66886
rect 36630 66824 36636 66836
rect 35820 66796 36636 66824
rect 1394 66688 1400 66700
rect 1355 66660 1400 66688
rect 1394 66648 1400 66660
rect 1452 66648 1458 66700
rect 34701 66691 34759 66697
rect 34701 66657 34713 66691
rect 34747 66688 34759 66691
rect 34790 66688 34796 66700
rect 34747 66660 34796 66688
rect 34747 66657 34759 66660
rect 34701 66651 34759 66657
rect 34790 66648 34796 66660
rect 34848 66648 34854 66700
rect 35342 66688 35348 66700
rect 35303 66660 35348 66688
rect 35342 66648 35348 66660
rect 35400 66648 35406 66700
rect 35820 66697 35848 66796
rect 36630 66784 36636 66796
rect 36688 66784 36694 66836
rect 36906 66784 36912 66836
rect 36964 66824 36970 66836
rect 38838 66824 38844 66836
rect 36964 66796 38844 66824
rect 36964 66784 36970 66796
rect 38838 66784 38844 66796
rect 38896 66784 38902 66836
rect 35989 66759 36047 66765
rect 35989 66725 36001 66759
rect 36035 66756 36047 66759
rect 36722 66756 36728 66768
rect 36035 66728 36728 66756
rect 36035 66725 36047 66728
rect 35989 66719 36047 66725
rect 36722 66716 36728 66728
rect 36780 66756 36786 66768
rect 37001 66759 37059 66765
rect 37001 66756 37013 66759
rect 36780 66728 37013 66756
rect 36780 66716 36786 66728
rect 37001 66725 37013 66728
rect 37047 66756 37059 66759
rect 37274 66756 37280 66768
rect 37047 66728 37280 66756
rect 37047 66725 37059 66728
rect 37001 66719 37059 66725
rect 37274 66716 37280 66728
rect 37332 66756 37338 66768
rect 37642 66756 37648 66768
rect 37332 66728 37648 66756
rect 37332 66716 37338 66728
rect 37642 66716 37648 66728
rect 37700 66716 37706 66768
rect 35805 66691 35863 66697
rect 35805 66657 35817 66691
rect 35851 66657 35863 66691
rect 35805 66651 35863 66657
rect 36081 66691 36139 66697
rect 36081 66657 36093 66691
rect 36127 66657 36139 66691
rect 36081 66651 36139 66657
rect 36096 66620 36124 66651
rect 36170 66648 36176 66700
rect 36228 66688 36234 66700
rect 36817 66691 36875 66697
rect 36228 66660 36273 66688
rect 36228 66648 36234 66660
rect 36817 66657 36829 66691
rect 36863 66688 36875 66691
rect 36906 66688 36912 66700
rect 36863 66660 36912 66688
rect 36863 66657 36875 66660
rect 36817 66651 36875 66657
rect 36906 66648 36912 66660
rect 36964 66648 36970 66700
rect 37090 66688 37096 66700
rect 37003 66660 37096 66688
rect 37090 66648 37096 66660
rect 37148 66648 37154 66700
rect 37182 66648 37188 66700
rect 37240 66688 37246 66700
rect 37240 66660 37285 66688
rect 37240 66648 37246 66660
rect 36262 66620 36268 66632
rect 36096 66592 36268 66620
rect 36262 66580 36268 66592
rect 36320 66620 36326 66632
rect 37108 66620 37136 66648
rect 36320 66592 37136 66620
rect 36320 66580 36326 66592
rect 31386 66512 31392 66564
rect 31444 66552 31450 66564
rect 36357 66555 36415 66561
rect 36357 66552 36369 66555
rect 31444 66524 36369 66552
rect 31444 66512 31450 66524
rect 36357 66521 36369 66524
rect 36403 66521 36415 66555
rect 36357 66515 36415 66521
rect 34514 66484 34520 66496
rect 34475 66456 34520 66484
rect 34514 66444 34520 66456
rect 34572 66444 34578 66496
rect 35161 66487 35219 66493
rect 35161 66453 35173 66487
rect 35207 66484 35219 66487
rect 36906 66484 36912 66496
rect 35207 66456 36912 66484
rect 35207 66453 35219 66456
rect 35161 66447 35219 66453
rect 36906 66444 36912 66456
rect 36964 66444 36970 66496
rect 37369 66487 37427 66493
rect 37369 66453 37381 66487
rect 37415 66484 37427 66487
rect 37826 66484 37832 66496
rect 37415 66456 37832 66484
rect 37415 66453 37427 66456
rect 37369 66447 37427 66453
rect 37826 66444 37832 66456
rect 37884 66444 37890 66496
rect 1104 66394 38824 66416
rect 1104 66342 4246 66394
rect 4298 66342 4310 66394
rect 4362 66342 4374 66394
rect 4426 66342 4438 66394
rect 4490 66342 34966 66394
rect 35018 66342 35030 66394
rect 35082 66342 35094 66394
rect 35146 66342 35158 66394
rect 35210 66342 38824 66394
rect 1104 66320 38824 66342
rect 38105 66215 38163 66221
rect 38105 66212 38117 66215
rect 31726 66184 38117 66212
rect 1394 66076 1400 66088
rect 1355 66048 1400 66076
rect 1394 66036 1400 66048
rect 1452 66036 1458 66088
rect 30282 65968 30288 66020
rect 30340 66008 30346 66020
rect 31726 66008 31754 66184
rect 38105 66181 38117 66184
rect 38151 66181 38163 66215
rect 38105 66175 38163 66181
rect 39022 66144 39028 66156
rect 37568 66116 39028 66144
rect 32953 66079 33011 66085
rect 32953 66045 32965 66079
rect 32999 66076 33011 66079
rect 33042 66076 33048 66088
rect 32999 66048 33048 66076
rect 32999 66045 33011 66048
rect 32953 66039 33011 66045
rect 33042 66036 33048 66048
rect 33100 66036 33106 66088
rect 35897 66079 35955 66085
rect 35897 66045 35909 66079
rect 35943 66076 35955 66079
rect 35986 66076 35992 66088
rect 35943 66048 35992 66076
rect 35943 66045 35955 66048
rect 35897 66039 35955 66045
rect 35986 66036 35992 66048
rect 36044 66076 36050 66088
rect 37568 66085 37596 66116
rect 39022 66104 39028 66116
rect 39080 66104 39086 66156
rect 36633 66079 36691 66085
rect 36633 66076 36645 66079
rect 36044 66048 36645 66076
rect 36044 66036 36050 66048
rect 36633 66045 36645 66048
rect 36679 66045 36691 66079
rect 36633 66039 36691 66045
rect 37553 66079 37611 66085
rect 37553 66045 37565 66079
rect 37599 66045 37611 66079
rect 37553 66039 37611 66045
rect 37921 66079 37979 66085
rect 37921 66045 37933 66079
rect 37967 66076 37979 66079
rect 38102 66076 38108 66088
rect 37967 66048 38108 66076
rect 37967 66045 37979 66048
rect 37921 66039 37979 66045
rect 38102 66036 38108 66048
rect 38160 66036 38166 66088
rect 30340 65980 31754 66008
rect 33137 66011 33195 66017
rect 30340 65968 30346 65980
rect 33137 65977 33149 66011
rect 33183 66008 33195 66011
rect 33594 66008 33600 66020
rect 33183 65980 33600 66008
rect 33183 65977 33195 65980
rect 33137 65971 33195 65977
rect 33594 65968 33600 65980
rect 33652 65968 33658 66020
rect 35802 65968 35808 66020
rect 35860 66008 35866 66020
rect 36817 66011 36875 66017
rect 36817 66008 36829 66011
rect 35860 65980 36829 66008
rect 35860 65968 35866 65980
rect 36817 65977 36829 65980
rect 36863 65977 36875 66011
rect 36817 65971 36875 65977
rect 37274 65968 37280 66020
rect 37332 66008 37338 66020
rect 37737 66011 37795 66017
rect 37737 66008 37749 66011
rect 37332 65980 37749 66008
rect 37332 65968 37338 65980
rect 37737 65977 37749 65980
rect 37783 65977 37795 66011
rect 37737 65971 37795 65977
rect 37829 66011 37887 66017
rect 37829 65977 37841 66011
rect 37875 65977 37887 66011
rect 37829 65971 37887 65977
rect 35989 65943 36047 65949
rect 35989 65909 36001 65943
rect 36035 65940 36047 65943
rect 36630 65940 36636 65952
rect 36035 65912 36636 65940
rect 36035 65909 36047 65912
rect 35989 65903 36047 65909
rect 36630 65900 36636 65912
rect 36688 65900 36694 65952
rect 37090 65900 37096 65952
rect 37148 65940 37154 65952
rect 37844 65940 37872 65971
rect 37148 65912 37872 65940
rect 37148 65900 37154 65912
rect 1104 65850 38824 65872
rect 1104 65798 19606 65850
rect 19658 65798 19670 65850
rect 19722 65798 19734 65850
rect 19786 65798 19798 65850
rect 19850 65798 38824 65850
rect 1104 65776 38824 65798
rect 34422 65696 34428 65748
rect 34480 65736 34486 65748
rect 38838 65736 38844 65748
rect 34480 65708 38844 65736
rect 34480 65696 34486 65708
rect 38838 65696 38844 65708
rect 38896 65696 38902 65748
rect 34514 65628 34520 65680
rect 34572 65668 34578 65680
rect 34572 65640 37252 65668
rect 34572 65628 34578 65640
rect 31754 65560 31760 65612
rect 31812 65600 31818 65612
rect 32766 65600 32772 65612
rect 31812 65572 32772 65600
rect 31812 65560 31818 65572
rect 32766 65560 32772 65572
rect 32824 65560 32830 65612
rect 32858 65560 32864 65612
rect 32916 65560 32922 65612
rect 33042 65560 33048 65612
rect 33100 65600 33106 65612
rect 33137 65603 33195 65609
rect 33137 65600 33149 65603
rect 33100 65572 33149 65600
rect 33100 65560 33106 65572
rect 33137 65569 33149 65572
rect 33183 65569 33195 65603
rect 35066 65600 35072 65612
rect 35027 65572 35072 65600
rect 33137 65563 33195 65569
rect 35066 65560 35072 65572
rect 35124 65560 35130 65612
rect 35710 65600 35716 65612
rect 35671 65572 35716 65600
rect 35710 65560 35716 65572
rect 35768 65560 35774 65612
rect 36357 65603 36415 65609
rect 36357 65569 36369 65603
rect 36403 65600 36415 65603
rect 36446 65600 36452 65612
rect 36403 65572 36452 65600
rect 36403 65569 36415 65572
rect 36357 65563 36415 65569
rect 36446 65560 36452 65572
rect 36504 65560 36510 65612
rect 36817 65603 36875 65609
rect 36817 65600 36829 65603
rect 36648 65572 36829 65600
rect 32030 65492 32036 65544
rect 32088 65532 32094 65544
rect 32674 65532 32680 65544
rect 32088 65504 32680 65532
rect 32088 65492 32094 65504
rect 32674 65492 32680 65504
rect 32732 65492 32738 65544
rect 32876 65408 32904 65560
rect 33318 65492 33324 65544
rect 33376 65532 33382 65544
rect 35526 65532 35532 65544
rect 33376 65504 35532 65532
rect 33376 65492 33382 65504
rect 35526 65492 35532 65504
rect 35584 65492 35590 65544
rect 33134 65424 33140 65476
rect 33192 65464 33198 65476
rect 34422 65464 34428 65476
rect 33192 65436 34428 65464
rect 33192 65424 33198 65436
rect 34422 65424 34428 65436
rect 34480 65424 34486 65476
rect 36648 65464 36676 65572
rect 36817 65569 36829 65572
rect 36863 65569 36875 65603
rect 36817 65563 36875 65569
rect 37001 65603 37059 65609
rect 37001 65569 37013 65603
rect 37047 65569 37059 65603
rect 37001 65563 37059 65569
rect 36722 65492 36728 65544
rect 36780 65532 36786 65544
rect 37016 65532 37044 65563
rect 37090 65560 37096 65612
rect 37148 65600 37154 65612
rect 37224 65609 37252 65640
rect 37642 65628 37648 65680
rect 37700 65668 37706 65680
rect 39390 65668 39396 65680
rect 37700 65640 39396 65668
rect 37700 65628 37706 65640
rect 39390 65628 39396 65640
rect 39448 65628 39454 65680
rect 37224 65603 37289 65609
rect 37148 65572 37193 65600
rect 37224 65572 37243 65603
rect 37148 65560 37154 65572
rect 37231 65569 37243 65572
rect 37277 65569 37289 65603
rect 37231 65563 37289 65569
rect 36780 65504 37044 65532
rect 36780 65492 36786 65504
rect 38562 65464 38568 65476
rect 36648 65436 38568 65464
rect 38562 65424 38568 65436
rect 38620 65424 38626 65476
rect 32858 65356 32864 65408
rect 32916 65356 32922 65408
rect 33229 65399 33287 65405
rect 33229 65365 33241 65399
rect 33275 65396 33287 65399
rect 34790 65396 34796 65408
rect 33275 65368 34796 65396
rect 33275 65365 33287 65368
rect 33229 65359 33287 65365
rect 34790 65356 34796 65368
rect 34848 65356 34854 65408
rect 34885 65399 34943 65405
rect 34885 65365 34897 65399
rect 34931 65396 34943 65399
rect 35434 65396 35440 65408
rect 34931 65368 35440 65396
rect 34931 65365 34943 65368
rect 34885 65359 34943 65365
rect 35434 65356 35440 65368
rect 35492 65356 35498 65408
rect 35526 65356 35532 65408
rect 35584 65396 35590 65408
rect 36170 65396 36176 65408
rect 35584 65368 35629 65396
rect 36131 65368 36176 65396
rect 35584 65356 35590 65368
rect 36170 65356 36176 65368
rect 36228 65356 36234 65408
rect 37369 65399 37427 65405
rect 37369 65365 37381 65399
rect 37415 65396 37427 65399
rect 39022 65396 39028 65408
rect 37415 65368 39028 65396
rect 37415 65365 37427 65368
rect 37369 65359 37427 65365
rect 39022 65356 39028 65368
rect 39080 65356 39086 65408
rect 1104 65306 38824 65328
rect 1104 65254 4246 65306
rect 4298 65254 4310 65306
rect 4362 65254 4374 65306
rect 4426 65254 4438 65306
rect 4490 65254 34966 65306
rect 35018 65254 35030 65306
rect 35082 65254 35094 65306
rect 35146 65254 35158 65306
rect 35210 65254 38824 65306
rect 1104 65232 38824 65254
rect 32953 65195 33011 65201
rect 32953 65161 32965 65195
rect 32999 65192 33011 65195
rect 34514 65192 34520 65204
rect 32999 65164 34520 65192
rect 32999 65161 33011 65164
rect 32953 65155 33011 65161
rect 34514 65152 34520 65164
rect 34572 65152 34578 65204
rect 35989 65195 36047 65201
rect 35989 65161 36001 65195
rect 36035 65192 36047 65195
rect 37182 65192 37188 65204
rect 36035 65164 37188 65192
rect 36035 65161 36047 65164
rect 35989 65155 36047 65161
rect 37182 65152 37188 65164
rect 37240 65152 37246 65204
rect 39666 65192 39672 65204
rect 37292 65164 39672 65192
rect 37093 65127 37151 65133
rect 37093 65124 37105 65127
rect 26206 65096 37105 65124
rect 26206 65068 26234 65096
rect 37093 65093 37105 65096
rect 37139 65093 37151 65127
rect 37093 65087 37151 65093
rect 26142 65016 26148 65068
rect 26200 65028 26234 65068
rect 26200 65016 26206 65028
rect 34606 65016 34612 65068
rect 34664 65056 34670 65068
rect 35158 65056 35164 65068
rect 34664 65028 35164 65056
rect 34664 65016 34670 65028
rect 35158 65016 35164 65028
rect 35216 65016 35222 65068
rect 37292 65056 37320 65164
rect 39666 65152 39672 65164
rect 39724 65152 39730 65204
rect 38105 65127 38163 65133
rect 38105 65093 38117 65127
rect 38151 65124 38163 65127
rect 39390 65124 39396 65136
rect 38151 65096 39396 65124
rect 38151 65093 38163 65096
rect 38105 65087 38163 65093
rect 39390 65084 39396 65096
rect 39448 65084 39454 65136
rect 39942 65056 39948 65068
rect 36556 65028 37320 65056
rect 37568 65028 39948 65056
rect 1394 64988 1400 65000
rect 1355 64960 1400 64988
rect 1394 64948 1400 64960
rect 1452 64948 1458 65000
rect 32861 64991 32919 64997
rect 32861 64957 32873 64991
rect 32907 64988 32919 64991
rect 33042 64988 33048 65000
rect 32907 64960 33048 64988
rect 32907 64957 32919 64960
rect 32861 64951 32919 64957
rect 33042 64948 33048 64960
rect 33100 64948 33106 65000
rect 34790 64988 34796 65000
rect 34751 64960 34796 64988
rect 34790 64948 34796 64960
rect 34848 64948 34854 65000
rect 35897 64991 35955 64997
rect 35897 64957 35909 64991
rect 35943 64988 35955 64991
rect 35986 64988 35992 65000
rect 35943 64960 35992 64988
rect 35943 64957 35955 64960
rect 35897 64951 35955 64957
rect 35986 64948 35992 64960
rect 36044 64948 36050 65000
rect 36556 64997 36584 65028
rect 36541 64991 36599 64997
rect 36541 64957 36553 64991
rect 36587 64957 36599 64991
rect 36541 64951 36599 64957
rect 36906 64948 36912 65000
rect 36964 64988 36970 65000
rect 37568 64997 37596 65028
rect 39942 65016 39948 65028
rect 40000 65016 40006 65068
rect 37553 64991 37611 64997
rect 36964 64960 37009 64988
rect 36964 64948 36970 64960
rect 37553 64957 37565 64991
rect 37599 64957 37611 64991
rect 37553 64951 37611 64957
rect 37921 64991 37979 64997
rect 37921 64957 37933 64991
rect 37967 64988 37979 64991
rect 38010 64988 38016 65000
rect 37967 64960 38016 64988
rect 37967 64957 37979 64960
rect 37921 64951 37979 64957
rect 38010 64948 38016 64960
rect 38068 64948 38074 65000
rect 32398 64880 32404 64932
rect 32456 64920 32462 64932
rect 32950 64920 32956 64932
rect 32456 64892 32956 64920
rect 32456 64880 32462 64892
rect 32950 64880 32956 64892
rect 33008 64880 33014 64932
rect 36722 64920 36728 64932
rect 36683 64892 36728 64920
rect 36722 64880 36728 64892
rect 36780 64880 36786 64932
rect 36817 64923 36875 64929
rect 36817 64889 36829 64923
rect 36863 64920 36875 64923
rect 37090 64920 37096 64932
rect 36863 64892 37096 64920
rect 36863 64889 36875 64892
rect 36817 64883 36875 64889
rect 37090 64880 37096 64892
rect 37148 64880 37154 64932
rect 37737 64923 37795 64929
rect 37737 64920 37749 64923
rect 37200 64892 37749 64920
rect 34606 64852 34612 64864
rect 34567 64824 34612 64852
rect 34606 64812 34612 64824
rect 34664 64812 34670 64864
rect 34790 64812 34796 64864
rect 34848 64852 34854 64864
rect 35342 64852 35348 64864
rect 34848 64824 35348 64852
rect 34848 64812 34854 64824
rect 35342 64812 35348 64824
rect 35400 64812 35406 64864
rect 36740 64852 36768 64880
rect 37200 64852 37228 64892
rect 37737 64889 37749 64892
rect 37783 64889 37795 64923
rect 37737 64883 37795 64889
rect 37829 64923 37887 64929
rect 37829 64889 37841 64923
rect 37875 64889 37887 64923
rect 37829 64883 37887 64889
rect 36740 64824 37228 64852
rect 37458 64812 37464 64864
rect 37516 64852 37522 64864
rect 37844 64852 37872 64883
rect 37516 64824 37872 64852
rect 37516 64812 37522 64824
rect 1104 64762 38824 64784
rect 1104 64710 19606 64762
rect 19658 64710 19670 64762
rect 19722 64710 19734 64762
rect 19786 64710 19798 64762
rect 19850 64710 38824 64762
rect 1104 64688 38824 64710
rect 35345 64651 35403 64657
rect 35345 64617 35357 64651
rect 35391 64648 35403 64651
rect 36262 64648 36268 64660
rect 35391 64620 36268 64648
rect 35391 64617 35403 64620
rect 35345 64611 35403 64617
rect 36262 64608 36268 64620
rect 36320 64608 36326 64660
rect 20162 64580 20168 64592
rect 20123 64552 20168 64580
rect 20162 64540 20168 64552
rect 20220 64540 20226 64592
rect 32490 64540 32496 64592
rect 32548 64580 32554 64592
rect 33137 64583 33195 64589
rect 33137 64580 33149 64583
rect 32548 64552 33149 64580
rect 32548 64540 32554 64552
rect 33137 64549 33149 64552
rect 33183 64549 33195 64583
rect 33137 64543 33195 64549
rect 35066 64540 35072 64592
rect 35124 64580 35130 64592
rect 36081 64583 36139 64589
rect 36081 64580 36093 64583
rect 35124 64552 35848 64580
rect 35124 64540 35130 64552
rect 1394 64512 1400 64524
rect 1355 64484 1400 64512
rect 1394 64472 1400 64484
rect 1452 64472 1458 64524
rect 31018 64472 31024 64524
rect 31076 64512 31082 64524
rect 31662 64512 31668 64524
rect 31076 64484 31668 64512
rect 31076 64472 31082 64484
rect 31662 64472 31668 64484
rect 31720 64472 31726 64524
rect 34146 64472 34152 64524
rect 34204 64512 34210 64524
rect 34701 64515 34759 64521
rect 34204 64484 34652 64512
rect 34204 64472 34210 64484
rect 3142 64336 3148 64388
rect 3200 64376 3206 64388
rect 28994 64376 29000 64388
rect 3200 64348 29000 64376
rect 3200 64336 3206 64348
rect 28994 64336 29000 64348
rect 29052 64336 29058 64388
rect 31849 64379 31907 64385
rect 31849 64345 31861 64379
rect 31895 64376 31907 64379
rect 34146 64376 34152 64388
rect 31895 64348 34152 64376
rect 31895 64345 31907 64348
rect 31849 64339 31907 64345
rect 34146 64336 34152 64348
rect 34204 64336 34210 64388
rect 34624 64376 34652 64484
rect 34701 64481 34713 64515
rect 34747 64481 34759 64515
rect 34701 64475 34759 64481
rect 34716 64444 34744 64475
rect 34882 64472 34888 64524
rect 34940 64512 34946 64524
rect 35820 64521 35848 64552
rect 35912 64552 36093 64580
rect 35161 64515 35219 64521
rect 35161 64512 35173 64515
rect 34940 64484 35173 64512
rect 34940 64472 34946 64484
rect 35161 64481 35173 64484
rect 35207 64481 35219 64515
rect 35161 64475 35219 64481
rect 35805 64515 35863 64521
rect 35805 64481 35817 64515
rect 35851 64481 35863 64515
rect 35805 64475 35863 64481
rect 35342 64444 35348 64456
rect 34716 64416 35348 64444
rect 35342 64404 35348 64416
rect 35400 64404 35406 64456
rect 35710 64376 35716 64388
rect 34624 64348 35716 64376
rect 35710 64336 35716 64348
rect 35768 64376 35774 64388
rect 35912 64376 35940 64552
rect 36081 64549 36093 64552
rect 36127 64549 36139 64583
rect 36081 64543 36139 64549
rect 36722 64540 36728 64592
rect 36780 64580 36786 64592
rect 37001 64583 37059 64589
rect 37001 64580 37013 64583
rect 36780 64552 37013 64580
rect 36780 64540 36786 64552
rect 37001 64549 37013 64552
rect 37047 64549 37059 64583
rect 37001 64543 37059 64549
rect 37090 64540 37096 64592
rect 37148 64580 37154 64592
rect 37458 64580 37464 64592
rect 37148 64552 37464 64580
rect 37148 64540 37154 64552
rect 37458 64540 37464 64552
rect 37516 64540 37522 64592
rect 35986 64472 35992 64524
rect 36044 64512 36050 64524
rect 36173 64515 36231 64521
rect 36044 64484 36089 64512
rect 36044 64472 36050 64484
rect 36173 64481 36185 64515
rect 36219 64481 36231 64515
rect 36173 64475 36231 64481
rect 36817 64515 36875 64521
rect 36817 64481 36829 64515
rect 36863 64512 36875 64515
rect 36906 64512 36912 64524
rect 36863 64484 36912 64512
rect 36863 64481 36875 64484
rect 36817 64475 36875 64481
rect 35768 64348 35940 64376
rect 35768 64336 35774 64348
rect 17310 64268 17316 64320
rect 17368 64308 17374 64320
rect 20257 64311 20315 64317
rect 20257 64308 20269 64311
rect 17368 64280 20269 64308
rect 17368 64268 17374 64280
rect 20257 64277 20269 64280
rect 20303 64277 20315 64311
rect 20257 64271 20315 64277
rect 33134 64268 33140 64320
rect 33192 64308 33198 64320
rect 33229 64311 33287 64317
rect 33229 64308 33241 64311
rect 33192 64280 33241 64308
rect 33192 64268 33198 64280
rect 33229 64277 33241 64280
rect 33275 64277 33287 64311
rect 33229 64271 33287 64277
rect 34517 64311 34575 64317
rect 34517 64277 34529 64311
rect 34563 64308 34575 64311
rect 36188 64308 36216 64475
rect 36906 64472 36912 64484
rect 36964 64472 36970 64524
rect 37185 64515 37243 64521
rect 37185 64481 37197 64515
rect 37231 64512 37243 64515
rect 37550 64512 37556 64524
rect 37231 64484 37556 64512
rect 37231 64481 37243 64484
rect 37185 64475 37243 64481
rect 37550 64472 37556 64484
rect 37608 64472 37614 64524
rect 36262 64404 36268 64456
rect 36320 64444 36326 64456
rect 37642 64444 37648 64456
rect 36320 64416 37648 64444
rect 36320 64404 36326 64416
rect 37642 64404 37648 64416
rect 37700 64404 37706 64456
rect 36354 64308 36360 64320
rect 34563 64280 36216 64308
rect 36315 64280 36360 64308
rect 34563 64277 34575 64280
rect 34517 64271 34575 64277
rect 36354 64268 36360 64280
rect 36412 64268 36418 64320
rect 37369 64311 37427 64317
rect 37369 64277 37381 64311
rect 37415 64308 37427 64311
rect 38562 64308 38568 64320
rect 37415 64280 38568 64308
rect 37415 64277 37427 64280
rect 37369 64271 37427 64277
rect 38562 64268 38568 64280
rect 38620 64268 38626 64320
rect 1104 64218 38824 64240
rect 1104 64166 4246 64218
rect 4298 64166 4310 64218
rect 4362 64166 4374 64218
rect 4426 64166 4438 64218
rect 4490 64166 34966 64218
rect 35018 64166 35030 64218
rect 35082 64166 35094 64218
rect 35146 64166 35158 64218
rect 35210 64166 38824 64218
rect 1104 64144 38824 64166
rect 37274 64104 37280 64116
rect 36648 64076 37280 64104
rect 36081 64039 36139 64045
rect 36081 64005 36093 64039
rect 36127 64036 36139 64039
rect 36648 64036 36676 64076
rect 37274 64064 37280 64076
rect 37332 64064 37338 64116
rect 37550 64064 37556 64116
rect 37608 64104 37614 64116
rect 39850 64104 39856 64116
rect 37608 64076 39856 64104
rect 37608 64064 37614 64076
rect 39850 64064 39856 64076
rect 39908 64064 39914 64116
rect 36127 64008 36676 64036
rect 36127 64005 36139 64008
rect 36081 63999 36139 64005
rect 39482 63968 39488 63980
rect 36740 63940 39488 63968
rect 34790 63900 34796 63912
rect 34751 63872 34796 63900
rect 34790 63860 34796 63872
rect 34848 63860 34854 63912
rect 34974 63860 34980 63912
rect 35032 63900 35038 63912
rect 35342 63900 35348 63912
rect 35032 63872 35348 63900
rect 35032 63860 35038 63872
rect 35342 63860 35348 63872
rect 35400 63900 35406 63912
rect 35802 63900 35808 63912
rect 35400 63872 35808 63900
rect 35400 63860 35406 63872
rect 35802 63860 35808 63872
rect 35860 63900 35866 63912
rect 35897 63903 35955 63909
rect 35897 63900 35909 63903
rect 35860 63872 35909 63900
rect 35860 63860 35866 63872
rect 35897 63869 35909 63872
rect 35943 63869 35955 63903
rect 35897 63863 35955 63869
rect 36541 63903 36599 63909
rect 36541 63869 36553 63903
rect 36587 63900 36599 63903
rect 36740 63900 36768 63940
rect 39482 63928 39488 63940
rect 39540 63928 39546 63980
rect 36906 63900 36912 63912
rect 36587 63872 36768 63900
rect 36867 63872 36912 63900
rect 36587 63869 36599 63872
rect 36541 63863 36599 63869
rect 36906 63860 36912 63872
rect 36964 63860 36970 63912
rect 37550 63900 37556 63912
rect 37511 63872 37556 63900
rect 37550 63860 37556 63872
rect 37608 63860 37614 63912
rect 37642 63860 37648 63912
rect 37700 63900 37706 63912
rect 37737 63903 37795 63909
rect 37737 63900 37749 63903
rect 37700 63872 37749 63900
rect 37700 63860 37706 63872
rect 37737 63869 37749 63872
rect 37783 63869 37795 63903
rect 37918 63900 37924 63912
rect 37879 63872 37924 63900
rect 37737 63863 37795 63869
rect 37918 63860 37924 63872
rect 37976 63860 37982 63912
rect 35986 63792 35992 63844
rect 36044 63832 36050 63844
rect 36725 63835 36783 63841
rect 36725 63832 36737 63835
rect 36044 63804 36737 63832
rect 36044 63792 36050 63804
rect 36725 63801 36737 63804
rect 36771 63801 36783 63835
rect 36725 63795 36783 63801
rect 36817 63835 36875 63841
rect 36817 63801 36829 63835
rect 36863 63801 36875 63835
rect 36817 63795 36875 63801
rect 34606 63764 34612 63776
rect 34567 63736 34612 63764
rect 34606 63724 34612 63736
rect 34664 63724 34670 63776
rect 35710 63724 35716 63776
rect 35768 63764 35774 63776
rect 36832 63764 36860 63795
rect 37458 63792 37464 63844
rect 37516 63832 37522 63844
rect 37829 63835 37887 63841
rect 37829 63832 37841 63835
rect 37516 63804 37841 63832
rect 37516 63792 37522 63804
rect 37829 63801 37841 63804
rect 37875 63801 37887 63835
rect 37829 63795 37887 63801
rect 38838 63792 38844 63844
rect 38896 63832 38902 63844
rect 38896 63804 38976 63832
rect 38896 63792 38902 63804
rect 37090 63764 37096 63776
rect 35768 63736 36860 63764
rect 37051 63736 37096 63764
rect 35768 63724 35774 63736
rect 37090 63724 37096 63736
rect 37148 63724 37154 63776
rect 38102 63764 38108 63776
rect 38063 63736 38108 63764
rect 38102 63724 38108 63736
rect 38160 63724 38166 63776
rect 1104 63674 38824 63696
rect 1104 63622 19606 63674
rect 19658 63622 19670 63674
rect 19722 63622 19734 63674
rect 19786 63622 19798 63674
rect 19850 63622 38824 63674
rect 38948 63640 38976 63804
rect 1104 63600 38824 63622
rect 38930 63588 38936 63640
rect 38988 63588 38994 63640
rect 34701 63563 34759 63569
rect 34701 63529 34713 63563
rect 34747 63560 34759 63563
rect 35802 63560 35808 63572
rect 34747 63532 35808 63560
rect 34747 63529 34759 63532
rect 34701 63523 34759 63529
rect 35802 63520 35808 63532
rect 35860 63520 35866 63572
rect 35986 63520 35992 63572
rect 36044 63560 36050 63572
rect 36446 63560 36452 63572
rect 36044 63532 36452 63560
rect 36044 63520 36050 63532
rect 36446 63520 36452 63532
rect 36504 63560 36510 63572
rect 36504 63532 37044 63560
rect 36504 63520 36510 63532
rect 1394 63424 1400 63436
rect 1355 63396 1400 63424
rect 1394 63384 1400 63396
rect 1452 63384 1458 63436
rect 34517 63427 34575 63433
rect 34517 63393 34529 63427
rect 34563 63424 34575 63427
rect 34974 63424 34980 63436
rect 34563 63396 34980 63424
rect 34563 63393 34575 63396
rect 34517 63387 34575 63393
rect 34974 63384 34980 63396
rect 35032 63384 35038 63436
rect 35158 63424 35164 63436
rect 35119 63396 35164 63424
rect 35158 63384 35164 63396
rect 35216 63424 35222 63436
rect 35526 63424 35532 63436
rect 35216 63396 35532 63424
rect 35216 63384 35222 63396
rect 35526 63384 35532 63396
rect 35584 63384 35590 63436
rect 35802 63424 35808 63436
rect 35763 63396 35808 63424
rect 35802 63384 35808 63396
rect 35860 63384 35866 63436
rect 36004 63433 36032 63520
rect 36081 63495 36139 63501
rect 36081 63461 36093 63495
rect 36127 63492 36139 63495
rect 36722 63492 36728 63504
rect 36127 63464 36728 63492
rect 36127 63461 36139 63464
rect 36081 63455 36139 63461
rect 35989 63427 36047 63433
rect 35989 63393 36001 63427
rect 36035 63393 36047 63427
rect 36170 63424 36176 63436
rect 36131 63396 36176 63424
rect 35989 63387 36047 63393
rect 36170 63384 36176 63396
rect 36228 63384 36234 63436
rect 35710 63316 35716 63368
rect 35768 63356 35774 63368
rect 36280 63356 36308 63464
rect 36722 63452 36728 63464
rect 36780 63492 36786 63504
rect 37016 63501 37044 63532
rect 37001 63495 37059 63501
rect 36780 63464 36952 63492
rect 36780 63452 36786 63464
rect 36817 63427 36875 63433
rect 36817 63393 36829 63427
rect 36863 63393 36875 63427
rect 36924 63424 36952 63464
rect 37001 63461 37013 63495
rect 37047 63461 37059 63495
rect 37001 63455 37059 63461
rect 37550 63452 37556 63504
rect 37608 63492 37614 63504
rect 38378 63492 38384 63504
rect 37608 63464 38384 63492
rect 37608 63452 37614 63464
rect 38378 63452 38384 63464
rect 38436 63452 38442 63504
rect 37093 63427 37151 63433
rect 37093 63424 37105 63427
rect 36924 63396 37105 63424
rect 36817 63387 36875 63393
rect 37093 63393 37105 63396
rect 37139 63393 37151 63427
rect 37093 63387 37151 63393
rect 37185 63427 37243 63433
rect 37185 63393 37197 63427
rect 37231 63424 37243 63427
rect 37274 63424 37280 63436
rect 37231 63396 37280 63424
rect 37231 63393 37243 63396
rect 37185 63387 37243 63393
rect 35768 63328 36308 63356
rect 36832 63356 36860 63387
rect 37274 63384 37280 63396
rect 37332 63384 37338 63436
rect 38746 63356 38752 63368
rect 36832 63328 38752 63356
rect 35768 63316 35774 63328
rect 38746 63316 38752 63328
rect 38804 63316 38810 63368
rect 37458 63288 37464 63300
rect 35728 63260 37464 63288
rect 35345 63223 35403 63229
rect 35345 63189 35357 63223
rect 35391 63220 35403 63223
rect 35728 63220 35756 63260
rect 37458 63248 37464 63260
rect 37516 63248 37522 63300
rect 35391 63192 35756 63220
rect 35391 63189 35403 63192
rect 35345 63183 35403 63189
rect 35802 63180 35808 63232
rect 35860 63220 35866 63232
rect 36357 63223 36415 63229
rect 36357 63220 36369 63223
rect 35860 63192 36369 63220
rect 35860 63180 35866 63192
rect 36357 63189 36369 63192
rect 36403 63189 36415 63223
rect 36357 63183 36415 63189
rect 37369 63223 37427 63229
rect 37369 63189 37381 63223
rect 37415 63220 37427 63223
rect 38286 63220 38292 63232
rect 37415 63192 38292 63220
rect 37415 63189 37427 63192
rect 37369 63183 37427 63189
rect 38286 63180 38292 63192
rect 38344 63180 38350 63232
rect 1104 63130 38824 63152
rect 1104 63078 4246 63130
rect 4298 63078 4310 63130
rect 4362 63078 4374 63130
rect 4426 63078 4438 63130
rect 4490 63078 34966 63130
rect 35018 63078 35030 63130
rect 35082 63078 35094 63130
rect 35146 63078 35158 63130
rect 35210 63078 38824 63130
rect 1104 63056 38824 63078
rect 36538 62976 36544 63028
rect 36596 63016 36602 63028
rect 36906 63016 36912 63028
rect 36596 62988 36912 63016
rect 36596 62976 36602 62988
rect 36906 62976 36912 62988
rect 36964 62976 36970 63028
rect 37274 62908 37280 62960
rect 37332 62948 37338 62960
rect 37550 62948 37556 62960
rect 37332 62920 37556 62948
rect 37332 62908 37338 62920
rect 32490 62840 32496 62892
rect 32548 62880 32554 62892
rect 32548 62852 32720 62880
rect 32548 62840 32554 62852
rect 1394 62812 1400 62824
rect 1355 62784 1400 62812
rect 1394 62772 1400 62784
rect 1452 62772 1458 62824
rect 31662 62772 31668 62824
rect 31720 62812 31726 62824
rect 32692 62821 32720 62852
rect 34606 62840 34612 62892
rect 34664 62880 34670 62892
rect 34664 62852 36400 62880
rect 34664 62840 34670 62852
rect 31849 62815 31907 62821
rect 31849 62812 31861 62815
rect 31720 62784 31861 62812
rect 31720 62772 31726 62784
rect 31849 62781 31861 62784
rect 31895 62781 31907 62815
rect 31849 62775 31907 62781
rect 32677 62815 32735 62821
rect 32677 62781 32689 62815
rect 32723 62781 32735 62815
rect 36078 62812 36084 62824
rect 36039 62784 36084 62812
rect 32677 62775 32735 62781
rect 36078 62772 36084 62784
rect 36136 62772 36142 62824
rect 36372 62812 36400 62852
rect 36630 62840 36636 62892
rect 36688 62880 36694 62892
rect 36688 62852 37320 62880
rect 36688 62840 36694 62852
rect 37292 62821 37320 62852
rect 37384 62821 37412 62920
rect 37550 62908 37556 62920
rect 37608 62908 37614 62960
rect 37645 62951 37703 62957
rect 37645 62917 37657 62951
rect 37691 62948 37703 62951
rect 38746 62948 38752 62960
rect 37691 62920 38752 62948
rect 37691 62917 37703 62920
rect 37645 62911 37703 62917
rect 38746 62908 38752 62920
rect 38804 62908 38810 62960
rect 36449 62815 36507 62821
rect 36449 62812 36461 62815
rect 36372 62784 36461 62812
rect 36449 62781 36461 62784
rect 36495 62781 36507 62815
rect 36449 62775 36507 62781
rect 37093 62815 37151 62821
rect 37093 62781 37105 62815
rect 37139 62781 37151 62815
rect 37093 62775 37151 62781
rect 37277 62815 37335 62821
rect 37277 62781 37289 62815
rect 37323 62781 37335 62815
rect 37277 62775 37335 62781
rect 37369 62815 37427 62821
rect 37369 62781 37381 62815
rect 37415 62781 37427 62815
rect 37369 62775 37427 62781
rect 32033 62747 32091 62753
rect 32033 62713 32045 62747
rect 32079 62744 32091 62747
rect 32490 62744 32496 62756
rect 32079 62716 32496 62744
rect 32079 62713 32091 62716
rect 32033 62707 32091 62713
rect 32490 62704 32496 62716
rect 32548 62704 32554 62756
rect 32861 62747 32919 62753
rect 32861 62713 32873 62747
rect 32907 62744 32919 62747
rect 33594 62744 33600 62756
rect 32907 62716 33600 62744
rect 32907 62713 32919 62716
rect 32861 62707 32919 62713
rect 33594 62704 33600 62716
rect 33652 62704 33658 62756
rect 36265 62747 36323 62753
rect 36265 62713 36277 62747
rect 36311 62713 36323 62747
rect 36265 62707 36323 62713
rect 36357 62747 36415 62753
rect 36357 62713 36369 62747
rect 36403 62744 36415 62747
rect 36722 62744 36728 62756
rect 36403 62716 36728 62744
rect 36403 62713 36415 62716
rect 36357 62707 36415 62713
rect 36280 62676 36308 62707
rect 36722 62704 36728 62716
rect 36780 62704 36786 62756
rect 36446 62676 36452 62688
rect 36280 62648 36452 62676
rect 36446 62636 36452 62648
rect 36504 62636 36510 62688
rect 36630 62676 36636 62688
rect 36591 62648 36636 62676
rect 36630 62636 36636 62648
rect 36688 62636 36694 62688
rect 37113 62676 37141 62775
rect 37458 62772 37464 62824
rect 37516 62821 37522 62824
rect 37516 62812 37524 62821
rect 37516 62784 37561 62812
rect 37516 62775 37524 62784
rect 37516 62772 37522 62775
rect 37642 62676 37648 62688
rect 37113 62648 37648 62676
rect 37642 62636 37648 62648
rect 37700 62636 37706 62688
rect 1104 62586 38824 62608
rect 1104 62534 19606 62586
rect 19658 62534 19670 62586
rect 19722 62534 19734 62586
rect 19786 62534 19798 62586
rect 19850 62534 38824 62586
rect 1104 62512 38824 62534
rect 35437 62475 35495 62481
rect 35437 62441 35449 62475
rect 35483 62472 35495 62475
rect 37458 62472 37464 62484
rect 35483 62444 37464 62472
rect 35483 62441 35495 62444
rect 35437 62435 35495 62441
rect 37458 62432 37464 62444
rect 37516 62432 37522 62484
rect 36538 62364 36544 62416
rect 36596 62404 36602 62416
rect 36909 62407 36967 62413
rect 36909 62404 36921 62407
rect 36596 62376 36921 62404
rect 36596 62364 36602 62376
rect 36909 62373 36921 62376
rect 36955 62404 36967 62407
rect 37274 62404 37280 62416
rect 36955 62376 37280 62404
rect 36955 62373 36967 62376
rect 36909 62367 36967 62373
rect 37274 62364 37280 62376
rect 37332 62364 37338 62416
rect 15378 62336 15384 62348
rect 15339 62308 15384 62336
rect 15378 62296 15384 62308
rect 15436 62296 15442 62348
rect 35621 62339 35679 62345
rect 35621 62305 35633 62339
rect 35667 62336 35679 62339
rect 35710 62336 35716 62348
rect 35667 62308 35716 62336
rect 35667 62305 35679 62308
rect 35621 62299 35679 62305
rect 35710 62296 35716 62308
rect 35768 62296 35774 62348
rect 36262 62336 36268 62348
rect 36223 62308 36268 62336
rect 36262 62296 36268 62308
rect 36320 62296 36326 62348
rect 36725 62339 36783 62345
rect 36725 62305 36737 62339
rect 36771 62336 36783 62339
rect 37001 62339 37059 62345
rect 36771 62308 36952 62336
rect 36771 62305 36783 62308
rect 36725 62299 36783 62305
rect 36081 62203 36139 62209
rect 36081 62169 36093 62203
rect 36127 62200 36139 62203
rect 36722 62200 36728 62212
rect 36127 62172 36728 62200
rect 36127 62169 36139 62172
rect 36081 62163 36139 62169
rect 36722 62160 36728 62172
rect 36780 62160 36786 62212
rect 36924 62200 36952 62308
rect 37001 62305 37013 62339
rect 37047 62305 37059 62339
rect 37001 62299 37059 62305
rect 37145 62339 37203 62345
rect 37145 62305 37157 62339
rect 37191 62336 37203 62339
rect 37458 62336 37464 62348
rect 37191 62308 37464 62336
rect 37191 62305 37203 62308
rect 37145 62299 37203 62305
rect 37016 62268 37044 62299
rect 37458 62296 37464 62308
rect 37516 62296 37522 62348
rect 37550 62268 37556 62280
rect 37016 62240 37556 62268
rect 37550 62228 37556 62240
rect 37608 62228 37614 62280
rect 39114 62200 39120 62212
rect 36924 62172 39120 62200
rect 39114 62160 39120 62172
rect 39172 62160 39178 62212
rect 3694 62092 3700 62144
rect 3752 62132 3758 62144
rect 15473 62135 15531 62141
rect 15473 62132 15485 62135
rect 3752 62104 15485 62132
rect 3752 62092 3758 62104
rect 15473 62101 15485 62104
rect 15519 62101 15531 62135
rect 15473 62095 15531 62101
rect 36170 62092 36176 62144
rect 36228 62132 36234 62144
rect 37277 62135 37335 62141
rect 37277 62132 37289 62135
rect 36228 62104 37289 62132
rect 36228 62092 36234 62104
rect 37277 62101 37289 62104
rect 37323 62101 37335 62135
rect 37277 62095 37335 62101
rect 1104 62042 38824 62064
rect 1104 61990 4246 62042
rect 4298 61990 4310 62042
rect 4362 61990 4374 62042
rect 4426 61990 4438 62042
rect 4490 61990 34966 62042
rect 35018 61990 35030 62042
rect 35082 61990 35094 62042
rect 35146 61990 35158 62042
rect 35210 61990 38824 62042
rect 1104 61968 38824 61990
rect 35805 61863 35863 61869
rect 35805 61829 35817 61863
rect 35851 61860 35863 61863
rect 37458 61860 37464 61872
rect 35851 61832 37464 61860
rect 35851 61829 35863 61832
rect 35805 61823 35863 61829
rect 37458 61820 37464 61832
rect 37516 61820 37522 61872
rect 37645 61863 37703 61869
rect 37645 61829 37657 61863
rect 37691 61860 37703 61863
rect 37734 61860 37740 61872
rect 37691 61832 37740 61860
rect 37691 61829 37703 61832
rect 37645 61823 37703 61829
rect 37734 61820 37740 61832
rect 37792 61820 37798 61872
rect 37366 61752 37372 61804
rect 37424 61752 37430 61804
rect 1394 61724 1400 61736
rect 1355 61696 1400 61724
rect 1394 61684 1400 61696
rect 1452 61684 1458 61736
rect 35802 61684 35808 61736
rect 35860 61724 35866 61736
rect 35989 61727 36047 61733
rect 35989 61724 36001 61727
rect 35860 61696 36001 61724
rect 35860 61684 35866 61696
rect 35989 61693 36001 61696
rect 36035 61693 36047 61727
rect 35989 61687 36047 61693
rect 36633 61727 36691 61733
rect 36633 61693 36645 61727
rect 36679 61724 36691 61727
rect 36722 61724 36728 61736
rect 36679 61696 36728 61724
rect 36679 61693 36691 61696
rect 36633 61687 36691 61693
rect 36722 61684 36728 61696
rect 36780 61684 36786 61736
rect 37093 61727 37151 61733
rect 37093 61693 37105 61727
rect 37139 61724 37151 61727
rect 37384 61724 37412 61752
rect 37139 61696 37412 61724
rect 37466 61727 37524 61733
rect 37139 61693 37151 61696
rect 37093 61687 37151 61693
rect 37466 61693 37478 61727
rect 37512 61724 37524 61727
rect 37512 61696 37688 61724
rect 37512 61693 37524 61696
rect 37466 61687 37524 61693
rect 35526 61616 35532 61668
rect 35584 61656 35590 61668
rect 36538 61656 36544 61668
rect 35584 61628 36544 61656
rect 35584 61616 35590 61628
rect 36538 61616 36544 61628
rect 36596 61616 36602 61668
rect 37274 61656 37280 61668
rect 37235 61628 37280 61656
rect 37274 61616 37280 61628
rect 37332 61616 37338 61668
rect 37369 61659 37427 61665
rect 37369 61625 37381 61659
rect 37415 61656 37427 61659
rect 37550 61656 37556 61668
rect 37415 61628 37556 61656
rect 37415 61625 37427 61628
rect 37369 61619 37427 61625
rect 37550 61616 37556 61628
rect 37608 61616 37614 61668
rect 36449 61591 36507 61597
rect 36449 61557 36461 61591
rect 36495 61588 36507 61591
rect 37660 61588 37688 61696
rect 36495 61560 37688 61588
rect 36495 61557 36507 61560
rect 36449 61551 36507 61557
rect 1104 61498 38824 61520
rect 1104 61446 19606 61498
rect 19658 61446 19670 61498
rect 19722 61446 19734 61498
rect 19786 61446 19798 61498
rect 19850 61446 38824 61498
rect 1104 61424 38824 61446
rect 35434 61344 35440 61396
rect 35492 61384 35498 61396
rect 36173 61387 36231 61393
rect 36173 61384 36185 61387
rect 35492 61356 36185 61384
rect 35492 61344 35498 61356
rect 36173 61353 36185 61356
rect 36219 61353 36231 61387
rect 37550 61384 37556 61396
rect 36173 61347 36231 61353
rect 36832 61356 37556 61384
rect 1394 61248 1400 61260
rect 1355 61220 1400 61248
rect 1394 61208 1400 61220
rect 1452 61208 1458 61260
rect 34882 61248 34888 61260
rect 34843 61220 34888 61248
rect 34882 61208 34888 61220
rect 34940 61208 34946 61260
rect 35526 61248 35532 61260
rect 35487 61220 35532 61248
rect 35526 61208 35532 61220
rect 35584 61208 35590 61260
rect 35989 61251 36047 61257
rect 35989 61217 36001 61251
rect 36035 61248 36047 61251
rect 36262 61248 36268 61260
rect 36035 61220 36268 61248
rect 36035 61217 36047 61220
rect 35989 61211 36047 61217
rect 36262 61208 36268 61220
rect 36320 61208 36326 61260
rect 36722 61248 36728 61260
rect 36683 61220 36728 61248
rect 36722 61208 36728 61220
rect 36780 61208 36786 61260
rect 36832 61248 36860 61356
rect 37550 61344 37556 61356
rect 37608 61344 37614 61396
rect 36909 61319 36967 61325
rect 36909 61285 36921 61319
rect 36955 61316 36967 61319
rect 37274 61316 37280 61328
rect 36955 61288 37280 61316
rect 36955 61285 36967 61288
rect 36909 61279 36967 61285
rect 37274 61276 37280 61288
rect 37332 61276 37338 61328
rect 37001 61251 37059 61257
rect 37001 61248 37013 61251
rect 36832 61220 37013 61248
rect 37001 61217 37013 61220
rect 37047 61217 37059 61251
rect 37001 61211 37059 61217
rect 37098 61251 37156 61257
rect 37098 61217 37110 61251
rect 37144 61217 37156 61251
rect 37098 61211 37156 61217
rect 37108 61180 37136 61211
rect 34716 61152 37136 61180
rect 34716 61121 34744 61152
rect 34701 61115 34759 61121
rect 34701 61081 34713 61115
rect 34747 61081 34759 61115
rect 37277 61115 37335 61121
rect 37277 61112 37289 61115
rect 34701 61075 34759 61081
rect 34808 61084 37289 61112
rect 33042 61004 33048 61056
rect 33100 61044 33106 61056
rect 34808 61044 34836 61084
rect 37277 61081 37289 61084
rect 37323 61081 37335 61115
rect 37277 61075 37335 61081
rect 35342 61044 35348 61056
rect 33100 61016 34836 61044
rect 35303 61016 35348 61044
rect 33100 61004 33106 61016
rect 35342 61004 35348 61016
rect 35400 61004 35406 61056
rect 36722 61004 36728 61056
rect 36780 61044 36786 61056
rect 39574 61044 39580 61056
rect 36780 61016 39580 61044
rect 36780 61004 36786 61016
rect 39574 61004 39580 61016
rect 39632 61004 39638 61056
rect 1104 60954 38824 60976
rect 1104 60902 4246 60954
rect 4298 60902 4310 60954
rect 4362 60902 4374 60954
rect 4426 60902 4438 60954
rect 4490 60902 34966 60954
rect 35018 60902 35030 60954
rect 35082 60902 35094 60954
rect 35146 60902 35158 60954
rect 35210 60902 38824 60954
rect 1104 60880 38824 60902
rect 28534 60732 28540 60784
rect 28592 60772 28598 60784
rect 34882 60772 34888 60784
rect 28592 60744 34888 60772
rect 28592 60732 28598 60744
rect 34882 60732 34888 60744
rect 34940 60732 34946 60784
rect 35158 60732 35164 60784
rect 35216 60772 35222 60784
rect 35526 60772 35532 60784
rect 35216 60744 35532 60772
rect 35216 60732 35222 60744
rect 35526 60732 35532 60744
rect 35584 60732 35590 60784
rect 37645 60775 37703 60781
rect 37645 60772 37657 60775
rect 35636 60744 37657 60772
rect 32674 60664 32680 60716
rect 32732 60704 32738 60716
rect 35636 60704 35664 60744
rect 37645 60741 37657 60744
rect 37691 60741 37703 60775
rect 37645 60735 37703 60741
rect 36538 60704 36544 60716
rect 32732 60676 35664 60704
rect 36280 60676 36544 60704
rect 32732 60664 32738 60676
rect 35250 60596 35256 60648
rect 35308 60636 35314 60648
rect 35526 60636 35532 60648
rect 35308 60608 35532 60636
rect 35308 60596 35314 60608
rect 35526 60596 35532 60608
rect 35584 60596 35590 60648
rect 35986 60636 35992 60648
rect 35947 60608 35992 60636
rect 35986 60596 35992 60608
rect 36044 60596 36050 60648
rect 36280 60645 36308 60676
rect 36538 60664 36544 60676
rect 36596 60704 36602 60716
rect 36722 60704 36728 60716
rect 36596 60676 36728 60704
rect 36596 60664 36602 60676
rect 36722 60664 36728 60676
rect 36780 60664 36786 60716
rect 36446 60645 36452 60648
rect 36265 60639 36323 60645
rect 36265 60605 36277 60639
rect 36311 60605 36323 60639
rect 36265 60599 36323 60605
rect 36409 60639 36452 60645
rect 36409 60605 36421 60639
rect 36409 60599 36452 60605
rect 36446 60596 36452 60599
rect 36504 60596 36510 60648
rect 36906 60596 36912 60648
rect 36964 60636 36970 60648
rect 37093 60639 37151 60645
rect 37093 60636 37105 60639
rect 36964 60608 37105 60636
rect 36964 60596 36970 60608
rect 37093 60605 37105 60608
rect 37139 60605 37151 60639
rect 37274 60636 37280 60648
rect 37235 60608 37280 60636
rect 37093 60599 37151 60605
rect 37274 60596 37280 60608
rect 37332 60596 37338 60648
rect 37458 60596 37464 60648
rect 37516 60645 37522 60648
rect 37516 60636 37524 60645
rect 37516 60608 37561 60636
rect 37516 60599 37524 60608
rect 37516 60596 37522 60599
rect 35434 60528 35440 60580
rect 35492 60568 35498 60580
rect 36173 60571 36231 60577
rect 36173 60568 36185 60571
rect 35492 60540 36185 60568
rect 35492 60528 35498 60540
rect 36173 60537 36185 60540
rect 36219 60537 36231 60571
rect 36173 60531 36231 60537
rect 37369 60571 37427 60577
rect 37369 60537 37381 60571
rect 37415 60568 37427 60571
rect 37550 60568 37556 60580
rect 37415 60540 37556 60568
rect 37415 60537 37427 60540
rect 37369 60531 37427 60537
rect 37550 60528 37556 60540
rect 37608 60528 37614 60580
rect 36538 60500 36544 60512
rect 36596 60509 36602 60512
rect 36507 60472 36544 60500
rect 36538 60460 36544 60472
rect 36596 60463 36607 60509
rect 36596 60460 36602 60463
rect 1104 60410 38824 60432
rect 1104 60358 19606 60410
rect 19658 60358 19670 60410
rect 19722 60358 19734 60410
rect 19786 60358 19798 60410
rect 19850 60358 38824 60410
rect 1104 60336 38824 60358
rect 33134 60256 33140 60308
rect 33192 60296 33198 60308
rect 33192 60268 33456 60296
rect 33192 60256 33198 60268
rect 33428 60237 33456 60268
rect 35342 60256 35348 60308
rect 35400 60296 35406 60308
rect 35400 60268 37504 60296
rect 35400 60256 35406 60268
rect 33413 60231 33471 60237
rect 33413 60197 33425 60231
rect 33459 60197 33471 60231
rect 33413 60191 33471 60197
rect 34514 60188 34520 60240
rect 34572 60228 34578 60240
rect 35897 60231 35955 60237
rect 35897 60228 35909 60231
rect 34572 60200 35909 60228
rect 34572 60188 34578 60200
rect 35897 60197 35909 60200
rect 35943 60228 35955 60231
rect 37002 60231 37060 60237
rect 37002 60228 37014 60231
rect 35943 60200 37014 60228
rect 35943 60197 35955 60200
rect 35897 60191 35955 60197
rect 37002 60197 37014 60200
rect 37048 60228 37060 60231
rect 37366 60228 37372 60240
rect 37048 60200 37372 60228
rect 37048 60197 37060 60200
rect 37002 60191 37060 60197
rect 37366 60188 37372 60200
rect 37424 60188 37430 60240
rect 1394 60160 1400 60172
rect 1355 60132 1400 60160
rect 1394 60120 1400 60132
rect 1452 60120 1458 60172
rect 16574 60120 16580 60172
rect 16632 60160 16638 60172
rect 33045 60163 33103 60169
rect 33045 60160 33057 60163
rect 16632 60132 33057 60160
rect 16632 60120 16638 60132
rect 33045 60129 33057 60132
rect 33091 60129 33103 60163
rect 33045 60123 33103 60129
rect 33193 60163 33251 60169
rect 33193 60129 33205 60163
rect 33239 60160 33251 60163
rect 33321 60163 33379 60169
rect 33239 60129 33272 60160
rect 33193 60123 33272 60129
rect 33321 60129 33333 60163
rect 33367 60129 33379 60163
rect 33321 60123 33379 60129
rect 33551 60163 33609 60169
rect 33551 60129 33563 60163
rect 33597 60160 33609 60163
rect 34054 60160 34060 60172
rect 33597 60132 34060 60160
rect 33597 60129 33609 60132
rect 33551 60123 33609 60129
rect 33244 60024 33272 60123
rect 33336 60092 33364 60123
rect 34054 60120 34060 60132
rect 34112 60120 34118 60172
rect 35158 60160 35164 60172
rect 35119 60132 35164 60160
rect 35158 60120 35164 60132
rect 35216 60120 35222 60172
rect 35618 60160 35624 60172
rect 35579 60132 35624 60160
rect 35618 60120 35624 60132
rect 35676 60120 35682 60172
rect 35805 60163 35863 60169
rect 35805 60129 35817 60163
rect 35851 60129 35863 60163
rect 35805 60123 35863 60129
rect 34146 60092 34152 60104
rect 33336 60064 34152 60092
rect 34146 60052 34152 60064
rect 34204 60052 34210 60104
rect 35820 60092 35848 60123
rect 35986 60120 35992 60172
rect 36044 60169 36050 60172
rect 36044 60160 36052 60169
rect 36745 60163 36803 60169
rect 36745 60160 36757 60163
rect 36044 60132 36089 60160
rect 36044 60123 36052 60132
rect 36740 60129 36757 60160
rect 36791 60129 36803 60163
rect 36740 60123 36803 60129
rect 36909 60163 36967 60169
rect 36909 60129 36921 60163
rect 36955 60129 36967 60163
rect 36909 60123 36967 60129
rect 37145 60163 37203 60169
rect 37145 60129 37157 60163
rect 37191 60160 37203 60163
rect 37476 60160 37504 60268
rect 37191 60132 37504 60160
rect 37191 60129 37203 60132
rect 37145 60123 37203 60129
rect 36044 60120 36050 60123
rect 35820 60064 36308 60092
rect 33778 60024 33784 60036
rect 33244 59996 33784 60024
rect 33778 59984 33784 59996
rect 33836 59984 33842 60036
rect 34514 59984 34520 60036
rect 34572 60024 34578 60036
rect 34882 60024 34888 60036
rect 34572 59996 34888 60024
rect 34572 59984 34578 59996
rect 34882 59984 34888 59996
rect 34940 59984 34946 60036
rect 35342 59984 35348 60036
rect 35400 60024 35406 60036
rect 36173 60027 36231 60033
rect 36173 60024 36185 60027
rect 35400 59996 36185 60024
rect 35400 59984 35406 59996
rect 36173 59993 36185 59996
rect 36219 59993 36231 60027
rect 36173 59987 36231 59993
rect 31662 59916 31668 59968
rect 31720 59956 31726 59968
rect 33689 59959 33747 59965
rect 33689 59956 33701 59959
rect 31720 59928 33701 59956
rect 31720 59916 31726 59928
rect 33689 59925 33701 59928
rect 33735 59925 33747 59959
rect 33689 59919 33747 59925
rect 34977 59959 35035 59965
rect 34977 59925 34989 59959
rect 35023 59956 35035 59959
rect 35802 59956 35808 59968
rect 35023 59928 35808 59956
rect 35023 59925 35035 59928
rect 34977 59919 35035 59925
rect 35802 59916 35808 59928
rect 35860 59916 35866 59968
rect 36280 59956 36308 60064
rect 36740 60024 36768 60123
rect 36924 60092 36952 60123
rect 37274 60092 37280 60104
rect 36924 60064 37280 60092
rect 37274 60052 37280 60064
rect 37332 60052 37338 60104
rect 39298 60024 39304 60036
rect 36740 59996 39304 60024
rect 39298 59984 39304 59996
rect 39356 59984 39362 60036
rect 37182 59956 37188 59968
rect 36280 59928 37188 59956
rect 37182 59916 37188 59928
rect 37240 59916 37246 59968
rect 37277 59959 37335 59965
rect 37277 59925 37289 59959
rect 37323 59956 37335 59959
rect 38654 59956 38660 59968
rect 37323 59928 38660 59956
rect 37323 59925 37335 59928
rect 37277 59919 37335 59925
rect 38654 59916 38660 59928
rect 38712 59916 38718 59968
rect 1104 59866 38824 59888
rect 1104 59814 4246 59866
rect 4298 59814 4310 59866
rect 4362 59814 4374 59866
rect 4426 59814 4438 59866
rect 4490 59814 34966 59866
rect 35018 59814 35030 59866
rect 35082 59814 35094 59866
rect 35146 59814 35158 59866
rect 35210 59814 38824 59866
rect 1104 59792 38824 59814
rect 31726 59724 33272 59752
rect 25682 59576 25688 59628
rect 25740 59616 25746 59628
rect 31726 59616 31754 59724
rect 25740 59588 31754 59616
rect 25740 59576 25746 59588
rect 33134 59576 33140 59628
rect 33192 59576 33198 59628
rect 33244 59616 33272 59724
rect 33594 59712 33600 59764
rect 33652 59752 33658 59764
rect 33870 59752 33876 59764
rect 33652 59724 33876 59752
rect 33652 59712 33658 59724
rect 33870 59712 33876 59724
rect 33928 59712 33934 59764
rect 34609 59755 34667 59761
rect 34609 59721 34621 59755
rect 34655 59752 34667 59755
rect 35986 59752 35992 59764
rect 34655 59724 35992 59752
rect 34655 59721 34667 59724
rect 34609 59715 34667 59721
rect 35986 59712 35992 59724
rect 36044 59712 36050 59764
rect 33318 59644 33324 59696
rect 33376 59684 33382 59696
rect 33376 59656 33824 59684
rect 33376 59644 33382 59656
rect 33244 59588 33364 59616
rect 1394 59548 1400 59560
rect 1355 59520 1400 59548
rect 1394 59508 1400 59520
rect 1452 59508 1458 59560
rect 31754 59508 31760 59560
rect 31812 59548 31818 59560
rect 32953 59551 33011 59557
rect 32953 59548 32965 59551
rect 31812 59520 32965 59548
rect 31812 59508 31818 59520
rect 32953 59517 32965 59520
rect 32999 59517 33011 59551
rect 33152 59548 33180 59576
rect 33336 59557 33364 59588
rect 33796 59557 33824 59656
rect 35618 59644 35624 59696
rect 35676 59684 35682 59696
rect 36541 59687 36599 59693
rect 36541 59684 36553 59687
rect 35676 59656 36553 59684
rect 35676 59644 35682 59656
rect 36541 59653 36553 59656
rect 36587 59653 36599 59687
rect 36541 59647 36599 59653
rect 37645 59687 37703 59693
rect 37645 59653 37657 59687
rect 37691 59684 37703 59687
rect 38378 59684 38384 59696
rect 37691 59656 38384 59684
rect 37691 59653 37703 59656
rect 37645 59647 37703 59653
rect 38378 59644 38384 59656
rect 38436 59644 38442 59696
rect 35802 59576 35808 59628
rect 35860 59616 35866 59628
rect 35860 59588 37228 59616
rect 35860 59576 35866 59588
rect 33229 59551 33287 59557
rect 33229 59548 33241 59551
rect 33152 59520 33241 59548
rect 32953 59511 33011 59517
rect 33229 59517 33241 59520
rect 33275 59517 33287 59551
rect 33229 59511 33287 59517
rect 33321 59551 33379 59557
rect 33321 59517 33333 59551
rect 33367 59517 33379 59551
rect 33321 59511 33379 59517
rect 33597 59551 33655 59557
rect 33597 59517 33609 59551
rect 33643 59517 33655 59551
rect 33597 59511 33655 59517
rect 33781 59551 33839 59557
rect 33781 59517 33793 59551
rect 33827 59517 33839 59551
rect 34790 59548 34796 59560
rect 34751 59520 34796 59548
rect 33781 59511 33839 59517
rect 30742 59440 30748 59492
rect 30800 59480 30806 59492
rect 32493 59483 32551 59489
rect 32493 59480 32505 59483
rect 30800 59452 32505 59480
rect 30800 59440 30806 59452
rect 32493 59449 32505 59452
rect 32539 59449 32551 59483
rect 32493 59443 32551 59449
rect 33244 59412 33272 59511
rect 33612 59480 33640 59511
rect 34790 59508 34796 59520
rect 34848 59508 34854 59560
rect 35989 59551 36047 59557
rect 35989 59517 36001 59551
rect 36035 59548 36047 59551
rect 36078 59548 36084 59560
rect 36035 59520 36084 59548
rect 36035 59517 36047 59520
rect 35989 59511 36047 59517
rect 36078 59508 36084 59520
rect 36136 59508 36142 59560
rect 36409 59551 36467 59557
rect 36409 59517 36421 59551
rect 36455 59548 36467 59551
rect 36722 59548 36728 59560
rect 36455 59520 36728 59548
rect 36455 59517 36467 59520
rect 36409 59511 36467 59517
rect 36722 59508 36728 59520
rect 36780 59508 36786 59560
rect 37093 59551 37151 59557
rect 37093 59517 37105 59551
rect 37139 59517 37151 59551
rect 37200 59548 37228 59588
rect 37466 59551 37524 59557
rect 37466 59548 37478 59551
rect 37200 59520 37478 59548
rect 37093 59511 37151 59517
rect 37466 59517 37478 59520
rect 37512 59517 37524 59551
rect 37466 59511 37524 59517
rect 34146 59480 34152 59492
rect 33612 59452 34152 59480
rect 34146 59440 34152 59452
rect 34204 59440 34210 59492
rect 35434 59440 35440 59492
rect 35492 59480 35498 59492
rect 36173 59483 36231 59489
rect 36173 59480 36185 59483
rect 35492 59452 36185 59480
rect 35492 59440 35498 59452
rect 36173 59449 36185 59452
rect 36219 59449 36231 59483
rect 36173 59443 36231 59449
rect 36265 59483 36323 59489
rect 36265 59449 36277 59483
rect 36311 59480 36323 59483
rect 36906 59480 36912 59492
rect 36311 59452 36912 59480
rect 36311 59449 36323 59452
rect 36265 59443 36323 59449
rect 36906 59440 36912 59452
rect 36964 59440 36970 59492
rect 33594 59412 33600 59424
rect 33244 59384 33600 59412
rect 33594 59372 33600 59384
rect 33652 59372 33658 59424
rect 37108 59412 37136 59511
rect 37182 59440 37188 59492
rect 37240 59480 37246 59492
rect 37277 59483 37335 59489
rect 37277 59480 37289 59483
rect 37240 59452 37289 59480
rect 37240 59440 37246 59452
rect 37277 59449 37289 59452
rect 37323 59449 37335 59483
rect 37277 59443 37335 59449
rect 37366 59440 37372 59492
rect 37424 59480 37430 59492
rect 37424 59452 37469 59480
rect 37424 59440 37430 59452
rect 38838 59412 38844 59424
rect 37108 59384 38844 59412
rect 38838 59372 38844 59384
rect 38896 59372 38902 59424
rect 1104 59322 38824 59344
rect 1104 59270 19606 59322
rect 19658 59270 19670 59322
rect 19722 59270 19734 59322
rect 19786 59270 19798 59322
rect 19850 59270 38824 59322
rect 1104 59248 38824 59270
rect 29638 59168 29644 59220
rect 29696 59208 29702 59220
rect 30098 59208 30104 59220
rect 29696 59180 30104 59208
rect 29696 59168 29702 59180
rect 30098 59168 30104 59180
rect 30156 59168 30162 59220
rect 34146 59208 34152 59220
rect 31680 59180 34152 59208
rect 31680 59149 31708 59180
rect 34146 59168 34152 59180
rect 34204 59168 34210 59220
rect 36722 59208 36728 59220
rect 35912 59180 36728 59208
rect 31665 59143 31723 59149
rect 31665 59109 31677 59143
rect 31711 59109 31723 59143
rect 31665 59103 31723 59109
rect 31757 59143 31815 59149
rect 31757 59109 31769 59143
rect 31803 59140 31815 59143
rect 33134 59140 33140 59152
rect 31803 59112 33140 59140
rect 31803 59109 31815 59112
rect 31757 59103 31815 59109
rect 33134 59100 33140 59112
rect 33192 59100 33198 59152
rect 35912 59149 35940 59180
rect 36722 59168 36728 59180
rect 36780 59168 36786 59220
rect 37182 59208 37188 59220
rect 36924 59180 37188 59208
rect 36924 59149 36952 59180
rect 37182 59168 37188 59180
rect 37240 59168 37246 59220
rect 35897 59143 35955 59149
rect 35897 59109 35909 59143
rect 35943 59109 35955 59143
rect 35897 59103 35955 59109
rect 36909 59143 36967 59149
rect 36909 59109 36921 59143
rect 36955 59109 36967 59143
rect 36909 59103 36967 59109
rect 37001 59143 37059 59149
rect 37001 59109 37013 59143
rect 37047 59140 37059 59143
rect 37366 59140 37372 59152
rect 37047 59112 37372 59140
rect 37047 59109 37059 59112
rect 37001 59103 37059 59109
rect 37366 59100 37372 59112
rect 37424 59100 37430 59152
rect 31389 59075 31447 59081
rect 31389 59072 31401 59075
rect 26206 59044 31401 59072
rect 25590 58964 25596 59016
rect 25648 59004 25654 59016
rect 26206 59004 26234 59044
rect 31389 59041 31401 59044
rect 31435 59041 31447 59075
rect 31389 59035 31447 59041
rect 31478 59032 31484 59084
rect 31536 59072 31542 59084
rect 31938 59081 31944 59084
rect 31895 59075 31944 59081
rect 31536 59044 31581 59072
rect 31536 59032 31542 59044
rect 31895 59041 31907 59075
rect 31941 59041 31944 59075
rect 31895 59035 31944 59041
rect 31938 59032 31944 59035
rect 31996 59032 32002 59084
rect 33505 59075 33563 59081
rect 33505 59041 33517 59075
rect 33551 59041 33563 59075
rect 33505 59035 33563 59041
rect 25648 58976 26234 59004
rect 33520 59004 33548 59035
rect 33594 59032 33600 59084
rect 33652 59072 33658 59084
rect 33873 59075 33931 59081
rect 33652 59044 33697 59072
rect 33652 59032 33658 59044
rect 33873 59041 33885 59075
rect 33919 59041 33931 59075
rect 34146 59072 34152 59084
rect 34107 59044 34152 59072
rect 33873 59035 33931 59041
rect 33778 59004 33784 59016
rect 33520 58976 33784 59004
rect 25648 58964 25654 58976
rect 33778 58964 33784 58976
rect 33836 58964 33842 59016
rect 30098 58896 30104 58948
rect 30156 58936 30162 58948
rect 33888 58936 33916 59035
rect 34146 59032 34152 59044
rect 34204 59032 34210 59084
rect 34330 59072 34336 59084
rect 34291 59044 34336 59072
rect 34330 59032 34336 59044
rect 34388 59032 34394 59084
rect 35434 59032 35440 59084
rect 35492 59072 35498 59084
rect 35621 59075 35679 59081
rect 35621 59072 35633 59075
rect 35492 59044 35633 59072
rect 35492 59032 35498 59044
rect 35621 59041 35633 59044
rect 35667 59041 35679 59075
rect 35621 59035 35679 59041
rect 35805 59075 35863 59081
rect 35805 59041 35817 59075
rect 35851 59041 35863 59075
rect 35986 59072 35992 59084
rect 36044 59081 36050 59084
rect 35952 59044 35992 59072
rect 35805 59035 35863 59041
rect 30156 58908 33916 58936
rect 35820 58936 35848 59035
rect 35986 59032 35992 59044
rect 36044 59035 36052 59081
rect 36725 59075 36783 59081
rect 36725 59041 36737 59075
rect 36771 59072 36783 59075
rect 36814 59072 36820 59084
rect 36771 59044 36820 59072
rect 36771 59041 36783 59044
rect 36725 59035 36783 59041
rect 36044 59032 36050 59035
rect 36814 59032 36820 59044
rect 36872 59032 36878 59084
rect 37145 59075 37203 59081
rect 37145 59041 37157 59075
rect 37191 59072 37203 59075
rect 37274 59072 37280 59084
rect 37191 59044 37280 59072
rect 37191 59041 37203 59044
rect 37145 59035 37203 59041
rect 37274 59032 37280 59044
rect 37332 59032 37338 59084
rect 37918 58936 37924 58948
rect 35820 58908 37924 58936
rect 30156 58896 30162 58908
rect 37918 58896 37924 58908
rect 37976 58896 37982 58948
rect 31018 58828 31024 58880
rect 31076 58868 31082 58880
rect 32033 58871 32091 58877
rect 32033 58868 32045 58871
rect 31076 58840 32045 58868
rect 31076 58828 31082 58840
rect 32033 58837 32045 58840
rect 32079 58837 32091 58871
rect 32033 58831 32091 58837
rect 32398 58828 32404 58880
rect 32456 58868 32462 58880
rect 33137 58871 33195 58877
rect 33137 58868 33149 58871
rect 32456 58840 33149 58868
rect 32456 58828 32462 58840
rect 33137 58837 33149 58840
rect 33183 58837 33195 58871
rect 36170 58868 36176 58880
rect 36131 58840 36176 58868
rect 33137 58831 33195 58837
rect 36170 58828 36176 58840
rect 36228 58828 36234 58880
rect 36722 58828 36728 58880
rect 36780 58868 36786 58880
rect 37277 58871 37335 58877
rect 37277 58868 37289 58871
rect 36780 58840 37289 58868
rect 36780 58828 36786 58840
rect 37277 58837 37289 58840
rect 37323 58837 37335 58871
rect 37277 58831 37335 58837
rect 1104 58778 38824 58800
rect 1104 58726 4246 58778
rect 4298 58726 4310 58778
rect 4362 58726 4374 58778
rect 4426 58726 4438 58778
rect 4490 58726 34966 58778
rect 35018 58726 35030 58778
rect 35082 58726 35094 58778
rect 35146 58726 35158 58778
rect 35210 58726 38824 58778
rect 1104 58704 38824 58726
rect 31202 58624 31208 58676
rect 31260 58664 31266 58676
rect 33778 58664 33784 58676
rect 31260 58636 33784 58664
rect 31260 58624 31266 58636
rect 33778 58624 33784 58636
rect 33836 58624 33842 58676
rect 36446 58664 36452 58676
rect 36407 58636 36452 58664
rect 36446 58624 36452 58636
rect 36504 58624 36510 58676
rect 37274 58664 37280 58676
rect 36556 58636 37280 58664
rect 31386 58556 31392 58608
rect 31444 58596 31450 58608
rect 34054 58596 34060 58608
rect 31444 58568 34060 58596
rect 31444 58556 31450 58568
rect 34054 58556 34060 58568
rect 34112 58556 34118 58608
rect 35805 58599 35863 58605
rect 35805 58565 35817 58599
rect 35851 58596 35863 58599
rect 36556 58596 36584 58636
rect 37274 58624 37280 58636
rect 37332 58624 37338 58676
rect 35851 58568 36584 58596
rect 35851 58565 35863 58568
rect 35805 58559 35863 58565
rect 36722 58556 36728 58608
rect 36780 58556 36786 58608
rect 37645 58599 37703 58605
rect 37645 58565 37657 58599
rect 37691 58596 37703 58599
rect 37826 58596 37832 58608
rect 37691 58568 37832 58596
rect 37691 58565 37703 58568
rect 37645 58559 37703 58565
rect 37826 58556 37832 58568
rect 37884 58556 37890 58608
rect 34146 58528 34152 58540
rect 26206 58500 33272 58528
rect 1394 58460 1400 58472
rect 1355 58432 1400 58460
rect 1394 58420 1400 58432
rect 1452 58420 1458 58472
rect 15654 58420 15660 58472
rect 15712 58460 15718 58472
rect 26206 58460 26234 58500
rect 32858 58460 32864 58472
rect 15712 58432 26234 58460
rect 32819 58432 32864 58460
rect 15712 58420 15718 58432
rect 32858 58420 32864 58432
rect 32916 58420 32922 58472
rect 33134 58460 33140 58472
rect 33095 58432 33140 58460
rect 33134 58420 33140 58432
rect 33192 58420 33198 58472
rect 33244 58469 33272 58500
rect 33520 58500 34152 58528
rect 33520 58469 33548 58500
rect 34146 58488 34152 58500
rect 34204 58488 34210 58540
rect 36740 58528 36768 58556
rect 36280 58500 36768 58528
rect 36280 58472 36308 58500
rect 33229 58463 33287 58469
rect 33229 58429 33241 58463
rect 33275 58429 33287 58463
rect 33229 58423 33287 58429
rect 33505 58463 33563 58469
rect 33505 58429 33517 58463
rect 33551 58429 33563 58463
rect 33505 58423 33563 58429
rect 33781 58463 33839 58469
rect 33781 58429 33793 58463
rect 33827 58460 33839 58463
rect 34790 58460 34796 58472
rect 33827 58432 34796 58460
rect 33827 58429 33839 58432
rect 33781 58423 33839 58429
rect 34790 58420 34796 58432
rect 34848 58420 34854 58472
rect 35802 58420 35808 58472
rect 35860 58460 35866 58472
rect 35989 58463 36047 58469
rect 35989 58460 36001 58463
rect 35860 58432 36001 58460
rect 35860 58420 35866 58432
rect 35989 58429 36001 58432
rect 36035 58429 36047 58463
rect 35989 58423 36047 58429
rect 36262 58420 36268 58472
rect 36320 58420 36326 58472
rect 36633 58463 36691 58469
rect 36633 58429 36645 58463
rect 36679 58460 36691 58463
rect 36722 58460 36728 58472
rect 36679 58432 36728 58460
rect 36679 58429 36691 58432
rect 36633 58423 36691 58429
rect 36722 58420 36728 58432
rect 36780 58420 36786 58472
rect 36998 58420 37004 58472
rect 37056 58460 37062 58472
rect 37093 58463 37151 58469
rect 37093 58460 37105 58463
rect 37056 58432 37105 58460
rect 37056 58420 37062 58432
rect 37093 58429 37105 58432
rect 37139 58429 37151 58463
rect 37093 58423 37151 58429
rect 37182 58420 37188 58472
rect 37240 58460 37246 58472
rect 37466 58463 37524 58469
rect 37466 58460 37478 58463
rect 37240 58432 37478 58460
rect 37240 58420 37246 58432
rect 37466 58429 37478 58432
rect 37512 58429 37524 58463
rect 37466 58423 37524 58429
rect 29730 58352 29736 58404
rect 29788 58392 29794 58404
rect 32401 58395 32459 58401
rect 32401 58392 32413 58395
rect 29788 58364 32413 58392
rect 29788 58352 29794 58364
rect 32401 58361 32413 58364
rect 32447 58361 32459 58395
rect 37274 58392 37280 58404
rect 37235 58364 37280 58392
rect 32401 58355 32459 58361
rect 37274 58352 37280 58364
rect 37332 58352 37338 58404
rect 37366 58352 37372 58404
rect 37424 58392 37430 58404
rect 37424 58364 37469 58392
rect 37424 58352 37430 58364
rect 29914 58284 29920 58336
rect 29972 58324 29978 58336
rect 33594 58324 33600 58336
rect 29972 58296 33600 58324
rect 29972 58284 29978 58296
rect 33594 58284 33600 58296
rect 33652 58284 33658 58336
rect 1104 58234 38824 58256
rect 1104 58182 19606 58234
rect 19658 58182 19670 58234
rect 19722 58182 19734 58234
rect 19786 58182 19798 58234
rect 19850 58182 38824 58234
rect 1104 58160 38824 58182
rect 18782 58080 18788 58132
rect 18840 58120 18846 58132
rect 30098 58120 30104 58132
rect 18840 58092 30104 58120
rect 18840 58080 18846 58092
rect 30098 58080 30104 58092
rect 30156 58080 30162 58132
rect 30190 58080 30196 58132
rect 30248 58120 30254 58132
rect 34054 58120 34060 58132
rect 30248 58092 34060 58120
rect 30248 58080 30254 58092
rect 34054 58080 34060 58092
rect 34112 58080 34118 58132
rect 36541 58123 36599 58129
rect 36541 58089 36553 58123
rect 36587 58120 36599 58123
rect 37182 58120 37188 58132
rect 36587 58092 37188 58120
rect 36587 58089 36599 58092
rect 36541 58083 36599 58089
rect 37182 58080 37188 58092
rect 37240 58080 37246 58132
rect 30282 58012 30288 58064
rect 30340 58052 30346 58064
rect 34330 58052 34336 58064
rect 30340 58024 34336 58052
rect 30340 58012 30346 58024
rect 34330 58012 34336 58024
rect 34388 58012 34394 58064
rect 35986 58012 35992 58064
rect 36044 58052 36050 58064
rect 37274 58052 37280 58064
rect 36044 58024 37280 58052
rect 36044 58012 36050 58024
rect 37274 58012 37280 58024
rect 37332 58012 37338 58064
rect 1394 57984 1400 57996
rect 1355 57956 1400 57984
rect 1394 57944 1400 57956
rect 1452 57944 1458 57996
rect 29638 57944 29644 57996
rect 29696 57984 29702 57996
rect 33318 57984 33324 57996
rect 29696 57956 33324 57984
rect 29696 57944 29702 57956
rect 33318 57944 33324 57956
rect 33376 57944 33382 57996
rect 36725 57987 36783 57993
rect 36725 57953 36737 57987
rect 36771 57984 36783 57987
rect 36814 57984 36820 57996
rect 36771 57956 36820 57984
rect 36771 57953 36783 57956
rect 36725 57947 36783 57953
rect 36814 57944 36820 57956
rect 36872 57944 36878 57996
rect 36906 57944 36912 57996
rect 36964 57984 36970 57996
rect 36964 57956 37136 57984
rect 36964 57944 36970 57956
rect 30466 57876 30472 57928
rect 30524 57916 30530 57928
rect 32030 57916 32036 57928
rect 30524 57888 32036 57916
rect 30524 57876 30530 57888
rect 32030 57876 32036 57888
rect 32088 57876 32094 57928
rect 37108 57848 37136 57956
rect 37182 57944 37188 57996
rect 37240 57984 37246 57996
rect 37369 57987 37427 57993
rect 37369 57984 37381 57987
rect 37240 57956 37381 57984
rect 37240 57944 37246 57956
rect 37369 57953 37381 57956
rect 37415 57953 37427 57987
rect 37369 57947 37427 57953
rect 37185 57851 37243 57857
rect 37185 57848 37197 57851
rect 37108 57820 37197 57848
rect 37185 57817 37197 57820
rect 37231 57817 37243 57851
rect 37185 57811 37243 57817
rect 1104 57690 38824 57712
rect 1104 57638 4246 57690
rect 4298 57638 4310 57690
rect 4362 57638 4374 57690
rect 4426 57638 4438 57690
rect 4490 57638 34966 57690
rect 35018 57638 35030 57690
rect 35082 57638 35094 57690
rect 35146 57638 35158 57690
rect 35210 57638 38824 57690
rect 1104 57616 38824 57638
rect 37274 57576 37280 57588
rect 37235 57548 37280 57576
rect 37274 57536 37280 57548
rect 37332 57536 37338 57588
rect 37458 57372 37464 57384
rect 37419 57344 37464 57372
rect 37458 57332 37464 57344
rect 37516 57332 37522 57384
rect 37918 57372 37924 57384
rect 37879 57344 37924 57372
rect 37918 57332 37924 57344
rect 37976 57332 37982 57384
rect 1104 57146 38824 57168
rect 1104 57094 19606 57146
rect 19658 57094 19670 57146
rect 19722 57094 19734 57146
rect 19786 57094 19798 57146
rect 19850 57094 38824 57146
rect 1104 57072 38824 57094
rect 1394 56896 1400 56908
rect 1355 56868 1400 56896
rect 1394 56856 1400 56868
rect 1452 56856 1458 56908
rect 31938 56652 31944 56704
rect 31996 56692 32002 56704
rect 37642 56692 37648 56704
rect 31996 56664 37648 56692
rect 31996 56652 32002 56664
rect 37642 56652 37648 56664
rect 37700 56652 37706 56704
rect 1104 56602 38824 56624
rect 1104 56550 4246 56602
rect 4298 56550 4310 56602
rect 4362 56550 4374 56602
rect 4426 56550 4438 56602
rect 4490 56550 34966 56602
rect 35018 56550 35030 56602
rect 35082 56550 35094 56602
rect 35146 56550 35158 56602
rect 35210 56550 38824 56602
rect 1104 56528 38824 56550
rect 15746 56488 15752 56500
rect 15707 56460 15752 56488
rect 15746 56448 15752 56460
rect 15804 56448 15810 56500
rect 16669 56491 16727 56497
rect 16669 56457 16681 56491
rect 16715 56488 16727 56491
rect 16850 56488 16856 56500
rect 16715 56460 16856 56488
rect 16715 56457 16727 56460
rect 16669 56451 16727 56457
rect 16850 56448 16856 56460
rect 16908 56448 16914 56500
rect 17589 56491 17647 56497
rect 17589 56457 17601 56491
rect 17635 56488 17647 56491
rect 17770 56488 17776 56500
rect 17635 56460 17776 56488
rect 17635 56457 17647 56460
rect 17589 56451 17647 56457
rect 17770 56448 17776 56460
rect 17828 56448 17834 56500
rect 33686 56352 33692 56364
rect 6886 56324 16528 56352
rect 1394 56284 1400 56296
rect 1355 56256 1400 56284
rect 1394 56244 1400 56256
rect 1452 56244 1458 56296
rect 2958 56176 2964 56228
rect 3016 56216 3022 56228
rect 6886 56216 6914 56324
rect 16500 56293 16528 56324
rect 33429 56324 33692 56352
rect 15381 56287 15439 56293
rect 15381 56253 15393 56287
rect 15427 56253 15439 56287
rect 15381 56247 15439 56253
rect 15565 56287 15623 56293
rect 15565 56253 15577 56287
rect 15611 56284 15623 56287
rect 16301 56287 16359 56293
rect 16301 56284 16313 56287
rect 15611 56256 16313 56284
rect 15611 56253 15623 56256
rect 15565 56247 15623 56253
rect 16301 56253 16313 56256
rect 16347 56253 16359 56287
rect 16301 56247 16359 56253
rect 16485 56287 16543 56293
rect 16485 56253 16497 56287
rect 16531 56253 16543 56287
rect 17310 56284 17316 56296
rect 16485 56247 16543 56253
rect 16960 56256 17316 56284
rect 3016 56188 6914 56216
rect 3016 56176 3022 56188
rect 6454 56108 6460 56160
rect 6512 56148 6518 56160
rect 15396 56148 15424 56247
rect 16316 56216 16344 56247
rect 16758 56216 16764 56228
rect 16316 56188 16764 56216
rect 16758 56176 16764 56188
rect 16816 56216 16822 56228
rect 16960 56216 16988 56256
rect 17310 56244 17316 56256
rect 17368 56244 17374 56296
rect 17405 56287 17463 56293
rect 17405 56253 17417 56287
rect 17451 56253 17463 56287
rect 33042 56284 33048 56296
rect 33003 56256 33048 56284
rect 17405 56247 17463 56253
rect 17420 56216 17448 56247
rect 33042 56244 33048 56256
rect 33100 56244 33106 56296
rect 33193 56287 33251 56293
rect 33193 56253 33205 56287
rect 33239 56284 33251 56287
rect 33429 56284 33457 56324
rect 33686 56312 33692 56324
rect 33744 56312 33750 56364
rect 34238 56312 34244 56364
rect 34296 56312 34302 56364
rect 33239 56256 33457 56284
rect 33551 56287 33609 56293
rect 33239 56253 33251 56256
rect 33193 56247 33251 56253
rect 33551 56253 33563 56287
rect 33597 56284 33609 56287
rect 34256 56284 34284 56312
rect 37458 56284 37464 56296
rect 33597 56256 34284 56284
rect 37419 56256 37464 56284
rect 33597 56253 33609 56256
rect 33551 56247 33609 56253
rect 37458 56244 37464 56256
rect 37516 56244 37522 56296
rect 37918 56284 37924 56296
rect 37879 56256 37924 56284
rect 37918 56244 37924 56256
rect 37976 56244 37982 56296
rect 16816 56188 16988 56216
rect 17052 56188 17448 56216
rect 16816 56176 16822 56188
rect 6512 56120 15424 56148
rect 6512 56108 6518 56120
rect 16850 56108 16856 56160
rect 16908 56148 16914 56160
rect 17052 56157 17080 56188
rect 32490 56176 32496 56228
rect 32548 56216 32554 56228
rect 33321 56219 33379 56225
rect 33321 56216 33333 56219
rect 32548 56188 33333 56216
rect 32548 56176 32554 56188
rect 33321 56185 33333 56188
rect 33367 56185 33379 56219
rect 33321 56179 33379 56185
rect 33413 56219 33471 56225
rect 33413 56185 33425 56219
rect 33459 56216 33471 56219
rect 33870 56216 33876 56228
rect 33459 56188 33876 56216
rect 33459 56185 33471 56188
rect 33413 56179 33471 56185
rect 33870 56176 33876 56188
rect 33928 56176 33934 56228
rect 17037 56151 17095 56157
rect 17037 56148 17049 56151
rect 16908 56120 17049 56148
rect 16908 56108 16914 56120
rect 17037 56117 17049 56120
rect 17083 56117 17095 56151
rect 17037 56111 17095 56117
rect 33689 56151 33747 56157
rect 33689 56117 33701 56151
rect 33735 56148 33747 56151
rect 34146 56148 34152 56160
rect 33735 56120 34152 56148
rect 33735 56117 33747 56120
rect 33689 56111 33747 56117
rect 34146 56108 34152 56120
rect 34204 56108 34210 56160
rect 37277 56151 37335 56157
rect 37277 56117 37289 56151
rect 37323 56148 37335 56151
rect 37550 56148 37556 56160
rect 37323 56120 37556 56148
rect 37323 56117 37335 56120
rect 37277 56111 37335 56117
rect 37550 56108 37556 56120
rect 37608 56108 37614 56160
rect 1104 56058 38824 56080
rect 1104 56006 19606 56058
rect 19658 56006 19670 56058
rect 19722 56006 19734 56058
rect 19786 56006 19798 56058
rect 19850 56006 38824 56058
rect 1104 55984 38824 56006
rect 2406 55904 2412 55956
rect 2464 55944 2470 55956
rect 16850 55944 16856 55956
rect 2464 55916 16856 55944
rect 2464 55904 2470 55916
rect 16850 55904 16856 55916
rect 16908 55904 16914 55956
rect 33502 55944 33508 55956
rect 33429 55916 33508 55944
rect 16022 55836 16028 55888
rect 16080 55876 16086 55888
rect 33042 55876 33048 55888
rect 16080 55848 33048 55876
rect 16080 55836 16086 55848
rect 33042 55836 33048 55848
rect 33100 55836 33106 55888
rect 17678 55768 17684 55820
rect 17736 55808 17742 55820
rect 33429 55817 33457 55916
rect 33502 55904 33508 55916
rect 33560 55904 33566 55956
rect 36446 55904 36452 55956
rect 36504 55944 36510 55956
rect 36998 55944 37004 55956
rect 36504 55916 37004 55944
rect 36504 55904 36510 55916
rect 36998 55904 37004 55916
rect 37056 55904 37062 55956
rect 33597 55879 33655 55885
rect 33597 55845 33609 55879
rect 33643 55876 33655 55879
rect 33870 55876 33876 55888
rect 33643 55848 33876 55876
rect 33643 55845 33655 55848
rect 33597 55839 33655 55845
rect 33870 55836 33876 55848
rect 33928 55836 33934 55888
rect 35250 55836 35256 55888
rect 35308 55876 35314 55888
rect 35802 55876 35808 55888
rect 35308 55848 35808 55876
rect 35308 55836 35314 55848
rect 35802 55836 35808 55848
rect 35860 55836 35866 55888
rect 36078 55836 36084 55888
rect 36136 55876 36142 55888
rect 36814 55876 36820 55888
rect 36136 55848 36820 55876
rect 36136 55836 36142 55848
rect 36814 55836 36820 55848
rect 36872 55836 36878 55888
rect 38470 55876 38476 55888
rect 37016 55848 38476 55876
rect 33229 55811 33287 55817
rect 33229 55808 33241 55811
rect 17736 55780 33241 55808
rect 17736 55768 17742 55780
rect 33229 55777 33241 55780
rect 33275 55777 33287 55811
rect 33229 55771 33287 55777
rect 33377 55811 33457 55817
rect 33377 55777 33389 55811
rect 33423 55780 33457 55811
rect 33505 55811 33563 55817
rect 33423 55777 33435 55780
rect 33377 55771 33435 55777
rect 33505 55777 33517 55811
rect 33551 55777 33563 55811
rect 33505 55771 33563 55777
rect 33735 55811 33793 55817
rect 33735 55777 33747 55811
rect 33781 55808 33793 55811
rect 37016 55808 37044 55848
rect 38470 55836 38476 55848
rect 38528 55836 38534 55888
rect 37182 55808 37188 55820
rect 33781 55780 37044 55808
rect 37143 55780 37188 55808
rect 33781 55777 33793 55780
rect 33735 55771 33793 55777
rect 32490 55700 32496 55752
rect 32548 55740 32554 55752
rect 32858 55740 32864 55752
rect 32548 55712 32864 55740
rect 32548 55700 32554 55712
rect 32858 55700 32864 55712
rect 32916 55740 32922 55752
rect 33520 55740 33548 55771
rect 37182 55768 37188 55780
rect 37240 55768 37246 55820
rect 32916 55712 33548 55740
rect 32916 55700 32922 55712
rect 35250 55700 35256 55752
rect 35308 55740 35314 55752
rect 35710 55740 35716 55752
rect 35308 55712 35716 55740
rect 35308 55700 35314 55712
rect 35710 55700 35716 55712
rect 35768 55700 35774 55752
rect 31938 55632 31944 55684
rect 31996 55672 32002 55684
rect 33873 55675 33931 55681
rect 33873 55672 33885 55675
rect 31996 55644 33885 55672
rect 31996 55632 32002 55644
rect 33873 55641 33885 55644
rect 33919 55641 33931 55675
rect 33873 55635 33931 55641
rect 32490 55564 32496 55616
rect 32548 55604 32554 55616
rect 32674 55604 32680 55616
rect 32548 55576 32680 55604
rect 32548 55564 32554 55576
rect 32674 55564 32680 55576
rect 32732 55564 32738 55616
rect 33134 55564 33140 55616
rect 33192 55604 33198 55616
rect 33594 55604 33600 55616
rect 33192 55576 33600 55604
rect 33192 55564 33198 55576
rect 33594 55564 33600 55576
rect 33652 55564 33658 55616
rect 1104 55514 38824 55536
rect 1104 55462 4246 55514
rect 4298 55462 4310 55514
rect 4362 55462 4374 55514
rect 4426 55462 4438 55514
rect 4490 55462 34966 55514
rect 35018 55462 35030 55514
rect 35082 55462 35094 55514
rect 35146 55462 35158 55514
rect 35210 55462 38824 55514
rect 1104 55440 38824 55462
rect 32858 55264 32864 55276
rect 32324 55236 32864 55264
rect 1394 55196 1400 55208
rect 1355 55168 1400 55196
rect 1394 55156 1400 55168
rect 1452 55156 1458 55208
rect 32214 55205 32220 55208
rect 32033 55199 32091 55205
rect 32033 55196 32045 55199
rect 26206 55168 32045 55196
rect 18506 55088 18512 55140
rect 18564 55128 18570 55140
rect 26206 55128 26234 55168
rect 32033 55165 32045 55168
rect 32079 55165 32091 55199
rect 32033 55159 32091 55165
rect 32181 55199 32220 55205
rect 32181 55165 32193 55199
rect 32181 55159 32220 55165
rect 32214 55156 32220 55159
rect 32272 55156 32278 55208
rect 32324 55205 32352 55236
rect 32858 55224 32864 55236
rect 32916 55224 32922 55276
rect 33502 55224 33508 55276
rect 33560 55264 33566 55276
rect 33870 55264 33876 55276
rect 33560 55236 33876 55264
rect 33560 55224 33566 55236
rect 32582 55205 32588 55208
rect 32309 55199 32367 55205
rect 32309 55165 32321 55199
rect 32355 55165 32367 55199
rect 32309 55159 32367 55165
rect 32539 55199 32588 55205
rect 32539 55165 32551 55199
rect 32585 55165 32588 55199
rect 32539 55159 32588 55165
rect 32582 55156 32588 55159
rect 32640 55156 32646 55208
rect 32674 55156 32680 55208
rect 32732 55196 32738 55208
rect 33410 55205 33416 55208
rect 33229 55199 33287 55205
rect 33229 55196 33241 55199
rect 32732 55168 33241 55196
rect 32732 55156 32738 55168
rect 33229 55165 33241 55168
rect 33275 55165 33287 55199
rect 33229 55159 33287 55165
rect 33377 55199 33416 55205
rect 33377 55165 33389 55199
rect 33377 55159 33416 55165
rect 33410 55156 33416 55159
rect 33468 55156 33474 55208
rect 33612 55205 33640 55236
rect 33870 55224 33876 55236
rect 33928 55224 33934 55276
rect 33597 55199 33655 55205
rect 33597 55165 33609 55199
rect 33643 55165 33655 55199
rect 33597 55159 33655 55165
rect 33735 55199 33793 55205
rect 33735 55165 33747 55199
rect 33781 55196 33793 55199
rect 33962 55196 33968 55208
rect 33781 55168 33968 55196
rect 33781 55165 33793 55168
rect 33735 55159 33793 55165
rect 18564 55100 26234 55128
rect 32401 55131 32459 55137
rect 18564 55088 18570 55100
rect 32401 55097 32413 55131
rect 32447 55128 32459 55131
rect 32447 55100 32812 55128
rect 32447 55097 32459 55100
rect 32401 55091 32459 55097
rect 31754 55020 31760 55072
rect 31812 55060 31818 55072
rect 32677 55063 32735 55069
rect 32677 55060 32689 55063
rect 31812 55032 32689 55060
rect 31812 55020 31818 55032
rect 32677 55029 32689 55032
rect 32723 55029 32735 55063
rect 32784 55060 32812 55100
rect 32858 55088 32864 55140
rect 32916 55128 32922 55140
rect 33505 55131 33563 55137
rect 33505 55128 33517 55131
rect 32916 55100 33517 55128
rect 32916 55088 32922 55100
rect 33505 55097 33517 55100
rect 33551 55097 33563 55131
rect 33505 55091 33563 55097
rect 33612 55060 33640 55159
rect 33962 55156 33968 55168
rect 34020 55156 34026 55208
rect 37458 55196 37464 55208
rect 37419 55168 37464 55196
rect 37458 55156 37464 55168
rect 37516 55156 37522 55208
rect 37918 55196 37924 55208
rect 37879 55168 37924 55196
rect 37918 55156 37924 55168
rect 37976 55156 37982 55208
rect 32784 55032 33640 55060
rect 32677 55023 32735 55029
rect 33686 55020 33692 55072
rect 33744 55060 33750 55072
rect 33873 55063 33931 55069
rect 33873 55060 33885 55063
rect 33744 55032 33885 55060
rect 33744 55020 33750 55032
rect 33873 55029 33885 55032
rect 33919 55029 33931 55063
rect 33873 55023 33931 55029
rect 37277 55063 37335 55069
rect 37277 55029 37289 55063
rect 37323 55060 37335 55063
rect 37366 55060 37372 55072
rect 37323 55032 37372 55060
rect 37323 55029 37335 55032
rect 37277 55023 37335 55029
rect 37366 55020 37372 55032
rect 37424 55020 37430 55072
rect 1104 54970 38824 54992
rect 1104 54918 19606 54970
rect 19658 54918 19670 54970
rect 19722 54918 19734 54970
rect 19786 54918 19798 54970
rect 19850 54918 38824 54970
rect 1104 54896 38824 54918
rect 33870 54816 33876 54868
rect 33928 54856 33934 54868
rect 34238 54856 34244 54868
rect 33928 54828 34244 54856
rect 33928 54816 33934 54828
rect 34238 54816 34244 54828
rect 34296 54816 34302 54868
rect 18690 54748 18696 54800
rect 18748 54788 18754 54800
rect 32674 54788 32680 54800
rect 18748 54760 32680 54788
rect 18748 54748 18754 54760
rect 32674 54748 32680 54760
rect 32732 54748 32738 54800
rect 34422 54788 34428 54800
rect 33336 54760 34428 54788
rect 1394 54720 1400 54732
rect 1355 54692 1400 54720
rect 1394 54680 1400 54692
rect 1452 54680 1458 54732
rect 29638 54680 29644 54732
rect 29696 54720 29702 54732
rect 33336 54729 33364 54760
rect 34422 54748 34428 54760
rect 34480 54748 34486 54800
rect 33137 54723 33195 54729
rect 33137 54720 33149 54723
rect 29696 54692 33149 54720
rect 29696 54680 29702 54692
rect 33137 54689 33149 54692
rect 33183 54689 33195 54723
rect 33137 54683 33195 54689
rect 33285 54723 33364 54729
rect 33285 54689 33297 54723
rect 33331 54692 33364 54723
rect 33413 54723 33471 54729
rect 33331 54689 33343 54692
rect 33285 54683 33343 54689
rect 33413 54689 33425 54723
rect 33459 54689 33471 54723
rect 33413 54683 33471 54689
rect 32858 54612 32864 54664
rect 32916 54652 32922 54664
rect 33428 54652 33456 54683
rect 33502 54680 33508 54732
rect 33560 54720 33566 54732
rect 33643 54723 33701 54729
rect 33560 54692 33605 54720
rect 33560 54680 33566 54692
rect 33643 54689 33655 54723
rect 33689 54720 33701 54723
rect 35526 54720 35532 54732
rect 33689 54692 35532 54720
rect 33689 54689 33701 54692
rect 33643 54683 33701 54689
rect 35526 54680 35532 54692
rect 35584 54680 35590 54732
rect 37182 54720 37188 54732
rect 37143 54692 37188 54720
rect 37182 54680 37188 54692
rect 37240 54680 37246 54732
rect 32916 54624 33456 54652
rect 32916 54612 32922 54624
rect 33410 54476 33416 54528
rect 33468 54516 33474 54528
rect 33781 54519 33839 54525
rect 33781 54516 33793 54519
rect 33468 54488 33793 54516
rect 33468 54476 33474 54488
rect 33781 54485 33793 54488
rect 33827 54485 33839 54519
rect 33781 54479 33839 54485
rect 1104 54426 38824 54448
rect 1104 54374 4246 54426
rect 4298 54374 4310 54426
rect 4362 54374 4374 54426
rect 4426 54374 4438 54426
rect 4490 54374 34966 54426
rect 35018 54374 35030 54426
rect 35082 54374 35094 54426
rect 35146 54374 35158 54426
rect 35210 54374 38824 54426
rect 1104 54352 38824 54374
rect 21542 54312 21548 54324
rect 21503 54284 21548 54312
rect 21542 54272 21548 54284
rect 21600 54272 21606 54324
rect 32122 54312 32128 54324
rect 32083 54284 32128 54312
rect 32122 54272 32128 54284
rect 32180 54272 32186 54324
rect 33226 54312 33232 54324
rect 33187 54284 33232 54312
rect 33226 54272 33232 54284
rect 33284 54272 33290 54324
rect 37553 54315 37611 54321
rect 37553 54281 37565 54315
rect 37599 54312 37611 54315
rect 38930 54312 38936 54324
rect 37599 54284 38936 54312
rect 37599 54281 37611 54284
rect 37553 54275 37611 54281
rect 38930 54272 38936 54284
rect 38988 54272 38994 54324
rect 32030 54204 32036 54256
rect 32088 54244 32094 54256
rect 34241 54247 34299 54253
rect 34241 54244 34253 54247
rect 32088 54216 34253 54244
rect 32088 54204 32094 54216
rect 34241 54213 34253 54216
rect 34287 54213 34299 54247
rect 34241 54207 34299 54213
rect 28166 54068 28172 54120
rect 28224 54108 28230 54120
rect 33137 54111 33195 54117
rect 33137 54108 33149 54111
rect 28224 54080 33149 54108
rect 28224 54068 28230 54080
rect 33137 54077 33149 54080
rect 33183 54077 33195 54111
rect 33137 54071 33195 54077
rect 7374 54000 7380 54052
rect 7432 54040 7438 54052
rect 21453 54043 21511 54049
rect 21453 54040 21465 54043
rect 7432 54012 21465 54040
rect 7432 54000 7438 54012
rect 21453 54009 21465 54012
rect 21499 54009 21511 54043
rect 21453 54003 21511 54009
rect 24394 54000 24400 54052
rect 24452 54040 24458 54052
rect 32033 54043 32091 54049
rect 32033 54040 32045 54043
rect 24452 54012 32045 54040
rect 24452 54000 24458 54012
rect 32033 54009 32045 54012
rect 32079 54009 32091 54043
rect 32033 54003 32091 54009
rect 34057 54043 34115 54049
rect 34057 54009 34069 54043
rect 34103 54009 34115 54043
rect 34057 54003 34115 54009
rect 37277 54043 37335 54049
rect 37277 54009 37289 54043
rect 37323 54040 37335 54043
rect 38194 54040 38200 54052
rect 37323 54012 38200 54040
rect 37323 54009 37335 54012
rect 37277 54003 37335 54009
rect 27706 53932 27712 53984
rect 27764 53972 27770 53984
rect 34072 53972 34100 54003
rect 38194 54000 38200 54012
rect 38252 54000 38258 54052
rect 27764 53944 34100 53972
rect 27764 53932 27770 53944
rect 1104 53882 38824 53904
rect 1104 53830 19606 53882
rect 19658 53830 19670 53882
rect 19722 53830 19734 53882
rect 19786 53830 19798 53882
rect 19850 53830 38824 53882
rect 1104 53808 38824 53830
rect 19334 53768 19340 53780
rect 19295 53740 19340 53768
rect 19334 53728 19340 53740
rect 19392 53728 19398 53780
rect 22922 53768 22928 53780
rect 22883 53740 22928 53768
rect 22922 53728 22928 53740
rect 22980 53728 22986 53780
rect 25038 53768 25044 53780
rect 24999 53740 25044 53768
rect 25038 53728 25044 53740
rect 25096 53728 25102 53780
rect 27982 53768 27988 53780
rect 27943 53740 27988 53768
rect 27982 53728 27988 53740
rect 28040 53728 28046 53780
rect 24949 53703 25007 53709
rect 24949 53700 24961 53703
rect 20732 53672 24961 53700
rect 1394 53632 1400 53644
rect 1355 53604 1400 53632
rect 1394 53592 1400 53604
rect 1452 53592 1458 53644
rect 3510 53592 3516 53644
rect 3568 53632 3574 53644
rect 19061 53635 19119 53641
rect 19061 53632 19073 53635
rect 3568 53604 19073 53632
rect 3568 53592 3574 53604
rect 19061 53601 19073 53604
rect 19107 53601 19119 53635
rect 19061 53595 19119 53601
rect 11238 53524 11244 53576
rect 11296 53564 11302 53576
rect 20732 53564 20760 53672
rect 24949 53669 24961 53672
rect 24995 53669 25007 53703
rect 24949 53663 25007 53669
rect 29365 53703 29423 53709
rect 29365 53669 29377 53703
rect 29411 53700 29423 53703
rect 29454 53700 29460 53712
rect 29411 53672 29460 53700
rect 29411 53669 29423 53672
rect 29365 53663 29423 53669
rect 29454 53660 29460 53672
rect 29512 53660 29518 53712
rect 22833 53635 22891 53641
rect 22833 53601 22845 53635
rect 22879 53601 22891 53635
rect 22833 53595 22891 53601
rect 11296 53536 20760 53564
rect 11296 53524 11302 53536
rect 9674 53456 9680 53508
rect 9732 53496 9738 53508
rect 22848 53496 22876 53595
rect 25038 53592 25044 53644
rect 25096 53632 25102 53644
rect 27893 53635 27951 53641
rect 27893 53632 27905 53635
rect 25096 53604 27905 53632
rect 25096 53592 25102 53604
rect 27893 53601 27905 53604
rect 27939 53601 27951 53635
rect 27893 53595 27951 53601
rect 28997 53635 29055 53641
rect 28997 53601 29009 53635
rect 29043 53601 29055 53635
rect 36722 53632 36728 53644
rect 36683 53604 36728 53632
rect 28997 53595 29055 53601
rect 9732 53468 22876 53496
rect 9732 53456 9738 53468
rect 19426 53388 19432 53440
rect 19484 53428 19490 53440
rect 29012 53428 29040 53595
rect 36722 53592 36728 53604
rect 36780 53592 36786 53644
rect 37182 53632 37188 53644
rect 37143 53604 37188 53632
rect 37182 53592 37188 53604
rect 37240 53592 37246 53644
rect 19484 53400 29040 53428
rect 19484 53388 19490 53400
rect 34238 53388 34244 53440
rect 34296 53428 34302 53440
rect 36541 53431 36599 53437
rect 36541 53428 36553 53431
rect 34296 53400 36553 53428
rect 34296 53388 34302 53400
rect 36541 53397 36553 53400
rect 36587 53397 36599 53431
rect 36541 53391 36599 53397
rect 1104 53338 38824 53360
rect 1104 53286 4246 53338
rect 4298 53286 4310 53338
rect 4362 53286 4374 53338
rect 4426 53286 4438 53338
rect 4490 53286 34966 53338
rect 35018 53286 35030 53338
rect 35082 53286 35094 53338
rect 35146 53286 35158 53338
rect 35210 53286 38824 53338
rect 1104 53264 38824 53286
rect 16482 53184 16488 53236
rect 16540 53224 16546 53236
rect 25038 53224 25044 53236
rect 16540 53196 25044 53224
rect 16540 53184 16546 53196
rect 25038 53184 25044 53196
rect 25096 53184 25102 53236
rect 38654 53116 38660 53168
rect 38712 53156 38718 53168
rect 38930 53156 38936 53168
rect 38712 53128 38936 53156
rect 38712 53116 38718 53128
rect 38930 53116 38936 53128
rect 38988 53116 38994 53168
rect 1394 53020 1400 53032
rect 1355 52992 1400 53020
rect 1394 52980 1400 52992
rect 1452 52980 1458 53032
rect 37274 53020 37280 53032
rect 37235 52992 37280 53020
rect 37274 52980 37280 52992
rect 37332 52980 37338 53032
rect 37918 53020 37924 53032
rect 37879 52992 37924 53020
rect 37918 52980 37924 52992
rect 37976 52980 37982 53032
rect 1104 52794 38824 52816
rect 1104 52742 19606 52794
rect 19658 52742 19670 52794
rect 19722 52742 19734 52794
rect 19786 52742 19798 52794
rect 19850 52742 38824 52794
rect 1104 52720 38824 52742
rect 1394 52544 1400 52556
rect 1355 52516 1400 52544
rect 1394 52504 1400 52516
rect 1452 52504 1458 52556
rect 32674 52368 32680 52420
rect 32732 52408 32738 52420
rect 36262 52408 36268 52420
rect 32732 52380 36268 52408
rect 32732 52368 32738 52380
rect 36262 52368 36268 52380
rect 36320 52368 36326 52420
rect 1104 52250 38824 52272
rect 1104 52198 4246 52250
rect 4298 52198 4310 52250
rect 4362 52198 4374 52250
rect 4426 52198 4438 52250
rect 4490 52198 34966 52250
rect 35018 52198 35030 52250
rect 35082 52198 35094 52250
rect 35146 52198 35158 52250
rect 35210 52198 38824 52250
rect 1104 52176 38824 52198
rect 33689 52071 33747 52077
rect 33689 52037 33701 52071
rect 33735 52068 33747 52071
rect 35526 52068 35532 52080
rect 33735 52040 35532 52068
rect 33735 52037 33747 52040
rect 33689 52031 33747 52037
rect 35526 52028 35532 52040
rect 35584 52028 35590 52080
rect 37550 52000 37556 52012
rect 35452 51972 37556 52000
rect 32950 51892 32956 51944
rect 33008 51932 33014 51944
rect 33045 51935 33103 51941
rect 33045 51932 33057 51935
rect 33008 51904 33057 51932
rect 33008 51892 33014 51904
rect 33045 51901 33057 51904
rect 33091 51901 33103 51935
rect 33045 51895 33103 51901
rect 33138 51935 33196 51941
rect 33138 51901 33150 51935
rect 33184 51901 33196 51935
rect 33138 51895 33196 51901
rect 33551 51935 33609 51941
rect 33551 51901 33563 51935
rect 33597 51932 33609 51935
rect 35452 51932 35480 51972
rect 37550 51960 37556 51972
rect 37608 51960 37614 52012
rect 37458 51932 37464 51944
rect 33597 51904 35480 51932
rect 37419 51904 37464 51932
rect 33597 51901 33609 51904
rect 33551 51895 33609 51901
rect 33152 51864 33180 51895
rect 37458 51892 37464 51904
rect 37516 51892 37522 51944
rect 37918 51932 37924 51944
rect 37879 51904 37924 51932
rect 37918 51892 37924 51904
rect 37976 51892 37982 51944
rect 32876 51836 33180 51864
rect 33321 51867 33379 51873
rect 32876 51808 32904 51836
rect 33321 51833 33333 51867
rect 33367 51833 33379 51867
rect 33321 51827 33379 51833
rect 33413 51867 33471 51873
rect 33413 51833 33425 51867
rect 33459 51864 33471 51867
rect 33459 51836 33640 51864
rect 33459 51833 33471 51836
rect 33413 51827 33471 51833
rect 32858 51796 32864 51808
rect 32819 51768 32864 51796
rect 32858 51756 32864 51768
rect 32916 51756 32922 51808
rect 33336 51796 33364 51827
rect 33612 51808 33640 51836
rect 38746 51824 38752 51876
rect 38804 51864 38810 51876
rect 38804 51836 38884 51864
rect 38804 51824 38810 51836
rect 33502 51796 33508 51808
rect 33336 51768 33508 51796
rect 33502 51756 33508 51768
rect 33560 51756 33566 51808
rect 33594 51756 33600 51808
rect 33652 51756 33658 51808
rect 35434 51756 35440 51808
rect 35492 51796 35498 51808
rect 37277 51799 37335 51805
rect 37277 51796 37289 51799
rect 35492 51768 37289 51796
rect 35492 51756 35498 51768
rect 37277 51765 37289 51768
rect 37323 51765 37335 51799
rect 37277 51759 37335 51765
rect 1104 51706 38824 51728
rect 1104 51654 19606 51706
rect 19658 51654 19670 51706
rect 19722 51654 19734 51706
rect 19786 51654 19798 51706
rect 19850 51654 38824 51706
rect 1104 51632 38824 51654
rect 33594 51552 33600 51604
rect 33652 51592 33658 51604
rect 33652 51564 33732 51592
rect 33652 51552 33658 51564
rect 33704 51533 33732 51564
rect 38746 51552 38752 51604
rect 38804 51592 38810 51604
rect 38856 51592 38884 51836
rect 38804 51564 38884 51592
rect 38804 51552 38810 51564
rect 33689 51527 33747 51533
rect 33689 51493 33701 51527
rect 33735 51493 33747 51527
rect 37366 51524 37372 51536
rect 33689 51487 33747 51493
rect 33842 51496 37372 51524
rect 1394 51456 1400 51468
rect 1355 51428 1400 51456
rect 1394 51416 1400 51428
rect 1452 51416 1458 51468
rect 33226 51416 33232 51468
rect 33284 51456 33290 51468
rect 33321 51459 33379 51465
rect 33321 51456 33333 51459
rect 33284 51428 33333 51456
rect 33284 51416 33290 51428
rect 33321 51425 33333 51428
rect 33367 51425 33379 51459
rect 33321 51419 33379 51425
rect 33414 51459 33472 51465
rect 33414 51425 33426 51459
rect 33460 51425 33472 51459
rect 33414 51419 33472 51425
rect 33429 51388 33457 51419
rect 33502 51416 33508 51468
rect 33560 51456 33566 51468
rect 33842 51465 33870 51496
rect 37366 51484 37372 51496
rect 37424 51484 37430 51536
rect 33597 51459 33655 51465
rect 33597 51456 33609 51459
rect 33560 51428 33609 51456
rect 33560 51416 33566 51428
rect 33597 51425 33609 51428
rect 33643 51425 33655 51459
rect 33597 51419 33655 51425
rect 33827 51459 33885 51465
rect 33827 51425 33839 51459
rect 33873 51425 33885 51459
rect 37182 51456 37188 51468
rect 37143 51428 37188 51456
rect 33827 51419 33885 51425
rect 37182 51416 37188 51428
rect 37240 51416 37246 51468
rect 33152 51360 33457 51388
rect 2314 51212 2320 51264
rect 2372 51252 2378 51264
rect 33152 51261 33180 51360
rect 33137 51255 33195 51261
rect 33137 51252 33149 51255
rect 2372 51224 33149 51252
rect 2372 51212 2378 51224
rect 33137 51221 33149 51224
rect 33183 51221 33195 51255
rect 33137 51215 33195 51221
rect 33965 51255 34023 51261
rect 33965 51221 33977 51255
rect 34011 51252 34023 51255
rect 34606 51252 34612 51264
rect 34011 51224 34612 51252
rect 34011 51221 34023 51224
rect 33965 51215 34023 51221
rect 34606 51212 34612 51224
rect 34664 51212 34670 51264
rect 1104 51162 38824 51184
rect 1104 51110 4246 51162
rect 4298 51110 4310 51162
rect 4362 51110 4374 51162
rect 4426 51110 4438 51162
rect 4490 51110 34966 51162
rect 35018 51110 35030 51162
rect 35082 51110 35094 51162
rect 35146 51110 35158 51162
rect 35210 51110 38824 51162
rect 1104 51088 38824 51110
rect 32582 50940 32588 50992
rect 32640 50980 32646 50992
rect 35618 50980 35624 50992
rect 32640 50952 35624 50980
rect 32640 50940 32646 50952
rect 35618 50940 35624 50952
rect 35676 50940 35682 50992
rect 33686 50872 33692 50924
rect 33744 50912 33750 50924
rect 34054 50912 34060 50924
rect 33744 50884 34060 50912
rect 33744 50872 33750 50884
rect 34054 50872 34060 50884
rect 34112 50872 34118 50924
rect 27522 50804 27528 50856
rect 27580 50844 27586 50856
rect 33321 50847 33379 50853
rect 33321 50844 33333 50847
rect 27580 50816 33333 50844
rect 27580 50804 27586 50816
rect 33321 50813 33333 50816
rect 33367 50813 33379 50847
rect 33321 50807 33379 50813
rect 33414 50847 33472 50853
rect 33414 50813 33426 50847
rect 33460 50813 33472 50847
rect 33414 50807 33472 50813
rect 1854 50776 1860 50788
rect 1815 50748 1860 50776
rect 1854 50736 1860 50748
rect 1912 50736 1918 50788
rect 33429 50776 33457 50807
rect 33502 50804 33508 50856
rect 33560 50853 33566 50856
rect 33560 50847 33609 50853
rect 33560 50813 33563 50847
rect 33597 50813 33609 50847
rect 33560 50807 33609 50813
rect 33805 50847 33863 50853
rect 33805 50813 33817 50847
rect 33851 50844 33863 50847
rect 34238 50844 34244 50856
rect 33851 50816 34244 50844
rect 33851 50813 33863 50816
rect 33805 50807 33863 50813
rect 33560 50804 33566 50807
rect 34238 50804 34244 50816
rect 34296 50804 34302 50856
rect 37458 50844 37464 50856
rect 37419 50816 37464 50844
rect 37458 50804 37464 50816
rect 37516 50804 37522 50856
rect 37918 50844 37924 50856
rect 37879 50816 37924 50844
rect 37918 50804 37924 50816
rect 37976 50804 37982 50856
rect 33336 50748 33457 50776
rect 33697 50779 33755 50785
rect 33336 50720 33364 50748
rect 33697 50745 33709 50779
rect 33743 50745 33755 50779
rect 33697 50739 33755 50745
rect 1949 50711 2007 50717
rect 1949 50677 1961 50711
rect 1995 50708 2007 50711
rect 32858 50708 32864 50720
rect 1995 50680 32864 50708
rect 1995 50677 2007 50680
rect 1949 50671 2007 50677
rect 32858 50668 32864 50680
rect 32916 50668 32922 50720
rect 33229 50711 33287 50717
rect 33229 50677 33241 50711
rect 33275 50708 33287 50711
rect 33318 50708 33324 50720
rect 33275 50680 33324 50708
rect 33275 50677 33287 50680
rect 33229 50671 33287 50677
rect 33318 50668 33324 50680
rect 33376 50668 33382 50720
rect 33594 50668 33600 50720
rect 33652 50708 33658 50720
rect 33704 50708 33732 50739
rect 33652 50680 33732 50708
rect 33965 50711 34023 50717
rect 33652 50668 33658 50680
rect 33965 50677 33977 50711
rect 34011 50708 34023 50711
rect 35802 50708 35808 50720
rect 34011 50680 35808 50708
rect 34011 50677 34023 50680
rect 33965 50671 34023 50677
rect 35802 50668 35808 50680
rect 35860 50668 35866 50720
rect 37277 50711 37335 50717
rect 37277 50677 37289 50711
rect 37323 50708 37335 50711
rect 37550 50708 37556 50720
rect 37323 50680 37556 50708
rect 37323 50677 37335 50680
rect 37277 50671 37335 50677
rect 37550 50668 37556 50680
rect 37608 50668 37614 50720
rect 1104 50618 38824 50640
rect 1104 50566 19606 50618
rect 19658 50566 19670 50618
rect 19722 50566 19734 50618
rect 19786 50566 19798 50618
rect 19850 50566 38824 50618
rect 1104 50544 38824 50566
rect 33686 50464 33692 50516
rect 33744 50464 33750 50516
rect 33597 50439 33655 50445
rect 33597 50405 33609 50439
rect 33643 50436 33655 50439
rect 33704 50436 33732 50464
rect 35434 50436 35440 50448
rect 33643 50408 33732 50436
rect 33842 50408 35440 50436
rect 33643 50405 33655 50408
rect 33597 50399 33655 50405
rect 3602 50328 3608 50380
rect 3660 50368 3666 50380
rect 28902 50368 28908 50380
rect 3660 50340 28908 50368
rect 3660 50328 3666 50340
rect 28902 50328 28908 50340
rect 28960 50328 28966 50380
rect 33134 50328 33140 50380
rect 33192 50368 33198 50380
rect 33842 50377 33870 50408
rect 35434 50396 35440 50408
rect 35492 50396 35498 50448
rect 33321 50371 33379 50377
rect 33321 50368 33333 50371
rect 33192 50340 33333 50368
rect 33192 50328 33198 50340
rect 33321 50337 33333 50340
rect 33367 50337 33379 50371
rect 33321 50331 33379 50337
rect 33414 50371 33472 50377
rect 33414 50337 33426 50371
rect 33460 50337 33472 50371
rect 33414 50331 33472 50337
rect 33702 50371 33760 50377
rect 33702 50337 33714 50371
rect 33748 50368 33760 50371
rect 33827 50371 33885 50377
rect 33748 50337 33778 50368
rect 33702 50331 33778 50337
rect 33827 50337 33839 50371
rect 33873 50337 33885 50371
rect 33827 50331 33885 50337
rect 24854 50260 24860 50312
rect 24912 50300 24918 50312
rect 33429 50300 33457 50331
rect 24912 50272 33457 50300
rect 24912 50260 24918 50272
rect 28721 50235 28779 50241
rect 28721 50201 28733 50235
rect 28767 50232 28779 50235
rect 28902 50232 28908 50244
rect 28767 50204 28908 50232
rect 28767 50201 28779 50204
rect 28721 50195 28779 50201
rect 28902 50192 28908 50204
rect 28960 50192 28966 50244
rect 29089 50235 29147 50241
rect 29089 50201 29101 50235
rect 29135 50232 29147 50235
rect 32122 50232 32128 50244
rect 29135 50204 32128 50232
rect 29135 50201 29147 50204
rect 29089 50195 29147 50201
rect 32122 50192 32128 50204
rect 32180 50232 32186 50244
rect 33594 50232 33600 50244
rect 32180 50204 33600 50232
rect 32180 50192 32186 50204
rect 33594 50192 33600 50204
rect 33652 50232 33658 50244
rect 33750 50232 33778 50331
rect 34514 50328 34520 50380
rect 34572 50368 34578 50380
rect 34609 50371 34667 50377
rect 34609 50368 34621 50371
rect 34572 50340 34621 50368
rect 34572 50328 34578 50340
rect 34609 50337 34621 50340
rect 34655 50337 34667 50371
rect 34609 50331 34667 50337
rect 34793 50235 34851 50241
rect 34793 50232 34805 50235
rect 33652 50204 33778 50232
rect 33888 50204 34805 50232
rect 33652 50192 33658 50204
rect 33502 50124 33508 50176
rect 33560 50164 33566 50176
rect 33686 50164 33692 50176
rect 33560 50136 33692 50164
rect 33560 50124 33566 50136
rect 33686 50124 33692 50136
rect 33744 50164 33750 50176
rect 33888 50164 33916 50204
rect 34793 50201 34805 50204
rect 34839 50201 34851 50235
rect 34793 50195 34851 50201
rect 33744 50136 33916 50164
rect 33965 50167 34023 50173
rect 33744 50124 33750 50136
rect 33965 50133 33977 50167
rect 34011 50164 34023 50167
rect 35618 50164 35624 50176
rect 34011 50136 35624 50164
rect 34011 50133 34023 50136
rect 33965 50127 34023 50133
rect 35618 50124 35624 50136
rect 35676 50124 35682 50176
rect 1104 50074 38824 50096
rect 1104 50022 4246 50074
rect 4298 50022 4310 50074
rect 4362 50022 4374 50074
rect 4426 50022 4438 50074
rect 4490 50022 34966 50074
rect 35018 50022 35030 50074
rect 35082 50022 35094 50074
rect 35146 50022 35158 50074
rect 35210 50022 38824 50074
rect 1104 50000 38824 50022
rect 2041 49895 2099 49901
rect 2041 49861 2053 49895
rect 2087 49892 2099 49895
rect 2314 49892 2320 49904
rect 2087 49864 2320 49892
rect 2087 49861 2099 49864
rect 2041 49855 2099 49861
rect 2314 49852 2320 49864
rect 2372 49852 2378 49904
rect 33502 49892 33508 49904
rect 32048 49864 33508 49892
rect 1854 49756 1860 49768
rect 1815 49728 1860 49756
rect 1854 49716 1860 49728
rect 1912 49716 1918 49768
rect 32048 49765 32076 49864
rect 33502 49852 33508 49864
rect 33560 49852 33566 49904
rect 32122 49784 32128 49836
rect 32180 49824 32186 49836
rect 32180 49796 32444 49824
rect 32180 49784 32186 49796
rect 32033 49759 32091 49765
rect 32033 49725 32045 49759
rect 32079 49725 32091 49759
rect 32214 49756 32220 49768
rect 32175 49728 32220 49756
rect 32033 49719 32091 49725
rect 32214 49716 32220 49728
rect 32272 49716 32278 49768
rect 32416 49765 32444 49796
rect 32401 49759 32459 49765
rect 32401 49725 32413 49759
rect 32447 49725 32459 49759
rect 32401 49719 32459 49725
rect 32677 49759 32735 49765
rect 32677 49725 32689 49759
rect 32723 49756 32735 49759
rect 32766 49756 32772 49768
rect 32723 49728 32772 49756
rect 32723 49725 32735 49728
rect 32677 49719 32735 49725
rect 32766 49716 32772 49728
rect 32824 49716 32830 49768
rect 34514 49716 34520 49768
rect 34572 49756 34578 49768
rect 34790 49756 34796 49768
rect 34572 49728 34796 49756
rect 34572 49716 34578 49728
rect 34790 49716 34796 49728
rect 34848 49716 34854 49768
rect 37918 49756 37924 49768
rect 37879 49728 37924 49756
rect 37918 49716 37924 49728
rect 37976 49716 37982 49768
rect 32030 49620 32036 49632
rect 31991 49592 32036 49620
rect 32030 49580 32036 49592
rect 32088 49580 32094 49632
rect 1104 49530 38824 49552
rect 1104 49478 19606 49530
rect 19658 49478 19670 49530
rect 19722 49478 19734 49530
rect 19786 49478 19798 49530
rect 19850 49478 38824 49530
rect 1104 49456 38824 49478
rect 1854 49280 1860 49292
rect 1815 49252 1860 49280
rect 1854 49240 1860 49252
rect 1912 49240 1918 49292
rect 37366 49280 37372 49292
rect 37327 49252 37372 49280
rect 37366 49240 37372 49252
rect 37424 49240 37430 49292
rect 2314 49172 2320 49224
rect 2372 49212 2378 49224
rect 24854 49212 24860 49224
rect 2372 49184 24860 49212
rect 2372 49172 2378 49184
rect 24854 49172 24860 49184
rect 24912 49172 24918 49224
rect 1949 49079 2007 49085
rect 1949 49045 1961 49079
rect 1995 49076 2007 49079
rect 33318 49076 33324 49088
rect 1995 49048 33324 49076
rect 1995 49045 2007 49048
rect 1949 49039 2007 49045
rect 33318 49036 33324 49048
rect 33376 49036 33382 49088
rect 34514 49036 34520 49088
rect 34572 49076 34578 49088
rect 37185 49079 37243 49085
rect 37185 49076 37197 49079
rect 34572 49048 37197 49076
rect 34572 49036 34578 49048
rect 37185 49045 37197 49048
rect 37231 49045 37243 49079
rect 37185 49039 37243 49045
rect 1104 48986 38824 49008
rect 1104 48934 4246 48986
rect 4298 48934 4310 48986
rect 4362 48934 4374 48986
rect 4426 48934 4438 48986
rect 4490 48934 34966 48986
rect 35018 48934 35030 48986
rect 35082 48934 35094 48986
rect 35146 48934 35158 48986
rect 35210 48934 38824 48986
rect 1104 48912 38824 48934
rect 29546 48804 29552 48816
rect 28092 48776 29552 48804
rect 16669 48671 16727 48677
rect 16669 48637 16681 48671
rect 16715 48668 16727 48671
rect 16758 48668 16764 48680
rect 16715 48640 16764 48668
rect 16715 48637 16727 48640
rect 16669 48631 16727 48637
rect 16758 48628 16764 48640
rect 16816 48628 16822 48680
rect 27614 48668 27620 48680
rect 27575 48640 27620 48668
rect 27614 48628 27620 48640
rect 27672 48628 27678 48680
rect 28092 48677 28120 48776
rect 29546 48764 29552 48776
rect 29604 48764 29610 48816
rect 32030 48736 32036 48748
rect 28368 48708 32036 48736
rect 28368 48677 28396 48708
rect 32030 48696 32036 48708
rect 32088 48696 32094 48748
rect 28077 48671 28135 48677
rect 28077 48637 28089 48671
rect 28123 48637 28135 48671
rect 28077 48631 28135 48637
rect 28353 48671 28411 48677
rect 28353 48637 28365 48671
rect 28399 48637 28411 48671
rect 28534 48668 28540 48680
rect 28495 48640 28540 48668
rect 28353 48631 28411 48637
rect 28534 48628 28540 48640
rect 28592 48628 28598 48680
rect 37274 48668 37280 48680
rect 37235 48640 37280 48668
rect 37274 48628 37280 48640
rect 37332 48628 37338 48680
rect 37918 48668 37924 48680
rect 37879 48640 37924 48668
rect 37918 48628 37924 48640
rect 37976 48628 37982 48680
rect 6638 48560 6644 48612
rect 6696 48600 6702 48612
rect 28813 48603 28871 48609
rect 28813 48600 28825 48603
rect 6696 48572 28825 48600
rect 6696 48560 6702 48572
rect 28813 48569 28825 48572
rect 28859 48569 28871 48603
rect 28813 48563 28871 48569
rect 16850 48532 16856 48544
rect 16811 48504 16856 48532
rect 16850 48492 16856 48504
rect 16908 48492 16914 48544
rect 1104 48442 38824 48464
rect 1104 48390 19606 48442
rect 19658 48390 19670 48442
rect 19722 48390 19734 48442
rect 19786 48390 19798 48442
rect 19850 48390 38824 48442
rect 1104 48368 38824 48390
rect 2041 48263 2099 48269
rect 2041 48229 2053 48263
rect 2087 48260 2099 48263
rect 2314 48260 2320 48272
rect 2087 48232 2320 48260
rect 2087 48229 2099 48232
rect 2041 48223 2099 48229
rect 2314 48220 2320 48232
rect 2372 48220 2378 48272
rect 1854 48192 1860 48204
rect 1815 48164 1860 48192
rect 1854 48152 1860 48164
rect 1912 48152 1918 48204
rect 37366 48192 37372 48204
rect 37327 48164 37372 48192
rect 37366 48152 37372 48164
rect 37424 48152 37430 48204
rect 34606 48084 34612 48136
rect 34664 48124 34670 48136
rect 35434 48124 35440 48136
rect 34664 48096 35440 48124
rect 34664 48084 34670 48096
rect 35434 48084 35440 48096
rect 35492 48084 35498 48136
rect 34606 47948 34612 48000
rect 34664 47988 34670 48000
rect 37185 47991 37243 47997
rect 37185 47988 37197 47991
rect 34664 47960 37197 47988
rect 34664 47948 34670 47960
rect 37185 47957 37197 47960
rect 37231 47957 37243 47991
rect 37185 47951 37243 47957
rect 1104 47898 38824 47920
rect 1104 47846 4246 47898
rect 4298 47846 4310 47898
rect 4362 47846 4374 47898
rect 4426 47846 4438 47898
rect 4490 47846 34966 47898
rect 35018 47846 35030 47898
rect 35082 47846 35094 47898
rect 35146 47846 35158 47898
rect 35210 47846 38824 47898
rect 1104 47824 38824 47846
rect 16758 47580 16764 47592
rect 16719 47552 16764 47580
rect 16758 47540 16764 47552
rect 16816 47540 16822 47592
rect 37274 47580 37280 47592
rect 37235 47552 37280 47580
rect 37274 47540 37280 47552
rect 37332 47540 37338 47592
rect 37918 47580 37924 47592
rect 37879 47552 37924 47580
rect 37918 47540 37924 47552
rect 37976 47540 37982 47592
rect 1854 47512 1860 47524
rect 1815 47484 1860 47512
rect 1854 47472 1860 47484
rect 1912 47472 1918 47524
rect 1946 47444 1952 47456
rect 1907 47416 1952 47444
rect 1946 47404 1952 47416
rect 2004 47404 2010 47456
rect 16945 47447 17003 47453
rect 16945 47413 16957 47447
rect 16991 47444 17003 47447
rect 17310 47444 17316 47456
rect 16991 47416 17316 47444
rect 16991 47413 17003 47416
rect 16945 47407 17003 47413
rect 17310 47404 17316 47416
rect 17368 47404 17374 47456
rect 1104 47354 38824 47376
rect 1104 47302 19606 47354
rect 19658 47302 19670 47354
rect 19722 47302 19734 47354
rect 19786 47302 19798 47354
rect 19850 47302 38824 47354
rect 1104 47280 38824 47302
rect 1946 47200 1952 47252
rect 2004 47240 2010 47252
rect 2004 47212 34100 47240
rect 2004 47200 2010 47212
rect 33962 47104 33968 47116
rect 33923 47076 33968 47104
rect 33962 47064 33968 47076
rect 34020 47064 34026 47116
rect 34072 47113 34100 47212
rect 34058 47107 34116 47113
rect 34058 47073 34070 47107
rect 34104 47073 34116 47107
rect 34238 47104 34244 47116
rect 34199 47076 34244 47104
rect 34058 47067 34116 47073
rect 34238 47064 34244 47076
rect 34296 47064 34302 47116
rect 34333 47107 34391 47113
rect 34333 47073 34345 47107
rect 34379 47073 34391 47107
rect 34333 47067 34391 47073
rect 34471 47107 34529 47113
rect 34471 47073 34483 47107
rect 34517 47104 34529 47107
rect 37550 47104 37556 47116
rect 34517 47076 37556 47104
rect 34517 47073 34529 47076
rect 34471 47067 34529 47073
rect 34348 47036 34376 47067
rect 37550 47064 37556 47076
rect 37608 47064 37614 47116
rect 34348 47008 34468 47036
rect 34440 46980 34468 47008
rect 34422 46928 34428 46980
rect 34480 46928 34486 46980
rect 34609 46971 34667 46977
rect 34609 46937 34621 46971
rect 34655 46968 34667 46971
rect 36078 46968 36084 46980
rect 34655 46940 36084 46968
rect 34655 46937 34667 46940
rect 34609 46931 34667 46937
rect 36078 46928 36084 46940
rect 36136 46928 36142 46980
rect 1104 46810 38824 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 34966 46810
rect 35018 46758 35030 46810
rect 35082 46758 35094 46810
rect 35146 46758 35158 46810
rect 35210 46758 38824 46810
rect 1104 46736 38824 46758
rect 34609 46631 34667 46637
rect 34609 46597 34621 46631
rect 34655 46628 34667 46631
rect 35342 46628 35348 46640
rect 34655 46600 35348 46628
rect 34655 46597 34667 46600
rect 34609 46591 34667 46597
rect 35342 46588 35348 46600
rect 35400 46588 35406 46640
rect 1854 46492 1860 46504
rect 1815 46464 1860 46492
rect 1854 46452 1860 46464
rect 1912 46452 1918 46504
rect 33778 46452 33784 46504
rect 33836 46492 33842 46504
rect 34514 46501 34520 46504
rect 33965 46495 34023 46501
rect 33965 46492 33977 46495
rect 33836 46464 33977 46492
rect 33836 46452 33842 46464
rect 33965 46461 33977 46464
rect 34011 46461 34023 46495
rect 33965 46455 34023 46461
rect 34058 46495 34116 46501
rect 34058 46461 34070 46495
rect 34104 46461 34116 46495
rect 34058 46455 34116 46461
rect 34471 46495 34520 46501
rect 34471 46461 34483 46495
rect 34517 46461 34520 46495
rect 34471 46455 34520 46461
rect 1949 46359 2007 46365
rect 1949 46325 1961 46359
rect 1995 46356 2007 46359
rect 34072 46356 34100 46455
rect 34514 46452 34520 46455
rect 34572 46452 34578 46504
rect 34790 46492 34796 46504
rect 34716 46464 34796 46492
rect 34238 46424 34244 46436
rect 34199 46396 34244 46424
rect 34238 46384 34244 46396
rect 34296 46384 34302 46436
rect 34333 46427 34391 46433
rect 34333 46393 34345 46427
rect 34379 46424 34391 46427
rect 34379 46396 34468 46424
rect 34379 46393 34391 46396
rect 34333 46387 34391 46393
rect 34440 46368 34468 46396
rect 1995 46328 34100 46356
rect 1995 46325 2007 46328
rect 1949 46319 2007 46325
rect 34422 46316 34428 46368
rect 34480 46316 34486 46368
rect 34514 46316 34520 46368
rect 34572 46356 34578 46368
rect 34716 46356 34744 46464
rect 34790 46452 34796 46464
rect 34848 46452 34854 46504
rect 37458 46492 37464 46504
rect 37419 46464 37464 46492
rect 37458 46452 37464 46464
rect 37516 46452 37522 46504
rect 37918 46492 37924 46504
rect 37879 46464 37924 46492
rect 37918 46452 37924 46464
rect 37976 46452 37982 46504
rect 34572 46328 34744 46356
rect 34572 46316 34578 46328
rect 34790 46316 34796 46368
rect 34848 46356 34854 46368
rect 37277 46359 37335 46365
rect 37277 46356 37289 46359
rect 34848 46328 37289 46356
rect 34848 46316 34854 46328
rect 37277 46325 37289 46328
rect 37323 46325 37335 46359
rect 37277 46319 37335 46325
rect 1104 46266 38824 46288
rect 1104 46214 19606 46266
rect 19658 46214 19670 46266
rect 19722 46214 19734 46266
rect 19786 46214 19798 46266
rect 19850 46214 38824 46266
rect 1104 46192 38824 46214
rect 34330 46152 34336 46164
rect 33980 46124 34336 46152
rect 1854 46016 1860 46028
rect 1815 45988 1860 46016
rect 1854 45976 1860 45988
rect 1912 45976 1918 46028
rect 33980 46025 34008 46124
rect 34330 46112 34336 46124
rect 34388 46112 34394 46164
rect 33965 46019 34023 46025
rect 33965 45985 33977 46019
rect 34011 45985 34023 46019
rect 33965 45979 34023 45985
rect 34058 46019 34116 46025
rect 34058 45985 34070 46019
rect 34104 45985 34116 46019
rect 34238 46016 34244 46028
rect 34199 45988 34244 46016
rect 34058 45979 34116 45985
rect 34072 45948 34100 45979
rect 34238 45976 34244 45988
rect 34296 45976 34302 46028
rect 34330 45976 34336 46028
rect 34388 46016 34394 46028
rect 34471 46019 34529 46025
rect 34388 45988 34433 46016
rect 34388 45976 34394 45988
rect 34471 45985 34483 46019
rect 34517 46016 34529 46019
rect 34606 46016 34612 46028
rect 34517 45988 34612 46016
rect 34517 45985 34529 45988
rect 34471 45979 34529 45985
rect 34606 45976 34612 45988
rect 34664 45976 34670 46028
rect 37182 46016 37188 46028
rect 37143 45988 37188 46016
rect 37182 45976 37188 45988
rect 37240 45976 37246 46028
rect 26206 45920 34100 45948
rect 1949 45815 2007 45821
rect 1949 45781 1961 45815
rect 1995 45812 2007 45815
rect 26206 45812 26234 45920
rect 30282 45840 30288 45892
rect 30340 45880 30346 45892
rect 34609 45883 34667 45889
rect 34609 45880 34621 45883
rect 30340 45852 34621 45880
rect 30340 45840 30346 45852
rect 34609 45849 34621 45852
rect 34655 45849 34667 45883
rect 34609 45843 34667 45849
rect 1995 45784 26234 45812
rect 1995 45781 2007 45784
rect 1949 45775 2007 45781
rect 1104 45722 38824 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 34966 45722
rect 35018 45670 35030 45722
rect 35082 45670 35094 45722
rect 35146 45670 35158 45722
rect 35210 45670 38824 45722
rect 1104 45648 38824 45670
rect 34609 45543 34667 45549
rect 34609 45509 34621 45543
rect 34655 45540 34667 45543
rect 36446 45540 36452 45552
rect 34655 45512 36452 45540
rect 34655 45509 34667 45512
rect 34609 45503 34667 45509
rect 36446 45500 36452 45512
rect 36504 45500 36510 45552
rect 35710 45472 35716 45484
rect 33980 45444 35716 45472
rect 33980 45413 34008 45444
rect 35710 45432 35716 45444
rect 35768 45432 35774 45484
rect 33965 45407 34023 45413
rect 33965 45373 33977 45407
rect 34011 45373 34023 45407
rect 33965 45367 34023 45373
rect 34054 45364 34060 45416
rect 34112 45404 34118 45416
rect 34471 45407 34529 45413
rect 34112 45376 34157 45404
rect 34112 45364 34118 45376
rect 34471 45373 34483 45407
rect 34517 45404 34529 45407
rect 34790 45404 34796 45416
rect 34517 45376 34796 45404
rect 34517 45373 34529 45376
rect 34471 45367 34529 45373
rect 34790 45364 34796 45376
rect 34848 45364 34854 45416
rect 37458 45404 37464 45416
rect 37419 45376 37464 45404
rect 37458 45364 37464 45376
rect 37516 45364 37522 45416
rect 37918 45404 37924 45416
rect 37879 45376 37924 45404
rect 37918 45364 37924 45376
rect 37976 45364 37982 45416
rect 34238 45336 34244 45348
rect 34199 45308 34244 45336
rect 34238 45296 34244 45308
rect 34296 45296 34302 45348
rect 34330 45296 34336 45348
rect 34388 45336 34394 45348
rect 34388 45308 34433 45336
rect 34388 45296 34394 45308
rect 34606 45296 34612 45348
rect 34664 45336 34670 45348
rect 35526 45336 35532 45348
rect 34664 45308 35532 45336
rect 34664 45296 34670 45308
rect 35526 45296 35532 45308
rect 35584 45296 35590 45348
rect 35710 45296 35716 45348
rect 35768 45336 35774 45348
rect 35894 45336 35900 45348
rect 35768 45308 35900 45336
rect 35768 45296 35774 45308
rect 35894 45296 35900 45308
rect 35952 45296 35958 45348
rect 34790 45228 34796 45280
rect 34848 45268 34854 45280
rect 37277 45271 37335 45277
rect 37277 45268 37289 45271
rect 34848 45240 37289 45268
rect 34848 45228 34854 45240
rect 37277 45237 37289 45240
rect 37323 45237 37335 45271
rect 37277 45231 37335 45237
rect 1104 45178 38824 45200
rect 1104 45126 19606 45178
rect 19658 45126 19670 45178
rect 19722 45126 19734 45178
rect 19786 45126 19798 45178
rect 19850 45126 38824 45178
rect 1104 45104 38824 45126
rect 33778 45024 33784 45076
rect 33836 45064 33842 45076
rect 39390 45064 39396 45076
rect 33836 45036 39396 45064
rect 33836 45024 33842 45036
rect 39390 45024 39396 45036
rect 39448 45024 39454 45076
rect 1854 44996 1860 45008
rect 1815 44968 1860 44996
rect 1854 44956 1860 44968
rect 1912 44956 1918 45008
rect 1949 44727 2007 44733
rect 1949 44693 1961 44727
rect 1995 44724 2007 44727
rect 34054 44724 34060 44736
rect 1995 44696 34060 44724
rect 1995 44693 2007 44696
rect 1949 44687 2007 44693
rect 34054 44684 34060 44696
rect 34112 44684 34118 44736
rect 1104 44634 38824 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 34966 44634
rect 35018 44582 35030 44634
rect 35082 44582 35094 44634
rect 35146 44582 35158 44634
rect 35210 44582 38824 44634
rect 1104 44560 38824 44582
rect 33410 44412 33416 44464
rect 33468 44452 33474 44464
rect 34054 44452 34060 44464
rect 33468 44424 34060 44452
rect 33468 44412 33474 44424
rect 34054 44412 34060 44424
rect 34112 44452 34118 44464
rect 34330 44452 34336 44464
rect 34112 44424 34336 44452
rect 34112 44412 34118 44424
rect 34330 44412 34336 44424
rect 34388 44412 34394 44464
rect 33686 44344 33692 44396
rect 33744 44384 33750 44396
rect 34238 44384 34244 44396
rect 33744 44356 34244 44384
rect 33744 44344 33750 44356
rect 33870 44316 33876 44328
rect 33831 44288 33876 44316
rect 33870 44276 33876 44288
rect 33928 44276 33934 44328
rect 34164 44325 34192 44356
rect 34238 44344 34244 44356
rect 34296 44344 34302 44396
rect 33966 44319 34024 44325
rect 33966 44285 33978 44319
rect 34012 44285 34024 44319
rect 33966 44279 34024 44285
rect 34149 44319 34207 44325
rect 34149 44285 34161 44319
rect 34195 44285 34207 44319
rect 34149 44279 34207 44285
rect 34379 44319 34437 44325
rect 34379 44285 34391 44319
rect 34425 44316 34437 44319
rect 34790 44316 34796 44328
rect 34425 44288 34796 44316
rect 34425 44285 34437 44288
rect 34379 44279 34437 44285
rect 1854 44248 1860 44260
rect 1815 44220 1860 44248
rect 1854 44208 1860 44220
rect 1912 44208 1918 44260
rect 1949 44183 2007 44189
rect 1949 44149 1961 44183
rect 1995 44180 2007 44183
rect 33980 44180 34008 44279
rect 34790 44276 34796 44288
rect 34848 44276 34854 44328
rect 37182 44276 37188 44328
rect 37240 44316 37246 44328
rect 37461 44319 37519 44325
rect 37461 44316 37473 44319
rect 37240 44288 37473 44316
rect 37240 44276 37246 44288
rect 37461 44285 37473 44288
rect 37507 44285 37519 44319
rect 37918 44316 37924 44328
rect 37879 44288 37924 44316
rect 37461 44279 37519 44285
rect 37918 44276 37924 44288
rect 37976 44276 37982 44328
rect 34054 44208 34060 44260
rect 34112 44248 34118 44260
rect 34241 44251 34299 44257
rect 34241 44248 34253 44251
rect 34112 44220 34253 44248
rect 34112 44208 34118 44220
rect 34241 44217 34253 44220
rect 34287 44217 34299 44251
rect 34241 44211 34299 44217
rect 1995 44152 34008 44180
rect 34517 44183 34575 44189
rect 1995 44149 2007 44152
rect 1949 44143 2007 44149
rect 34517 44149 34529 44183
rect 34563 44180 34575 44183
rect 36722 44180 36728 44192
rect 34563 44152 36728 44180
rect 34563 44149 34575 44152
rect 34517 44143 34575 44149
rect 36722 44140 36728 44152
rect 36780 44140 36786 44192
rect 37274 44180 37280 44192
rect 37235 44152 37280 44180
rect 37274 44140 37280 44152
rect 37332 44140 37338 44192
rect 1104 44090 38824 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 38824 44090
rect 1104 44016 38824 44038
rect 33962 43936 33968 43988
rect 34020 43976 34026 43988
rect 34238 43976 34244 43988
rect 34020 43948 34244 43976
rect 34020 43936 34026 43948
rect 34238 43936 34244 43948
rect 34296 43936 34302 43988
rect 37182 43840 37188 43852
rect 37143 43812 37188 43840
rect 37182 43800 37188 43812
rect 37240 43800 37246 43852
rect 1104 43546 38824 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 38824 43546
rect 1104 43472 38824 43494
rect 15654 43432 15660 43444
rect 15615 43404 15660 43432
rect 15654 43392 15660 43404
rect 15712 43392 15718 43444
rect 16298 43392 16304 43444
rect 16356 43432 16362 43444
rect 25682 43432 25688 43444
rect 16356 43404 25688 43432
rect 16356 43392 16362 43404
rect 25682 43392 25688 43404
rect 25740 43392 25746 43444
rect 16577 43367 16635 43373
rect 16577 43333 16589 43367
rect 16623 43364 16635 43367
rect 18782 43364 18788 43376
rect 16623 43336 18788 43364
rect 16623 43333 16635 43336
rect 16577 43327 16635 43333
rect 18782 43324 18788 43336
rect 18840 43324 18846 43376
rect 15289 43299 15347 43305
rect 15289 43265 15301 43299
rect 15335 43296 15347 43299
rect 16209 43299 16267 43305
rect 16209 43296 16221 43299
rect 15335 43268 16221 43296
rect 15335 43265 15347 43268
rect 15289 43259 15347 43265
rect 16209 43265 16221 43268
rect 16255 43296 16267 43299
rect 16850 43296 16856 43308
rect 16255 43268 16856 43296
rect 16255 43265 16267 43268
rect 16209 43259 16267 43265
rect 16850 43256 16856 43268
rect 16908 43256 16914 43308
rect 1854 43228 1860 43240
rect 1815 43200 1860 43228
rect 1854 43188 1860 43200
rect 1912 43188 1918 43240
rect 15470 43228 15476 43240
rect 15431 43200 15476 43228
rect 15470 43188 15476 43200
rect 15528 43188 15534 43240
rect 16390 43228 16396 43240
rect 16351 43200 16396 43228
rect 16390 43188 16396 43200
rect 16448 43188 16454 43240
rect 37918 43228 37924 43240
rect 37879 43200 37924 43228
rect 37918 43188 37924 43200
rect 37976 43188 37982 43240
rect 1946 43092 1952 43104
rect 1907 43064 1952 43092
rect 1946 43052 1952 43064
rect 2004 43052 2010 43104
rect 1104 43002 38824 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 38824 43002
rect 1104 42928 38824 42950
rect 1946 42848 1952 42900
rect 2004 42888 2010 42900
rect 24854 42888 24860 42900
rect 2004 42860 24860 42888
rect 2004 42848 2010 42860
rect 24854 42848 24860 42860
rect 24912 42848 24918 42900
rect 1854 42752 1860 42764
rect 1815 42724 1860 42752
rect 1854 42712 1860 42724
rect 1912 42712 1918 42764
rect 16114 42752 16120 42764
rect 16075 42724 16120 42752
rect 16114 42712 16120 42724
rect 16172 42712 16178 42764
rect 16298 42752 16304 42764
rect 16259 42724 16304 42752
rect 16298 42712 16304 42724
rect 16356 42712 16362 42764
rect 17494 42752 17500 42764
rect 17455 42724 17500 42752
rect 17494 42712 17500 42724
rect 17552 42712 17558 42764
rect 17681 42755 17739 42761
rect 17681 42721 17693 42755
rect 17727 42752 17739 42755
rect 25590 42752 25596 42764
rect 17727 42724 25596 42752
rect 17727 42721 17739 42724
rect 17681 42715 17739 42721
rect 25590 42712 25596 42724
rect 25648 42712 25654 42764
rect 33042 42712 33048 42764
rect 33100 42752 33106 42764
rect 36814 42752 36820 42764
rect 33100 42724 36820 42752
rect 33100 42712 33106 42724
rect 36814 42712 36820 42724
rect 36872 42712 36878 42764
rect 37366 42752 37372 42764
rect 37327 42724 37372 42752
rect 37366 42712 37372 42724
rect 37424 42712 37430 42764
rect 15933 42687 15991 42693
rect 15933 42653 15945 42687
rect 15979 42684 15991 42687
rect 16850 42684 16856 42696
rect 15979 42656 16856 42684
rect 15979 42653 15991 42656
rect 15933 42647 15991 42653
rect 16850 42644 16856 42656
rect 16908 42684 16914 42696
rect 17313 42687 17371 42693
rect 17313 42684 17325 42687
rect 16908 42656 17325 42684
rect 16908 42644 16914 42656
rect 17313 42653 17325 42656
rect 17359 42653 17371 42687
rect 17313 42647 17371 42653
rect 33870 42616 33876 42628
rect 6886 42588 33876 42616
rect 1949 42551 2007 42557
rect 1949 42517 1961 42551
rect 1995 42548 2007 42551
rect 6886 42548 6914 42588
rect 33870 42576 33876 42588
rect 33928 42576 33934 42628
rect 1995 42520 6914 42548
rect 1995 42517 2007 42520
rect 1949 42511 2007 42517
rect 34422 42508 34428 42560
rect 34480 42548 34486 42560
rect 37185 42551 37243 42557
rect 37185 42548 37197 42551
rect 34480 42520 37197 42548
rect 34480 42508 34486 42520
rect 37185 42517 37197 42520
rect 37231 42517 37243 42551
rect 37185 42511 37243 42517
rect 1104 42458 38824 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 38824 42458
rect 1104 42384 38824 42406
rect 16574 42304 16580 42356
rect 16632 42344 16638 42356
rect 16632 42316 16677 42344
rect 16632 42304 16638 42316
rect 37274 42304 37280 42356
rect 37332 42304 37338 42356
rect 16209 42211 16267 42217
rect 16209 42177 16221 42211
rect 16255 42208 16267 42211
rect 16850 42208 16856 42220
rect 16255 42180 16856 42208
rect 16255 42177 16267 42180
rect 16209 42171 16267 42177
rect 16850 42168 16856 42180
rect 16908 42168 16914 42220
rect 37292 42208 37320 42304
rect 35820 42180 37320 42208
rect 16298 42100 16304 42152
rect 16356 42140 16362 42152
rect 16393 42143 16451 42149
rect 16393 42140 16405 42143
rect 16356 42112 16405 42140
rect 16356 42100 16362 42112
rect 16393 42109 16405 42112
rect 16439 42109 16451 42143
rect 16393 42103 16451 42109
rect 24854 42100 24860 42152
rect 24912 42140 24918 42152
rect 33778 42140 33784 42152
rect 24912 42112 26234 42140
rect 33739 42112 33784 42140
rect 24912 42100 24918 42112
rect 26206 42072 26234 42112
rect 33778 42100 33784 42112
rect 33836 42100 33842 42152
rect 33874 42143 33932 42149
rect 33874 42109 33886 42143
rect 33920 42109 33932 42143
rect 33874 42103 33932 42109
rect 33888 42072 33916 42103
rect 33962 42100 33968 42152
rect 34020 42140 34026 42152
rect 34149 42143 34207 42149
rect 34149 42140 34161 42143
rect 34020 42112 34161 42140
rect 34020 42100 34026 42112
rect 34149 42109 34161 42112
rect 34195 42109 34207 42143
rect 34149 42103 34207 42109
rect 34287 42143 34345 42149
rect 34287 42109 34299 42143
rect 34333 42140 34345 42143
rect 35820 42140 35848 42180
rect 37274 42140 37280 42152
rect 34333 42112 35848 42140
rect 37235 42112 37280 42140
rect 34333 42109 34345 42112
rect 34287 42103 34345 42109
rect 37274 42100 37280 42112
rect 37332 42100 37338 42152
rect 37918 42140 37924 42152
rect 37879 42112 37924 42140
rect 37918 42100 37924 42112
rect 37976 42100 37982 42152
rect 34054 42072 34060 42084
rect 26206 42044 33916 42072
rect 34015 42044 34060 42072
rect 34054 42032 34060 42044
rect 34112 42032 34118 42084
rect 34330 41964 34336 42016
rect 34388 42004 34394 42016
rect 34425 42007 34483 42013
rect 34425 42004 34437 42007
rect 34388 41976 34437 42004
rect 34388 41964 34394 41976
rect 34425 41973 34437 41976
rect 34471 41973 34483 42007
rect 34425 41967 34483 41973
rect 1104 41914 38824 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 38824 41914
rect 1104 41840 38824 41862
rect 1854 41732 1860 41744
rect 1815 41704 1860 41732
rect 1854 41692 1860 41704
rect 1912 41692 1918 41744
rect 34054 41732 34060 41744
rect 33967 41704 34060 41732
rect 34054 41692 34060 41704
rect 34112 41692 34118 41744
rect 33781 41667 33839 41673
rect 33781 41633 33793 41667
rect 33827 41633 33839 41667
rect 33781 41627 33839 41633
rect 2041 41531 2099 41537
rect 2041 41497 2053 41531
rect 2087 41528 2099 41531
rect 2682 41528 2688 41540
rect 2087 41500 2688 41528
rect 2087 41497 2099 41500
rect 2041 41491 2099 41497
rect 2682 41488 2688 41500
rect 2740 41488 2746 41540
rect 30926 41420 30932 41472
rect 30984 41460 30990 41472
rect 32398 41460 32404 41472
rect 30984 41432 32404 41460
rect 30984 41420 30990 41432
rect 32398 41420 32404 41432
rect 32456 41420 32462 41472
rect 33796 41460 33824 41627
rect 33870 41624 33876 41676
rect 33928 41664 33934 41676
rect 33928 41636 33973 41664
rect 33928 41624 33934 41636
rect 34073 41596 34101 41692
rect 34149 41667 34207 41673
rect 34149 41633 34161 41667
rect 34195 41633 34207 41667
rect 34149 41627 34207 41633
rect 34287 41667 34345 41673
rect 34287 41633 34299 41667
rect 34333 41664 34345 41667
rect 34422 41664 34428 41676
rect 34333 41636 34428 41664
rect 34333 41633 34345 41636
rect 34287 41627 34345 41633
rect 33888 41568 34101 41596
rect 33888 41540 33916 41568
rect 33870 41488 33876 41540
rect 33928 41488 33934 41540
rect 34054 41488 34060 41540
rect 34112 41528 34118 41540
rect 34164 41528 34192 41627
rect 34422 41624 34428 41636
rect 34480 41624 34486 41676
rect 37182 41624 37188 41676
rect 37240 41664 37246 41676
rect 37369 41667 37427 41673
rect 37369 41664 37381 41667
rect 37240 41636 37381 41664
rect 37240 41624 37246 41636
rect 37369 41633 37381 41636
rect 37415 41633 37427 41667
rect 37369 41627 37427 41633
rect 39022 41596 39028 41608
rect 34112 41500 34192 41528
rect 34348 41568 39028 41596
rect 34112 41488 34118 41500
rect 34348 41460 34376 41568
rect 39022 41556 39028 41568
rect 39080 41556 39086 41608
rect 35250 41488 35256 41540
rect 35308 41528 35314 41540
rect 37185 41531 37243 41537
rect 37185 41528 37197 41531
rect 35308 41500 37197 41528
rect 35308 41488 35314 41500
rect 37185 41497 37197 41500
rect 37231 41497 37243 41531
rect 37185 41491 37243 41497
rect 33796 41432 34376 41460
rect 34425 41463 34483 41469
rect 34425 41429 34437 41463
rect 34471 41460 34483 41463
rect 35894 41460 35900 41472
rect 34471 41432 35900 41460
rect 34471 41429 34483 41432
rect 34425 41423 34483 41429
rect 35894 41420 35900 41432
rect 35952 41420 35958 41472
rect 1104 41370 38824 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 38824 41370
rect 1104 41296 38824 41318
rect 26142 41080 26148 41132
rect 26200 41120 26206 41132
rect 26200 41092 31754 41120
rect 26200 41080 26206 41092
rect 2682 41012 2688 41064
rect 2740 41052 2746 41064
rect 31726 41052 31754 41092
rect 33689 41055 33747 41061
rect 33689 41052 33701 41055
rect 2740 41024 26234 41052
rect 31726 41024 33701 41052
rect 2740 41012 2746 41024
rect 1854 40984 1860 40996
rect 1815 40956 1860 40984
rect 1854 40944 1860 40956
rect 1912 40944 1918 40996
rect 2041 40987 2099 40993
rect 2041 40953 2053 40987
rect 2087 40984 2099 40987
rect 2590 40984 2596 40996
rect 2087 40956 2596 40984
rect 2087 40953 2099 40956
rect 2041 40947 2099 40953
rect 2590 40944 2596 40956
rect 2648 40944 2654 40996
rect 26206 40984 26234 41024
rect 33689 41021 33701 41024
rect 33735 41021 33747 41055
rect 33689 41015 33747 41021
rect 33782 41055 33840 41061
rect 33782 41021 33794 41055
rect 33828 41021 33840 41055
rect 33782 41015 33840 41021
rect 33796 40984 33824 41015
rect 33870 41012 33876 41064
rect 33928 41052 33934 41064
rect 33965 41055 34023 41061
rect 33965 41052 33977 41055
rect 33928 41024 33977 41052
rect 33928 41012 33934 41024
rect 33965 41021 33977 41024
rect 34011 41021 34023 41055
rect 33965 41015 34023 41021
rect 34195 41055 34253 41061
rect 34195 41021 34207 41055
rect 34241 41052 34253 41055
rect 35250 41052 35256 41064
rect 34241 41024 35256 41052
rect 34241 41021 34253 41024
rect 34195 41015 34253 41021
rect 35250 41012 35256 41024
rect 35308 41012 35314 41064
rect 37274 41052 37280 41064
rect 37235 41024 37280 41052
rect 37274 41012 37280 41024
rect 37332 41012 37338 41064
rect 37918 41052 37924 41064
rect 37879 41024 37924 41052
rect 37918 41012 37924 41024
rect 37976 41012 37982 41064
rect 34054 40984 34060 40996
rect 26206 40956 33824 40984
rect 34015 40956 34060 40984
rect 34054 40944 34060 40956
rect 34112 40944 34118 40996
rect 34333 40919 34391 40925
rect 34333 40885 34345 40919
rect 34379 40916 34391 40919
rect 35434 40916 35440 40928
rect 34379 40888 35440 40916
rect 34379 40885 34391 40888
rect 34333 40879 34391 40885
rect 35434 40876 35440 40888
rect 35492 40876 35498 40928
rect 1104 40826 38824 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 38824 40826
rect 1104 40752 38824 40774
rect 1854 40576 1860 40588
rect 1815 40548 1860 40576
rect 1854 40536 1860 40548
rect 1912 40536 1918 40588
rect 17218 40536 17224 40588
rect 17276 40576 17282 40588
rect 17497 40579 17555 40585
rect 17497 40576 17509 40579
rect 17276 40548 17509 40576
rect 17276 40536 17282 40548
rect 17497 40545 17509 40548
rect 17543 40545 17555 40579
rect 17497 40539 17555 40545
rect 17310 40508 17316 40520
rect 17271 40480 17316 40508
rect 17310 40468 17316 40480
rect 17368 40468 17374 40520
rect 2041 40443 2099 40449
rect 2041 40409 2053 40443
rect 2087 40440 2099 40443
rect 2682 40440 2688 40452
rect 2087 40412 2688 40440
rect 2087 40409 2099 40412
rect 2041 40403 2099 40409
rect 2682 40400 2688 40412
rect 2740 40400 2746 40452
rect 17681 40375 17739 40381
rect 17681 40341 17693 40375
rect 17727 40372 17739 40375
rect 29638 40372 29644 40384
rect 17727 40344 29644 40372
rect 17727 40341 17739 40344
rect 17681 40335 17739 40341
rect 29638 40332 29644 40344
rect 29696 40332 29702 40384
rect 36170 40332 36176 40384
rect 36228 40372 36234 40384
rect 36814 40372 36820 40384
rect 36228 40344 36820 40372
rect 36228 40332 36234 40344
rect 36814 40332 36820 40344
rect 36872 40332 36878 40384
rect 1104 40282 38824 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 38824 40282
rect 1104 40208 38824 40230
rect 17678 40168 17684 40180
rect 17639 40140 17684 40168
rect 17678 40128 17684 40140
rect 17736 40128 17742 40180
rect 17310 40060 17316 40112
rect 17368 40100 17374 40112
rect 17368 40072 17816 40100
rect 17368 40060 17374 40072
rect 2590 39992 2596 40044
rect 2648 40032 2654 40044
rect 2648 40004 6914 40032
rect 2648 39992 2654 40004
rect 6886 39828 6914 40004
rect 9122 39992 9128 40044
rect 9180 40032 9186 40044
rect 16022 40032 16028 40044
rect 9180 40004 15884 40032
rect 15983 40004 16028 40032
rect 9180 39992 9186 40004
rect 15856 39973 15884 40004
rect 16022 39992 16028 40004
rect 16080 39992 16086 40044
rect 16485 40035 16543 40041
rect 16485 40032 16497 40035
rect 16224 40004 16497 40032
rect 15749 39967 15807 39973
rect 15749 39933 15761 39967
rect 15795 39933 15807 39967
rect 15749 39927 15807 39933
rect 15841 39967 15899 39973
rect 15841 39933 15853 39967
rect 15887 39933 15899 39967
rect 15841 39927 15899 39933
rect 15764 39896 15792 39927
rect 16224 39896 16252 40004
rect 16485 40001 16497 40004
rect 16531 40032 16543 40035
rect 16853 40035 16911 40041
rect 16531 40004 16804 40032
rect 16531 40001 16543 40004
rect 16485 39995 16543 40001
rect 16666 39964 16672 39976
rect 16627 39936 16672 39964
rect 16666 39924 16672 39936
rect 16724 39924 16730 39976
rect 16776 39964 16804 40004
rect 16853 40001 16865 40035
rect 16899 40032 16911 40035
rect 17788 40032 17816 40072
rect 36170 40060 36176 40112
rect 36228 40100 36234 40112
rect 36630 40100 36636 40112
rect 36228 40072 36636 40100
rect 36228 40060 36234 40072
rect 36630 40060 36636 40072
rect 36688 40060 36694 40112
rect 18141 40035 18199 40041
rect 18141 40032 18153 40035
rect 16899 40004 17632 40032
rect 17788 40004 18153 40032
rect 16899 40001 16911 40004
rect 16853 39995 16911 40001
rect 17310 39964 17316 39976
rect 16776 39936 17316 39964
rect 17310 39924 17316 39936
rect 17368 39924 17374 39976
rect 17497 39967 17555 39973
rect 17497 39933 17509 39967
rect 17543 39933 17555 39967
rect 17497 39927 17555 39933
rect 15764 39868 16252 39896
rect 16546 39868 17080 39896
rect 16546 39828 16574 39868
rect 6886 39800 16574 39828
rect 17052 39828 17080 39868
rect 17126 39856 17132 39908
rect 17184 39896 17190 39908
rect 17512 39896 17540 39927
rect 17184 39868 17540 39896
rect 17604 39896 17632 40004
rect 18141 40001 18153 40004
rect 18187 40001 18199 40035
rect 18506 40032 18512 40044
rect 18467 40004 18512 40032
rect 18141 39995 18199 40001
rect 18506 39992 18512 40004
rect 18564 39992 18570 40044
rect 38102 40032 38108 40044
rect 33704 40004 38108 40032
rect 18322 39964 18328 39976
rect 18283 39936 18328 39964
rect 18322 39924 18328 39936
rect 18380 39924 18386 39976
rect 33704 39973 33732 40004
rect 38102 39992 38108 40004
rect 38160 39992 38166 40044
rect 33689 39967 33747 39973
rect 33689 39933 33701 39967
rect 33735 39933 33747 39967
rect 33689 39927 33747 39933
rect 33782 39967 33840 39973
rect 33782 39933 33794 39967
rect 33828 39933 33840 39967
rect 33782 39927 33840 39933
rect 18690 39896 18696 39908
rect 17604 39868 18696 39896
rect 17184 39856 17190 39868
rect 18690 39856 18696 39868
rect 18748 39856 18754 39908
rect 33796 39828 33824 39927
rect 33870 39924 33876 39976
rect 33928 39964 33934 39976
rect 33965 39967 34023 39973
rect 33965 39964 33977 39967
rect 33928 39936 33977 39964
rect 33928 39924 33934 39936
rect 33965 39933 33977 39936
rect 34011 39933 34023 39967
rect 33965 39927 34023 39933
rect 34195 39967 34253 39973
rect 34195 39933 34207 39967
rect 34241 39964 34253 39967
rect 37458 39964 37464 39976
rect 34241 39936 37320 39964
rect 37419 39936 37464 39964
rect 34241 39933 34253 39936
rect 34195 39927 34253 39933
rect 34054 39896 34060 39908
rect 34015 39868 34060 39896
rect 34054 39856 34060 39868
rect 34112 39856 34118 39908
rect 17052 39800 33824 39828
rect 34333 39831 34391 39837
rect 34333 39797 34345 39831
rect 34379 39828 34391 39831
rect 36630 39828 36636 39840
rect 34379 39800 36636 39828
rect 34379 39797 34391 39800
rect 34333 39791 34391 39797
rect 36630 39788 36636 39800
rect 36688 39788 36694 39840
rect 37292 39837 37320 39936
rect 37458 39924 37464 39936
rect 37516 39924 37522 39976
rect 37918 39964 37924 39976
rect 37879 39936 37924 39964
rect 37918 39924 37924 39936
rect 37976 39924 37982 39976
rect 37277 39831 37335 39837
rect 37277 39797 37289 39831
rect 37323 39797 37335 39831
rect 37277 39791 37335 39797
rect 1104 39738 38824 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 38824 39738
rect 1104 39664 38824 39686
rect 26206 39528 33824 39556
rect 1854 39488 1860 39500
rect 1815 39460 1860 39488
rect 1854 39448 1860 39460
rect 1912 39448 1918 39500
rect 2682 39448 2688 39500
rect 2740 39488 2746 39500
rect 26206 39488 26234 39528
rect 33796 39497 33824 39528
rect 33870 39516 33876 39568
rect 33928 39556 33934 39568
rect 33965 39559 34023 39565
rect 33965 39556 33977 39559
rect 33928 39528 33977 39556
rect 33928 39516 33934 39528
rect 33965 39525 33977 39528
rect 34011 39525 34023 39559
rect 33965 39519 34023 39525
rect 2740 39460 26234 39488
rect 33689 39491 33747 39497
rect 2740 39448 2746 39460
rect 33689 39457 33701 39491
rect 33735 39457 33747 39491
rect 33689 39451 33747 39457
rect 33782 39491 33840 39497
rect 33782 39457 33794 39491
rect 33828 39457 33840 39491
rect 34054 39488 34060 39500
rect 34015 39460 34060 39488
rect 33782 39451 33840 39457
rect 33704 39420 33732 39451
rect 34054 39448 34060 39460
rect 34112 39448 34118 39500
rect 34195 39491 34253 39497
rect 34195 39457 34207 39491
rect 34241 39488 34253 39491
rect 37274 39488 37280 39500
rect 34241 39460 37280 39488
rect 34241 39457 34253 39460
rect 34195 39451 34253 39457
rect 37274 39448 37280 39460
rect 37332 39448 37338 39500
rect 38562 39420 38568 39432
rect 33704 39392 38568 39420
rect 38562 39380 38568 39392
rect 38620 39380 38626 39432
rect 2041 39355 2099 39361
rect 2041 39321 2053 39355
rect 2087 39352 2099 39355
rect 2682 39352 2688 39364
rect 2087 39324 2688 39352
rect 2087 39321 2099 39324
rect 2041 39315 2099 39321
rect 2682 39312 2688 39324
rect 2740 39312 2746 39364
rect 34333 39287 34391 39293
rect 34333 39253 34345 39287
rect 34379 39284 34391 39287
rect 34422 39284 34428 39296
rect 34379 39256 34428 39284
rect 34379 39253 34391 39256
rect 34333 39247 34391 39253
rect 34422 39244 34428 39256
rect 34480 39244 34486 39296
rect 1104 39194 38824 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 38824 39194
rect 1104 39120 38824 39142
rect 37274 39080 37280 39092
rect 37235 39052 37280 39080
rect 37274 39040 37280 39052
rect 37332 39040 37338 39092
rect 37458 38876 37464 38888
rect 37419 38848 37464 38876
rect 37458 38836 37464 38848
rect 37516 38836 37522 38888
rect 37918 38876 37924 38888
rect 37879 38848 37924 38876
rect 37918 38836 37924 38848
rect 37976 38836 37982 38888
rect 1854 38808 1860 38820
rect 1815 38780 1860 38808
rect 1854 38768 1860 38780
rect 1912 38768 1918 38820
rect 2041 38811 2099 38817
rect 2041 38777 2053 38811
rect 2087 38808 2099 38811
rect 2590 38808 2596 38820
rect 2087 38780 2596 38808
rect 2087 38777 2099 38780
rect 2041 38771 2099 38777
rect 2590 38768 2596 38780
rect 2648 38768 2654 38820
rect 32766 38700 32772 38752
rect 32824 38740 32830 38752
rect 35802 38740 35808 38752
rect 32824 38712 35808 38740
rect 32824 38700 32830 38712
rect 35802 38700 35808 38712
rect 35860 38700 35866 38752
rect 1104 38650 38824 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 38824 38650
rect 1104 38576 38824 38598
rect 33686 38496 33692 38548
rect 33744 38536 33750 38548
rect 34057 38539 34115 38545
rect 34057 38536 34069 38539
rect 33744 38508 34069 38536
rect 33744 38496 33750 38508
rect 34057 38505 34069 38508
rect 34103 38505 34115 38539
rect 34057 38499 34115 38505
rect 34330 38496 34336 38548
rect 34388 38536 34394 38548
rect 34790 38536 34796 38548
rect 34388 38508 34796 38536
rect 34388 38496 34394 38508
rect 34790 38496 34796 38508
rect 34848 38496 34854 38548
rect 28902 38428 28908 38480
rect 28960 38468 28966 38480
rect 28997 38471 29055 38477
rect 28997 38468 29009 38471
rect 28960 38440 29009 38468
rect 28960 38428 28966 38440
rect 28997 38437 29009 38440
rect 29043 38437 29055 38471
rect 33410 38468 33416 38480
rect 33371 38440 33416 38468
rect 28997 38431 29055 38437
rect 33410 38428 33416 38440
rect 33468 38428 33474 38480
rect 33502 38428 33508 38480
rect 33560 38468 33566 38480
rect 36354 38468 36360 38480
rect 33560 38440 36360 38468
rect 33560 38428 33566 38440
rect 36354 38428 36360 38440
rect 36412 38428 36418 38480
rect 33229 38403 33287 38409
rect 33229 38369 33241 38403
rect 33275 38400 33287 38403
rect 33778 38400 33784 38412
rect 33275 38372 33784 38400
rect 33275 38369 33287 38372
rect 33229 38363 33287 38369
rect 33778 38360 33784 38372
rect 33836 38360 33842 38412
rect 33965 38403 34023 38409
rect 33965 38369 33977 38403
rect 34011 38400 34023 38403
rect 34330 38400 34336 38412
rect 34011 38372 34336 38400
rect 34011 38369 34023 38372
rect 33965 38363 34023 38369
rect 34330 38360 34336 38372
rect 34388 38360 34394 38412
rect 34514 38360 34520 38412
rect 34572 38400 34578 38412
rect 34609 38403 34667 38409
rect 34609 38400 34621 38403
rect 34572 38372 34621 38400
rect 34572 38360 34578 38372
rect 34609 38369 34621 38372
rect 34655 38369 34667 38403
rect 37182 38400 37188 38412
rect 37143 38372 37188 38400
rect 34609 38363 34667 38369
rect 37182 38360 37188 38372
rect 37240 38360 37246 38412
rect 29181 38267 29239 38273
rect 29181 38233 29193 38267
rect 29227 38264 29239 38267
rect 33686 38264 33692 38276
rect 29227 38236 33692 38264
rect 29227 38233 29239 38236
rect 29181 38227 29239 38233
rect 33686 38224 33692 38236
rect 33744 38224 33750 38276
rect 33594 38156 33600 38208
rect 33652 38196 33658 38208
rect 34793 38199 34851 38205
rect 34793 38196 34805 38199
rect 33652 38168 34805 38196
rect 33652 38156 33658 38168
rect 34793 38165 34805 38168
rect 34839 38165 34851 38199
rect 34793 38159 34851 38165
rect 1104 38106 38824 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 38824 38106
rect 1104 38032 38824 38054
rect 37090 37856 37096 37868
rect 33336 37828 37096 37856
rect 1854 37788 1860 37800
rect 1815 37760 1860 37788
rect 1854 37748 1860 37760
rect 1912 37748 1918 37800
rect 33336 37797 33364 37828
rect 37090 37816 37096 37828
rect 37148 37816 37154 37868
rect 33321 37791 33379 37797
rect 33321 37757 33333 37791
rect 33367 37757 33379 37791
rect 33321 37751 33379 37757
rect 33414 37791 33472 37797
rect 33414 37757 33426 37791
rect 33460 37757 33472 37791
rect 33594 37788 33600 37800
rect 33555 37760 33600 37788
rect 33414 37751 33472 37757
rect 2041 37723 2099 37729
rect 2041 37689 2053 37723
rect 2087 37720 2099 37723
rect 4062 37720 4068 37732
rect 2087 37692 4068 37720
rect 2087 37689 2099 37692
rect 2041 37683 2099 37689
rect 4062 37680 4068 37692
rect 4120 37680 4126 37732
rect 33428 37720 33456 37751
rect 33594 37748 33600 37760
rect 33652 37748 33658 37800
rect 33686 37748 33692 37800
rect 33744 37788 33750 37800
rect 33827 37791 33885 37797
rect 33744 37760 33789 37788
rect 33744 37748 33750 37760
rect 33827 37757 33839 37791
rect 33873 37788 33885 37791
rect 37182 37788 37188 37800
rect 33873 37760 37188 37788
rect 33873 37757 33885 37760
rect 33827 37751 33885 37757
rect 37182 37748 37188 37760
rect 37240 37748 37246 37800
rect 37918 37788 37924 37800
rect 37879 37760 37924 37788
rect 37918 37748 37924 37760
rect 37976 37748 37982 37800
rect 33152 37692 33456 37720
rect 2682 37612 2688 37664
rect 2740 37652 2746 37664
rect 33152 37661 33180 37692
rect 33137 37655 33195 37661
rect 33137 37652 33149 37655
rect 2740 37624 33149 37652
rect 2740 37612 2746 37624
rect 33137 37621 33149 37624
rect 33183 37621 33195 37655
rect 33137 37615 33195 37621
rect 33965 37655 34023 37661
rect 33965 37621 33977 37655
rect 34011 37652 34023 37655
rect 34054 37652 34060 37664
rect 34011 37624 34060 37652
rect 34011 37621 34023 37624
rect 33965 37615 34023 37621
rect 34054 37612 34060 37624
rect 34112 37612 34118 37664
rect 1104 37562 38824 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 38824 37562
rect 1104 37488 38824 37510
rect 34514 37408 34520 37460
rect 34572 37408 34578 37460
rect 37182 37448 37188 37460
rect 37143 37420 37188 37448
rect 37182 37408 37188 37420
rect 37240 37408 37246 37460
rect 1854 37312 1860 37324
rect 1815 37284 1860 37312
rect 1854 37272 1860 37284
rect 1912 37272 1918 37324
rect 2041 37315 2099 37321
rect 2041 37281 2053 37315
rect 2087 37312 2099 37315
rect 2682 37312 2688 37324
rect 2087 37284 2688 37312
rect 2087 37281 2099 37284
rect 2041 37275 2099 37281
rect 2682 37272 2688 37284
rect 2740 37272 2746 37324
rect 34532 37312 34560 37408
rect 37366 37312 37372 37324
rect 34440 37284 34560 37312
rect 37327 37284 37372 37312
rect 34440 37256 34468 37284
rect 37366 37272 37372 37284
rect 37424 37272 37430 37324
rect 34422 37204 34428 37256
rect 34480 37204 34486 37256
rect 1104 37018 38824 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 38824 37018
rect 1104 36944 38824 36966
rect 33870 36864 33876 36916
rect 33928 36904 33934 36916
rect 34517 36907 34575 36913
rect 34517 36904 34529 36907
rect 33928 36876 34529 36904
rect 33928 36864 33934 36876
rect 34517 36873 34529 36876
rect 34563 36873 34575 36907
rect 34517 36867 34575 36873
rect 36354 36864 36360 36916
rect 36412 36904 36418 36916
rect 36538 36904 36544 36916
rect 36412 36876 36544 36904
rect 36412 36864 36418 36876
rect 36538 36864 36544 36876
rect 36596 36864 36602 36916
rect 38286 36836 38292 36848
rect 33244 36808 38292 36836
rect 33244 36709 33272 36808
rect 38286 36796 38292 36808
rect 38344 36796 38350 36848
rect 33594 36768 33600 36780
rect 33520 36740 33600 36768
rect 33520 36709 33548 36740
rect 33594 36728 33600 36740
rect 33652 36728 33658 36780
rect 33229 36703 33287 36709
rect 33229 36669 33241 36703
rect 33275 36669 33287 36703
rect 33229 36663 33287 36669
rect 33322 36703 33380 36709
rect 33322 36669 33334 36703
rect 33368 36669 33380 36703
rect 33322 36663 33380 36669
rect 33505 36703 33563 36709
rect 33505 36669 33517 36703
rect 33551 36669 33563 36703
rect 33505 36663 33563 36669
rect 33735 36703 33793 36709
rect 33735 36669 33747 36703
rect 33781 36700 33793 36703
rect 37090 36700 37096 36712
rect 33781 36672 37096 36700
rect 33781 36669 33793 36672
rect 33735 36663 33793 36669
rect 33336 36632 33364 36663
rect 37090 36660 37096 36672
rect 37148 36660 37154 36712
rect 37274 36700 37280 36712
rect 37235 36672 37280 36700
rect 37274 36660 37280 36672
rect 37332 36660 37338 36712
rect 37918 36700 37924 36712
rect 37879 36672 37924 36700
rect 37918 36660 37924 36672
rect 37976 36660 37982 36712
rect 33152 36604 33364 36632
rect 33597 36635 33655 36641
rect 2590 36524 2596 36576
rect 2648 36564 2654 36576
rect 33152 36573 33180 36604
rect 33597 36601 33609 36635
rect 33643 36632 33655 36635
rect 33643 36604 33732 36632
rect 33643 36601 33655 36604
rect 33597 36595 33655 36601
rect 33704 36576 33732 36604
rect 34330 36592 34336 36644
rect 34388 36632 34394 36644
rect 34425 36635 34483 36641
rect 34425 36632 34437 36635
rect 34388 36604 34437 36632
rect 34388 36592 34394 36604
rect 34425 36601 34437 36604
rect 34471 36601 34483 36635
rect 34425 36595 34483 36601
rect 33137 36567 33195 36573
rect 33137 36564 33149 36567
rect 2648 36536 33149 36564
rect 2648 36524 2654 36536
rect 33137 36533 33149 36536
rect 33183 36533 33195 36567
rect 33137 36527 33195 36533
rect 33686 36524 33692 36576
rect 33744 36524 33750 36576
rect 33870 36564 33876 36576
rect 33831 36536 33876 36564
rect 33870 36524 33876 36536
rect 33928 36524 33934 36576
rect 1104 36474 38824 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 38824 36474
rect 1104 36400 38824 36422
rect 28813 36363 28871 36369
rect 28813 36329 28825 36363
rect 28859 36360 28871 36363
rect 32398 36360 32404 36372
rect 28859 36332 32404 36360
rect 28859 36329 28871 36332
rect 28813 36323 28871 36329
rect 32398 36320 32404 36332
rect 32456 36320 32462 36372
rect 33594 36360 33600 36372
rect 33520 36332 33600 36360
rect 4062 36252 4068 36304
rect 4120 36292 4126 36304
rect 28718 36292 28724 36304
rect 4120 36264 26234 36292
rect 28631 36264 28724 36292
rect 4120 36252 4126 36264
rect 1854 36224 1860 36236
rect 1815 36196 1860 36224
rect 1854 36184 1860 36196
rect 1912 36184 1918 36236
rect 26206 36224 26234 36264
rect 28718 36252 28724 36264
rect 28776 36292 28782 36304
rect 28902 36292 28908 36304
rect 28776 36264 28908 36292
rect 28776 36252 28782 36264
rect 28902 36252 28908 36264
rect 28960 36252 28966 36304
rect 33520 36301 33548 36332
rect 33594 36320 33600 36332
rect 33652 36320 33658 36372
rect 33686 36320 33692 36372
rect 33744 36320 33750 36372
rect 33962 36320 33968 36372
rect 34020 36360 34026 36372
rect 34517 36363 34575 36369
rect 34517 36360 34529 36363
rect 34020 36332 34529 36360
rect 34020 36320 34026 36332
rect 34517 36329 34529 36332
rect 34563 36329 34575 36363
rect 34517 36323 34575 36329
rect 37090 36320 37096 36372
rect 37148 36360 37154 36372
rect 37185 36363 37243 36369
rect 37185 36360 37197 36363
rect 37148 36332 37197 36360
rect 37148 36320 37154 36332
rect 37185 36329 37197 36332
rect 37231 36329 37243 36363
rect 37185 36323 37243 36329
rect 33505 36295 33563 36301
rect 33152 36264 33364 36292
rect 33152 36233 33180 36264
rect 33336 36233 33364 36264
rect 33505 36261 33517 36295
rect 33551 36261 33563 36295
rect 33704 36292 33732 36320
rect 33505 36255 33563 36261
rect 33612 36264 33732 36292
rect 33612 36233 33640 36264
rect 33870 36252 33876 36304
rect 33928 36292 33934 36304
rect 34698 36292 34704 36304
rect 33928 36264 34704 36292
rect 33928 36252 33934 36264
rect 34698 36252 34704 36264
rect 34756 36252 34762 36304
rect 33137 36227 33195 36233
rect 33137 36224 33149 36227
rect 26206 36196 33149 36224
rect 33137 36193 33149 36196
rect 33183 36193 33195 36227
rect 33137 36187 33195 36193
rect 33229 36227 33287 36233
rect 33229 36193 33241 36227
rect 33275 36193 33287 36227
rect 33229 36187 33287 36193
rect 33322 36227 33380 36233
rect 33322 36193 33334 36227
rect 33368 36193 33380 36227
rect 33322 36187 33380 36193
rect 33597 36227 33655 36233
rect 33597 36193 33609 36227
rect 33643 36193 33655 36227
rect 33597 36187 33655 36193
rect 33735 36227 33793 36233
rect 33735 36193 33747 36227
rect 33781 36224 33793 36227
rect 33962 36224 33968 36236
rect 33781 36196 33968 36224
rect 33781 36193 33793 36196
rect 33735 36187 33793 36193
rect 33244 36156 33272 36187
rect 33962 36184 33968 36196
rect 34020 36184 34026 36236
rect 34425 36227 34483 36233
rect 34425 36193 34437 36227
rect 34471 36224 34483 36227
rect 34882 36224 34888 36236
rect 34471 36196 34888 36224
rect 34471 36193 34483 36196
rect 34425 36187 34483 36193
rect 34882 36184 34888 36196
rect 34940 36184 34946 36236
rect 37366 36224 37372 36236
rect 37327 36196 37372 36224
rect 37366 36184 37372 36196
rect 37424 36184 37430 36236
rect 33502 36156 33508 36168
rect 33244 36128 33508 36156
rect 33502 36116 33508 36128
rect 33560 36116 33566 36168
rect 35342 36116 35348 36168
rect 35400 36156 35406 36168
rect 36262 36156 36268 36168
rect 35400 36128 36268 36156
rect 35400 36116 35406 36128
rect 36262 36116 36268 36128
rect 36320 36116 36326 36168
rect 2041 36091 2099 36097
rect 2041 36057 2053 36091
rect 2087 36088 2099 36091
rect 2682 36088 2688 36100
rect 2087 36060 2688 36088
rect 2087 36057 2099 36060
rect 2041 36051 2099 36057
rect 2682 36048 2688 36060
rect 2740 36048 2746 36100
rect 33873 36023 33931 36029
rect 33873 35989 33885 36023
rect 33919 36020 33931 36023
rect 35342 36020 35348 36032
rect 33919 35992 35348 36020
rect 33919 35989 33931 35992
rect 33873 35983 33931 35989
rect 35342 35980 35348 35992
rect 35400 35980 35406 36032
rect 1104 35930 38824 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 38824 35930
rect 1104 35856 38824 35878
rect 33134 35776 33140 35828
rect 33192 35816 33198 35828
rect 36170 35816 36176 35828
rect 33192 35788 36176 35816
rect 33192 35776 33198 35788
rect 36170 35776 36176 35788
rect 36228 35776 36234 35828
rect 35250 35748 35256 35760
rect 33244 35720 35256 35748
rect 2590 35572 2596 35624
rect 2648 35612 2654 35624
rect 33244 35621 33272 35720
rect 35250 35708 35256 35720
rect 35308 35708 35314 35760
rect 33594 35640 33600 35692
rect 33652 35640 33658 35692
rect 33137 35615 33195 35621
rect 33137 35612 33149 35615
rect 2648 35584 33149 35612
rect 2648 35572 2654 35584
rect 33137 35581 33149 35584
rect 33183 35581 33195 35615
rect 33137 35575 33195 35581
rect 33229 35615 33287 35621
rect 33229 35581 33241 35615
rect 33275 35581 33287 35615
rect 33229 35575 33287 35581
rect 33322 35615 33380 35621
rect 33322 35581 33334 35615
rect 33368 35581 33380 35615
rect 33322 35575 33380 35581
rect 33505 35615 33563 35621
rect 33505 35581 33517 35615
rect 33551 35612 33563 35615
rect 33612 35612 33640 35640
rect 33551 35584 33640 35612
rect 33735 35615 33793 35621
rect 33551 35581 33563 35584
rect 33505 35575 33563 35581
rect 33735 35581 33747 35615
rect 33781 35612 33793 35615
rect 36170 35612 36176 35624
rect 33781 35584 36176 35612
rect 33781 35581 33793 35584
rect 33735 35575 33793 35581
rect 1854 35544 1860 35556
rect 1815 35516 1860 35544
rect 1854 35504 1860 35516
rect 1912 35504 1918 35556
rect 2041 35547 2099 35553
rect 2041 35513 2053 35547
rect 2087 35544 2099 35547
rect 2406 35544 2412 35556
rect 2087 35516 2412 35544
rect 2087 35513 2099 35516
rect 2041 35507 2099 35513
rect 2406 35504 2412 35516
rect 2464 35504 2470 35556
rect 28718 35504 28724 35556
rect 28776 35544 28782 35556
rect 28813 35547 28871 35553
rect 28813 35544 28825 35547
rect 28776 35516 28825 35544
rect 28776 35504 28782 35516
rect 28813 35513 28825 35516
rect 28859 35513 28871 35547
rect 28813 35507 28871 35513
rect 28997 35547 29055 35553
rect 28997 35513 29009 35547
rect 29043 35513 29055 35547
rect 33152 35544 33180 35575
rect 33336 35544 33364 35575
rect 36170 35572 36176 35584
rect 36228 35572 36234 35624
rect 37274 35612 37280 35624
rect 37235 35584 37280 35612
rect 37274 35572 37280 35584
rect 37332 35572 37338 35624
rect 37918 35612 37924 35624
rect 37879 35584 37924 35612
rect 37918 35572 37924 35584
rect 37976 35572 37982 35624
rect 33152 35516 33364 35544
rect 33597 35547 33655 35553
rect 28997 35507 29055 35513
rect 33597 35513 33609 35547
rect 33643 35513 33655 35547
rect 34422 35544 34428 35556
rect 34383 35516 34428 35544
rect 33597 35507 33655 35513
rect 29012 35476 29040 35507
rect 33410 35476 33416 35488
rect 29012 35448 33416 35476
rect 33410 35436 33416 35448
rect 33468 35436 33474 35488
rect 33502 35436 33508 35488
rect 33560 35476 33566 35488
rect 33612 35476 33640 35507
rect 34422 35504 34428 35516
rect 34480 35504 34486 35556
rect 33686 35476 33692 35488
rect 33560 35448 33692 35476
rect 33560 35436 33566 35448
rect 33686 35436 33692 35448
rect 33744 35436 33750 35488
rect 33870 35476 33876 35488
rect 33831 35448 33876 35476
rect 33870 35436 33876 35448
rect 33928 35436 33934 35488
rect 34330 35436 34336 35488
rect 34388 35476 34394 35488
rect 34517 35479 34575 35485
rect 34517 35476 34529 35479
rect 34388 35448 34529 35476
rect 34388 35436 34394 35448
rect 34517 35445 34529 35448
rect 34563 35445 34575 35479
rect 34517 35439 34575 35445
rect 1104 35386 38824 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 38824 35386
rect 1104 35312 38824 35334
rect 33594 35232 33600 35284
rect 33652 35232 33658 35284
rect 33413 35207 33471 35213
rect 33413 35173 33425 35207
rect 33459 35204 33471 35207
rect 33612 35204 33640 35232
rect 33459 35176 33640 35204
rect 33459 35173 33471 35176
rect 33413 35167 33471 35173
rect 33778 35164 33784 35216
rect 33836 35204 33842 35216
rect 34333 35207 34391 35213
rect 34333 35204 34345 35207
rect 33836 35176 34345 35204
rect 33836 35164 33842 35176
rect 34333 35173 34345 35176
rect 34379 35204 34391 35207
rect 34422 35204 34428 35216
rect 34379 35176 34428 35204
rect 34379 35173 34391 35176
rect 34333 35167 34391 35173
rect 34422 35164 34428 35176
rect 34480 35164 34486 35216
rect 33134 35136 33140 35148
rect 33095 35108 33140 35136
rect 33134 35096 33140 35108
rect 33192 35096 33198 35148
rect 33230 35139 33288 35145
rect 33230 35105 33242 35139
rect 33276 35105 33288 35139
rect 33502 35136 33508 35148
rect 33463 35108 33508 35136
rect 33230 35099 33288 35105
rect 33244 35068 33272 35099
rect 33502 35096 33508 35108
rect 33560 35096 33566 35148
rect 33643 35139 33701 35145
rect 33643 35105 33655 35139
rect 33689 35136 33701 35139
rect 33689 35108 34284 35136
rect 33689 35105 33701 35108
rect 33643 35099 33701 35105
rect 32968 35040 33272 35068
rect 2682 34892 2688 34944
rect 2740 34932 2746 34944
rect 32968 34941 32996 35040
rect 33870 35028 33876 35080
rect 33928 35028 33934 35080
rect 34256 35068 34284 35108
rect 37090 35068 37096 35080
rect 34256 35040 37096 35068
rect 37090 35028 37096 35040
rect 37148 35028 37154 35080
rect 33686 34960 33692 35012
rect 33744 35000 33750 35012
rect 33888 35000 33916 35028
rect 33744 34972 33916 35000
rect 33744 34960 33750 34972
rect 32953 34935 33011 34941
rect 32953 34932 32965 34935
rect 2740 34904 32965 34932
rect 2740 34892 2746 34904
rect 32953 34901 32965 34904
rect 32999 34901 33011 34935
rect 32953 34895 33011 34901
rect 33781 34935 33839 34941
rect 33781 34901 33793 34935
rect 33827 34932 33839 34935
rect 33870 34932 33876 34944
rect 33827 34904 33876 34932
rect 33827 34901 33839 34904
rect 33781 34895 33839 34901
rect 33870 34892 33876 34904
rect 33928 34892 33934 34944
rect 34422 34932 34428 34944
rect 34383 34904 34428 34932
rect 34422 34892 34428 34904
rect 34480 34892 34486 34944
rect 1104 34842 38824 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 38824 34842
rect 1104 34768 38824 34790
rect 33962 34688 33968 34740
rect 34020 34728 34026 34740
rect 37277 34731 37335 34737
rect 37277 34728 37289 34731
rect 34020 34700 37289 34728
rect 34020 34688 34026 34700
rect 37277 34697 37289 34700
rect 37323 34697 37335 34731
rect 37277 34691 37335 34697
rect 2041 34527 2099 34533
rect 2041 34493 2053 34527
rect 2087 34524 2099 34527
rect 2590 34524 2596 34536
rect 2087 34496 2596 34524
rect 2087 34493 2099 34496
rect 2041 34487 2099 34493
rect 2590 34484 2596 34496
rect 2648 34484 2654 34536
rect 37458 34524 37464 34536
rect 37419 34496 37464 34524
rect 37458 34484 37464 34496
rect 37516 34484 37522 34536
rect 37918 34524 37924 34536
rect 37879 34496 37924 34524
rect 37918 34484 37924 34496
rect 37976 34484 37982 34536
rect 1854 34456 1860 34468
rect 1815 34428 1860 34456
rect 1854 34416 1860 34428
rect 1912 34416 1918 34468
rect 1104 34298 38824 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 38824 34298
rect 1104 34224 38824 34246
rect 1854 34048 1860 34060
rect 1815 34020 1860 34048
rect 1854 34008 1860 34020
rect 1912 34008 1918 34060
rect 2041 33915 2099 33921
rect 2041 33881 2053 33915
rect 2087 33912 2099 33915
rect 2682 33912 2688 33924
rect 2087 33884 2688 33912
rect 2087 33881 2099 33884
rect 2041 33875 2099 33881
rect 2682 33872 2688 33884
rect 2740 33872 2746 33924
rect 35802 33804 35808 33856
rect 35860 33844 35866 33856
rect 36538 33844 36544 33856
rect 35860 33816 36544 33844
rect 35860 33804 35866 33816
rect 36538 33804 36544 33816
rect 36596 33804 36602 33856
rect 1104 33754 38824 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 38824 33754
rect 1104 33680 38824 33702
rect 36170 33600 36176 33652
rect 36228 33640 36234 33652
rect 37277 33643 37335 33649
rect 37277 33640 37289 33643
rect 36228 33612 37289 33640
rect 36228 33600 36234 33612
rect 37277 33609 37289 33612
rect 37323 33609 37335 33643
rect 37277 33603 37335 33609
rect 36170 33464 36176 33516
rect 36228 33504 36234 33516
rect 36354 33504 36360 33516
rect 36228 33476 36360 33504
rect 36228 33464 36234 33476
rect 36354 33464 36360 33476
rect 36412 33464 36418 33516
rect 28718 33436 28724 33448
rect 28679 33408 28724 33436
rect 28718 33396 28724 33408
rect 28776 33396 28782 33448
rect 33689 33439 33747 33445
rect 33689 33405 33701 33439
rect 33735 33436 33747 33439
rect 33778 33436 33784 33448
rect 33735 33408 33784 33436
rect 33735 33405 33747 33408
rect 33689 33399 33747 33405
rect 33778 33396 33784 33408
rect 33836 33396 33842 33448
rect 37458 33436 37464 33448
rect 37419 33408 37464 33436
rect 37458 33396 37464 33408
rect 37516 33396 37522 33448
rect 37918 33436 37924 33448
rect 37879 33408 37924 33436
rect 37918 33396 37924 33408
rect 37976 33396 37982 33448
rect 28905 33371 28963 33377
rect 28905 33337 28917 33371
rect 28951 33368 28963 33371
rect 33134 33368 33140 33380
rect 28951 33340 33140 33368
rect 28951 33337 28963 33340
rect 28905 33331 28963 33337
rect 33134 33328 33140 33340
rect 33192 33328 33198 33380
rect 32858 33260 32864 33312
rect 32916 33300 32922 33312
rect 33781 33303 33839 33309
rect 33781 33300 33793 33303
rect 32916 33272 33793 33300
rect 32916 33260 32922 33272
rect 33781 33269 33793 33272
rect 33827 33269 33839 33303
rect 33781 33263 33839 33269
rect 1104 33210 38824 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 38824 33210
rect 1104 33136 38824 33158
rect 1854 33028 1860 33040
rect 1815 33000 1860 33028
rect 1854 32988 1860 33000
rect 1912 32988 1918 33040
rect 32398 32988 32404 33040
rect 32456 33028 32462 33040
rect 36814 33028 36820 33040
rect 32456 33000 36820 33028
rect 32456 32988 32462 33000
rect 36814 32988 36820 33000
rect 36872 32988 36878 33040
rect 34698 32920 34704 32972
rect 34756 32960 34762 32972
rect 35802 32960 35808 32972
rect 34756 32932 35808 32960
rect 34756 32920 34762 32932
rect 35802 32920 35808 32932
rect 35860 32920 35866 32972
rect 37182 32960 37188 32972
rect 37143 32932 37188 32960
rect 37182 32920 37188 32932
rect 37240 32920 37246 32972
rect 1946 32756 1952 32768
rect 1907 32728 1952 32756
rect 1946 32716 1952 32728
rect 2004 32716 2010 32768
rect 1104 32666 38824 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 38824 32666
rect 1104 32592 38824 32614
rect 2406 32512 2412 32564
rect 2464 32552 2470 32564
rect 32861 32555 32919 32561
rect 32861 32552 32873 32555
rect 2464 32524 32873 32552
rect 2464 32512 2470 32524
rect 32861 32521 32873 32524
rect 32907 32521 32919 32555
rect 32861 32515 32919 32521
rect 32876 32416 32904 32515
rect 34422 32416 34428 32428
rect 32876 32388 33180 32416
rect 33152 32357 33180 32388
rect 33336 32388 34428 32416
rect 33336 32360 33364 32388
rect 34422 32376 34428 32388
rect 34480 32376 34486 32428
rect 33045 32351 33103 32357
rect 33045 32317 33057 32351
rect 33091 32317 33103 32351
rect 33045 32311 33103 32317
rect 33138 32351 33196 32357
rect 33138 32317 33150 32351
rect 33184 32317 33196 32351
rect 33318 32348 33324 32360
rect 33231 32320 33324 32348
rect 33138 32311 33196 32317
rect 1854 32280 1860 32292
rect 1815 32252 1860 32280
rect 1854 32240 1860 32252
rect 1912 32240 1918 32292
rect 2041 32283 2099 32289
rect 2041 32249 2053 32283
rect 2087 32280 2099 32283
rect 2406 32280 2412 32292
rect 2087 32252 2412 32280
rect 2087 32249 2099 32252
rect 2041 32243 2099 32249
rect 2406 32240 2412 32252
rect 2464 32240 2470 32292
rect 33060 32280 33088 32311
rect 33318 32308 33324 32320
rect 33376 32308 33382 32360
rect 33410 32308 33416 32360
rect 33468 32348 33474 32360
rect 33551 32351 33609 32357
rect 33468 32320 33513 32348
rect 33468 32308 33474 32320
rect 33551 32317 33563 32351
rect 33597 32348 33609 32351
rect 37182 32348 37188 32360
rect 33597 32320 37188 32348
rect 33597 32317 33609 32320
rect 33551 32311 33609 32317
rect 37182 32308 37188 32320
rect 37240 32308 37246 32360
rect 37918 32348 37924 32360
rect 37879 32320 37924 32348
rect 37918 32308 37924 32320
rect 37976 32308 37982 32360
rect 38746 32280 38752 32292
rect 33060 32252 38752 32280
rect 38746 32240 38752 32252
rect 38804 32240 38810 32292
rect 33689 32215 33747 32221
rect 33689 32181 33701 32215
rect 33735 32212 33747 32215
rect 35342 32212 35348 32224
rect 33735 32184 35348 32212
rect 33735 32181 33747 32184
rect 33689 32175 33747 32181
rect 35342 32172 35348 32184
rect 35400 32172 35406 32224
rect 1104 32122 38824 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 38824 32122
rect 1104 32048 38824 32070
rect 33689 32011 33747 32017
rect 33689 31977 33701 32011
rect 33735 32008 33747 32011
rect 33962 32008 33968 32020
rect 33735 31980 33968 32008
rect 33735 31977 33747 31980
rect 33689 31971 33747 31977
rect 33962 31968 33968 31980
rect 34020 31968 34026 32020
rect 37090 31968 37096 32020
rect 37148 32008 37154 32020
rect 37185 32011 37243 32017
rect 37185 32008 37197 32011
rect 37148 31980 37197 32008
rect 37148 31968 37154 31980
rect 37185 31977 37197 31980
rect 37231 31977 37243 32011
rect 37185 31971 37243 31977
rect 33318 31940 33324 31952
rect 33279 31912 33324 31940
rect 33318 31900 33324 31912
rect 33376 31900 33382 31952
rect 33410 31900 33416 31952
rect 33468 31940 33474 31952
rect 33468 31912 33513 31940
rect 33468 31900 33474 31912
rect 33042 31872 33048 31884
rect 33003 31844 33048 31872
rect 33042 31832 33048 31844
rect 33100 31832 33106 31884
rect 33138 31875 33196 31881
rect 33138 31841 33150 31875
rect 33184 31841 33196 31875
rect 33138 31835 33196 31841
rect 33551 31875 33609 31881
rect 33551 31841 33563 31875
rect 33597 31872 33609 31875
rect 36814 31872 36820 31884
rect 33597 31844 36820 31872
rect 33597 31841 33609 31844
rect 33551 31835 33609 31841
rect 2590 31764 2596 31816
rect 2648 31804 2654 31816
rect 32861 31807 32919 31813
rect 32861 31804 32873 31807
rect 2648 31776 32873 31804
rect 2648 31764 2654 31776
rect 32861 31773 32873 31776
rect 32907 31804 32919 31807
rect 33152 31804 33180 31835
rect 36814 31832 36820 31844
rect 36872 31832 36878 31884
rect 37366 31872 37372 31884
rect 37327 31844 37372 31872
rect 37366 31832 37372 31844
rect 37424 31832 37430 31884
rect 32907 31776 33180 31804
rect 32907 31773 32919 31776
rect 32861 31767 32919 31773
rect 36630 31764 36636 31816
rect 36688 31804 36694 31816
rect 37090 31804 37096 31816
rect 36688 31776 37096 31804
rect 36688 31764 36694 31776
rect 37090 31764 37096 31776
rect 37148 31764 37154 31816
rect 35526 31696 35532 31748
rect 35584 31736 35590 31748
rect 35584 31708 36400 31736
rect 35584 31696 35590 31708
rect 36372 31680 36400 31708
rect 36354 31628 36360 31680
rect 36412 31628 36418 31680
rect 1104 31578 38824 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 38824 31578
rect 1104 31504 38824 31526
rect 33318 31424 33324 31476
rect 33376 31464 33382 31476
rect 33502 31464 33508 31476
rect 33376 31436 33508 31464
rect 33376 31424 33382 31436
rect 33502 31424 33508 31436
rect 33560 31424 33566 31476
rect 33686 31424 33692 31476
rect 33744 31464 33750 31476
rect 35526 31464 35532 31476
rect 33744 31436 35532 31464
rect 33744 31424 33750 31436
rect 35526 31424 35532 31436
rect 35584 31424 35590 31476
rect 37734 31464 37740 31476
rect 36648 31436 37740 31464
rect 36648 31396 36676 31436
rect 37734 31424 37740 31436
rect 37792 31424 37798 31476
rect 32968 31368 36676 31396
rect 1854 31260 1860 31272
rect 1815 31232 1860 31260
rect 1854 31220 1860 31232
rect 1912 31220 1918 31272
rect 2682 31220 2688 31272
rect 2740 31260 2746 31272
rect 32968 31269 32996 31368
rect 36722 31356 36728 31408
rect 36780 31396 36786 31408
rect 36906 31396 36912 31408
rect 36780 31368 36912 31396
rect 36780 31356 36786 31368
rect 36906 31356 36912 31368
rect 36964 31356 36970 31408
rect 32769 31263 32827 31269
rect 32769 31260 32781 31263
rect 2740 31232 32781 31260
rect 2740 31220 2746 31232
rect 32769 31229 32781 31232
rect 32815 31229 32827 31263
rect 32769 31223 32827 31229
rect 32953 31263 33011 31269
rect 32953 31229 32965 31263
rect 32999 31229 33011 31263
rect 32953 31223 33011 31229
rect 33046 31263 33104 31269
rect 33046 31229 33058 31263
rect 33092 31229 33104 31263
rect 33318 31260 33324 31272
rect 33279 31232 33324 31260
rect 33046 31223 33104 31229
rect 2041 31195 2099 31201
rect 2041 31161 2053 31195
rect 2087 31192 2099 31195
rect 2590 31192 2596 31204
rect 2087 31164 2596 31192
rect 2087 31161 2099 31164
rect 2041 31155 2099 31161
rect 2590 31152 2596 31164
rect 2648 31152 2654 31204
rect 32784 31192 32812 31223
rect 33060 31192 33088 31223
rect 33318 31220 33324 31232
rect 33376 31220 33382 31272
rect 33459 31263 33517 31269
rect 33459 31229 33471 31263
rect 33505 31260 33517 31263
rect 36906 31260 36912 31272
rect 33505 31232 36912 31260
rect 33505 31229 33517 31232
rect 33459 31223 33517 31229
rect 36906 31220 36912 31232
rect 36964 31220 36970 31272
rect 37274 31260 37280 31272
rect 37235 31232 37280 31260
rect 37274 31220 37280 31232
rect 37332 31220 37338 31272
rect 37918 31260 37924 31272
rect 37879 31232 37924 31260
rect 37918 31220 37924 31232
rect 37976 31220 37982 31272
rect 32784 31164 33088 31192
rect 33229 31195 33287 31201
rect 33229 31161 33241 31195
rect 33275 31161 33287 31195
rect 33229 31155 33287 31161
rect 33244 31124 33272 31155
rect 33318 31124 33324 31136
rect 33231 31096 33324 31124
rect 33318 31084 33324 31096
rect 33376 31124 33382 31136
rect 33502 31124 33508 31136
rect 33376 31096 33508 31124
rect 33376 31084 33382 31096
rect 33502 31084 33508 31096
rect 33560 31084 33566 31136
rect 33597 31127 33655 31133
rect 33597 31093 33609 31127
rect 33643 31124 33655 31127
rect 33778 31124 33784 31136
rect 33643 31096 33784 31124
rect 33643 31093 33655 31096
rect 33597 31087 33655 31093
rect 33778 31084 33784 31096
rect 33836 31084 33842 31136
rect 34054 31084 34060 31136
rect 34112 31124 34118 31136
rect 34606 31124 34612 31136
rect 34112 31096 34612 31124
rect 34112 31084 34118 31096
rect 34606 31084 34612 31096
rect 34664 31084 34670 31136
rect 1104 31034 38824 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 38824 31034
rect 1104 30960 38824 30982
rect 37182 30920 37188 30932
rect 37143 30892 37188 30920
rect 37182 30880 37188 30892
rect 37240 30880 37246 30932
rect 33410 30852 33416 30864
rect 33371 30824 33416 30852
rect 33410 30812 33416 30824
rect 33468 30812 33474 30864
rect 1854 30784 1860 30796
rect 1815 30756 1860 30784
rect 1854 30744 1860 30756
rect 1912 30744 1918 30796
rect 32950 30744 32956 30796
rect 33008 30784 33014 30796
rect 33045 30787 33103 30793
rect 33045 30784 33057 30787
rect 33008 30756 33057 30784
rect 33008 30744 33014 30756
rect 33045 30753 33057 30756
rect 33091 30753 33103 30787
rect 33045 30747 33103 30753
rect 33138 30787 33196 30793
rect 33138 30753 33150 30787
rect 33184 30753 33196 30787
rect 33318 30784 33324 30796
rect 33279 30756 33324 30784
rect 33138 30747 33196 30753
rect 1946 30676 1952 30728
rect 2004 30716 2010 30728
rect 33153 30716 33181 30747
rect 33318 30744 33324 30756
rect 33376 30744 33382 30796
rect 33551 30787 33609 30793
rect 33551 30753 33563 30787
rect 33597 30784 33609 30787
rect 36630 30784 36636 30796
rect 33597 30756 36636 30784
rect 33597 30753 33609 30756
rect 33551 30747 33609 30753
rect 36630 30744 36636 30756
rect 36688 30744 36694 30796
rect 37366 30784 37372 30796
rect 37327 30756 37372 30784
rect 37366 30744 37372 30756
rect 37424 30744 37430 30796
rect 2004 30688 6914 30716
rect 2004 30676 2010 30688
rect 1946 30580 1952 30592
rect 1907 30552 1952 30580
rect 1946 30540 1952 30552
rect 2004 30540 2010 30592
rect 6886 30580 6914 30688
rect 32876 30688 33181 30716
rect 32876 30589 32904 30688
rect 32861 30583 32919 30589
rect 32861 30580 32873 30583
rect 6886 30552 32873 30580
rect 32861 30549 32873 30552
rect 32907 30549 32919 30583
rect 32861 30543 32919 30549
rect 33689 30583 33747 30589
rect 33689 30549 33701 30583
rect 33735 30580 33747 30583
rect 34422 30580 34428 30592
rect 33735 30552 34428 30580
rect 33735 30549 33747 30552
rect 33689 30543 33747 30549
rect 34422 30540 34428 30552
rect 34480 30540 34486 30592
rect 1104 30490 38824 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 38824 30490
rect 1104 30416 38824 30438
rect 1946 30336 1952 30388
rect 2004 30376 2010 30388
rect 27522 30376 27528 30388
rect 2004 30348 27528 30376
rect 2004 30336 2010 30348
rect 27522 30336 27528 30348
rect 27580 30336 27586 30388
rect 33318 30308 33324 30320
rect 33153 30280 33324 30308
rect 32490 30132 32496 30184
rect 32548 30172 32554 30184
rect 33153 30181 33181 30280
rect 33318 30268 33324 30280
rect 33376 30268 33382 30320
rect 33410 30268 33416 30320
rect 33468 30268 33474 30320
rect 33428 30240 33456 30268
rect 33244 30212 33456 30240
rect 33244 30181 33272 30212
rect 32861 30175 32919 30181
rect 32861 30172 32873 30175
rect 32548 30144 32873 30172
rect 32548 30132 32554 30144
rect 32861 30141 32873 30144
rect 32907 30141 32919 30175
rect 32861 30135 32919 30141
rect 32954 30175 33012 30181
rect 32954 30141 32966 30175
rect 33000 30141 33012 30175
rect 32954 30135 33012 30141
rect 33137 30175 33195 30181
rect 33137 30141 33149 30175
rect 33183 30141 33195 30175
rect 33137 30135 33195 30141
rect 33229 30175 33287 30181
rect 33229 30141 33241 30175
rect 33275 30141 33287 30175
rect 33229 30135 33287 30141
rect 33367 30175 33425 30181
rect 33367 30141 33379 30175
rect 33413 30172 33425 30175
rect 37274 30172 37280 30184
rect 33413 30144 37136 30172
rect 37235 30144 37280 30172
rect 33413 30141 33425 30144
rect 33367 30135 33425 30141
rect 32968 30104 32996 30135
rect 32692 30076 32996 30104
rect 2406 29996 2412 30048
rect 2464 30036 2470 30048
rect 32692 30045 32720 30076
rect 32677 30039 32735 30045
rect 32677 30036 32689 30039
rect 2464 30008 32689 30036
rect 2464 29996 2470 30008
rect 32677 30005 32689 30008
rect 32723 30005 32735 30039
rect 32677 29999 32735 30005
rect 33505 30039 33563 30045
rect 33505 30005 33517 30039
rect 33551 30036 33563 30039
rect 33870 30036 33876 30048
rect 33551 30008 33876 30036
rect 33551 30005 33563 30008
rect 33505 29999 33563 30005
rect 33870 29996 33876 30008
rect 33928 29996 33934 30048
rect 37108 30036 37136 30144
rect 37274 30132 37280 30144
rect 37332 30132 37338 30184
rect 37918 30172 37924 30184
rect 37879 30144 37924 30172
rect 37918 30132 37924 30144
rect 37976 30132 37982 30184
rect 37274 30036 37280 30048
rect 37108 30008 37280 30036
rect 37274 29996 37280 30008
rect 37332 29996 37338 30048
rect 1104 29946 38824 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 38824 29946
rect 1104 29872 38824 29894
rect 1854 29764 1860 29776
rect 1815 29736 1860 29764
rect 1854 29724 1860 29736
rect 1912 29724 1918 29776
rect 2041 29563 2099 29569
rect 2041 29529 2053 29563
rect 2087 29560 2099 29563
rect 2682 29560 2688 29572
rect 2087 29532 2688 29560
rect 2087 29529 2099 29532
rect 2041 29523 2099 29529
rect 2682 29520 2688 29532
rect 2740 29520 2746 29572
rect 1104 29402 38824 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 38824 29402
rect 1104 29328 38824 29350
rect 36814 29248 36820 29300
rect 36872 29288 36878 29300
rect 37277 29291 37335 29297
rect 37277 29288 37289 29291
rect 36872 29260 37289 29288
rect 36872 29248 36878 29260
rect 37277 29257 37289 29260
rect 37323 29257 37335 29291
rect 37277 29251 37335 29257
rect 34422 29180 34428 29232
rect 34480 29220 34486 29232
rect 34882 29220 34888 29232
rect 34480 29192 34888 29220
rect 34480 29180 34486 29192
rect 34882 29180 34888 29192
rect 34940 29180 34946 29232
rect 1854 29084 1860 29096
rect 1815 29056 1860 29084
rect 1854 29044 1860 29056
rect 1912 29044 1918 29096
rect 37458 29084 37464 29096
rect 37419 29056 37464 29084
rect 37458 29044 37464 29056
rect 37516 29044 37522 29096
rect 37918 29084 37924 29096
rect 37879 29056 37924 29084
rect 37918 29044 37924 29056
rect 37976 29044 37982 29096
rect 2041 29019 2099 29025
rect 2041 28985 2053 29019
rect 2087 29016 2099 29019
rect 4062 29016 4068 29028
rect 2087 28988 4068 29016
rect 2087 28985 2099 28988
rect 2041 28979 2099 28985
rect 4062 28976 4068 28988
rect 4120 28976 4126 29028
rect 36354 28976 36360 29028
rect 36412 29016 36418 29028
rect 36814 29016 36820 29028
rect 36412 28988 36820 29016
rect 36412 28976 36418 28988
rect 36814 28976 36820 28988
rect 36872 28976 36878 29028
rect 1104 28858 38824 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 38824 28858
rect 1104 28784 38824 28806
rect 32490 28704 32496 28756
rect 32548 28744 32554 28756
rect 37826 28744 37832 28756
rect 32548 28716 37832 28744
rect 32548 28704 32554 28716
rect 37826 28704 37832 28716
rect 37884 28704 37890 28756
rect 34882 28432 34888 28484
rect 34940 28472 34946 28484
rect 38470 28472 38476 28484
rect 34940 28444 38476 28472
rect 34940 28432 34946 28444
rect 38470 28432 38476 28444
rect 38528 28432 38534 28484
rect 33042 28364 33048 28416
rect 33100 28404 33106 28416
rect 38378 28404 38384 28416
rect 33100 28376 38384 28404
rect 33100 28364 33106 28376
rect 38378 28364 38384 28376
rect 38436 28364 38442 28416
rect 1104 28314 38824 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 38824 28314
rect 1104 28240 38824 28262
rect 36906 28160 36912 28212
rect 36964 28200 36970 28212
rect 37277 28203 37335 28209
rect 37277 28200 37289 28203
rect 36964 28172 37289 28200
rect 36964 28160 36970 28172
rect 37277 28169 37289 28172
rect 37323 28169 37335 28203
rect 37277 28163 37335 28169
rect 2590 28024 2596 28076
rect 2648 28064 2654 28076
rect 32585 28067 32643 28073
rect 32585 28064 32597 28067
rect 2648 28036 32597 28064
rect 2648 28024 2654 28036
rect 32585 28033 32597 28036
rect 32631 28064 32643 28067
rect 32631 28036 32904 28064
rect 32631 28033 32643 28036
rect 32585 28027 32643 28033
rect 1854 27996 1860 28008
rect 1815 27968 1860 27996
rect 1854 27956 1860 27968
rect 1912 27956 1918 28008
rect 26789 27999 26847 28005
rect 26789 27965 26801 27999
rect 26835 27965 26847 27999
rect 26789 27959 26847 27965
rect 26881 27999 26939 28005
rect 26881 27965 26893 27999
rect 26927 27996 26939 27999
rect 26970 27996 26976 28008
rect 26927 27968 26976 27996
rect 26927 27965 26939 27968
rect 26881 27959 26939 27965
rect 2041 27931 2099 27937
rect 2041 27897 2053 27931
rect 2087 27928 2099 27931
rect 2406 27928 2412 27940
rect 2087 27900 2412 27928
rect 2087 27897 2099 27900
rect 2041 27891 2099 27897
rect 2406 27888 2412 27900
rect 2464 27888 2470 27940
rect 26804 27860 26832 27959
rect 26970 27956 26976 27968
rect 27028 27956 27034 28008
rect 27065 27999 27123 28005
rect 27065 27965 27077 27999
rect 27111 27996 27123 27999
rect 27154 27996 27160 28008
rect 27111 27968 27160 27996
rect 27111 27965 27123 27968
rect 27065 27959 27123 27965
rect 27154 27956 27160 27968
rect 27212 27956 27218 28008
rect 27525 27999 27583 28005
rect 27525 27965 27537 27999
rect 27571 27996 27583 27999
rect 27798 27996 27804 28008
rect 27571 27968 27804 27996
rect 27571 27965 27583 27968
rect 27525 27959 27583 27965
rect 27798 27956 27804 27968
rect 27856 27996 27862 28008
rect 28534 27996 28540 28008
rect 27856 27968 28540 27996
rect 27856 27956 27862 27968
rect 28534 27956 28540 27968
rect 28592 27956 28598 28008
rect 32876 28005 32904 28036
rect 32769 27999 32827 28005
rect 32769 27965 32781 27999
rect 32815 27965 32827 27999
rect 32769 27959 32827 27965
rect 32862 27999 32920 28005
rect 32862 27965 32874 27999
rect 32908 27965 32920 27999
rect 33134 27996 33140 28008
rect 33095 27968 33140 27996
rect 32862 27959 32920 27965
rect 26878 27860 26884 27872
rect 26804 27832 26884 27860
rect 26878 27820 26884 27832
rect 26936 27820 26942 27872
rect 32784 27860 32812 27959
rect 33134 27956 33140 27968
rect 33192 27956 33198 28008
rect 33275 27999 33333 28005
rect 33275 27965 33287 27999
rect 33321 27996 33333 27999
rect 36906 27996 36912 28008
rect 33321 27968 36912 27996
rect 33321 27965 33333 27968
rect 33275 27959 33333 27965
rect 36906 27956 36912 27968
rect 36964 27956 36970 28008
rect 37458 27996 37464 28008
rect 37419 27968 37464 27996
rect 37458 27956 37464 27968
rect 37516 27956 37522 28008
rect 37921 27999 37979 28005
rect 37921 27965 37933 27999
rect 37967 27996 37979 27999
rect 38010 27996 38016 28008
rect 37967 27968 38016 27996
rect 37967 27965 37979 27968
rect 37921 27959 37979 27965
rect 38010 27956 38016 27968
rect 38068 27956 38074 28008
rect 32950 27888 32956 27940
rect 33008 27928 33014 27940
rect 33045 27931 33103 27937
rect 33045 27928 33057 27931
rect 33008 27900 33057 27928
rect 33008 27888 33014 27900
rect 33045 27897 33057 27900
rect 33091 27897 33103 27931
rect 38930 27928 38936 27940
rect 33045 27891 33103 27897
rect 33336 27900 38936 27928
rect 33336 27860 33364 27900
rect 38930 27888 38936 27900
rect 38988 27888 38994 27940
rect 32784 27832 33364 27860
rect 33413 27863 33471 27869
rect 33413 27829 33425 27863
rect 33459 27860 33471 27863
rect 33502 27860 33508 27872
rect 33459 27832 33508 27860
rect 33459 27829 33471 27832
rect 33413 27823 33471 27829
rect 33502 27820 33508 27832
rect 33560 27820 33566 27872
rect 33594 27820 33600 27872
rect 33652 27860 33658 27872
rect 34146 27860 34152 27872
rect 33652 27832 34152 27860
rect 33652 27820 33658 27832
rect 34146 27820 34152 27832
rect 34204 27820 34210 27872
rect 1104 27770 38824 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 38824 27770
rect 1104 27696 38824 27718
rect 33134 27616 33140 27668
rect 33192 27656 33198 27668
rect 33192 27628 33456 27656
rect 33192 27616 33198 27628
rect 27801 27591 27859 27597
rect 27801 27557 27813 27591
rect 27847 27557 27859 27591
rect 27801 27551 27859 27557
rect 1854 27520 1860 27532
rect 1815 27492 1860 27520
rect 1854 27480 1860 27492
rect 1912 27480 1918 27532
rect 27816 27520 27844 27551
rect 27982 27548 27988 27600
rect 28040 27597 28046 27600
rect 28040 27591 28064 27597
rect 28052 27557 28064 27591
rect 28040 27551 28064 27557
rect 28040 27548 28046 27551
rect 32950 27548 32956 27600
rect 33008 27588 33014 27600
rect 33428 27597 33456 27628
rect 33594 27616 33600 27668
rect 33652 27656 33658 27668
rect 33689 27659 33747 27665
rect 33689 27656 33701 27659
rect 33652 27628 33701 27656
rect 33652 27616 33658 27628
rect 33689 27625 33701 27628
rect 33735 27625 33747 27659
rect 33689 27619 33747 27625
rect 33321 27591 33379 27597
rect 33321 27588 33333 27591
rect 33008 27560 33333 27588
rect 33008 27548 33014 27560
rect 33321 27557 33333 27560
rect 33367 27557 33379 27591
rect 33321 27551 33379 27557
rect 33413 27591 33471 27597
rect 33413 27557 33425 27591
rect 33459 27557 33471 27591
rect 33413 27551 33471 27557
rect 35618 27548 35624 27600
rect 35676 27588 35682 27600
rect 36354 27588 36360 27600
rect 35676 27560 36360 27588
rect 35676 27548 35682 27560
rect 36354 27548 36360 27560
rect 36412 27548 36418 27600
rect 37458 27588 37464 27600
rect 36740 27560 37464 27588
rect 28534 27520 28540 27532
rect 27816 27492 28540 27520
rect 28534 27480 28540 27492
rect 28592 27480 28598 27532
rect 33042 27520 33048 27532
rect 33003 27492 33048 27520
rect 33042 27480 33048 27492
rect 33100 27480 33106 27532
rect 33138 27523 33196 27529
rect 33138 27489 33150 27523
rect 33184 27489 33196 27523
rect 33138 27483 33196 27489
rect 33551 27523 33609 27529
rect 33551 27489 33563 27523
rect 33597 27520 33609 27523
rect 36740 27520 36768 27560
rect 37458 27548 37464 27560
rect 37516 27548 37522 27600
rect 37182 27520 37188 27532
rect 33597 27492 36768 27520
rect 37143 27492 37188 27520
rect 33597 27489 33609 27492
rect 33551 27483 33609 27489
rect 27522 27412 27528 27464
rect 27580 27452 27586 27464
rect 32861 27455 32919 27461
rect 32861 27452 32873 27455
rect 27580 27424 32873 27452
rect 27580 27412 27586 27424
rect 32861 27421 32873 27424
rect 32907 27452 32919 27455
rect 33153 27452 33181 27483
rect 37182 27480 37188 27492
rect 37240 27480 37246 27532
rect 32907 27424 33181 27452
rect 32907 27421 32919 27424
rect 32861 27415 32919 27421
rect 34238 27412 34244 27464
rect 34296 27452 34302 27464
rect 34422 27452 34428 27464
rect 34296 27424 34428 27452
rect 34296 27412 34302 27424
rect 34422 27412 34428 27424
rect 34480 27412 34486 27464
rect 6886 27356 30236 27384
rect 1949 27319 2007 27325
rect 1949 27285 1961 27319
rect 1995 27316 2007 27319
rect 6886 27316 6914 27356
rect 1995 27288 6914 27316
rect 1995 27285 2007 27288
rect 1949 27279 2007 27285
rect 27798 27276 27804 27328
rect 27856 27316 27862 27328
rect 27985 27319 28043 27325
rect 27985 27316 27997 27319
rect 27856 27288 27997 27316
rect 27856 27276 27862 27288
rect 27985 27285 27997 27288
rect 28031 27285 28043 27319
rect 27985 27279 28043 27285
rect 28074 27276 28080 27328
rect 28132 27316 28138 27328
rect 28169 27319 28227 27325
rect 28169 27316 28181 27319
rect 28132 27288 28181 27316
rect 28132 27276 28138 27288
rect 28169 27285 28181 27288
rect 28215 27285 28227 27319
rect 30208 27316 30236 27356
rect 34238 27316 34244 27328
rect 30208 27288 34244 27316
rect 28169 27279 28227 27285
rect 34238 27276 34244 27288
rect 34296 27276 34302 27328
rect 1104 27226 38824 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 38824 27226
rect 1104 27152 38824 27174
rect 26789 27115 26847 27121
rect 26789 27081 26801 27115
rect 26835 27112 26847 27115
rect 27982 27112 27988 27124
rect 26835 27084 27988 27112
rect 26835 27081 26847 27084
rect 26789 27075 26847 27081
rect 27982 27072 27988 27084
rect 28040 27072 28046 27124
rect 31846 27112 31852 27124
rect 30484 27084 31432 27112
rect 31807 27084 31852 27112
rect 30484 27044 30512 27084
rect 6886 27016 30512 27044
rect 31404 27044 31432 27084
rect 31846 27072 31852 27084
rect 31904 27072 31910 27124
rect 32585 27047 32643 27053
rect 32585 27044 32597 27047
rect 31404 27016 32597 27044
rect 2682 26936 2688 26988
rect 2740 26976 2746 26988
rect 6886 26976 6914 27016
rect 32585 27013 32597 27016
rect 32631 27013 32643 27047
rect 32585 27007 32643 27013
rect 2740 26948 6914 26976
rect 25317 26979 25375 26985
rect 2740 26936 2746 26948
rect 25317 26945 25329 26979
rect 25363 26976 25375 26979
rect 26878 26976 26884 26988
rect 25363 26948 26884 26976
rect 25363 26945 25375 26948
rect 25317 26939 25375 26945
rect 26878 26936 26884 26948
rect 26936 26936 26942 26988
rect 29914 26936 29920 26988
rect 29972 26976 29978 26988
rect 30745 26979 30803 26985
rect 30745 26976 30757 26979
rect 29972 26948 30757 26976
rect 29972 26936 29978 26948
rect 30745 26945 30757 26948
rect 30791 26945 30803 26979
rect 32600 26976 32628 27007
rect 36906 27004 36912 27056
rect 36964 27044 36970 27056
rect 37182 27044 37188 27056
rect 36964 27016 37188 27044
rect 36964 27004 36970 27016
rect 37182 27004 37188 27016
rect 37240 27004 37246 27056
rect 32600 26948 32904 26976
rect 30745 26939 30803 26945
rect 9582 26868 9588 26920
rect 9640 26908 9646 26920
rect 25225 26911 25283 26917
rect 25225 26908 25237 26911
rect 9640 26880 25237 26908
rect 9640 26868 9646 26880
rect 25225 26877 25237 26880
rect 25271 26908 25283 26911
rect 25406 26908 25412 26920
rect 25271 26880 25412 26908
rect 25271 26877 25283 26880
rect 25225 26871 25283 26877
rect 25406 26868 25412 26880
rect 25464 26868 25470 26920
rect 26605 26911 26663 26917
rect 26605 26877 26617 26911
rect 26651 26877 26663 26911
rect 26605 26871 26663 26877
rect 26697 26911 26755 26917
rect 26697 26877 26709 26911
rect 26743 26908 26755 26911
rect 26970 26908 26976 26920
rect 26743 26880 26976 26908
rect 26743 26877 26755 26880
rect 26697 26871 26755 26877
rect 1854 26840 1860 26852
rect 1815 26812 1860 26840
rect 1854 26800 1860 26812
rect 1912 26800 1918 26852
rect 2041 26843 2099 26849
rect 2041 26809 2053 26843
rect 2087 26840 2099 26843
rect 2590 26840 2596 26852
rect 2087 26812 2596 26840
rect 2087 26809 2099 26812
rect 2041 26803 2099 26809
rect 2590 26800 2596 26812
rect 2648 26800 2654 26852
rect 26620 26840 26648 26871
rect 26970 26868 26976 26880
rect 27028 26908 27034 26920
rect 27522 26908 27528 26920
rect 27028 26880 27528 26908
rect 27028 26868 27034 26880
rect 27522 26868 27528 26880
rect 27580 26868 27586 26920
rect 30469 26911 30527 26917
rect 30469 26877 30481 26911
rect 30515 26908 30527 26911
rect 31386 26908 31392 26920
rect 30515 26880 31392 26908
rect 30515 26877 30527 26880
rect 30469 26871 30527 26877
rect 31386 26868 31392 26880
rect 31444 26868 31450 26920
rect 32766 26908 32772 26920
rect 32727 26880 32772 26908
rect 32766 26868 32772 26880
rect 32824 26868 32830 26920
rect 32876 26917 32904 26948
rect 32862 26911 32920 26917
rect 32862 26877 32874 26911
rect 32908 26877 32920 26911
rect 33134 26908 33140 26920
rect 33095 26880 33140 26908
rect 32862 26871 32920 26877
rect 33134 26868 33140 26880
rect 33192 26868 33198 26920
rect 33275 26911 33333 26917
rect 33275 26877 33287 26911
rect 33321 26908 33333 26911
rect 37550 26908 37556 26920
rect 33321 26880 37556 26908
rect 33321 26877 33333 26880
rect 33275 26871 33333 26877
rect 37550 26868 37556 26880
rect 37608 26868 37614 26920
rect 37918 26908 37924 26920
rect 37879 26880 37924 26908
rect 37918 26868 37924 26880
rect 37976 26868 37982 26920
rect 27154 26840 27160 26852
rect 26620 26812 27160 26840
rect 27154 26800 27160 26812
rect 27212 26800 27218 26852
rect 32950 26800 32956 26852
rect 33008 26840 33014 26852
rect 33045 26843 33103 26849
rect 33045 26840 33057 26843
rect 33008 26812 33057 26840
rect 33008 26800 33014 26812
rect 33045 26809 33057 26812
rect 33091 26809 33103 26843
rect 33045 26803 33103 26809
rect 32766 26732 32772 26784
rect 32824 26772 32830 26784
rect 33413 26775 33471 26781
rect 33413 26772 33425 26775
rect 32824 26744 33425 26772
rect 32824 26732 32830 26744
rect 33413 26741 33425 26744
rect 33459 26741 33471 26775
rect 33413 26735 33471 26741
rect 1104 26682 38824 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 38824 26682
rect 1104 26608 38824 26630
rect 4062 26528 4068 26580
rect 4120 26568 4126 26580
rect 32861 26571 32919 26577
rect 32861 26568 32873 26571
rect 4120 26540 32873 26568
rect 4120 26528 4126 26540
rect 32861 26537 32873 26540
rect 32907 26537 32919 26571
rect 32861 26531 32919 26537
rect 32876 26500 32904 26531
rect 33134 26528 33140 26580
rect 33192 26568 33198 26580
rect 33192 26540 33456 26568
rect 33192 26528 33198 26540
rect 33428 26509 33456 26540
rect 33566 26540 36584 26568
rect 33413 26503 33471 26509
rect 32876 26472 33181 26500
rect 25317 26435 25375 26441
rect 25317 26401 25329 26435
rect 25363 26432 25375 26435
rect 28074 26432 28080 26444
rect 25363 26404 28080 26432
rect 25363 26401 25375 26404
rect 25317 26395 25375 26401
rect 28074 26392 28080 26404
rect 28132 26392 28138 26444
rect 32674 26392 32680 26444
rect 32732 26432 32738 26444
rect 33153 26441 33181 26472
rect 33413 26469 33425 26503
rect 33459 26469 33471 26503
rect 33413 26463 33471 26469
rect 33566 26441 33594 26540
rect 36170 26500 36176 26512
rect 34164 26472 36176 26500
rect 34164 26441 34192 26472
rect 36170 26460 36176 26472
rect 36228 26460 36234 26512
rect 36556 26500 36584 26540
rect 36630 26528 36636 26580
rect 36688 26568 36694 26580
rect 37185 26571 37243 26577
rect 37185 26568 37197 26571
rect 36688 26540 37197 26568
rect 36688 26528 36694 26540
rect 37185 26537 37197 26540
rect 37231 26537 37243 26571
rect 37185 26531 37243 26537
rect 37826 26500 37832 26512
rect 36556 26472 37832 26500
rect 37826 26460 37832 26472
rect 37884 26460 37890 26512
rect 33045 26435 33103 26441
rect 33045 26432 33057 26435
rect 32732 26404 33057 26432
rect 32732 26392 32738 26404
rect 33045 26401 33057 26404
rect 33091 26401 33103 26435
rect 33045 26395 33103 26401
rect 33138 26435 33196 26441
rect 33138 26401 33150 26435
rect 33184 26401 33196 26435
rect 33138 26395 33196 26401
rect 33321 26435 33379 26441
rect 33321 26401 33333 26435
rect 33367 26401 33379 26435
rect 33321 26395 33379 26401
rect 33551 26435 33609 26441
rect 33551 26401 33563 26435
rect 33597 26401 33609 26435
rect 33551 26395 33609 26401
rect 34149 26435 34207 26441
rect 34149 26401 34161 26435
rect 34195 26401 34207 26435
rect 34149 26395 34207 26401
rect 25041 26367 25099 26373
rect 25041 26333 25053 26367
rect 25087 26364 25099 26367
rect 25222 26364 25228 26376
rect 25087 26336 25228 26364
rect 25087 26333 25099 26336
rect 25041 26327 25099 26333
rect 25222 26324 25228 26336
rect 25280 26324 25286 26376
rect 25406 26324 25412 26376
rect 25464 26364 25470 26376
rect 26050 26364 26056 26376
rect 25464 26336 26056 26364
rect 25464 26324 25470 26336
rect 26050 26324 26056 26336
rect 26108 26364 26114 26376
rect 26421 26367 26479 26373
rect 26421 26364 26433 26367
rect 26108 26336 26433 26364
rect 26108 26324 26114 26336
rect 26421 26333 26433 26336
rect 26467 26333 26479 26367
rect 26421 26327 26479 26333
rect 32950 26324 32956 26376
rect 33008 26364 33014 26376
rect 33336 26364 33364 26395
rect 34238 26392 34244 26444
rect 34296 26432 34302 26444
rect 34425 26435 34483 26441
rect 34296 26404 34341 26432
rect 34296 26392 34302 26404
rect 34425 26401 34437 26435
rect 34471 26401 34483 26435
rect 34425 26395 34483 26401
rect 34517 26435 34575 26441
rect 34517 26401 34529 26435
rect 34563 26401 34575 26435
rect 34517 26395 34575 26401
rect 34655 26435 34713 26441
rect 34655 26401 34667 26435
rect 34701 26432 34713 26435
rect 37366 26432 37372 26444
rect 34701 26404 37228 26432
rect 37327 26404 37372 26432
rect 34701 26401 34713 26404
rect 34655 26395 34713 26401
rect 34330 26364 34336 26376
rect 33008 26336 33364 26364
rect 33796 26336 34336 26364
rect 33008 26324 33014 26336
rect 33410 26256 33416 26308
rect 33468 26296 33474 26308
rect 33689 26299 33747 26305
rect 33689 26296 33701 26299
rect 33468 26268 33701 26296
rect 33468 26256 33474 26268
rect 33689 26265 33701 26268
rect 33735 26265 33747 26299
rect 33689 26259 33747 26265
rect 33318 26188 33324 26240
rect 33376 26228 33382 26240
rect 33796 26228 33824 26336
rect 34330 26324 34336 26336
rect 34388 26364 34394 26376
rect 34440 26364 34468 26395
rect 34388 26336 34468 26364
rect 34388 26324 34394 26336
rect 34146 26256 34152 26308
rect 34204 26296 34210 26308
rect 34532 26296 34560 26395
rect 34790 26324 34796 26376
rect 34848 26324 34854 26376
rect 37200 26364 37228 26404
rect 37366 26392 37372 26404
rect 37424 26392 37430 26444
rect 38654 26364 38660 26376
rect 37200 26336 38660 26364
rect 38654 26324 38660 26336
rect 38712 26324 38718 26376
rect 34204 26268 34560 26296
rect 34204 26256 34210 26268
rect 34606 26256 34612 26308
rect 34664 26296 34670 26308
rect 34808 26296 34836 26324
rect 34664 26268 34836 26296
rect 34664 26256 34670 26268
rect 34790 26228 34796 26240
rect 33376 26200 33824 26228
rect 34751 26200 34796 26228
rect 33376 26188 33382 26200
rect 34790 26188 34796 26200
rect 34848 26188 34854 26240
rect 1104 26138 38824 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 38824 26138
rect 1104 26064 38824 26086
rect 32306 25916 32312 25968
rect 32364 25956 32370 25968
rect 32674 25956 32680 25968
rect 32364 25928 32680 25956
rect 32364 25916 32370 25928
rect 32674 25916 32680 25928
rect 32732 25916 32738 25968
rect 33042 25916 33048 25968
rect 33100 25956 33106 25968
rect 33413 25959 33471 25965
rect 33413 25956 33425 25959
rect 33100 25928 33425 25956
rect 33100 25916 33106 25928
rect 33413 25925 33425 25928
rect 33459 25925 33471 25959
rect 33413 25919 33471 25925
rect 34440 25928 36032 25956
rect 34440 25900 34468 25928
rect 32214 25848 32220 25900
rect 32272 25888 32278 25900
rect 34422 25888 34428 25900
rect 32272 25860 34428 25888
rect 32272 25848 32278 25860
rect 34422 25848 34428 25860
rect 34480 25848 34486 25900
rect 1854 25820 1860 25832
rect 1815 25792 1860 25820
rect 1854 25780 1860 25792
rect 1912 25780 1918 25832
rect 32490 25780 32496 25832
rect 32548 25820 32554 25832
rect 32769 25823 32827 25829
rect 32769 25820 32781 25823
rect 32548 25792 32781 25820
rect 32548 25780 32554 25792
rect 32769 25789 32781 25792
rect 32815 25789 32827 25823
rect 32769 25783 32827 25789
rect 32862 25823 32920 25829
rect 32862 25789 32874 25823
rect 32908 25789 32920 25823
rect 33134 25820 33140 25832
rect 33095 25792 33140 25820
rect 32862 25783 32920 25789
rect 2041 25755 2099 25761
rect 2041 25721 2053 25755
rect 2087 25752 2099 25755
rect 2682 25752 2688 25764
rect 2087 25724 2688 25752
rect 2087 25721 2099 25724
rect 2041 25715 2099 25721
rect 2682 25712 2688 25724
rect 2740 25712 2746 25764
rect 32876 25752 32904 25783
rect 33134 25780 33140 25792
rect 33192 25780 33198 25832
rect 33275 25823 33333 25829
rect 33275 25789 33287 25823
rect 33321 25820 33333 25823
rect 34974 25820 34980 25832
rect 33321 25792 34980 25820
rect 33321 25789 33333 25792
rect 33275 25783 33333 25789
rect 34974 25780 34980 25792
rect 35032 25780 35038 25832
rect 36004 25829 36032 25928
rect 35897 25823 35955 25829
rect 35897 25789 35909 25823
rect 35943 25789 35955 25823
rect 35897 25783 35955 25789
rect 35989 25823 36047 25829
rect 35989 25789 36001 25823
rect 36035 25789 36047 25823
rect 36170 25820 36176 25832
rect 36131 25792 36176 25820
rect 35989 25783 36047 25789
rect 32600 25724 32904 25752
rect 2406 25644 2412 25696
rect 2464 25684 2470 25696
rect 32600 25693 32628 25724
rect 32950 25712 32956 25764
rect 33008 25752 33014 25764
rect 33045 25755 33103 25761
rect 33045 25752 33057 25755
rect 33008 25724 33057 25752
rect 33008 25712 33014 25724
rect 33045 25721 33057 25724
rect 33091 25721 33103 25755
rect 33045 25715 33103 25721
rect 35158 25712 35164 25764
rect 35216 25752 35222 25764
rect 35912 25752 35940 25783
rect 36170 25780 36176 25792
rect 36228 25780 36234 25832
rect 36265 25823 36323 25829
rect 36265 25789 36277 25823
rect 36311 25820 36323 25823
rect 36354 25820 36360 25832
rect 36311 25792 36360 25820
rect 36311 25789 36323 25792
rect 36265 25783 36323 25789
rect 36354 25780 36360 25792
rect 36412 25780 36418 25832
rect 37274 25820 37280 25832
rect 37235 25792 37280 25820
rect 37274 25780 37280 25792
rect 37332 25780 37338 25832
rect 37918 25820 37924 25832
rect 37879 25792 37924 25820
rect 37918 25780 37924 25792
rect 37976 25780 37982 25832
rect 36630 25752 36636 25764
rect 35216 25724 35848 25752
rect 35912 25724 36636 25752
rect 35216 25712 35222 25724
rect 32585 25687 32643 25693
rect 32585 25684 32597 25687
rect 2464 25656 32597 25684
rect 2464 25644 2470 25656
rect 32585 25653 32597 25656
rect 32631 25653 32643 25687
rect 32585 25647 32643 25653
rect 35618 25644 35624 25696
rect 35676 25684 35682 25696
rect 35713 25687 35771 25693
rect 35713 25684 35725 25687
rect 35676 25656 35725 25684
rect 35676 25644 35682 25656
rect 35713 25653 35725 25656
rect 35759 25653 35771 25687
rect 35820 25684 35848 25724
rect 36630 25712 36636 25724
rect 36688 25712 36694 25764
rect 36906 25712 36912 25764
rect 36964 25752 36970 25764
rect 37090 25752 37096 25764
rect 36964 25724 37096 25752
rect 36964 25712 36970 25724
rect 37090 25712 37096 25724
rect 37148 25712 37154 25764
rect 38378 25684 38384 25696
rect 35820 25656 38384 25684
rect 35713 25647 35771 25653
rect 38378 25644 38384 25656
rect 38436 25644 38442 25696
rect 1104 25594 38824 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 38824 25594
rect 1104 25520 38824 25542
rect 37366 25480 37372 25492
rect 35360 25452 37228 25480
rect 37327 25452 37372 25480
rect 32950 25372 32956 25424
rect 33008 25412 33014 25424
rect 33318 25412 33324 25424
rect 33008 25384 33324 25412
rect 33008 25372 33014 25384
rect 33318 25372 33324 25384
rect 33376 25372 33382 25424
rect 33413 25415 33471 25421
rect 33413 25381 33425 25415
rect 33459 25412 33471 25415
rect 34238 25412 34244 25424
rect 33459 25384 34244 25412
rect 33459 25381 33471 25384
rect 33413 25375 33471 25381
rect 34238 25372 34244 25384
rect 34296 25372 34302 25424
rect 35158 25412 35164 25424
rect 34348 25384 35164 25412
rect 1854 25344 1860 25356
rect 1815 25316 1860 25344
rect 1854 25304 1860 25316
rect 1912 25304 1918 25356
rect 32582 25304 32588 25356
rect 32640 25344 32646 25356
rect 33045 25347 33103 25353
rect 33045 25344 33057 25347
rect 32640 25316 33057 25344
rect 32640 25304 32646 25316
rect 33045 25313 33057 25316
rect 33091 25313 33103 25347
rect 33045 25307 33103 25313
rect 33138 25347 33196 25353
rect 33138 25313 33150 25347
rect 33184 25313 33196 25347
rect 33138 25307 33196 25313
rect 33551 25347 33609 25353
rect 33551 25313 33563 25347
rect 33597 25344 33609 25347
rect 34146 25344 34152 25356
rect 33597 25316 34152 25344
rect 33597 25313 33609 25316
rect 33551 25307 33609 25313
rect 2133 25279 2191 25285
rect 2133 25245 2145 25279
rect 2179 25276 2191 25279
rect 10318 25276 10324 25288
rect 2179 25248 10324 25276
rect 2179 25245 2191 25248
rect 2133 25239 2191 25245
rect 10318 25236 10324 25248
rect 10376 25236 10382 25288
rect 33153 25276 33181 25307
rect 34146 25304 34152 25316
rect 34204 25304 34210 25356
rect 34348 25353 34376 25384
rect 35158 25372 35164 25384
rect 35216 25372 35222 25424
rect 34333 25347 34391 25353
rect 34333 25313 34345 25347
rect 34379 25313 34391 25347
rect 34333 25307 34391 25313
rect 34422 25304 34428 25356
rect 34480 25344 34486 25356
rect 34609 25347 34667 25353
rect 34480 25316 34525 25344
rect 34480 25304 34486 25316
rect 34609 25313 34621 25347
rect 34655 25313 34667 25347
rect 34609 25307 34667 25313
rect 34624 25276 34652 25307
rect 34698 25304 34704 25356
rect 34756 25344 34762 25356
rect 35360 25353 35388 25452
rect 35452 25384 36492 25412
rect 35452 25353 35480 25384
rect 35345 25347 35403 25353
rect 34756 25316 34801 25344
rect 34756 25304 34762 25316
rect 35345 25313 35357 25347
rect 35391 25313 35403 25347
rect 35345 25307 35403 25313
rect 35437 25347 35495 25353
rect 35437 25313 35449 25347
rect 35483 25313 35495 25347
rect 35437 25307 35495 25313
rect 35621 25347 35679 25353
rect 35621 25313 35633 25347
rect 35667 25313 35679 25347
rect 35621 25307 35679 25313
rect 35452 25276 35480 25307
rect 32876 25248 33181 25276
rect 33244 25248 34652 25276
rect 35360 25248 35480 25276
rect 35636 25276 35664 25307
rect 35710 25304 35716 25356
rect 35768 25344 35774 25356
rect 36354 25344 36360 25356
rect 35768 25316 35813 25344
rect 36315 25316 36360 25344
rect 35768 25304 35774 25316
rect 36354 25304 36360 25316
rect 36412 25304 36418 25356
rect 36464 25353 36492 25384
rect 36538 25372 36544 25424
rect 36596 25412 36602 25424
rect 37200 25412 37228 25452
rect 37366 25440 37372 25452
rect 37424 25440 37430 25492
rect 38746 25412 38752 25424
rect 36596 25384 36768 25412
rect 37200 25384 38752 25412
rect 36596 25372 36602 25384
rect 36740 25353 36768 25384
rect 38746 25372 38752 25384
rect 38804 25372 38810 25424
rect 36449 25347 36507 25353
rect 36449 25313 36461 25347
rect 36495 25313 36507 25347
rect 36449 25307 36507 25313
rect 36633 25347 36691 25353
rect 36633 25313 36645 25347
rect 36679 25313 36691 25347
rect 36633 25307 36691 25313
rect 36725 25347 36783 25353
rect 36725 25313 36737 25347
rect 36771 25313 36783 25347
rect 37182 25344 37188 25356
rect 37143 25316 37188 25344
rect 36725 25307 36783 25313
rect 35636 25248 35756 25276
rect 2590 25100 2596 25152
rect 2648 25140 2654 25152
rect 32876 25149 32904 25248
rect 33134 25168 33140 25220
rect 33192 25208 33198 25220
rect 33244 25208 33272 25248
rect 33192 25180 33272 25208
rect 33192 25168 33198 25180
rect 33318 25168 33324 25220
rect 33376 25208 33382 25220
rect 34149 25211 34207 25217
rect 34149 25208 34161 25211
rect 33376 25180 34161 25208
rect 33376 25168 33382 25180
rect 34149 25177 34161 25180
rect 34195 25177 34207 25211
rect 34149 25171 34207 25177
rect 34422 25168 34428 25220
rect 34480 25208 34486 25220
rect 35360 25208 35388 25248
rect 35728 25220 35756 25248
rect 35894 25236 35900 25288
rect 35952 25276 35958 25288
rect 36538 25276 36544 25288
rect 35952 25248 36544 25276
rect 35952 25236 35958 25248
rect 36538 25236 36544 25248
rect 36596 25236 36602 25288
rect 34480 25180 35388 25208
rect 34480 25168 34486 25180
rect 35710 25168 35716 25220
rect 35768 25208 35774 25220
rect 36648 25208 36676 25307
rect 37182 25304 37188 25316
rect 37240 25304 37246 25356
rect 35768 25180 36676 25208
rect 35768 25168 35774 25180
rect 32861 25143 32919 25149
rect 32861 25140 32873 25143
rect 2648 25112 32873 25140
rect 2648 25100 2654 25112
rect 32861 25109 32873 25112
rect 32907 25109 32919 25143
rect 32861 25103 32919 25109
rect 33689 25143 33747 25149
rect 33689 25109 33701 25143
rect 33735 25140 33747 25143
rect 34238 25140 34244 25152
rect 33735 25112 34244 25140
rect 33735 25109 33747 25112
rect 33689 25103 33747 25109
rect 34238 25100 34244 25112
rect 34296 25100 34302 25152
rect 34514 25100 34520 25152
rect 34572 25140 34578 25152
rect 35161 25143 35219 25149
rect 35161 25140 35173 25143
rect 34572 25112 35173 25140
rect 34572 25100 34578 25112
rect 35161 25109 35173 25112
rect 35207 25109 35219 25143
rect 35161 25103 35219 25109
rect 35894 25100 35900 25152
rect 35952 25140 35958 25152
rect 36173 25143 36231 25149
rect 36173 25140 36185 25143
rect 35952 25112 36185 25140
rect 35952 25100 35958 25112
rect 36173 25109 36185 25112
rect 36219 25109 36231 25143
rect 36173 25103 36231 25109
rect 1104 25050 38824 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 38824 25050
rect 1104 24976 38824 24998
rect 32858 24828 32864 24880
rect 32916 24868 32922 24880
rect 33686 24868 33692 24880
rect 32916 24840 33692 24868
rect 32916 24828 32922 24840
rect 33686 24828 33692 24840
rect 33744 24828 33750 24880
rect 35710 24828 35716 24880
rect 35768 24868 35774 24880
rect 36170 24868 36176 24880
rect 35768 24840 36176 24868
rect 35768 24828 35774 24840
rect 27154 24800 27160 24812
rect 27115 24772 27160 24800
rect 27154 24760 27160 24772
rect 27212 24760 27218 24812
rect 34146 24800 34152 24812
rect 33244 24772 34152 24800
rect 27065 24735 27123 24741
rect 27065 24701 27077 24735
rect 27111 24732 27123 24735
rect 27614 24732 27620 24744
rect 27111 24704 27620 24732
rect 27111 24701 27123 24704
rect 27065 24695 27123 24701
rect 27614 24692 27620 24704
rect 27672 24692 27678 24744
rect 27709 24735 27767 24741
rect 27709 24701 27721 24735
rect 27755 24732 27767 24735
rect 27890 24732 27896 24744
rect 27755 24704 27896 24732
rect 27755 24701 27767 24704
rect 27709 24695 27767 24701
rect 27890 24692 27896 24704
rect 27948 24692 27954 24744
rect 32398 24692 32404 24744
rect 32456 24732 32462 24744
rect 32861 24735 32919 24741
rect 32861 24732 32873 24735
rect 32456 24704 32873 24732
rect 32456 24692 32462 24704
rect 32861 24701 32873 24704
rect 32907 24701 32919 24735
rect 32861 24695 32919 24701
rect 32950 24692 32956 24744
rect 33008 24732 33014 24744
rect 33244 24741 33272 24772
rect 34146 24760 34152 24772
rect 34204 24760 34210 24812
rect 35820 24772 36032 24800
rect 33229 24735 33287 24741
rect 33008 24704 33053 24732
rect 33008 24692 33014 24704
rect 33229 24701 33241 24735
rect 33275 24701 33287 24735
rect 33229 24695 33287 24701
rect 33367 24735 33425 24741
rect 33367 24701 33379 24735
rect 33413 24732 33425 24735
rect 33686 24732 33692 24744
rect 33413 24704 33692 24732
rect 33413 24701 33425 24704
rect 33367 24695 33425 24701
rect 33686 24692 33692 24704
rect 33744 24692 33750 24744
rect 2682 24624 2688 24676
rect 2740 24664 2746 24676
rect 32677 24667 32735 24673
rect 32677 24664 32689 24667
rect 2740 24636 32689 24664
rect 2740 24624 2746 24636
rect 32677 24633 32689 24636
rect 32723 24664 32735 24667
rect 33137 24667 33195 24673
rect 33137 24664 33149 24667
rect 32723 24636 33149 24664
rect 32723 24633 32735 24636
rect 32677 24627 32735 24633
rect 33137 24633 33149 24636
rect 33183 24633 33195 24667
rect 33137 24627 33195 24633
rect 34514 24624 34520 24676
rect 34572 24664 34578 24676
rect 35250 24664 35256 24676
rect 34572 24636 35256 24664
rect 34572 24624 34578 24636
rect 35250 24624 35256 24636
rect 35308 24624 35314 24676
rect 27522 24556 27528 24608
rect 27580 24596 27586 24608
rect 27801 24599 27859 24605
rect 27801 24596 27813 24599
rect 27580 24568 27813 24596
rect 27580 24556 27586 24568
rect 27801 24565 27813 24568
rect 27847 24565 27859 24599
rect 27801 24559 27859 24565
rect 32582 24556 32588 24608
rect 32640 24596 32646 24608
rect 33505 24599 33563 24605
rect 33505 24596 33517 24599
rect 32640 24568 33517 24596
rect 32640 24556 32646 24568
rect 33505 24565 33517 24568
rect 33551 24565 33563 24599
rect 33505 24559 33563 24565
rect 34146 24556 34152 24608
rect 34204 24596 34210 24608
rect 35713 24599 35771 24605
rect 35713 24596 35725 24599
rect 34204 24568 35725 24596
rect 34204 24556 34210 24568
rect 35713 24565 35725 24568
rect 35759 24565 35771 24599
rect 35820 24596 35848 24772
rect 36004 24741 36032 24772
rect 35897 24735 35955 24741
rect 35897 24701 35909 24735
rect 35943 24701 35955 24735
rect 35897 24695 35955 24701
rect 35989 24735 36047 24741
rect 35989 24701 36001 24735
rect 36035 24701 36047 24735
rect 36088 24732 36116 24840
rect 36170 24828 36176 24840
rect 36228 24828 36234 24880
rect 36173 24735 36231 24741
rect 36173 24732 36185 24735
rect 36088 24704 36185 24732
rect 35989 24695 36047 24701
rect 36173 24701 36185 24704
rect 36219 24701 36231 24735
rect 36173 24695 36231 24701
rect 35912 24664 35940 24695
rect 36262 24692 36268 24744
rect 36320 24732 36326 24744
rect 37274 24732 37280 24744
rect 36320 24704 36365 24732
rect 37235 24704 37280 24732
rect 36320 24692 36326 24704
rect 37274 24692 37280 24704
rect 37332 24692 37338 24744
rect 37918 24732 37924 24744
rect 37879 24704 37924 24732
rect 37918 24692 37924 24704
rect 37976 24692 37982 24744
rect 37090 24664 37096 24676
rect 35912 24636 37096 24664
rect 37090 24624 37096 24636
rect 37148 24624 37154 24676
rect 36170 24596 36176 24608
rect 35820 24568 36176 24596
rect 35713 24559 35771 24565
rect 36170 24556 36176 24568
rect 36228 24556 36234 24608
rect 36262 24556 36268 24608
rect 36320 24596 36326 24608
rect 36814 24596 36820 24608
rect 36320 24568 36820 24596
rect 36320 24556 36326 24568
rect 36814 24556 36820 24568
rect 36872 24556 36878 24608
rect 1104 24506 38824 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 38824 24506
rect 1104 24432 38824 24454
rect 28905 24395 28963 24401
rect 28905 24361 28917 24395
rect 28951 24392 28963 24395
rect 29914 24392 29920 24404
rect 28951 24364 29920 24392
rect 28951 24361 28963 24364
rect 28905 24355 28963 24361
rect 29914 24352 29920 24364
rect 29972 24352 29978 24404
rect 34238 24352 34244 24404
rect 34296 24392 34302 24404
rect 35250 24392 35256 24404
rect 34296 24364 35256 24392
rect 34296 24352 34302 24364
rect 35250 24352 35256 24364
rect 35308 24352 35314 24404
rect 37182 24392 37188 24404
rect 37143 24364 37188 24392
rect 37182 24352 37188 24364
rect 37240 24352 37246 24404
rect 27614 24284 27620 24336
rect 27672 24324 27678 24336
rect 29457 24327 29515 24333
rect 27672 24296 28396 24324
rect 27672 24284 27678 24296
rect 1854 24256 1860 24268
rect 1815 24228 1860 24256
rect 1854 24216 1860 24228
rect 1912 24216 1918 24268
rect 27154 24216 27160 24268
rect 27212 24256 27218 24268
rect 28368 24265 28396 24296
rect 29457 24293 29469 24327
rect 29503 24324 29515 24327
rect 31846 24324 31852 24336
rect 29503 24296 31852 24324
rect 29503 24293 29515 24296
rect 29457 24287 29515 24293
rect 31846 24284 31852 24296
rect 31904 24284 31910 24336
rect 32398 24284 32404 24336
rect 32456 24324 32462 24336
rect 38286 24324 38292 24336
rect 32456 24296 33640 24324
rect 32456 24284 32462 24296
rect 27985 24259 28043 24265
rect 27985 24256 27997 24259
rect 27212 24228 27997 24256
rect 27212 24216 27218 24228
rect 27985 24225 27997 24228
rect 28031 24225 28043 24259
rect 27985 24219 28043 24225
rect 28077 24259 28135 24265
rect 28077 24225 28089 24259
rect 28123 24225 28135 24259
rect 28077 24219 28135 24225
rect 28353 24259 28411 24265
rect 28353 24225 28365 24259
rect 28399 24225 28411 24259
rect 28353 24219 28411 24225
rect 27890 24148 27896 24200
rect 27948 24188 27954 24200
rect 28092 24188 28120 24219
rect 28626 24216 28632 24268
rect 28684 24256 28690 24268
rect 29181 24259 29239 24265
rect 29181 24256 29193 24259
rect 28684 24228 29193 24256
rect 28684 24216 28690 24228
rect 29181 24225 29193 24228
rect 29227 24225 29239 24259
rect 29181 24219 29239 24225
rect 32950 24216 32956 24268
rect 33008 24256 33014 24268
rect 33612 24265 33640 24296
rect 35544 24296 38292 24324
rect 35544 24265 35572 24296
rect 38286 24284 38292 24296
rect 38344 24284 38350 24336
rect 33229 24259 33287 24265
rect 33229 24256 33241 24259
rect 33008 24228 33241 24256
rect 33008 24216 33014 24228
rect 33229 24225 33241 24228
rect 33275 24225 33287 24259
rect 33229 24219 33287 24225
rect 33321 24259 33379 24265
rect 33321 24225 33333 24259
rect 33367 24225 33379 24259
rect 33321 24219 33379 24225
rect 33597 24259 33655 24265
rect 33597 24225 33609 24259
rect 33643 24225 33655 24259
rect 33597 24219 33655 24225
rect 35529 24259 35587 24265
rect 35529 24225 35541 24259
rect 35575 24225 35587 24259
rect 35529 24219 35587 24225
rect 35621 24259 35679 24265
rect 35621 24225 35633 24259
rect 35667 24225 35679 24259
rect 35621 24219 35679 24225
rect 29086 24188 29092 24200
rect 27948 24160 28120 24188
rect 28999 24160 29092 24188
rect 27948 24148 27954 24160
rect 29086 24148 29092 24160
rect 29144 24188 29150 24200
rect 29549 24191 29607 24197
rect 29549 24188 29561 24191
rect 29144 24160 29561 24188
rect 29144 24148 29150 24160
rect 29549 24157 29561 24160
rect 29595 24188 29607 24191
rect 33134 24188 33140 24200
rect 29595 24160 33140 24188
rect 29595 24157 29607 24160
rect 29549 24151 29607 24157
rect 33134 24148 33140 24160
rect 33192 24148 33198 24200
rect 33336 24188 33364 24219
rect 35345 24191 35403 24197
rect 35345 24188 35357 24191
rect 33336 24160 35357 24188
rect 35345 24157 35357 24160
rect 35391 24157 35403 24191
rect 35636 24188 35664 24219
rect 35710 24216 35716 24268
rect 35768 24256 35774 24268
rect 35805 24259 35863 24265
rect 35805 24256 35817 24259
rect 35768 24228 35817 24256
rect 35768 24216 35774 24228
rect 35805 24225 35817 24228
rect 35851 24225 35863 24259
rect 35805 24219 35863 24225
rect 35897 24259 35955 24265
rect 35897 24225 35909 24259
rect 35943 24256 35955 24259
rect 36078 24256 36084 24268
rect 35943 24228 36084 24256
rect 35943 24225 35955 24228
rect 35897 24219 35955 24225
rect 36078 24216 36084 24228
rect 36136 24216 36142 24268
rect 37366 24256 37372 24268
rect 37327 24228 37372 24256
rect 37366 24216 37372 24228
rect 37424 24216 37430 24268
rect 35636 24160 36124 24188
rect 35345 24151 35403 24157
rect 36096 24132 36124 24160
rect 27522 24080 27528 24132
rect 27580 24120 27586 24132
rect 28261 24123 28319 24129
rect 28261 24120 28273 24123
rect 27580 24092 28273 24120
rect 27580 24080 27586 24092
rect 28261 24089 28273 24092
rect 28307 24089 28319 24123
rect 28261 24083 28319 24089
rect 32122 24080 32128 24132
rect 32180 24120 32186 24132
rect 33505 24123 33563 24129
rect 33505 24120 33517 24123
rect 32180 24092 33517 24120
rect 32180 24080 32186 24092
rect 33505 24089 33517 24092
rect 33551 24089 33563 24123
rect 33505 24083 33563 24089
rect 34330 24080 34336 24132
rect 34388 24120 34394 24132
rect 35158 24120 35164 24132
rect 34388 24092 35164 24120
rect 34388 24080 34394 24092
rect 35158 24080 35164 24092
rect 35216 24080 35222 24132
rect 36078 24080 36084 24132
rect 36136 24080 36142 24132
rect 2133 24055 2191 24061
rect 2133 24021 2145 24055
rect 2179 24052 2191 24055
rect 20990 24052 20996 24064
rect 2179 24024 20996 24052
rect 2179 24021 2191 24024
rect 2133 24015 2191 24021
rect 20990 24012 20996 24024
rect 21048 24012 21054 24064
rect 27246 24012 27252 24064
rect 27304 24052 27310 24064
rect 27801 24055 27859 24061
rect 27801 24052 27813 24055
rect 27304 24024 27813 24052
rect 27304 24012 27310 24024
rect 27801 24021 27813 24024
rect 27847 24021 27859 24055
rect 27801 24015 27859 24021
rect 31938 24012 31944 24064
rect 31996 24052 32002 24064
rect 33045 24055 33103 24061
rect 33045 24052 33057 24055
rect 31996 24024 33057 24052
rect 31996 24012 32002 24024
rect 33045 24021 33057 24024
rect 33091 24021 33103 24055
rect 33045 24015 33103 24021
rect 33686 24012 33692 24064
rect 33744 24052 33750 24064
rect 38010 24052 38016 24064
rect 33744 24024 38016 24052
rect 33744 24012 33750 24024
rect 38010 24012 38016 24024
rect 38068 24012 38074 24064
rect 1104 23962 38824 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 38824 23962
rect 1104 23888 38824 23910
rect 2133 23851 2191 23857
rect 2133 23817 2145 23851
rect 2179 23848 2191 23851
rect 9030 23848 9036 23860
rect 2179 23820 9036 23848
rect 2179 23817 2191 23820
rect 2133 23811 2191 23817
rect 9030 23808 9036 23820
rect 9088 23808 9094 23860
rect 31846 23808 31852 23860
rect 31904 23848 31910 23860
rect 34422 23848 34428 23860
rect 31904 23820 34428 23848
rect 31904 23808 31910 23820
rect 34422 23808 34428 23820
rect 34480 23808 34486 23860
rect 35710 23808 35716 23860
rect 35768 23848 35774 23860
rect 37182 23848 37188 23860
rect 35768 23820 37188 23848
rect 35768 23808 35774 23820
rect 37182 23808 37188 23820
rect 37240 23808 37246 23860
rect 28534 23740 28540 23792
rect 28592 23780 28598 23792
rect 32950 23780 32956 23792
rect 28592 23752 32956 23780
rect 28592 23740 28598 23752
rect 32950 23740 32956 23752
rect 33008 23780 33014 23792
rect 33008 23752 33548 23780
rect 33008 23740 33014 23752
rect 28718 23672 28724 23724
rect 28776 23712 28782 23724
rect 28776 23684 31754 23712
rect 28776 23672 28782 23684
rect 27246 23644 27252 23656
rect 27207 23616 27252 23644
rect 27246 23604 27252 23616
rect 27304 23604 27310 23656
rect 27433 23647 27491 23653
rect 27433 23613 27445 23647
rect 27479 23613 27491 23647
rect 27890 23644 27896 23656
rect 27851 23616 27896 23644
rect 27433 23607 27491 23613
rect 1854 23576 1860 23588
rect 1815 23548 1860 23576
rect 1854 23536 1860 23548
rect 1912 23536 1918 23588
rect 26142 23536 26148 23588
rect 26200 23576 26206 23588
rect 27448 23576 27476 23607
rect 27890 23604 27896 23616
rect 27948 23604 27954 23656
rect 28077 23647 28135 23653
rect 28077 23613 28089 23647
rect 28123 23644 28135 23647
rect 29086 23644 29092 23656
rect 28123 23616 29092 23644
rect 28123 23613 28135 23616
rect 28077 23607 28135 23613
rect 28092 23576 28120 23607
rect 29086 23604 29092 23616
rect 29144 23604 29150 23656
rect 31726 23644 31754 23684
rect 33321 23647 33379 23653
rect 33321 23644 33333 23647
rect 31726 23616 33333 23644
rect 33321 23613 33333 23616
rect 33367 23613 33379 23647
rect 33321 23607 33379 23613
rect 33413 23647 33471 23653
rect 33413 23613 33425 23647
rect 33459 23613 33471 23647
rect 33520 23644 33548 23752
rect 35894 23740 35900 23792
rect 35952 23740 35958 23792
rect 33597 23715 33655 23721
rect 33597 23681 33609 23715
rect 33643 23712 33655 23715
rect 34238 23712 34244 23724
rect 33643 23684 34244 23712
rect 33643 23681 33655 23684
rect 33597 23675 33655 23681
rect 34238 23672 34244 23684
rect 34296 23672 34302 23724
rect 34974 23672 34980 23724
rect 35032 23712 35038 23724
rect 35912 23712 35940 23740
rect 36078 23712 36084 23724
rect 35032 23684 35940 23712
rect 36004 23684 36084 23712
rect 35032 23672 35038 23684
rect 33689 23647 33747 23653
rect 33689 23644 33701 23647
rect 33520 23616 33701 23644
rect 33413 23607 33471 23613
rect 33689 23613 33701 23616
rect 33735 23613 33747 23647
rect 33689 23607 33747 23613
rect 26200 23548 28120 23576
rect 33428 23576 33456 23607
rect 35250 23604 35256 23656
rect 35308 23644 35314 23656
rect 36004 23653 36032 23684
rect 36078 23672 36084 23684
rect 36136 23672 36142 23724
rect 35897 23647 35955 23653
rect 35308 23616 35848 23644
rect 35308 23604 35314 23616
rect 35618 23576 35624 23588
rect 33428 23548 35624 23576
rect 26200 23536 26206 23548
rect 35618 23536 35624 23548
rect 35676 23536 35682 23588
rect 26694 23468 26700 23520
rect 26752 23508 26758 23520
rect 27341 23511 27399 23517
rect 27341 23508 27353 23511
rect 26752 23480 27353 23508
rect 26752 23468 26758 23480
rect 27341 23477 27353 23480
rect 27387 23477 27399 23511
rect 27982 23508 27988 23520
rect 27943 23480 27988 23508
rect 27341 23471 27399 23477
rect 27982 23468 27988 23480
rect 28040 23468 28046 23520
rect 33134 23508 33140 23520
rect 33095 23480 33140 23508
rect 33134 23468 33140 23480
rect 33192 23468 33198 23520
rect 35710 23508 35716 23520
rect 35671 23480 35716 23508
rect 35710 23468 35716 23480
rect 35768 23468 35774 23520
rect 35820 23508 35848 23616
rect 35897 23613 35909 23647
rect 35943 23613 35955 23647
rect 35897 23607 35955 23613
rect 35989 23647 36047 23653
rect 35989 23613 36001 23647
rect 36035 23613 36047 23647
rect 36170 23644 36176 23656
rect 36131 23616 36176 23644
rect 35989 23607 36047 23613
rect 35912 23576 35940 23607
rect 36170 23604 36176 23616
rect 36228 23604 36234 23656
rect 36265 23647 36323 23653
rect 36265 23613 36277 23647
rect 36311 23644 36323 23647
rect 36446 23644 36452 23656
rect 36311 23616 36452 23644
rect 36311 23613 36323 23616
rect 36265 23607 36323 23613
rect 36446 23604 36452 23616
rect 36504 23604 36510 23656
rect 37274 23644 37280 23656
rect 37235 23616 37280 23644
rect 37274 23604 37280 23616
rect 37332 23604 37338 23656
rect 37918 23644 37924 23656
rect 37879 23616 37924 23644
rect 37918 23604 37924 23616
rect 37976 23604 37982 23656
rect 36814 23576 36820 23588
rect 35912 23548 36820 23576
rect 36814 23536 36820 23548
rect 36872 23536 36878 23588
rect 35894 23508 35900 23520
rect 35820 23480 35900 23508
rect 35894 23468 35900 23480
rect 35952 23468 35958 23520
rect 1104 23418 38824 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 38824 23418
rect 1104 23344 38824 23366
rect 27890 23264 27896 23316
rect 27948 23304 27954 23316
rect 29181 23307 29239 23313
rect 29181 23304 29193 23307
rect 27948 23276 29193 23304
rect 27948 23264 27954 23276
rect 29181 23273 29193 23276
rect 29227 23273 29239 23307
rect 29181 23267 29239 23273
rect 30282 23264 30288 23316
rect 30340 23304 30346 23316
rect 30340 23276 35848 23304
rect 30340 23264 30346 23276
rect 27982 23196 27988 23248
rect 28040 23245 28046 23248
rect 28040 23239 28104 23245
rect 28040 23205 28058 23239
rect 28092 23205 28104 23239
rect 28040 23199 28104 23205
rect 28040 23196 28046 23199
rect 32490 23196 32496 23248
rect 32548 23236 32554 23248
rect 34146 23236 34152 23248
rect 32548 23208 34152 23236
rect 32548 23196 32554 23208
rect 34146 23196 34152 23208
rect 34204 23196 34210 23248
rect 34974 23236 34980 23248
rect 34348 23208 34980 23236
rect 28350 23128 28356 23180
rect 28408 23168 28414 23180
rect 33229 23171 33287 23177
rect 33229 23168 33241 23171
rect 28408 23140 33241 23168
rect 28408 23128 28414 23140
rect 33229 23137 33241 23140
rect 33275 23137 33287 23171
rect 33229 23131 33287 23137
rect 33318 23128 33324 23180
rect 33376 23168 33382 23180
rect 33597 23171 33655 23177
rect 33376 23140 33421 23168
rect 33376 23128 33382 23140
rect 33597 23137 33609 23171
rect 33643 23137 33655 23171
rect 33597 23131 33655 23137
rect 27430 23060 27436 23112
rect 27488 23100 27494 23112
rect 27801 23103 27859 23109
rect 27801 23100 27813 23103
rect 27488 23072 27813 23100
rect 27488 23060 27494 23072
rect 27801 23069 27813 23072
rect 27847 23069 27859 23103
rect 27801 23063 27859 23069
rect 32950 23060 32956 23112
rect 33008 23100 33014 23112
rect 33612 23100 33640 23131
rect 33686 23128 33692 23180
rect 33744 23168 33750 23180
rect 34348 23177 34376 23208
rect 34974 23196 34980 23208
rect 35032 23196 35038 23248
rect 34241 23171 34299 23177
rect 34241 23168 34253 23171
rect 33744 23140 34253 23168
rect 33744 23128 33750 23140
rect 34241 23137 34253 23140
rect 34287 23137 34299 23171
rect 34241 23131 34299 23137
rect 34333 23171 34391 23177
rect 34333 23137 34345 23171
rect 34379 23137 34391 23171
rect 34606 23168 34612 23180
rect 34567 23140 34612 23168
rect 34333 23131 34391 23137
rect 34606 23128 34612 23140
rect 34664 23128 34670 23180
rect 35820 23177 35848 23276
rect 35437 23171 35495 23177
rect 35437 23137 35449 23171
rect 35483 23137 35495 23171
rect 35437 23131 35495 23137
rect 35529 23171 35587 23177
rect 35529 23137 35541 23171
rect 35575 23137 35587 23171
rect 35529 23131 35587 23137
rect 35713 23171 35771 23177
rect 35713 23137 35725 23171
rect 35759 23137 35771 23171
rect 35713 23131 35771 23137
rect 35805 23171 35863 23177
rect 35805 23137 35817 23171
rect 35851 23137 35863 23171
rect 35805 23131 35863 23137
rect 33008 23072 33640 23100
rect 33008 23060 33014 23072
rect 33336 23044 33364 23072
rect 31478 23032 31484 23044
rect 28736 23004 31484 23032
rect 27798 22924 27804 22976
rect 27856 22964 27862 22976
rect 28736 22964 28764 23004
rect 31478 22992 31484 23004
rect 31536 22992 31542 23044
rect 33318 22992 33324 23044
rect 33376 22992 33382 23044
rect 33505 23035 33563 23041
rect 33505 23001 33517 23035
rect 33551 23032 33563 23035
rect 34517 23035 34575 23041
rect 33551 23004 33732 23032
rect 33551 23001 33563 23004
rect 33505 22995 33563 23001
rect 33704 22976 33732 23004
rect 34517 23001 34529 23035
rect 34563 23032 34575 23035
rect 35342 23032 35348 23044
rect 34563 23004 35348 23032
rect 34563 23001 34575 23004
rect 34517 22995 34575 23001
rect 35342 22992 35348 23004
rect 35400 22992 35406 23044
rect 27856 22936 28764 22964
rect 27856 22924 27862 22936
rect 32950 22924 32956 22976
rect 33008 22964 33014 22976
rect 33045 22967 33103 22973
rect 33045 22964 33057 22967
rect 33008 22936 33057 22964
rect 33008 22924 33014 22936
rect 33045 22933 33057 22936
rect 33091 22933 33103 22967
rect 33045 22927 33103 22933
rect 33686 22924 33692 22976
rect 33744 22924 33750 22976
rect 33870 22924 33876 22976
rect 33928 22964 33934 22976
rect 34057 22967 34115 22973
rect 34057 22964 34069 22967
rect 33928 22936 34069 22964
rect 33928 22924 33934 22936
rect 34057 22933 34069 22936
rect 34103 22933 34115 22967
rect 34057 22927 34115 22933
rect 34606 22924 34612 22976
rect 34664 22964 34670 22976
rect 35253 22967 35311 22973
rect 35253 22964 35265 22967
rect 34664 22936 35265 22964
rect 34664 22924 34670 22936
rect 35253 22933 35265 22936
rect 35299 22933 35311 22967
rect 35452 22964 35480 23131
rect 35544 23032 35572 23131
rect 35728 23100 35756 23131
rect 36170 23100 36176 23112
rect 35728 23072 36176 23100
rect 36170 23060 36176 23072
rect 36228 23060 36234 23112
rect 36078 23032 36084 23044
rect 35544 23004 36084 23032
rect 36078 22992 36084 23004
rect 36136 22992 36142 23044
rect 37366 22964 37372 22976
rect 35452 22936 37372 22964
rect 35253 22927 35311 22933
rect 37366 22924 37372 22936
rect 37424 22924 37430 22976
rect 1104 22874 38824 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 38824 22874
rect 1104 22800 38824 22822
rect 27430 22760 27436 22772
rect 26436 22732 27436 22760
rect 26436 22633 26464 22732
rect 27430 22720 27436 22732
rect 27488 22720 27494 22772
rect 32214 22720 32220 22772
rect 32272 22760 32278 22772
rect 32309 22763 32367 22769
rect 32309 22760 32321 22763
rect 32272 22732 32321 22760
rect 32272 22720 32278 22732
rect 32309 22729 32321 22732
rect 32355 22729 32367 22763
rect 32309 22723 32367 22729
rect 32416 22732 33088 22760
rect 31846 22652 31852 22704
rect 31904 22692 31910 22704
rect 32416 22692 32444 22732
rect 31904 22664 32444 22692
rect 31904 22652 31910 22664
rect 32490 22652 32496 22704
rect 32548 22652 32554 22704
rect 26421 22627 26479 22633
rect 26421 22593 26433 22627
rect 26467 22593 26479 22627
rect 32508 22624 32536 22652
rect 26421 22587 26479 22593
rect 32140 22596 32536 22624
rect 1854 22556 1860 22568
rect 1815 22528 1860 22556
rect 1854 22516 1860 22528
rect 1912 22516 1918 22568
rect 26694 22565 26700 22568
rect 26688 22556 26700 22565
rect 26655 22528 26700 22556
rect 26688 22519 26700 22528
rect 26694 22516 26700 22519
rect 26752 22516 26758 22568
rect 31846 22516 31852 22568
rect 31904 22516 31910 22568
rect 32030 22556 32036 22568
rect 31991 22528 32036 22556
rect 32030 22516 32036 22528
rect 32088 22516 32094 22568
rect 32140 22565 32168 22596
rect 32674 22584 32680 22636
rect 32732 22584 32738 22636
rect 33060 22624 33088 22732
rect 33888 22732 35112 22760
rect 33321 22695 33379 22701
rect 33321 22661 33333 22695
rect 33367 22692 33379 22695
rect 33888 22692 33916 22732
rect 35084 22704 35112 22732
rect 36538 22720 36544 22772
rect 36596 22760 36602 22772
rect 37458 22760 37464 22772
rect 36596 22732 36860 22760
rect 37419 22732 37464 22760
rect 36596 22720 36602 22732
rect 34054 22692 34060 22704
rect 33367 22664 33916 22692
rect 33980 22664 34060 22692
rect 33367 22661 33379 22664
rect 33321 22655 33379 22661
rect 33060 22596 33180 22624
rect 32125 22559 32183 22565
rect 32125 22525 32137 22559
rect 32171 22525 32183 22559
rect 32125 22519 32183 22525
rect 32401 22559 32459 22565
rect 32401 22525 32413 22559
rect 32447 22556 32459 22559
rect 32490 22556 32496 22568
rect 32447 22528 32496 22556
rect 32447 22525 32459 22528
rect 32401 22519 32459 22525
rect 32490 22516 32496 22528
rect 32548 22516 32554 22568
rect 32692 22556 32720 22584
rect 33152 22565 33180 22596
rect 33045 22559 33103 22565
rect 33045 22556 33057 22559
rect 32692 22528 33057 22556
rect 33045 22525 33057 22528
rect 33091 22525 33103 22559
rect 33045 22519 33103 22525
rect 33137 22559 33195 22565
rect 33137 22525 33149 22559
rect 33183 22525 33195 22559
rect 33137 22519 33195 22525
rect 33318 22516 33324 22568
rect 33376 22565 33382 22568
rect 33376 22559 33425 22565
rect 33376 22525 33379 22559
rect 33413 22525 33425 22559
rect 33980 22556 34008 22664
rect 34054 22652 34060 22664
rect 34112 22652 34118 22704
rect 34146 22652 34152 22704
rect 34204 22692 34210 22704
rect 34204 22664 34285 22692
rect 34204 22652 34210 22664
rect 34257 22624 34285 22664
rect 35066 22652 35072 22704
rect 35124 22652 35130 22704
rect 35710 22652 35716 22704
rect 35768 22652 35774 22704
rect 34333 22627 34391 22633
rect 34333 22624 34345 22627
rect 34257 22596 34345 22624
rect 34333 22593 34345 22596
rect 34379 22593 34391 22627
rect 35728 22624 35756 22652
rect 36078 22624 36084 22636
rect 34333 22587 34391 22593
rect 34900 22596 35756 22624
rect 35991 22596 36084 22624
rect 34058 22559 34116 22565
rect 34058 22556 34070 22559
rect 33980 22528 34070 22556
rect 33376 22519 33425 22525
rect 34058 22525 34070 22528
rect 34104 22525 34116 22559
rect 34058 22519 34116 22525
rect 34149 22559 34207 22565
rect 34149 22525 34161 22559
rect 34195 22525 34207 22559
rect 34149 22519 34207 22525
rect 33376 22516 33382 22519
rect 31864 22488 31892 22516
rect 34164 22488 34192 22519
rect 34422 22516 34428 22568
rect 34480 22556 34486 22568
rect 34480 22528 34525 22556
rect 34480 22516 34486 22528
rect 34900 22488 34928 22596
rect 35250 22516 35256 22568
rect 35308 22556 35314 22568
rect 35710 22556 35716 22568
rect 35308 22528 35716 22556
rect 35308 22516 35314 22528
rect 35710 22516 35716 22528
rect 35768 22516 35774 22568
rect 36004 22565 36032 22596
rect 36078 22584 36084 22596
rect 36136 22624 36142 22636
rect 36538 22624 36544 22636
rect 36136 22596 36544 22624
rect 36136 22584 36142 22596
rect 36538 22584 36544 22596
rect 36596 22584 36602 22636
rect 35897 22559 35955 22565
rect 35897 22525 35909 22559
rect 35943 22525 35955 22559
rect 35897 22519 35955 22525
rect 35989 22559 36047 22565
rect 35989 22525 36001 22559
rect 36035 22525 36047 22559
rect 36170 22556 36176 22568
rect 36131 22528 36176 22556
rect 35989 22519 36047 22525
rect 31864 22460 32996 22488
rect 34164 22460 34928 22488
rect 35912 22488 35940 22519
rect 36170 22516 36176 22528
rect 36228 22516 36234 22568
rect 36265 22559 36323 22565
rect 36265 22525 36277 22559
rect 36311 22556 36323 22559
rect 36722 22556 36728 22568
rect 36311 22528 36728 22556
rect 36311 22525 36323 22528
rect 36265 22519 36323 22525
rect 36722 22516 36728 22528
rect 36780 22516 36786 22568
rect 36446 22488 36452 22500
rect 35912 22460 36452 22488
rect 2133 22423 2191 22429
rect 2133 22389 2145 22423
rect 2179 22420 2191 22423
rect 14550 22420 14556 22432
rect 2179 22392 14556 22420
rect 2179 22389 2191 22392
rect 2133 22383 2191 22389
rect 14550 22380 14556 22392
rect 14608 22380 14614 22432
rect 27614 22380 27620 22432
rect 27672 22420 27678 22432
rect 27801 22423 27859 22429
rect 27801 22420 27813 22423
rect 27672 22392 27813 22420
rect 27672 22380 27678 22392
rect 27801 22389 27813 22392
rect 27847 22389 27859 22423
rect 27801 22383 27859 22389
rect 31849 22423 31907 22429
rect 31849 22389 31861 22423
rect 31895 22420 31907 22423
rect 32398 22420 32404 22432
rect 31895 22392 32404 22420
rect 31895 22389 31907 22392
rect 31849 22383 31907 22389
rect 32398 22380 32404 22392
rect 32456 22380 32462 22432
rect 32858 22420 32864 22432
rect 32819 22392 32864 22420
rect 32858 22380 32864 22392
rect 32916 22380 32922 22432
rect 32968 22420 32996 22460
rect 36446 22448 36452 22460
rect 36504 22448 36510 22500
rect 33873 22423 33931 22429
rect 33873 22420 33885 22423
rect 32968 22392 33885 22420
rect 33873 22389 33885 22392
rect 33919 22389 33931 22423
rect 33873 22383 33931 22389
rect 34330 22380 34336 22432
rect 34388 22420 34394 22432
rect 34698 22420 34704 22432
rect 34388 22392 34704 22420
rect 34388 22380 34394 22392
rect 34698 22380 34704 22392
rect 34756 22380 34762 22432
rect 34882 22380 34888 22432
rect 34940 22420 34946 22432
rect 35713 22423 35771 22429
rect 35713 22420 35725 22423
rect 34940 22392 35725 22420
rect 34940 22380 34946 22392
rect 35713 22389 35725 22392
rect 35759 22389 35771 22423
rect 35713 22383 35771 22389
rect 36722 22380 36728 22432
rect 36780 22420 36786 22432
rect 36832 22420 36860 22732
rect 37458 22720 37464 22732
rect 37516 22720 37522 22772
rect 37274 22556 37280 22568
rect 37235 22528 37280 22556
rect 37274 22516 37280 22528
rect 37332 22516 37338 22568
rect 37918 22556 37924 22568
rect 37879 22528 37924 22556
rect 37918 22516 37924 22528
rect 37976 22516 37982 22568
rect 36780 22392 36860 22420
rect 36780 22380 36786 22392
rect 1104 22330 38824 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 38824 22330
rect 1104 22256 38824 22278
rect 36078 22216 36084 22228
rect 35360 22188 36084 22216
rect 1854 22148 1860 22160
rect 1815 22120 1860 22148
rect 1854 22108 1860 22120
rect 1912 22108 1918 22160
rect 32490 22108 32496 22160
rect 32548 22148 32554 22160
rect 34422 22148 34428 22160
rect 32548 22120 34428 22148
rect 32548 22108 32554 22120
rect 33226 22080 33232 22092
rect 33187 22052 33232 22080
rect 33226 22040 33232 22052
rect 33284 22040 33290 22092
rect 33612 22089 33640 22120
rect 34422 22108 34428 22120
rect 34480 22108 34486 22160
rect 33321 22083 33379 22089
rect 33321 22049 33333 22083
rect 33367 22049 33379 22083
rect 33321 22043 33379 22049
rect 33597 22083 33655 22089
rect 33597 22049 33609 22083
rect 33643 22049 33655 22083
rect 34606 22080 34612 22092
rect 33597 22043 33655 22049
rect 33704 22052 34612 22080
rect 30374 21972 30380 22024
rect 30432 22012 30438 22024
rect 30558 22012 30564 22024
rect 30432 21984 30564 22012
rect 30432 21972 30438 21984
rect 30558 21972 30564 21984
rect 30616 21972 30622 22024
rect 33336 22012 33364 22043
rect 33704 22012 33732 22052
rect 34606 22040 34612 22052
rect 34664 22040 34670 22092
rect 35066 22080 35072 22092
rect 35027 22052 35072 22080
rect 35066 22040 35072 22052
rect 35124 22040 35130 22092
rect 35360 22089 35388 22188
rect 36078 22176 36084 22188
rect 36136 22216 36142 22228
rect 36136 22188 36400 22216
rect 36136 22176 36142 22188
rect 36096 22120 36308 22148
rect 35161 22083 35219 22089
rect 35161 22049 35173 22083
rect 35207 22049 35219 22083
rect 35161 22043 35219 22049
rect 35345 22083 35403 22089
rect 35345 22049 35357 22083
rect 35391 22049 35403 22083
rect 35345 22043 35403 22049
rect 35437 22083 35495 22089
rect 35437 22049 35449 22083
rect 35483 22080 35495 22083
rect 35618 22080 35624 22092
rect 35483 22052 35624 22080
rect 35483 22049 35495 22052
rect 35437 22043 35495 22049
rect 34885 22015 34943 22021
rect 34885 22012 34897 22015
rect 33336 21984 33732 22012
rect 34670 21984 34897 22012
rect 34670 21956 34698 21984
rect 34885 21981 34897 21984
rect 34931 21981 34943 22015
rect 34885 21975 34943 21981
rect 32122 21904 32128 21956
rect 32180 21944 32186 21956
rect 34054 21944 34060 21956
rect 32180 21916 34060 21944
rect 32180 21904 32186 21916
rect 34054 21904 34060 21916
rect 34112 21904 34118 21956
rect 34606 21904 34612 21956
rect 34664 21916 34698 21956
rect 35176 21944 35204 22043
rect 35618 22040 35624 22052
rect 35676 22040 35682 22092
rect 36096 22089 36124 22120
rect 36081 22083 36139 22089
rect 36081 22049 36093 22083
rect 36127 22049 36139 22083
rect 36081 22043 36139 22049
rect 36173 22083 36231 22089
rect 36173 22049 36185 22083
rect 36219 22049 36231 22083
rect 36173 22043 36231 22049
rect 36188 21956 36216 22043
rect 36280 22012 36308 22120
rect 36372 22089 36400 22188
rect 36357 22083 36415 22089
rect 36357 22049 36369 22083
rect 36403 22049 36415 22083
rect 36357 22043 36415 22049
rect 36449 22083 36507 22089
rect 36449 22049 36461 22083
rect 36495 22080 36507 22083
rect 36722 22080 36728 22092
rect 36495 22052 36728 22080
rect 36495 22049 36507 22052
rect 36449 22043 36507 22049
rect 36722 22040 36728 22052
rect 36780 22040 36786 22092
rect 38562 22012 38568 22024
rect 36280 21984 38568 22012
rect 38562 21972 38568 21984
rect 38620 21972 38626 22024
rect 35176 21916 36032 21944
rect 34664 21904 34670 21916
rect 1949 21879 2007 21885
rect 1949 21845 1961 21879
rect 1995 21876 2007 21879
rect 16666 21876 16672 21888
rect 1995 21848 16672 21876
rect 1995 21845 2007 21848
rect 1949 21839 2007 21845
rect 16666 21836 16672 21848
rect 16724 21836 16730 21888
rect 33042 21876 33048 21888
rect 33003 21848 33048 21876
rect 33042 21836 33048 21848
rect 33100 21836 33106 21888
rect 33505 21879 33563 21885
rect 33505 21845 33517 21879
rect 33551 21876 33563 21879
rect 33686 21876 33692 21888
rect 33551 21848 33692 21876
rect 33551 21845 33563 21848
rect 33505 21839 33563 21845
rect 33686 21836 33692 21848
rect 33744 21836 33750 21888
rect 35894 21876 35900 21888
rect 35855 21848 35900 21876
rect 35894 21836 35900 21848
rect 35952 21836 35958 21888
rect 36004 21876 36032 21916
rect 36170 21904 36176 21956
rect 36228 21904 36234 21956
rect 36188 21876 36216 21904
rect 36004 21848 36216 21876
rect 1104 21786 38824 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 38824 21786
rect 1104 21712 38824 21734
rect 31386 21632 31392 21684
rect 31444 21672 31450 21684
rect 32677 21675 32735 21681
rect 32677 21672 32689 21675
rect 31444 21644 32689 21672
rect 31444 21632 31450 21644
rect 31680 21400 31708 21644
rect 32677 21641 32689 21644
rect 32723 21672 32735 21675
rect 32766 21672 32772 21684
rect 32723 21644 32772 21672
rect 32723 21641 32735 21644
rect 32677 21635 32735 21641
rect 32766 21632 32772 21644
rect 32824 21632 32830 21684
rect 37461 21675 37519 21681
rect 37461 21641 37473 21675
rect 37507 21672 37519 21675
rect 37550 21672 37556 21684
rect 37507 21644 37556 21672
rect 37507 21641 37519 21644
rect 37461 21635 37519 21641
rect 37550 21632 37556 21644
rect 37608 21632 37614 21684
rect 32306 21564 32312 21616
rect 32364 21604 32370 21616
rect 34606 21604 34612 21616
rect 32364 21576 34612 21604
rect 32364 21564 32370 21576
rect 34606 21564 34612 21576
rect 34664 21564 34670 21616
rect 37182 21604 37188 21616
rect 35176 21576 37188 21604
rect 32030 21496 32036 21548
rect 32088 21536 32094 21548
rect 32125 21539 32183 21545
rect 32125 21536 32137 21539
rect 32088 21508 32137 21536
rect 32088 21496 32094 21508
rect 32125 21505 32137 21508
rect 32171 21505 32183 21539
rect 32125 21499 32183 21505
rect 34333 21539 34391 21545
rect 34333 21505 34345 21539
rect 34379 21536 34391 21539
rect 35176 21536 35204 21576
rect 37182 21564 37188 21576
rect 37240 21564 37246 21616
rect 34379 21508 35204 21536
rect 34379 21505 34391 21508
rect 34333 21499 34391 21505
rect 35250 21496 35256 21548
rect 35308 21536 35314 21548
rect 38470 21536 38476 21548
rect 35308 21508 38476 21536
rect 35308 21496 35314 21508
rect 38470 21496 38476 21508
rect 38528 21496 38534 21548
rect 31754 21428 31760 21480
rect 31812 21468 31818 21480
rect 31849 21471 31907 21477
rect 31849 21468 31861 21471
rect 31812 21440 31861 21468
rect 31812 21428 31818 21440
rect 31849 21437 31861 21440
rect 31895 21437 31907 21471
rect 31849 21431 31907 21437
rect 31941 21471 31999 21477
rect 31941 21437 31953 21471
rect 31987 21437 31999 21471
rect 32214 21468 32220 21480
rect 32175 21440 32220 21468
rect 31941 21431 31999 21437
rect 31956 21400 31984 21431
rect 32214 21428 32220 21440
rect 32272 21428 32278 21480
rect 32490 21428 32496 21480
rect 32548 21468 32554 21480
rect 32861 21471 32919 21477
rect 32861 21468 32873 21471
rect 32548 21440 32873 21468
rect 32548 21428 32554 21440
rect 32861 21437 32873 21440
rect 32907 21437 32919 21471
rect 37274 21468 37280 21480
rect 37235 21440 37280 21468
rect 32861 21431 32919 21437
rect 37274 21428 37280 21440
rect 37332 21428 37338 21480
rect 37918 21468 37924 21480
rect 37879 21440 37924 21468
rect 37918 21428 37924 21440
rect 37976 21428 37982 21480
rect 34054 21400 34060 21412
rect 31680 21372 31800 21400
rect 31956 21372 34060 21400
rect 31772 21344 31800 21372
rect 34054 21360 34060 21372
rect 34112 21360 34118 21412
rect 34149 21403 34207 21409
rect 34149 21369 34161 21403
rect 34195 21400 34207 21403
rect 36722 21400 36728 21412
rect 34195 21372 36728 21400
rect 34195 21369 34207 21372
rect 34149 21363 34207 21369
rect 36722 21360 36728 21372
rect 36780 21360 36786 21412
rect 31478 21292 31484 21344
rect 31536 21332 31542 21344
rect 31665 21335 31723 21341
rect 31665 21332 31677 21335
rect 31536 21304 31677 21332
rect 31536 21292 31542 21304
rect 31665 21301 31677 21304
rect 31711 21301 31723 21335
rect 31665 21295 31723 21301
rect 31754 21292 31760 21344
rect 31812 21292 31818 21344
rect 33318 21292 33324 21344
rect 33376 21332 33382 21344
rect 34330 21332 34336 21344
rect 33376 21304 34336 21332
rect 33376 21292 33382 21304
rect 34330 21292 34336 21304
rect 34388 21292 34394 21344
rect 1104 21242 38824 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 38824 21242
rect 1104 21168 38824 21190
rect 35894 21128 35900 21140
rect 30576 21100 35900 21128
rect 1854 20992 1860 21004
rect 1815 20964 1860 20992
rect 1854 20952 1860 20964
rect 1912 20952 1918 21004
rect 30576 21001 30604 21100
rect 35894 21088 35900 21100
rect 35952 21088 35958 21140
rect 31662 21060 31668 21072
rect 31496 21032 31668 21060
rect 30469 20995 30527 21001
rect 30469 20961 30481 20995
rect 30515 20961 30527 20995
rect 30469 20955 30527 20961
rect 30561 20995 30619 21001
rect 30561 20961 30573 20995
rect 30607 20961 30619 20995
rect 30561 20955 30619 20961
rect 30837 20995 30895 21001
rect 30837 20961 30849 20995
rect 30883 20992 30895 20995
rect 31386 20992 31392 21004
rect 30883 20964 31392 20992
rect 30883 20961 30895 20964
rect 30837 20955 30895 20961
rect 30484 20924 30512 20955
rect 31386 20952 31392 20964
rect 31444 20952 31450 21004
rect 31496 21001 31524 21032
rect 31662 21020 31668 21032
rect 31720 21020 31726 21072
rect 32306 21060 32312 21072
rect 31772 21032 32312 21060
rect 31481 20995 31539 21001
rect 31481 20961 31493 20995
rect 31527 20961 31539 20995
rect 31481 20955 31539 20961
rect 31573 20995 31631 21001
rect 31573 20961 31585 20995
rect 31619 20992 31631 20995
rect 31772 20992 31800 21032
rect 32306 21020 32312 21032
rect 32364 21020 32370 21072
rect 33134 21020 33140 21072
rect 33192 21060 33198 21072
rect 33290 21063 33348 21069
rect 33290 21060 33302 21063
rect 33192 21032 33302 21060
rect 33192 21020 33198 21032
rect 33290 21029 33302 21032
rect 33336 21029 33348 21063
rect 33290 21023 33348 21029
rect 35360 21032 36400 21060
rect 35360 21004 35388 21032
rect 31619 20964 31800 20992
rect 31849 20995 31907 21001
rect 31619 20961 31631 20964
rect 31573 20955 31631 20961
rect 31849 20961 31861 20995
rect 31895 20992 31907 20995
rect 32214 20992 32220 21004
rect 31895 20964 32220 20992
rect 31895 20961 31907 20964
rect 31849 20955 31907 20961
rect 32214 20952 32220 20964
rect 32272 20952 32278 21004
rect 32490 20992 32496 21004
rect 32324 20964 32496 20992
rect 31018 20924 31024 20936
rect 30484 20896 31024 20924
rect 31018 20884 31024 20896
rect 31076 20884 31082 20936
rect 32324 20868 32352 20964
rect 32490 20952 32496 20964
rect 32548 20952 32554 21004
rect 32766 20952 32772 21004
rect 32824 20992 32830 21004
rect 33045 20995 33103 21001
rect 33045 20992 33057 20995
rect 32824 20964 33057 20992
rect 32824 20952 32830 20964
rect 33045 20961 33057 20964
rect 33091 20961 33103 20995
rect 33045 20955 33103 20961
rect 35069 20995 35127 21001
rect 35069 20961 35081 20995
rect 35115 20961 35127 20995
rect 35069 20955 35127 20961
rect 35161 20995 35219 21001
rect 35161 20961 35173 20995
rect 35207 20961 35219 20995
rect 35342 20992 35348 21004
rect 35255 20964 35348 20992
rect 35161 20955 35219 20961
rect 30466 20816 30472 20868
rect 30524 20856 30530 20868
rect 31297 20859 31355 20865
rect 31297 20856 31309 20859
rect 30524 20828 31309 20856
rect 30524 20816 30530 20828
rect 31297 20825 31309 20828
rect 31343 20825 31355 20859
rect 31297 20819 31355 20825
rect 31386 20816 31392 20868
rect 31444 20856 31450 20868
rect 32214 20856 32220 20868
rect 31444 20828 32220 20856
rect 31444 20816 31450 20828
rect 32214 20816 32220 20828
rect 32272 20816 32278 20868
rect 32306 20816 32312 20868
rect 32364 20816 32370 20868
rect 1949 20791 2007 20797
rect 1949 20757 1961 20791
rect 1995 20788 2007 20791
rect 17126 20788 17132 20800
rect 1995 20760 17132 20788
rect 1995 20757 2007 20760
rect 1949 20751 2007 20757
rect 17126 20748 17132 20760
rect 17184 20748 17190 20800
rect 30282 20788 30288 20800
rect 30243 20760 30288 20788
rect 30282 20748 30288 20760
rect 30340 20748 30346 20800
rect 30745 20791 30803 20797
rect 30745 20757 30757 20791
rect 30791 20788 30803 20791
rect 31018 20788 31024 20800
rect 30791 20760 31024 20788
rect 30791 20757 30803 20760
rect 30745 20751 30803 20757
rect 31018 20748 31024 20760
rect 31076 20748 31082 20800
rect 31754 20748 31760 20800
rect 31812 20788 31818 20800
rect 31812 20760 31857 20788
rect 31812 20748 31818 20760
rect 32490 20748 32496 20800
rect 32548 20788 32554 20800
rect 32950 20788 32956 20800
rect 32548 20760 32956 20788
rect 32548 20748 32554 20760
rect 32950 20748 32956 20760
rect 33008 20748 33014 20800
rect 34238 20748 34244 20800
rect 34296 20788 34302 20800
rect 34425 20791 34483 20797
rect 34425 20788 34437 20791
rect 34296 20760 34437 20788
rect 34296 20748 34302 20760
rect 34425 20757 34437 20760
rect 34471 20757 34483 20791
rect 34425 20751 34483 20757
rect 34514 20748 34520 20800
rect 34572 20788 34578 20800
rect 34885 20791 34943 20797
rect 34885 20788 34897 20791
rect 34572 20760 34897 20788
rect 34572 20748 34578 20760
rect 34885 20757 34897 20760
rect 34931 20757 34943 20791
rect 35084 20788 35112 20955
rect 35176 20924 35204 20955
rect 35342 20952 35348 20964
rect 35400 20952 35406 21004
rect 35434 20952 35440 21004
rect 35492 20992 35498 21004
rect 36081 20995 36139 21001
rect 35492 20964 35537 20992
rect 35492 20952 35498 20964
rect 36081 20961 36093 20995
rect 36127 20961 36139 20995
rect 36081 20955 36139 20961
rect 36096 20924 36124 20955
rect 36170 20952 36176 21004
rect 36228 20992 36234 21004
rect 36372 21001 36400 21032
rect 36357 20995 36415 21001
rect 36228 20964 36273 20992
rect 36228 20952 36234 20964
rect 36357 20961 36369 20995
rect 36403 20961 36415 20995
rect 36357 20955 36415 20961
rect 36449 20995 36507 21001
rect 36449 20961 36461 20995
rect 36495 20992 36507 20995
rect 36906 20992 36912 21004
rect 36495 20964 36912 20992
rect 36495 20961 36507 20964
rect 36449 20955 36507 20961
rect 36906 20952 36912 20964
rect 36964 20952 36970 21004
rect 37182 20992 37188 21004
rect 37143 20964 37188 20992
rect 37182 20952 37188 20964
rect 37240 20952 37246 21004
rect 38470 20924 38476 20936
rect 35176 20896 36032 20924
rect 36096 20896 38476 20924
rect 35894 20856 35900 20868
rect 35855 20828 35900 20856
rect 35894 20816 35900 20828
rect 35952 20816 35958 20868
rect 36004 20856 36032 20896
rect 38470 20884 38476 20896
rect 38528 20884 38534 20936
rect 36170 20856 36176 20868
rect 36004 20828 36176 20856
rect 36170 20816 36176 20828
rect 36228 20816 36234 20868
rect 37458 20788 37464 20800
rect 35084 20760 37464 20788
rect 34885 20751 34943 20757
rect 37458 20748 37464 20760
rect 37516 20748 37522 20800
rect 1104 20698 38824 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 38824 20698
rect 1104 20624 38824 20646
rect 27154 20544 27160 20596
rect 27212 20584 27218 20596
rect 27249 20587 27307 20593
rect 27249 20584 27261 20587
rect 27212 20556 27261 20584
rect 27212 20544 27218 20556
rect 27249 20553 27261 20556
rect 27295 20584 27307 20587
rect 27430 20584 27436 20596
rect 27295 20556 27436 20584
rect 27295 20553 27307 20556
rect 27249 20547 27307 20553
rect 27430 20544 27436 20556
rect 27488 20544 27494 20596
rect 34514 20584 34520 20596
rect 31036 20556 34520 20584
rect 28077 20519 28135 20525
rect 28077 20485 28089 20519
rect 28123 20516 28135 20519
rect 29546 20516 29552 20528
rect 28123 20488 29552 20516
rect 28123 20485 28135 20488
rect 28077 20479 28135 20485
rect 29546 20476 29552 20488
rect 29604 20476 29610 20528
rect 30926 20516 30932 20528
rect 30852 20488 30932 20516
rect 27430 20380 27436 20392
rect 27391 20352 27436 20380
rect 27430 20340 27436 20352
rect 27488 20340 27494 20392
rect 27890 20380 27896 20392
rect 27803 20352 27896 20380
rect 27890 20340 27896 20352
rect 27948 20380 27954 20392
rect 27948 20352 28396 20380
rect 27948 20340 27954 20352
rect 1854 20312 1860 20324
rect 1815 20284 1860 20312
rect 1854 20272 1860 20284
rect 1912 20272 1918 20324
rect 28368 20312 28396 20352
rect 28534 20340 28540 20392
rect 28592 20380 28598 20392
rect 30852 20389 30880 20488
rect 30926 20476 30932 20488
rect 30984 20476 30990 20528
rect 30837 20383 30895 20389
rect 28592 20352 28856 20380
rect 28592 20340 28598 20352
rect 28828 20324 28856 20352
rect 30837 20349 30849 20383
rect 30883 20349 30895 20383
rect 30837 20343 30895 20349
rect 30929 20383 30987 20389
rect 30929 20349 30941 20383
rect 30975 20380 30987 20383
rect 31036 20380 31064 20556
rect 34514 20544 34520 20556
rect 34572 20544 34578 20596
rect 31113 20519 31171 20525
rect 31113 20485 31125 20519
rect 31159 20516 31171 20519
rect 31202 20516 31208 20528
rect 31159 20488 31208 20516
rect 31159 20485 31171 20488
rect 31113 20479 31171 20485
rect 31202 20476 31208 20488
rect 31260 20476 31266 20528
rect 33226 20476 33232 20528
rect 33284 20516 33290 20528
rect 33689 20519 33747 20525
rect 33689 20516 33701 20519
rect 33284 20488 33701 20516
rect 33284 20476 33290 20488
rect 33689 20485 33701 20488
rect 33735 20485 33747 20519
rect 33689 20479 33747 20485
rect 35989 20519 36047 20525
rect 35989 20485 36001 20519
rect 36035 20516 36047 20519
rect 36078 20516 36084 20528
rect 36035 20488 36084 20516
rect 36035 20485 36047 20488
rect 35989 20479 36047 20485
rect 36078 20476 36084 20488
rect 36136 20476 36142 20528
rect 31662 20448 31668 20460
rect 31623 20420 31668 20448
rect 31662 20408 31668 20420
rect 31720 20408 31726 20460
rect 34238 20448 34244 20460
rect 33244 20420 34244 20448
rect 30975 20352 31064 20380
rect 31205 20383 31263 20389
rect 30975 20349 30987 20352
rect 30929 20343 30987 20349
rect 31205 20349 31217 20383
rect 31251 20380 31263 20383
rect 31386 20380 31392 20392
rect 31251 20352 31392 20380
rect 31251 20349 31263 20352
rect 31205 20343 31263 20349
rect 31386 20340 31392 20352
rect 31444 20340 31450 20392
rect 28629 20315 28687 20321
rect 28629 20312 28641 20315
rect 28368 20284 28641 20312
rect 28629 20281 28641 20284
rect 28675 20281 28687 20315
rect 28810 20312 28816 20324
rect 28771 20284 28816 20312
rect 28629 20275 28687 20281
rect 1949 20247 2007 20253
rect 1949 20213 1961 20247
rect 1995 20244 2007 20247
rect 17218 20244 17224 20256
rect 1995 20216 17224 20244
rect 1995 20213 2007 20216
rect 1949 20207 2007 20213
rect 17218 20204 17224 20216
rect 17276 20204 17282 20256
rect 23566 20204 23572 20256
rect 23624 20244 23630 20256
rect 25498 20244 25504 20256
rect 23624 20216 25504 20244
rect 23624 20204 23630 20216
rect 25498 20204 25504 20216
rect 25556 20204 25562 20256
rect 28644 20244 28672 20275
rect 28810 20272 28816 20284
rect 28868 20272 28874 20324
rect 31680 20312 31708 20408
rect 33244 20392 33272 20420
rect 34238 20408 34244 20420
rect 34296 20408 34302 20460
rect 36170 20448 36176 20460
rect 34532 20420 36176 20448
rect 31938 20389 31944 20392
rect 31932 20343 31944 20389
rect 31996 20380 32002 20392
rect 31996 20352 32032 20380
rect 31938 20340 31944 20343
rect 31996 20340 32002 20352
rect 33226 20340 33232 20392
rect 33284 20340 33290 20392
rect 34532 20389 34560 20420
rect 36170 20408 36176 20420
rect 36228 20408 36234 20460
rect 33505 20383 33563 20389
rect 33505 20349 33517 20383
rect 33551 20349 33563 20383
rect 33505 20343 33563 20349
rect 34425 20383 34483 20389
rect 34425 20349 34437 20383
rect 34471 20349 34483 20383
rect 34425 20343 34483 20349
rect 34517 20383 34575 20389
rect 34517 20349 34529 20383
rect 34563 20349 34575 20383
rect 34517 20343 34575 20349
rect 34660 20383 34718 20389
rect 34660 20349 34672 20383
rect 34706 20349 34718 20383
rect 34790 20380 34796 20392
rect 34751 20352 34796 20380
rect 34660 20343 34718 20349
rect 32214 20312 32220 20324
rect 31680 20284 32220 20312
rect 32214 20272 32220 20284
rect 32272 20272 32278 20324
rect 29454 20244 29460 20256
rect 28644 20216 29460 20244
rect 29454 20204 29460 20216
rect 29512 20204 29518 20256
rect 30374 20204 30380 20256
rect 30432 20244 30438 20256
rect 30653 20247 30711 20253
rect 30653 20244 30665 20247
rect 30432 20216 30665 20244
rect 30432 20204 30438 20216
rect 30653 20213 30665 20216
rect 30699 20213 30711 20247
rect 30653 20207 30711 20213
rect 31386 20204 31392 20256
rect 31444 20244 31450 20256
rect 31662 20244 31668 20256
rect 31444 20216 31668 20244
rect 31444 20204 31450 20216
rect 31662 20204 31668 20216
rect 31720 20204 31726 20256
rect 31938 20204 31944 20256
rect 31996 20244 32002 20256
rect 32306 20244 32312 20256
rect 31996 20216 32312 20244
rect 31996 20204 32002 20216
rect 32306 20204 32312 20216
rect 32364 20204 32370 20256
rect 32766 20204 32772 20256
rect 32824 20244 32830 20256
rect 33045 20247 33103 20253
rect 33045 20244 33057 20247
rect 32824 20216 33057 20244
rect 32824 20204 32830 20216
rect 33045 20213 33057 20216
rect 33091 20213 33103 20247
rect 33045 20207 33103 20213
rect 33318 20204 33324 20256
rect 33376 20244 33382 20256
rect 33520 20244 33548 20343
rect 34238 20244 34244 20256
rect 33376 20216 33548 20244
rect 34199 20216 34244 20244
rect 33376 20204 33382 20216
rect 34238 20204 34244 20216
rect 34296 20204 34302 20256
rect 34440 20244 34468 20343
rect 34675 20312 34703 20343
rect 34790 20340 34796 20352
rect 34848 20340 34854 20392
rect 35805 20383 35863 20389
rect 35805 20349 35817 20383
rect 35851 20380 35863 20383
rect 36078 20380 36084 20392
rect 35851 20352 36084 20380
rect 35851 20349 35863 20352
rect 35805 20343 35863 20349
rect 36078 20340 36084 20352
rect 36136 20380 36142 20392
rect 36722 20380 36728 20392
rect 36136 20352 36728 20380
rect 36136 20340 36142 20352
rect 36722 20340 36728 20352
rect 36780 20340 36786 20392
rect 37918 20380 37924 20392
rect 37879 20352 37924 20380
rect 37918 20340 37924 20352
rect 37976 20340 37982 20392
rect 35342 20312 35348 20324
rect 34675 20284 35348 20312
rect 35342 20272 35348 20284
rect 35400 20272 35406 20324
rect 34790 20244 34796 20256
rect 34440 20216 34796 20244
rect 34790 20204 34796 20216
rect 34848 20204 34854 20256
rect 1104 20154 38824 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 38824 20154
rect 1104 20080 38824 20102
rect 34885 20043 34943 20049
rect 34885 20040 34897 20043
rect 28828 20012 34897 20040
rect 26050 19972 26056 19984
rect 25792 19944 26056 19972
rect 25792 19916 25820 19944
rect 26050 19932 26056 19944
rect 26108 19932 26114 19984
rect 25685 19907 25743 19913
rect 25685 19873 25697 19907
rect 25731 19904 25743 19907
rect 25774 19904 25780 19916
rect 25731 19876 25780 19904
rect 25731 19873 25743 19876
rect 25685 19867 25743 19873
rect 25774 19864 25780 19876
rect 25832 19864 25838 19916
rect 25961 19907 26019 19913
rect 25961 19873 25973 19907
rect 26007 19904 26019 19907
rect 27614 19904 27620 19916
rect 26007 19876 27620 19904
rect 26007 19873 26019 19876
rect 25961 19867 26019 19873
rect 27614 19864 27620 19876
rect 27672 19864 27678 19916
rect 27890 19904 27896 19916
rect 27851 19876 27896 19904
rect 27890 19864 27896 19876
rect 27948 19864 27954 19916
rect 28258 19864 28264 19916
rect 28316 19904 28322 19916
rect 28828 19913 28856 20012
rect 34885 20009 34897 20012
rect 34931 20009 34943 20043
rect 34885 20003 34943 20009
rect 37369 20043 37427 20049
rect 37369 20009 37381 20043
rect 37415 20040 37427 20043
rect 37826 20040 37832 20052
rect 37415 20012 37832 20040
rect 37415 20009 37427 20012
rect 37369 20003 37427 20009
rect 37826 20000 37832 20012
rect 37884 20000 37890 20052
rect 29638 19972 29644 19984
rect 29104 19944 29644 19972
rect 29104 19913 29132 19944
rect 29638 19932 29644 19944
rect 29696 19932 29702 19984
rect 34238 19972 34244 19984
rect 29840 19944 34244 19972
rect 28721 19907 28779 19913
rect 28721 19904 28733 19907
rect 28316 19876 28733 19904
rect 28316 19864 28322 19876
rect 28721 19873 28733 19876
rect 28767 19873 28779 19907
rect 28721 19867 28779 19873
rect 28813 19907 28871 19913
rect 28813 19873 28825 19907
rect 28859 19873 28871 19907
rect 29089 19907 29147 19913
rect 29089 19904 29101 19907
rect 28813 19867 28871 19873
rect 28920 19876 29101 19904
rect 26421 19839 26479 19845
rect 26421 19805 26433 19839
rect 26467 19836 26479 19839
rect 26970 19836 26976 19848
rect 26467 19808 26976 19836
rect 26467 19805 26479 19808
rect 26421 19799 26479 19805
rect 26970 19796 26976 19808
rect 27028 19796 27034 19848
rect 28920 19836 28948 19876
rect 29089 19873 29101 19876
rect 29135 19873 29147 19907
rect 29730 19904 29736 19916
rect 29691 19876 29736 19904
rect 29089 19867 29147 19873
rect 29730 19864 29736 19876
rect 29788 19864 29794 19916
rect 29840 19913 29868 19944
rect 34238 19932 34244 19944
rect 34296 19932 34302 19984
rect 34514 19932 34520 19984
rect 34572 19932 34578 19984
rect 36173 19975 36231 19981
rect 35084 19944 36124 19972
rect 29825 19907 29883 19913
rect 29825 19873 29837 19907
rect 29871 19873 29883 19907
rect 29825 19867 29883 19873
rect 30101 19907 30159 19913
rect 30101 19873 30113 19907
rect 30147 19873 30159 19907
rect 30742 19904 30748 19916
rect 30703 19876 30748 19904
rect 30101 19867 30159 19873
rect 28092 19808 28948 19836
rect 25777 19771 25835 19777
rect 25777 19737 25789 19771
rect 25823 19768 25835 19771
rect 27522 19768 27528 19780
rect 25823 19740 27528 19768
rect 25823 19737 25835 19740
rect 25777 19731 25835 19737
rect 27522 19728 27528 19740
rect 27580 19728 27586 19780
rect 28092 19777 28120 19808
rect 28994 19796 29000 19848
rect 29052 19836 29058 19848
rect 29549 19839 29607 19845
rect 29549 19836 29561 19839
rect 29052 19808 29561 19836
rect 29052 19796 29058 19808
rect 29549 19805 29561 19808
rect 29595 19805 29607 19839
rect 29549 19799 29607 19805
rect 29638 19796 29644 19848
rect 29696 19836 29702 19848
rect 30116 19836 30144 19867
rect 30742 19864 30748 19876
rect 30800 19864 30806 19916
rect 30837 19907 30895 19913
rect 30837 19873 30849 19907
rect 30883 19904 30895 19907
rect 30926 19904 30932 19916
rect 30883 19876 30932 19904
rect 30883 19873 30895 19876
rect 30837 19867 30895 19873
rect 30926 19864 30932 19876
rect 30984 19864 30990 19916
rect 31113 19907 31171 19913
rect 31113 19873 31125 19907
rect 31159 19904 31171 19907
rect 31386 19904 31392 19916
rect 31159 19876 31392 19904
rect 31159 19873 31171 19876
rect 31113 19867 31171 19873
rect 31386 19864 31392 19876
rect 31444 19864 31450 19916
rect 31573 19907 31631 19913
rect 31573 19873 31585 19907
rect 31619 19873 31631 19907
rect 31573 19867 31631 19873
rect 29696 19808 30144 19836
rect 29696 19796 29702 19808
rect 28077 19771 28135 19777
rect 28077 19737 28089 19771
rect 28123 19737 28135 19771
rect 28077 19731 28135 19737
rect 28902 19728 28908 19780
rect 28960 19768 28966 19780
rect 30009 19771 30067 19777
rect 30009 19768 30021 19771
rect 28960 19740 30021 19768
rect 28960 19728 28966 19740
rect 30009 19737 30021 19740
rect 30055 19737 30067 19771
rect 31588 19768 31616 19867
rect 32214 19864 32220 19916
rect 32272 19904 32278 19916
rect 33045 19907 33103 19913
rect 33045 19904 33057 19907
rect 32272 19876 33057 19904
rect 32272 19864 32278 19876
rect 33045 19873 33057 19876
rect 33091 19873 33103 19907
rect 33045 19867 33103 19873
rect 33312 19907 33370 19913
rect 33312 19873 33324 19907
rect 33358 19904 33370 19907
rect 33870 19904 33876 19916
rect 33358 19876 33876 19904
rect 33358 19873 33370 19876
rect 33312 19867 33370 19873
rect 33870 19864 33876 19876
rect 33928 19864 33934 19916
rect 34532 19904 34560 19932
rect 35084 19913 35112 19944
rect 34440 19876 34560 19904
rect 35069 19907 35127 19913
rect 30009 19731 30067 19737
rect 30116 19740 31616 19768
rect 28534 19700 28540 19712
rect 28495 19672 28540 19700
rect 28534 19660 28540 19672
rect 28592 19660 28598 19712
rect 28626 19660 28632 19712
rect 28684 19700 28690 19712
rect 28997 19703 29055 19709
rect 28997 19700 29009 19703
rect 28684 19672 29009 19700
rect 28684 19660 28690 19672
rect 28997 19669 29009 19672
rect 29043 19669 29055 19703
rect 28997 19663 29055 19669
rect 29454 19660 29460 19712
rect 29512 19700 29518 19712
rect 29730 19700 29736 19712
rect 29512 19672 29736 19700
rect 29512 19660 29518 19672
rect 29730 19660 29736 19672
rect 29788 19700 29794 19712
rect 30116 19700 30144 19740
rect 31662 19728 31668 19780
rect 31720 19768 31726 19780
rect 34440 19777 34468 19876
rect 35069 19873 35081 19907
rect 35115 19873 35127 19907
rect 35069 19867 35127 19873
rect 35161 19907 35219 19913
rect 35161 19873 35173 19907
rect 35207 19873 35219 19907
rect 35342 19904 35348 19916
rect 35303 19876 35348 19904
rect 35161 19867 35219 19873
rect 34514 19796 34520 19848
rect 34572 19836 34578 19848
rect 35176 19836 35204 19867
rect 35342 19864 35348 19876
rect 35400 19864 35406 19916
rect 35437 19907 35495 19913
rect 35437 19873 35449 19907
rect 35483 19904 35495 19907
rect 35802 19904 35808 19916
rect 35483 19876 35808 19904
rect 35483 19873 35495 19876
rect 35437 19867 35495 19873
rect 35802 19864 35808 19876
rect 35860 19864 35866 19916
rect 35894 19864 35900 19916
rect 35952 19904 35958 19916
rect 35989 19907 36047 19913
rect 35989 19904 36001 19907
rect 35952 19876 36001 19904
rect 35952 19864 35958 19876
rect 35989 19873 36001 19876
rect 36035 19873 36047 19907
rect 35989 19867 36047 19873
rect 34572 19808 35204 19836
rect 36096 19836 36124 19944
rect 36173 19941 36185 19975
rect 36219 19972 36231 19975
rect 36538 19972 36544 19984
rect 36219 19944 36544 19972
rect 36219 19941 36231 19944
rect 36173 19935 36231 19941
rect 36538 19932 36544 19944
rect 36596 19932 36602 19984
rect 37182 19904 37188 19916
rect 37143 19876 37188 19904
rect 37182 19864 37188 19876
rect 37240 19864 37246 19916
rect 37826 19836 37832 19848
rect 36096 19808 37832 19836
rect 34572 19796 34578 19808
rect 37826 19796 37832 19808
rect 37884 19796 37890 19848
rect 31757 19771 31815 19777
rect 31757 19768 31769 19771
rect 31720 19740 31769 19768
rect 31720 19728 31726 19740
rect 31757 19737 31769 19740
rect 31803 19737 31815 19771
rect 31757 19731 31815 19737
rect 34425 19771 34483 19777
rect 34425 19737 34437 19771
rect 34471 19737 34483 19771
rect 34425 19731 34483 19737
rect 30558 19700 30564 19712
rect 29788 19672 30144 19700
rect 30519 19672 30564 19700
rect 29788 19660 29794 19672
rect 30558 19660 30564 19672
rect 30616 19660 30622 19712
rect 31018 19700 31024 19712
rect 30979 19672 31024 19700
rect 31018 19660 31024 19672
rect 31076 19660 31082 19712
rect 32858 19660 32864 19712
rect 32916 19700 32922 19712
rect 33226 19700 33232 19712
rect 32916 19672 33232 19700
rect 32916 19660 32922 19672
rect 33226 19660 33232 19672
rect 33284 19660 33290 19712
rect 1104 19610 38824 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 38824 19610
rect 1104 19536 38824 19558
rect 24121 19499 24179 19505
rect 24121 19465 24133 19499
rect 24167 19496 24179 19499
rect 26786 19496 26792 19508
rect 24167 19468 26792 19496
rect 24167 19465 24179 19468
rect 24121 19459 24179 19465
rect 26786 19456 26792 19468
rect 26844 19456 26850 19508
rect 27062 19496 27068 19508
rect 27023 19468 27068 19496
rect 27062 19456 27068 19468
rect 27120 19456 27126 19508
rect 27430 19456 27436 19508
rect 27488 19496 27494 19508
rect 31938 19496 31944 19508
rect 27488 19468 31944 19496
rect 27488 19456 27494 19468
rect 31938 19456 31944 19468
rect 31996 19456 32002 19508
rect 31662 19388 31668 19440
rect 31720 19428 31726 19440
rect 31849 19431 31907 19437
rect 31849 19428 31861 19431
rect 31720 19400 31861 19428
rect 31720 19388 31726 19400
rect 31849 19397 31861 19400
rect 31895 19428 31907 19431
rect 32122 19428 32128 19440
rect 31895 19400 32128 19428
rect 31895 19397 31907 19400
rect 31849 19391 31907 19397
rect 32122 19388 32128 19400
rect 32180 19388 32186 19440
rect 35066 19388 35072 19440
rect 35124 19428 35130 19440
rect 36078 19428 36084 19440
rect 35124 19400 36084 19428
rect 35124 19388 35130 19400
rect 26605 19363 26663 19369
rect 25976 19332 26280 19360
rect 1854 19292 1860 19304
rect 1815 19264 1860 19292
rect 1854 19252 1860 19264
rect 1912 19252 1918 19304
rect 23937 19295 23995 19301
rect 23937 19261 23949 19295
rect 23983 19261 23995 19295
rect 24118 19292 24124 19304
rect 24079 19264 24124 19292
rect 23937 19255 23995 19261
rect 2041 19227 2099 19233
rect 2041 19193 2053 19227
rect 2087 19224 2099 19227
rect 9122 19224 9128 19236
rect 2087 19196 9128 19224
rect 2087 19193 2099 19196
rect 2041 19187 2099 19193
rect 9122 19184 9128 19196
rect 9180 19184 9186 19236
rect 23952 19224 23980 19255
rect 24118 19252 24124 19264
rect 24176 19252 24182 19304
rect 25976 19292 26004 19332
rect 26252 19304 26280 19332
rect 26605 19329 26617 19363
rect 26651 19360 26663 19363
rect 27338 19360 27344 19372
rect 26651 19332 27344 19360
rect 26651 19329 26663 19332
rect 26605 19323 26663 19329
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 32214 19320 32220 19372
rect 32272 19360 32278 19372
rect 32309 19363 32367 19369
rect 32309 19360 32321 19363
rect 32272 19332 32321 19360
rect 32272 19320 32278 19332
rect 32309 19329 32321 19332
rect 32355 19329 32367 19363
rect 32309 19323 32367 19329
rect 34348 19332 34928 19360
rect 26142 19292 26148 19304
rect 25792 19264 26004 19292
rect 26103 19264 26148 19292
rect 25792 19224 25820 19264
rect 26142 19252 26148 19264
rect 26200 19252 26206 19304
rect 26234 19252 26240 19304
rect 26292 19252 26298 19304
rect 26970 19292 26976 19304
rect 26931 19264 26976 19292
rect 26970 19252 26976 19264
rect 27028 19252 27034 19304
rect 30098 19252 30104 19304
rect 30156 19292 30162 19304
rect 30469 19295 30527 19301
rect 30469 19292 30481 19295
rect 30156 19264 30481 19292
rect 30156 19252 30162 19264
rect 30469 19261 30481 19264
rect 30515 19261 30527 19295
rect 30469 19255 30527 19261
rect 30736 19295 30794 19301
rect 30736 19261 30748 19295
rect 30782 19292 30794 19295
rect 31846 19292 31852 19304
rect 30782 19264 31852 19292
rect 30782 19261 30794 19264
rect 30736 19255 30794 19261
rect 31846 19252 31852 19264
rect 31904 19252 31910 19304
rect 34348 19301 34376 19332
rect 34514 19301 34520 19304
rect 34149 19295 34207 19301
rect 34149 19292 34161 19295
rect 32508 19264 34161 19292
rect 25958 19224 25964 19236
rect 23952 19196 25820 19224
rect 25919 19196 25964 19224
rect 25958 19184 25964 19196
rect 26016 19184 26022 19236
rect 26050 19184 26056 19236
rect 26108 19224 26114 19236
rect 27801 19227 27859 19233
rect 27801 19224 27813 19227
rect 26108 19196 27813 19224
rect 26108 19184 26114 19196
rect 27801 19193 27813 19196
rect 27847 19193 27859 19227
rect 27801 19187 27859 19193
rect 27890 19184 27896 19236
rect 27948 19224 27954 19236
rect 27948 19196 28994 19224
rect 27948 19184 27954 19196
rect 24305 19159 24363 19165
rect 24305 19125 24317 19159
rect 24351 19156 24363 19159
rect 28442 19156 28448 19168
rect 24351 19128 28448 19156
rect 24351 19125 24363 19128
rect 24305 19119 24363 19125
rect 28442 19116 28448 19128
rect 28500 19116 28506 19168
rect 28966 19156 28994 19196
rect 29454 19184 29460 19236
rect 29512 19224 29518 19236
rect 32508 19224 32536 19264
rect 34149 19261 34161 19264
rect 34195 19261 34207 19295
rect 34149 19255 34207 19261
rect 34336 19295 34394 19301
rect 34336 19261 34348 19295
rect 34382 19261 34394 19295
rect 34336 19255 34394 19261
rect 34471 19295 34520 19301
rect 34471 19261 34483 19295
rect 34517 19261 34520 19295
rect 34471 19255 34520 19261
rect 34514 19252 34520 19255
rect 34572 19252 34578 19304
rect 34609 19295 34667 19301
rect 34609 19261 34621 19295
rect 34655 19261 34667 19295
rect 34609 19255 34667 19261
rect 29512 19196 32536 19224
rect 32576 19227 32634 19233
rect 29512 19184 29518 19196
rect 32576 19193 32588 19227
rect 32622 19224 32634 19227
rect 33042 19224 33048 19236
rect 32622 19196 33048 19224
rect 32622 19193 32634 19196
rect 32576 19187 32634 19193
rect 33042 19184 33048 19196
rect 33100 19184 33106 19236
rect 34624 19224 34652 19255
rect 34698 19252 34704 19304
rect 34756 19292 34762 19304
rect 34900 19292 34928 19332
rect 35158 19292 35164 19304
rect 34756 19264 34801 19292
rect 34900 19264 35164 19292
rect 34756 19252 34762 19264
rect 35158 19252 35164 19264
rect 35216 19252 35222 19304
rect 35728 19301 35756 19400
rect 36078 19388 36084 19400
rect 36136 19388 36142 19440
rect 35713 19295 35771 19301
rect 35713 19261 35725 19295
rect 35759 19261 35771 19295
rect 37274 19292 37280 19304
rect 37235 19264 37280 19292
rect 35713 19255 35771 19261
rect 37274 19252 37280 19264
rect 37332 19252 37338 19304
rect 37918 19292 37924 19304
rect 37879 19264 37924 19292
rect 37918 19252 37924 19264
rect 37976 19252 37982 19304
rect 34624 19196 35388 19224
rect 35360 19168 35388 19196
rect 29273 19159 29331 19165
rect 29273 19156 29285 19159
rect 28966 19128 29285 19156
rect 29273 19125 29285 19128
rect 29319 19156 29331 19159
rect 31386 19156 31392 19168
rect 29319 19128 31392 19156
rect 29319 19125 29331 19128
rect 29273 19119 29331 19125
rect 31386 19116 31392 19128
rect 31444 19116 31450 19168
rect 33686 19156 33692 19168
rect 33647 19128 33692 19156
rect 33686 19116 33692 19128
rect 33744 19116 33750 19168
rect 35342 19116 35348 19168
rect 35400 19156 35406 19168
rect 35897 19159 35955 19165
rect 35897 19156 35909 19159
rect 35400 19128 35909 19156
rect 35400 19116 35406 19128
rect 35897 19125 35909 19128
rect 35943 19125 35955 19159
rect 35897 19119 35955 19125
rect 1104 19066 38824 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 38824 19066
rect 1104 18992 38824 19014
rect 24118 18912 24124 18964
rect 24176 18952 24182 18964
rect 28350 18952 28356 18964
rect 24176 18924 28356 18952
rect 24176 18912 24182 18924
rect 28350 18912 28356 18924
rect 28408 18912 28414 18964
rect 29273 18955 29331 18961
rect 29273 18921 29285 18955
rect 29319 18952 29331 18955
rect 30745 18955 30803 18961
rect 30745 18952 30757 18955
rect 29319 18924 30757 18952
rect 29319 18921 29331 18924
rect 29273 18915 29331 18921
rect 30745 18921 30757 18924
rect 30791 18952 30803 18955
rect 31754 18952 31760 18964
rect 30791 18924 31760 18952
rect 30791 18921 30803 18924
rect 30745 18915 30803 18921
rect 31754 18912 31760 18924
rect 31812 18912 31818 18964
rect 31938 18952 31944 18964
rect 31899 18924 31944 18952
rect 31938 18912 31944 18924
rect 31996 18912 32002 18964
rect 33134 18952 33140 18964
rect 32877 18924 33140 18952
rect 24305 18887 24363 18893
rect 24305 18853 24317 18887
rect 24351 18884 24363 18887
rect 25498 18884 25504 18896
rect 24351 18856 25504 18884
rect 24351 18853 24363 18856
rect 24305 18847 24363 18853
rect 25498 18844 25504 18856
rect 25556 18844 25562 18896
rect 29632 18887 29690 18893
rect 26436 18856 28580 18884
rect 1854 18816 1860 18828
rect 1815 18788 1860 18816
rect 1854 18776 1860 18788
rect 1912 18776 1918 18828
rect 26050 18816 26056 18828
rect 22066 18788 26056 18816
rect 1302 18708 1308 18760
rect 1360 18748 1366 18760
rect 22066 18748 22094 18788
rect 26050 18776 26056 18788
rect 26108 18776 26114 18828
rect 26326 18816 26332 18828
rect 26287 18788 26332 18816
rect 26326 18776 26332 18788
rect 26384 18776 26390 18828
rect 26436 18825 26464 18856
rect 26421 18819 26479 18825
rect 26421 18785 26433 18819
rect 26467 18785 26479 18819
rect 26421 18779 26479 18785
rect 26602 18776 26608 18828
rect 26660 18816 26666 18828
rect 26697 18819 26755 18825
rect 26697 18816 26709 18819
rect 26660 18788 26709 18816
rect 26660 18776 26666 18788
rect 26697 18785 26709 18788
rect 26743 18785 26755 18819
rect 26697 18779 26755 18785
rect 26878 18776 26884 18828
rect 26936 18816 26942 18828
rect 27801 18819 27859 18825
rect 27801 18816 27813 18819
rect 26936 18788 27813 18816
rect 26936 18776 26942 18788
rect 27801 18785 27813 18788
rect 27847 18785 27859 18819
rect 28074 18816 28080 18828
rect 28035 18788 28080 18816
rect 27801 18779 27859 18785
rect 28074 18776 28080 18788
rect 28132 18776 28138 18828
rect 28261 18819 28319 18825
rect 28261 18785 28273 18819
rect 28307 18785 28319 18819
rect 28442 18816 28448 18828
rect 28403 18788 28448 18816
rect 28261 18779 28319 18785
rect 24670 18748 24676 18760
rect 1360 18720 22094 18748
rect 24631 18720 24676 18748
rect 1360 18708 1366 18720
rect 24670 18708 24676 18720
rect 24728 18708 24734 18760
rect 25041 18751 25099 18757
rect 25041 18717 25053 18751
rect 25087 18748 25099 18751
rect 28276 18748 28304 18779
rect 28442 18776 28448 18788
rect 28500 18776 28506 18828
rect 28552 18816 28580 18856
rect 29632 18853 29644 18887
rect 29678 18884 29690 18887
rect 30466 18884 30472 18896
rect 29678 18856 30472 18884
rect 29678 18853 29690 18856
rect 29632 18847 29690 18853
rect 30466 18844 30472 18856
rect 30524 18844 30530 18896
rect 31481 18887 31539 18893
rect 31481 18853 31493 18887
rect 31527 18884 31539 18887
rect 32877 18884 32905 18924
rect 33134 18912 33140 18924
rect 33192 18912 33198 18964
rect 34146 18912 34152 18964
rect 34204 18952 34210 18964
rect 34425 18955 34483 18961
rect 34425 18952 34437 18955
rect 34204 18924 34437 18952
rect 34204 18912 34210 18924
rect 34425 18921 34437 18924
rect 34471 18921 34483 18955
rect 34425 18915 34483 18921
rect 34882 18912 34888 18964
rect 34940 18952 34946 18964
rect 36078 18952 36084 18964
rect 34940 18924 36084 18952
rect 34940 18912 34946 18924
rect 36078 18912 36084 18924
rect 36136 18912 36142 18964
rect 37369 18955 37427 18961
rect 37369 18921 37381 18955
rect 37415 18952 37427 18955
rect 37734 18952 37740 18964
rect 37415 18924 37740 18952
rect 37415 18921 37427 18924
rect 37369 18915 37427 18921
rect 37734 18912 37740 18924
rect 37792 18912 37798 18964
rect 31527 18856 32905 18884
rect 31527 18853 31539 18856
rect 31481 18847 31539 18853
rect 32950 18844 32956 18896
rect 33008 18884 33014 18896
rect 33290 18887 33348 18893
rect 33290 18884 33302 18887
rect 33008 18856 33302 18884
rect 33008 18844 33014 18856
rect 33290 18853 33302 18856
rect 33336 18853 33348 18887
rect 33290 18847 33348 18853
rect 34514 18844 34520 18896
rect 34572 18884 34578 18896
rect 34698 18884 34704 18896
rect 34572 18856 34704 18884
rect 34572 18844 34578 18856
rect 34698 18844 34704 18856
rect 34756 18884 34762 18896
rect 34756 18856 35204 18884
rect 34756 18844 34762 18856
rect 29914 18816 29920 18828
rect 28552 18788 29920 18816
rect 29914 18776 29920 18788
rect 29972 18776 29978 18828
rect 30190 18776 30196 18828
rect 30248 18816 30254 18828
rect 31297 18819 31355 18825
rect 30248 18788 30512 18816
rect 30248 18776 30254 18788
rect 30484 18760 30512 18788
rect 31297 18785 31309 18819
rect 31343 18785 31355 18819
rect 31297 18779 31355 18785
rect 25087 18720 26556 18748
rect 25087 18717 25099 18720
rect 25041 18711 25099 18717
rect 24470 18683 24528 18689
rect 24470 18649 24482 18683
rect 24516 18680 24528 18683
rect 26528 18680 26556 18720
rect 26896 18720 28304 18748
rect 28629 18751 28687 18757
rect 26896 18680 26924 18720
rect 28629 18717 28641 18751
rect 28675 18748 28687 18751
rect 28718 18748 28724 18760
rect 28675 18720 28724 18748
rect 28675 18717 28687 18720
rect 28629 18711 28687 18717
rect 28718 18708 28724 18720
rect 28776 18708 28782 18760
rect 29365 18751 29423 18757
rect 29365 18717 29377 18751
rect 29411 18717 29423 18751
rect 29365 18711 29423 18717
rect 24516 18652 26464 18680
rect 26528 18652 26924 18680
rect 24516 18649 24528 18652
rect 24470 18643 24528 18649
rect 26436 18624 26464 18652
rect 27154 18640 27160 18692
rect 27212 18680 27218 18692
rect 29380 18680 29408 18711
rect 30466 18708 30472 18760
rect 30524 18708 30530 18760
rect 27212 18652 29408 18680
rect 31312 18680 31340 18779
rect 31386 18776 31392 18828
rect 31444 18816 31450 18828
rect 32125 18819 32183 18825
rect 32125 18816 32137 18819
rect 31444 18788 32137 18816
rect 31444 18776 31450 18788
rect 32125 18785 32137 18788
rect 32171 18785 32183 18819
rect 32125 18779 32183 18785
rect 32214 18776 32220 18828
rect 32272 18816 32278 18828
rect 33045 18819 33103 18825
rect 33045 18816 33057 18819
rect 32272 18788 33057 18816
rect 32272 18776 32278 18788
rect 33045 18785 33057 18788
rect 33091 18785 33103 18819
rect 34054 18816 34060 18828
rect 33045 18779 33103 18785
rect 33153 18788 34060 18816
rect 32674 18708 32680 18760
rect 32732 18748 32738 18760
rect 33153 18748 33181 18788
rect 34054 18776 34060 18788
rect 34112 18776 34118 18828
rect 35176 18825 35204 18856
rect 35894 18844 35900 18896
rect 35952 18884 35958 18896
rect 35989 18887 36047 18893
rect 35989 18884 36001 18887
rect 35952 18856 36001 18884
rect 35952 18844 35958 18856
rect 35989 18853 36001 18856
rect 36035 18853 36047 18887
rect 36170 18884 36176 18896
rect 36131 18856 36176 18884
rect 35989 18847 36047 18853
rect 36170 18844 36176 18856
rect 36228 18844 36234 18896
rect 35069 18819 35127 18825
rect 35069 18785 35081 18819
rect 35115 18785 35127 18819
rect 35069 18779 35127 18785
rect 35161 18819 35219 18825
rect 35161 18785 35173 18819
rect 35207 18785 35219 18819
rect 35342 18816 35348 18828
rect 35303 18788 35348 18816
rect 35161 18779 35219 18785
rect 32732 18720 33181 18748
rect 35084 18748 35112 18779
rect 35342 18776 35348 18788
rect 35400 18776 35406 18828
rect 35437 18819 35495 18825
rect 35437 18785 35449 18819
rect 35483 18816 35495 18819
rect 35526 18816 35532 18828
rect 35483 18788 35532 18816
rect 35483 18785 35495 18788
rect 35437 18779 35495 18785
rect 35526 18776 35532 18788
rect 35584 18776 35590 18828
rect 37182 18816 37188 18828
rect 37143 18788 37188 18816
rect 37182 18776 37188 18788
rect 37240 18776 37246 18828
rect 36906 18748 36912 18760
rect 35084 18720 36912 18748
rect 32732 18708 32738 18720
rect 36906 18708 36912 18720
rect 36964 18708 36970 18760
rect 31312 18652 31524 18680
rect 27212 18640 27218 18652
rect 1949 18615 2007 18621
rect 1949 18581 1961 18615
rect 1995 18612 2007 18615
rect 18322 18612 18328 18624
rect 1995 18584 18328 18612
rect 1995 18581 2007 18584
rect 1949 18575 2007 18581
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 24581 18615 24639 18621
rect 24581 18581 24593 18615
rect 24627 18612 24639 18615
rect 24762 18612 24768 18624
rect 24627 18584 24768 18612
rect 24627 18581 24639 18584
rect 24581 18575 24639 18581
rect 24762 18572 24768 18584
rect 24820 18572 24826 18624
rect 24946 18572 24952 18624
rect 25004 18612 25010 18624
rect 26145 18615 26203 18621
rect 26145 18612 26157 18615
rect 25004 18584 26157 18612
rect 25004 18572 25010 18584
rect 26145 18581 26157 18584
rect 26191 18581 26203 18615
rect 26145 18575 26203 18581
rect 26418 18572 26424 18624
rect 26476 18572 26482 18624
rect 26602 18612 26608 18624
rect 26563 18584 26608 18612
rect 26602 18572 26608 18584
rect 26660 18572 26666 18624
rect 27246 18572 27252 18624
rect 27304 18612 27310 18624
rect 29273 18615 29331 18621
rect 29273 18612 29285 18615
rect 27304 18584 29285 18612
rect 27304 18572 27310 18584
rect 29273 18581 29285 18584
rect 29319 18581 29331 18615
rect 29380 18612 29408 18652
rect 30098 18612 30104 18624
rect 29380 18584 30104 18612
rect 29273 18575 29331 18581
rect 30098 18572 30104 18584
rect 30156 18572 30162 18624
rect 30926 18572 30932 18624
rect 30984 18612 30990 18624
rect 31386 18612 31392 18624
rect 30984 18584 31392 18612
rect 30984 18572 30990 18584
rect 31386 18572 31392 18584
rect 31444 18572 31450 18624
rect 31496 18612 31524 18652
rect 34054 18640 34060 18692
rect 34112 18680 34118 18692
rect 34885 18683 34943 18689
rect 34885 18680 34897 18683
rect 34112 18652 34897 18680
rect 34112 18640 34118 18652
rect 34885 18649 34897 18652
rect 34931 18649 34943 18683
rect 34885 18643 34943 18649
rect 35158 18640 35164 18692
rect 35216 18680 35222 18692
rect 35216 18652 35480 18680
rect 35216 18640 35222 18652
rect 35452 18624 35480 18652
rect 31938 18612 31944 18624
rect 31496 18584 31944 18612
rect 31938 18572 31944 18584
rect 31996 18572 32002 18624
rect 35434 18572 35440 18624
rect 35492 18572 35498 18624
rect 35802 18572 35808 18624
rect 35860 18612 35866 18624
rect 37550 18612 37556 18624
rect 35860 18584 37556 18612
rect 35860 18572 35866 18584
rect 37550 18572 37556 18584
rect 37608 18572 37614 18624
rect 1104 18522 38824 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 38824 18522
rect 1104 18448 38824 18470
rect 26418 18368 26424 18420
rect 26476 18408 26482 18420
rect 26605 18411 26663 18417
rect 26605 18408 26617 18411
rect 26476 18380 26617 18408
rect 26476 18368 26482 18380
rect 26605 18377 26617 18380
rect 26651 18377 26663 18411
rect 26605 18371 26663 18377
rect 28350 18368 28356 18420
rect 28408 18408 28414 18420
rect 28445 18411 28503 18417
rect 28445 18408 28457 18411
rect 28408 18380 28457 18408
rect 28408 18368 28414 18380
rect 28445 18377 28457 18380
rect 28491 18377 28503 18411
rect 31938 18408 31944 18420
rect 28445 18371 28503 18377
rect 28966 18380 31944 18408
rect 28258 18300 28264 18352
rect 28316 18340 28322 18352
rect 28966 18340 28994 18380
rect 31938 18368 31944 18380
rect 31996 18368 32002 18420
rect 28316 18312 28994 18340
rect 29457 18343 29515 18349
rect 28316 18300 28322 18312
rect 29457 18309 29469 18343
rect 29503 18340 29515 18343
rect 29546 18340 29552 18352
rect 29503 18312 29552 18340
rect 29503 18309 29515 18312
rect 29457 18303 29515 18309
rect 29546 18300 29552 18312
rect 29604 18300 29610 18352
rect 32214 18340 32220 18352
rect 31726 18312 32220 18340
rect 25222 18272 25228 18284
rect 25183 18244 25228 18272
rect 25222 18232 25228 18244
rect 25280 18232 25286 18284
rect 29362 18272 29368 18284
rect 29196 18244 29368 18272
rect 26602 18204 26608 18216
rect 25332 18176 26608 18204
rect 23382 18096 23388 18148
rect 23440 18136 23446 18148
rect 25332 18136 25360 18176
rect 26602 18164 26608 18176
rect 26660 18164 26666 18216
rect 27065 18207 27123 18213
rect 27065 18173 27077 18207
rect 27111 18204 27123 18207
rect 27154 18204 27160 18216
rect 27111 18176 27160 18204
rect 27111 18173 27123 18176
rect 27065 18167 27123 18173
rect 27154 18164 27160 18176
rect 27212 18164 27218 18216
rect 27614 18164 27620 18216
rect 27672 18204 27678 18216
rect 28718 18204 28724 18216
rect 27672 18176 28724 18204
rect 27672 18164 27678 18176
rect 28718 18164 28724 18176
rect 28776 18164 28782 18216
rect 29196 18213 29224 18244
rect 29362 18232 29368 18244
rect 29420 18232 29426 18284
rect 29181 18207 29239 18213
rect 29181 18173 29193 18207
rect 29227 18173 29239 18207
rect 29181 18167 29239 18173
rect 29273 18207 29331 18213
rect 29273 18173 29285 18207
rect 29319 18173 29331 18207
rect 29273 18167 29331 18173
rect 29549 18207 29607 18213
rect 29549 18173 29561 18207
rect 29595 18204 29607 18207
rect 29638 18204 29644 18216
rect 29595 18176 29644 18204
rect 29595 18173 29607 18176
rect 29549 18167 29607 18173
rect 25498 18145 25504 18148
rect 25492 18136 25504 18145
rect 23440 18108 25360 18136
rect 25459 18108 25504 18136
rect 23440 18096 23446 18108
rect 25492 18099 25504 18108
rect 25498 18096 25504 18099
rect 25556 18096 25562 18148
rect 26786 18096 26792 18148
rect 26844 18136 26850 18148
rect 27310 18139 27368 18145
rect 27310 18136 27322 18139
rect 26844 18108 27322 18136
rect 26844 18096 26850 18108
rect 27310 18105 27322 18108
rect 27356 18136 27368 18139
rect 27430 18136 27436 18148
rect 27356 18108 27436 18136
rect 27356 18105 27368 18108
rect 27310 18099 27368 18105
rect 27430 18096 27436 18108
rect 27488 18096 27494 18148
rect 29288 18136 29316 18167
rect 29638 18164 29644 18176
rect 29696 18164 29702 18216
rect 30469 18207 30527 18213
rect 30469 18173 30481 18207
rect 30515 18204 30527 18207
rect 31726 18204 31754 18312
rect 32214 18300 32220 18312
rect 32272 18340 32278 18352
rect 32272 18312 32352 18340
rect 32272 18300 32278 18312
rect 32324 18281 32352 18312
rect 33318 18300 33324 18352
rect 33376 18340 33382 18352
rect 33870 18340 33876 18352
rect 33376 18312 33876 18340
rect 33376 18300 33382 18312
rect 33870 18300 33876 18312
rect 33928 18300 33934 18352
rect 34698 18340 34704 18352
rect 34440 18312 34704 18340
rect 32309 18275 32367 18281
rect 32309 18241 32321 18275
rect 32355 18241 32367 18275
rect 32309 18235 32367 18241
rect 30515 18176 31754 18204
rect 30515 18173 30527 18176
rect 30469 18167 30527 18173
rect 32398 18164 32404 18216
rect 32456 18204 32462 18216
rect 32565 18207 32623 18213
rect 32565 18204 32577 18207
rect 32456 18176 32577 18204
rect 32456 18164 32462 18176
rect 32565 18173 32577 18176
rect 32611 18173 32623 18207
rect 32565 18167 32623 18173
rect 33870 18164 33876 18216
rect 33928 18204 33934 18216
rect 34440 18213 34468 18312
rect 34698 18300 34704 18312
rect 34756 18300 34762 18352
rect 35897 18343 35955 18349
rect 35897 18309 35909 18343
rect 35943 18309 35955 18343
rect 35897 18303 35955 18309
rect 35342 18272 35348 18284
rect 34624 18244 35348 18272
rect 34333 18207 34391 18213
rect 34333 18204 34345 18207
rect 33928 18176 34345 18204
rect 33928 18164 33934 18176
rect 34333 18173 34345 18176
rect 34379 18173 34391 18207
rect 34333 18167 34391 18173
rect 34425 18207 34483 18213
rect 34425 18173 34437 18207
rect 34471 18173 34483 18207
rect 34425 18167 34483 18173
rect 29454 18136 29460 18148
rect 29288 18108 29460 18136
rect 29454 18096 29460 18108
rect 29512 18096 29518 18148
rect 30736 18139 30794 18145
rect 30736 18105 30748 18139
rect 30782 18136 30794 18139
rect 30782 18108 30880 18136
rect 30782 18105 30794 18108
rect 30736 18099 30794 18105
rect 23842 18028 23848 18080
rect 23900 18068 23906 18080
rect 28074 18068 28080 18080
rect 23900 18040 28080 18068
rect 23900 18028 23906 18040
rect 28074 18028 28080 18040
rect 28132 18028 28138 18080
rect 28997 18071 29055 18077
rect 28997 18037 29009 18071
rect 29043 18068 29055 18071
rect 29086 18068 29092 18080
rect 29043 18040 29092 18068
rect 29043 18037 29055 18040
rect 28997 18031 29055 18037
rect 29086 18028 29092 18040
rect 29144 18028 29150 18080
rect 30852 18068 30880 18108
rect 30926 18096 30932 18148
rect 30984 18136 30990 18148
rect 34149 18139 34207 18145
rect 34149 18136 34161 18139
rect 30984 18108 34161 18136
rect 30984 18096 30990 18108
rect 34149 18105 34161 18108
rect 34195 18105 34207 18139
rect 34440 18136 34468 18167
rect 34514 18164 34520 18216
rect 34572 18204 34578 18216
rect 34624 18213 34652 18244
rect 35342 18232 35348 18244
rect 35400 18272 35406 18284
rect 35912 18272 35940 18303
rect 35400 18244 35940 18272
rect 35400 18232 35406 18244
rect 34609 18207 34667 18213
rect 34609 18204 34621 18207
rect 34572 18176 34621 18204
rect 34572 18164 34578 18176
rect 34609 18173 34621 18176
rect 34655 18173 34667 18207
rect 34609 18167 34667 18173
rect 34698 18164 34704 18216
rect 34756 18204 34762 18216
rect 34756 18176 34801 18204
rect 34756 18164 34762 18176
rect 34882 18164 34888 18216
rect 34940 18204 34946 18216
rect 35713 18207 35771 18213
rect 35713 18204 35725 18207
rect 34940 18176 35725 18204
rect 34940 18164 34946 18176
rect 35713 18173 35725 18176
rect 35759 18173 35771 18207
rect 37274 18204 37280 18216
rect 37235 18176 37280 18204
rect 35713 18167 35771 18173
rect 37274 18164 37280 18176
rect 37332 18164 37338 18216
rect 37918 18204 37924 18216
rect 37879 18176 37924 18204
rect 37918 18164 37924 18176
rect 37976 18164 37982 18216
rect 34440 18108 34744 18136
rect 34149 18099 34207 18105
rect 34716 18080 34744 18108
rect 31478 18068 31484 18080
rect 30852 18040 31484 18068
rect 31478 18028 31484 18040
rect 31536 18028 31542 18080
rect 31849 18071 31907 18077
rect 31849 18037 31861 18071
rect 31895 18068 31907 18071
rect 32030 18068 32036 18080
rect 31895 18040 32036 18068
rect 31895 18037 31907 18040
rect 31849 18031 31907 18037
rect 32030 18028 32036 18040
rect 32088 18028 32094 18080
rect 32582 18028 32588 18080
rect 32640 18068 32646 18080
rect 33042 18068 33048 18080
rect 32640 18040 33048 18068
rect 32640 18028 32646 18040
rect 33042 18028 33048 18040
rect 33100 18068 33106 18080
rect 33689 18071 33747 18077
rect 33689 18068 33701 18071
rect 33100 18040 33701 18068
rect 33100 18028 33106 18040
rect 33689 18037 33701 18040
rect 33735 18037 33747 18071
rect 33689 18031 33747 18037
rect 34698 18028 34704 18080
rect 34756 18028 34762 18080
rect 1104 17978 38824 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 38824 17978
rect 1104 17904 38824 17926
rect 24762 17824 24768 17876
rect 24820 17864 24826 17876
rect 26789 17867 26847 17873
rect 26789 17864 26801 17867
rect 24820 17836 26801 17864
rect 24820 17824 24826 17836
rect 26789 17833 26801 17836
rect 26835 17833 26847 17867
rect 26789 17827 26847 17833
rect 28258 17824 28264 17876
rect 28316 17864 28322 17876
rect 28902 17864 28908 17876
rect 28316 17836 28908 17864
rect 28316 17824 28322 17836
rect 28902 17824 28908 17836
rect 28960 17864 28966 17876
rect 29181 17867 29239 17873
rect 29181 17864 29193 17867
rect 28960 17836 29193 17864
rect 28960 17824 28966 17836
rect 29181 17833 29193 17836
rect 29227 17833 29239 17867
rect 29181 17827 29239 17833
rect 29362 17824 29368 17876
rect 29420 17864 29426 17876
rect 31481 17867 31539 17873
rect 31481 17864 31493 17867
rect 29420 17836 31493 17864
rect 29420 17824 29426 17836
rect 31481 17833 31493 17836
rect 31527 17833 31539 17867
rect 34054 17864 34060 17876
rect 31481 17827 31539 17833
rect 31956 17836 34060 17864
rect 1854 17796 1860 17808
rect 1815 17768 1860 17796
rect 1854 17756 1860 17768
rect 1912 17756 1918 17808
rect 23842 17805 23848 17808
rect 23836 17796 23848 17805
rect 23803 17768 23848 17796
rect 23836 17759 23848 17768
rect 23842 17756 23848 17759
rect 23900 17756 23906 17808
rect 23934 17756 23940 17808
rect 23992 17796 23998 17808
rect 25222 17796 25228 17808
rect 23992 17768 25228 17796
rect 23992 17756 23998 17768
rect 25222 17756 25228 17768
rect 25280 17756 25286 17808
rect 25676 17799 25734 17805
rect 25676 17796 25688 17799
rect 25608 17768 25688 17796
rect 23569 17731 23627 17737
rect 23569 17697 23581 17731
rect 23615 17728 23627 17731
rect 23952 17728 23980 17756
rect 25608 17728 25636 17768
rect 25676 17765 25688 17768
rect 25722 17796 25734 17799
rect 26878 17796 26884 17808
rect 25722 17768 26884 17796
rect 25722 17765 25734 17768
rect 25676 17759 25734 17765
rect 26878 17756 26884 17768
rect 26936 17756 26942 17808
rect 28068 17799 28126 17805
rect 28068 17765 28080 17799
rect 28114 17796 28126 17799
rect 28994 17796 29000 17808
rect 28114 17768 29000 17796
rect 28114 17765 28126 17768
rect 28068 17759 28126 17765
rect 28994 17756 29000 17768
rect 29052 17756 29058 17808
rect 29908 17799 29966 17805
rect 29908 17765 29920 17799
rect 29954 17796 29966 17799
rect 30374 17796 30380 17808
rect 29954 17768 30380 17796
rect 29954 17765 29966 17768
rect 29908 17759 29966 17765
rect 30374 17756 30380 17768
rect 30432 17756 30438 17808
rect 31846 17796 31852 17808
rect 30484 17768 31852 17796
rect 30484 17728 30512 17768
rect 31846 17756 31852 17768
rect 31904 17756 31910 17808
rect 23615 17700 23980 17728
rect 24964 17700 25636 17728
rect 26436 17700 30512 17728
rect 23615 17697 23627 17700
rect 23569 17691 23627 17697
rect 24964 17601 24992 17700
rect 25222 17620 25228 17672
rect 25280 17660 25286 17672
rect 25409 17663 25467 17669
rect 25409 17660 25421 17663
rect 25280 17632 25421 17660
rect 25280 17620 25286 17632
rect 25409 17629 25421 17632
rect 25455 17629 25467 17663
rect 25409 17623 25467 17629
rect 24949 17595 25007 17601
rect 24949 17561 24961 17595
rect 24995 17561 25007 17595
rect 24949 17555 25007 17561
rect 1949 17527 2007 17533
rect 1949 17493 1961 17527
rect 1995 17524 2007 17527
rect 16298 17524 16304 17536
rect 1995 17496 16304 17524
rect 1995 17493 2007 17496
rect 1949 17487 2007 17493
rect 16298 17484 16304 17496
rect 16356 17484 16362 17536
rect 24302 17484 24308 17536
rect 24360 17524 24366 17536
rect 26436 17524 26464 17700
rect 30742 17688 30748 17740
rect 30800 17728 30806 17740
rect 31665 17731 31723 17737
rect 31665 17728 31677 17731
rect 30800 17700 31677 17728
rect 30800 17688 30806 17700
rect 31665 17697 31677 17700
rect 31711 17697 31723 17731
rect 31665 17691 31723 17697
rect 31757 17731 31815 17737
rect 31757 17697 31769 17731
rect 31803 17728 31815 17731
rect 31956 17728 31984 17836
rect 34054 17824 34060 17836
rect 34112 17824 34118 17876
rect 34422 17864 34428 17876
rect 34383 17836 34428 17864
rect 34422 17824 34428 17836
rect 34480 17824 34486 17876
rect 32490 17756 32496 17808
rect 32548 17796 32554 17808
rect 33290 17799 33348 17805
rect 33290 17796 33302 17799
rect 32548 17768 33302 17796
rect 32548 17756 32554 17768
rect 33290 17765 33302 17768
rect 33336 17765 33348 17799
rect 33290 17759 33348 17765
rect 34606 17756 34612 17808
rect 34664 17796 34670 17808
rect 34664 17768 35204 17796
rect 34664 17756 34670 17768
rect 31803 17700 31984 17728
rect 32033 17731 32091 17737
rect 31803 17697 31815 17700
rect 31757 17691 31815 17697
rect 32033 17697 32045 17731
rect 32079 17697 32091 17731
rect 32033 17691 32091 17697
rect 27154 17620 27160 17672
rect 27212 17660 27218 17672
rect 27798 17660 27804 17672
rect 27212 17632 27804 17660
rect 27212 17620 27218 17632
rect 27798 17620 27804 17632
rect 27856 17620 27862 17672
rect 29641 17663 29699 17669
rect 29641 17660 29653 17663
rect 28828 17632 29653 17660
rect 24360 17496 26464 17524
rect 24360 17484 24366 17496
rect 27798 17484 27804 17536
rect 27856 17524 27862 17536
rect 28828 17524 28856 17632
rect 29641 17629 29653 17632
rect 29687 17629 29699 17663
rect 32048 17660 32076 17691
rect 32214 17688 32220 17740
rect 32272 17728 32278 17740
rect 33045 17731 33103 17737
rect 33045 17728 33057 17731
rect 32272 17700 33057 17728
rect 32272 17688 32278 17700
rect 33045 17697 33057 17700
rect 33091 17697 33103 17731
rect 33045 17691 33103 17697
rect 33134 17688 33140 17740
rect 33192 17728 33198 17740
rect 34882 17728 34888 17740
rect 33192 17700 34888 17728
rect 33192 17688 33198 17700
rect 34882 17688 34888 17700
rect 34940 17688 34946 17740
rect 35066 17728 35072 17740
rect 35027 17700 35072 17728
rect 35066 17688 35072 17700
rect 35124 17688 35130 17740
rect 35176 17737 35204 17768
rect 35161 17731 35219 17737
rect 35161 17697 35173 17731
rect 35207 17697 35219 17731
rect 35357 17731 35415 17737
rect 35357 17728 35369 17731
rect 35161 17691 35219 17697
rect 35268 17700 35369 17728
rect 29641 17623 29699 17629
rect 30668 17632 32076 17660
rect 27856 17496 28856 17524
rect 27856 17484 27862 17496
rect 29638 17484 29644 17536
rect 29696 17524 29702 17536
rect 30668 17524 30696 17632
rect 34514 17620 34520 17672
rect 34572 17660 34578 17672
rect 35268 17660 35296 17700
rect 35357 17697 35369 17700
rect 35403 17697 35415 17731
rect 35357 17691 35415 17697
rect 35447 17731 35505 17737
rect 35447 17697 35459 17731
rect 35493 17728 35505 17731
rect 35710 17728 35716 17740
rect 35493 17700 35716 17728
rect 35493 17697 35505 17700
rect 35447 17691 35505 17697
rect 35710 17688 35716 17700
rect 35768 17688 35774 17740
rect 34572 17632 35296 17660
rect 34572 17620 34578 17632
rect 31386 17552 31392 17604
rect 31444 17592 31450 17604
rect 34885 17595 34943 17601
rect 34885 17592 34897 17595
rect 31444 17564 33088 17592
rect 31444 17552 31450 17564
rect 29696 17496 30696 17524
rect 29696 17484 29702 17496
rect 30742 17484 30748 17536
rect 30800 17524 30806 17536
rect 31021 17527 31079 17533
rect 31021 17524 31033 17527
rect 30800 17496 31033 17524
rect 30800 17484 30806 17496
rect 31021 17493 31033 17496
rect 31067 17524 31079 17527
rect 31202 17524 31208 17536
rect 31067 17496 31208 17524
rect 31067 17493 31079 17496
rect 31021 17487 31079 17493
rect 31202 17484 31208 17496
rect 31260 17484 31266 17536
rect 31754 17484 31760 17536
rect 31812 17524 31818 17536
rect 31941 17527 31999 17533
rect 31941 17524 31953 17527
rect 31812 17496 31953 17524
rect 31812 17484 31818 17496
rect 31941 17493 31953 17496
rect 31987 17493 31999 17527
rect 33060 17524 33088 17564
rect 33980 17564 34897 17592
rect 33980 17524 34008 17564
rect 34885 17561 34897 17564
rect 34931 17561 34943 17595
rect 34885 17555 34943 17561
rect 35066 17552 35072 17604
rect 35124 17592 35130 17604
rect 35342 17592 35348 17604
rect 35124 17564 35348 17592
rect 35124 17552 35130 17564
rect 35342 17552 35348 17564
rect 35400 17552 35406 17604
rect 33060 17496 34008 17524
rect 31941 17487 31999 17493
rect 1104 17434 38824 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 38824 17434
rect 1104 17360 38824 17382
rect 24670 17280 24676 17332
rect 24728 17320 24734 17332
rect 26605 17323 26663 17329
rect 26605 17320 26617 17323
rect 24728 17292 26617 17320
rect 24728 17280 24734 17292
rect 26605 17289 26617 17292
rect 26651 17289 26663 17323
rect 26605 17283 26663 17289
rect 27430 17280 27436 17332
rect 27488 17320 27494 17332
rect 28445 17323 28503 17329
rect 28445 17320 28457 17323
rect 27488 17292 28457 17320
rect 27488 17280 27494 17292
rect 28445 17289 28457 17292
rect 28491 17289 28503 17323
rect 28445 17283 28503 17289
rect 28552 17292 31432 17320
rect 25222 17184 25228 17196
rect 25183 17156 25228 17184
rect 25222 17144 25228 17156
rect 25280 17144 25286 17196
rect 24305 17119 24363 17125
rect 24305 17085 24317 17119
rect 24351 17116 24363 17119
rect 25130 17116 25136 17128
rect 24351 17088 25136 17116
rect 24351 17085 24363 17088
rect 24305 17079 24363 17085
rect 25130 17076 25136 17088
rect 25188 17076 25194 17128
rect 25958 17076 25964 17128
rect 26016 17116 26022 17128
rect 27065 17119 27123 17125
rect 27065 17116 27077 17119
rect 26016 17088 27077 17116
rect 26016 17076 26022 17088
rect 27065 17085 27077 17088
rect 27111 17085 27123 17119
rect 27065 17079 27123 17085
rect 27154 17076 27160 17128
rect 27212 17116 27218 17128
rect 28552 17116 28580 17292
rect 29270 17252 29276 17264
rect 29196 17224 29276 17252
rect 28994 17116 29000 17128
rect 27212 17088 28580 17116
rect 27212 17076 27218 17088
rect 28966 17076 29000 17116
rect 29052 17076 29058 17128
rect 29196 17125 29224 17224
rect 29270 17212 29276 17224
rect 29328 17212 29334 17264
rect 31404 17252 31432 17292
rect 31478 17280 31484 17332
rect 31536 17320 31542 17332
rect 31849 17323 31907 17329
rect 31849 17320 31861 17323
rect 31536 17292 31861 17320
rect 31536 17280 31542 17292
rect 31849 17289 31861 17292
rect 31895 17289 31907 17323
rect 31849 17283 31907 17289
rect 37461 17323 37519 17329
rect 37461 17289 37473 17323
rect 37507 17320 37519 17323
rect 38654 17320 38660 17332
rect 37507 17292 38660 17320
rect 37507 17289 37519 17292
rect 37461 17283 37519 17289
rect 38654 17280 38660 17292
rect 38712 17280 38718 17332
rect 31404 17224 31754 17252
rect 29454 17184 29460 17196
rect 29415 17156 29460 17184
rect 29454 17144 29460 17156
rect 29512 17144 29518 17196
rect 29181 17119 29239 17125
rect 29181 17085 29193 17119
rect 29227 17085 29239 17119
rect 29181 17079 29239 17085
rect 29319 17119 29377 17125
rect 29319 17085 29331 17119
rect 29365 17085 29377 17119
rect 29319 17079 29377 17085
rect 29549 17119 29607 17125
rect 29549 17085 29561 17119
rect 29595 17116 29607 17119
rect 29638 17116 29644 17128
rect 29595 17088 29644 17116
rect 29595 17085 29607 17088
rect 29549 17079 29607 17085
rect 1854 17048 1860 17060
rect 1815 17020 1860 17048
rect 1854 17008 1860 17020
rect 1912 17008 1918 17060
rect 24118 17048 24124 17060
rect 24079 17020 24124 17048
rect 24118 17008 24124 17020
rect 24176 17008 24182 17060
rect 24762 17008 24768 17060
rect 24820 17048 24826 17060
rect 25470 17051 25528 17057
rect 25470 17048 25482 17051
rect 24820 17020 25482 17048
rect 24820 17008 24826 17020
rect 25470 17017 25482 17020
rect 25516 17017 25528 17051
rect 25470 17011 25528 17017
rect 26418 17008 26424 17060
rect 26476 17048 26482 17060
rect 27310 17051 27368 17057
rect 27310 17048 27322 17051
rect 26476 17020 27322 17048
rect 26476 17008 26482 17020
rect 27310 17017 27322 17020
rect 27356 17017 27368 17051
rect 28966 17048 28994 17076
rect 27310 17011 27368 17017
rect 27448 17020 28994 17048
rect 1949 16983 2007 16989
rect 1949 16949 1961 16983
rect 1995 16980 2007 16983
rect 17494 16980 17500 16992
rect 1995 16952 17500 16980
rect 1995 16949 2007 16952
rect 1949 16943 2007 16949
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 24854 16940 24860 16992
rect 24912 16980 24918 16992
rect 27448 16980 27476 17020
rect 28994 16980 29000 16992
rect 24912 16952 27476 16980
rect 28955 16952 29000 16980
rect 24912 16940 24918 16952
rect 28994 16940 29000 16952
rect 29052 16940 29058 16992
rect 29334 16980 29362 17079
rect 29638 17076 29644 17088
rect 29696 17076 29702 17128
rect 30374 17076 30380 17128
rect 30432 17116 30438 17128
rect 30469 17119 30527 17125
rect 30469 17116 30481 17119
rect 30432 17088 30481 17116
rect 30432 17076 30438 17088
rect 30469 17085 30481 17088
rect 30515 17116 30527 17119
rect 31202 17116 31208 17128
rect 30515 17088 31208 17116
rect 30515 17085 30527 17088
rect 30469 17079 30527 17085
rect 31202 17076 31208 17088
rect 31260 17076 31266 17128
rect 30282 17008 30288 17060
rect 30340 17048 30346 17060
rect 30714 17051 30772 17057
rect 30714 17048 30726 17051
rect 30340 17020 30726 17048
rect 30340 17008 30346 17020
rect 30714 17017 30726 17020
rect 30760 17017 30772 17051
rect 30714 17011 30772 17017
rect 30926 16980 30932 16992
rect 29334 16952 30932 16980
rect 30926 16940 30932 16952
rect 30984 16940 30990 16992
rect 31726 16980 31754 17224
rect 36538 17212 36544 17264
rect 36596 17252 36602 17264
rect 37090 17252 37096 17264
rect 36596 17224 37096 17252
rect 36596 17212 36602 17224
rect 37090 17212 37096 17224
rect 37148 17212 37154 17264
rect 32122 17144 32128 17196
rect 32180 17184 32186 17196
rect 33781 17187 33839 17193
rect 33781 17184 33793 17187
rect 32180 17156 33793 17184
rect 32180 17144 32186 17156
rect 33781 17153 33793 17156
rect 33827 17153 33839 17187
rect 34514 17184 34520 17196
rect 33781 17147 33839 17153
rect 34256 17156 34520 17184
rect 32306 17116 32312 17128
rect 32267 17088 32312 17116
rect 32306 17076 32312 17088
rect 32364 17076 32370 17128
rect 33965 17119 34023 17125
rect 33965 17085 33977 17119
rect 34011 17085 34023 17119
rect 33965 17079 34023 17085
rect 34057 17119 34115 17125
rect 34057 17085 34069 17119
rect 34103 17085 34115 17119
rect 34057 17079 34115 17085
rect 31846 17008 31852 17060
rect 31904 17048 31910 17060
rect 33042 17048 33048 17060
rect 31904 17020 33048 17048
rect 31904 17008 31910 17020
rect 33042 17008 33048 17020
rect 33100 17008 33106 17060
rect 32493 16983 32551 16989
rect 32493 16980 32505 16983
rect 31726 16952 32505 16980
rect 32493 16949 32505 16952
rect 32539 16949 32551 16983
rect 33980 16980 34008 17079
rect 34072 17048 34100 17079
rect 34146 17076 34152 17128
rect 34204 17116 34210 17128
rect 34256 17125 34284 17156
rect 34514 17144 34520 17156
rect 34572 17144 34578 17196
rect 36630 17144 36636 17196
rect 36688 17184 36694 17196
rect 36814 17184 36820 17196
rect 36688 17156 36820 17184
rect 36688 17144 36694 17156
rect 36814 17144 36820 17156
rect 36872 17144 36878 17196
rect 34241 17119 34299 17125
rect 34241 17116 34253 17119
rect 34204 17088 34253 17116
rect 34204 17076 34210 17088
rect 34241 17085 34253 17088
rect 34287 17085 34299 17119
rect 34241 17079 34299 17085
rect 34330 17076 34336 17128
rect 34388 17116 34394 17128
rect 37274 17116 37280 17128
rect 34388 17088 34433 17116
rect 37235 17088 37280 17116
rect 34388 17076 34394 17088
rect 37274 17076 37280 17088
rect 37332 17076 37338 17128
rect 37918 17116 37924 17128
rect 37879 17088 37924 17116
rect 37918 17076 37924 17088
rect 37976 17076 37982 17128
rect 34698 17048 34704 17060
rect 34072 17020 34704 17048
rect 34698 17008 34704 17020
rect 34756 17008 34762 17060
rect 37550 16980 37556 16992
rect 33980 16952 37556 16980
rect 32493 16943 32551 16949
rect 37550 16940 37556 16952
rect 37608 16940 37614 16992
rect 1104 16890 38824 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 38824 16890
rect 1104 16816 38824 16838
rect 23584 16748 25452 16776
rect 23584 16649 23612 16748
rect 24670 16668 24676 16720
rect 24728 16708 24734 16720
rect 25286 16711 25344 16717
rect 25286 16708 25298 16711
rect 24728 16680 25298 16708
rect 24728 16668 24734 16680
rect 25286 16677 25298 16680
rect 25332 16677 25344 16711
rect 25286 16671 25344 16677
rect 23569 16643 23627 16649
rect 23569 16609 23581 16643
rect 23615 16609 23627 16643
rect 24026 16640 24032 16652
rect 23987 16612 24032 16640
rect 23569 16603 23627 16609
rect 24026 16600 24032 16612
rect 24084 16600 24090 16652
rect 24210 16640 24216 16652
rect 24171 16612 24216 16640
rect 24210 16600 24216 16612
rect 24268 16600 24274 16652
rect 24302 16600 24308 16652
rect 24360 16640 24366 16652
rect 24581 16643 24639 16649
rect 24360 16612 24405 16640
rect 24360 16600 24366 16612
rect 24581 16609 24593 16643
rect 24627 16640 24639 16643
rect 24854 16640 24860 16652
rect 24627 16612 24860 16640
rect 24627 16609 24639 16612
rect 24581 16603 24639 16609
rect 24854 16600 24860 16612
rect 24912 16600 24918 16652
rect 25424 16640 25452 16748
rect 25498 16736 25504 16788
rect 25556 16776 25562 16788
rect 26421 16779 26479 16785
rect 26421 16776 26433 16779
rect 25556 16748 26433 16776
rect 25556 16736 25562 16748
rect 26421 16745 26433 16748
rect 26467 16745 26479 16779
rect 29181 16779 29239 16785
rect 29181 16776 29193 16779
rect 26421 16739 26479 16745
rect 26620 16748 29193 16776
rect 26234 16668 26240 16720
rect 26292 16708 26298 16720
rect 26620 16708 26648 16748
rect 29181 16745 29193 16748
rect 29227 16745 29239 16779
rect 29181 16739 29239 16745
rect 29270 16736 29276 16788
rect 29328 16776 29334 16788
rect 31018 16776 31024 16788
rect 29328 16748 30696 16776
rect 30979 16748 31024 16776
rect 29328 16736 29334 16748
rect 27890 16708 27896 16720
rect 26292 16680 26648 16708
rect 27632 16680 27896 16708
rect 26292 16668 26298 16680
rect 27632 16640 27660 16680
rect 27890 16668 27896 16680
rect 27948 16668 27954 16720
rect 28068 16711 28126 16717
rect 28068 16677 28080 16711
rect 28114 16708 28126 16711
rect 28350 16708 28356 16720
rect 28114 16680 28356 16708
rect 28114 16677 28126 16680
rect 28068 16671 28126 16677
rect 28350 16668 28356 16680
rect 28408 16668 28414 16720
rect 29908 16711 29966 16717
rect 29908 16677 29920 16711
rect 29954 16708 29966 16711
rect 30558 16708 30564 16720
rect 29954 16680 30564 16708
rect 29954 16677 29966 16680
rect 29908 16671 29966 16677
rect 30558 16668 30564 16680
rect 30616 16668 30622 16720
rect 30668 16708 30696 16748
rect 31018 16736 31024 16748
rect 31076 16736 31082 16788
rect 31202 16736 31208 16788
rect 31260 16776 31266 16788
rect 32214 16776 32220 16788
rect 31260 16748 32220 16776
rect 31260 16736 31266 16748
rect 32214 16736 32220 16748
rect 32272 16736 32278 16788
rect 34606 16776 34612 16788
rect 33796 16748 34612 16776
rect 31481 16711 31539 16717
rect 31481 16708 31493 16711
rect 30668 16680 31493 16708
rect 31481 16677 31493 16680
rect 31527 16677 31539 16711
rect 31481 16671 31539 16677
rect 31772 16680 32536 16708
rect 27798 16640 27804 16652
rect 25424 16612 27660 16640
rect 27759 16612 27804 16640
rect 27798 16600 27804 16612
rect 27856 16600 27862 16652
rect 29641 16643 29699 16649
rect 29641 16609 29653 16643
rect 29687 16640 29699 16643
rect 30374 16640 30380 16652
rect 29687 16612 30380 16640
rect 29687 16609 29699 16612
rect 29641 16603 29699 16609
rect 30374 16600 30380 16612
rect 30432 16600 30438 16652
rect 31570 16600 31576 16652
rect 31628 16640 31634 16652
rect 31772 16649 31800 16680
rect 31665 16643 31723 16649
rect 31665 16640 31677 16643
rect 31628 16612 31677 16640
rect 31628 16600 31634 16612
rect 31665 16609 31677 16612
rect 31711 16609 31723 16643
rect 31665 16603 31723 16609
rect 31757 16643 31815 16649
rect 31757 16609 31769 16643
rect 31803 16609 31815 16643
rect 31757 16603 31815 16609
rect 32033 16643 32091 16649
rect 32033 16609 32045 16643
rect 32079 16609 32091 16643
rect 32306 16640 32312 16652
rect 32033 16603 32091 16609
rect 32140 16612 32312 16640
rect 25038 16572 25044 16584
rect 24999 16544 25044 16572
rect 25038 16532 25044 16544
rect 25096 16532 25102 16584
rect 31202 16532 31208 16584
rect 31260 16572 31266 16584
rect 32048 16572 32076 16603
rect 31260 16544 32076 16572
rect 31260 16532 31266 16544
rect 23474 16464 23480 16516
rect 23532 16504 23538 16516
rect 24118 16504 24124 16516
rect 23532 16476 24124 16504
rect 23532 16464 23538 16476
rect 24118 16464 24124 16476
rect 24176 16504 24182 16516
rect 32140 16504 32168 16612
rect 32306 16600 32312 16612
rect 32364 16600 32370 16652
rect 24176 16476 24799 16504
rect 24176 16464 24182 16476
rect 22922 16396 22928 16448
rect 22980 16436 22986 16448
rect 23385 16439 23443 16445
rect 23385 16436 23397 16439
rect 22980 16408 23397 16436
rect 22980 16396 22986 16408
rect 23385 16405 23397 16408
rect 23431 16405 23443 16439
rect 23385 16399 23443 16405
rect 24489 16439 24547 16445
rect 24489 16405 24501 16439
rect 24535 16436 24547 16439
rect 24670 16436 24676 16448
rect 24535 16408 24676 16436
rect 24535 16405 24547 16408
rect 24489 16399 24547 16405
rect 24670 16396 24676 16408
rect 24728 16396 24734 16448
rect 24771 16436 24799 16476
rect 31726 16476 32168 16504
rect 28718 16436 28724 16448
rect 24771 16408 28724 16436
rect 28718 16396 28724 16408
rect 28776 16396 28782 16448
rect 29638 16396 29644 16448
rect 29696 16436 29702 16448
rect 31726 16436 31754 16476
rect 31938 16436 31944 16448
rect 29696 16408 31754 16436
rect 31899 16408 31944 16436
rect 29696 16396 29702 16408
rect 31938 16396 31944 16408
rect 31996 16396 32002 16448
rect 32508 16436 32536 16680
rect 33318 16668 33324 16720
rect 33376 16708 33382 16720
rect 33796 16708 33824 16748
rect 34606 16736 34612 16748
rect 34664 16736 34670 16788
rect 35710 16736 35716 16788
rect 35768 16776 35774 16788
rect 36078 16776 36084 16788
rect 35768 16748 36084 16776
rect 35768 16736 35774 16748
rect 36078 16736 36084 16748
rect 36136 16736 36142 16788
rect 34146 16708 34152 16720
rect 33376 16680 33824 16708
rect 33376 16668 33382 16680
rect 33796 16649 33824 16680
rect 33980 16680 34152 16708
rect 33980 16649 34008 16680
rect 34146 16668 34152 16680
rect 34204 16668 34210 16720
rect 34624 16708 34652 16736
rect 34624 16680 34836 16708
rect 33689 16643 33747 16649
rect 33689 16609 33701 16643
rect 33735 16609 33747 16643
rect 33689 16603 33747 16609
rect 33781 16643 33839 16649
rect 33781 16609 33793 16643
rect 33827 16609 33839 16643
rect 33781 16603 33839 16609
rect 33965 16643 34023 16649
rect 33965 16609 33977 16643
rect 34011 16609 34023 16643
rect 33965 16603 34023 16609
rect 34057 16643 34115 16649
rect 34057 16609 34069 16643
rect 34103 16640 34115 16643
rect 34330 16640 34336 16652
rect 34103 16612 34336 16640
rect 34103 16609 34115 16612
rect 34057 16603 34115 16609
rect 33704 16572 33732 16603
rect 34330 16600 34336 16612
rect 34388 16600 34394 16652
rect 34606 16600 34612 16652
rect 34664 16640 34670 16652
rect 34808 16649 34836 16680
rect 34701 16643 34759 16649
rect 34701 16640 34713 16643
rect 34664 16612 34713 16640
rect 34664 16600 34670 16612
rect 34701 16609 34713 16612
rect 34747 16609 34759 16643
rect 34701 16603 34759 16609
rect 34793 16643 34851 16649
rect 34793 16609 34805 16643
rect 34839 16609 34851 16643
rect 34793 16603 34851 16609
rect 34977 16643 35035 16649
rect 34977 16609 34989 16643
rect 35023 16609 35035 16643
rect 34977 16603 35035 16609
rect 35069 16643 35127 16649
rect 35069 16609 35081 16643
rect 35115 16640 35127 16643
rect 35250 16640 35256 16652
rect 35115 16612 35256 16640
rect 35115 16609 35127 16612
rect 35069 16603 35127 16609
rect 34146 16572 34152 16584
rect 33704 16544 34152 16572
rect 34146 16532 34152 16544
rect 34204 16532 34210 16584
rect 34517 16575 34575 16581
rect 34517 16572 34529 16575
rect 34256 16544 34529 16572
rect 32582 16464 32588 16516
rect 32640 16504 32646 16516
rect 33505 16507 33563 16513
rect 33505 16504 33517 16507
rect 32640 16476 33517 16504
rect 32640 16464 32646 16476
rect 33505 16473 33517 16476
rect 33551 16473 33563 16507
rect 33505 16467 33563 16473
rect 34256 16436 34284 16544
rect 34517 16541 34529 16544
rect 34563 16541 34575 16575
rect 34517 16535 34575 16541
rect 32508 16408 34284 16436
rect 34606 16396 34612 16448
rect 34664 16436 34670 16448
rect 34992 16436 35020 16603
rect 35250 16600 35256 16612
rect 35308 16600 35314 16652
rect 34664 16408 35020 16436
rect 34664 16396 34670 16408
rect 1104 16346 38824 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 38824 16346
rect 1104 16272 38824 16294
rect 23842 16192 23848 16244
rect 23900 16232 23906 16244
rect 23937 16235 23995 16241
rect 23937 16232 23949 16235
rect 23900 16204 23949 16232
rect 23900 16192 23906 16204
rect 23937 16201 23949 16204
rect 23983 16201 23995 16235
rect 25958 16232 25964 16244
rect 23937 16195 23995 16201
rect 25608 16204 25964 16232
rect 25038 16056 25044 16108
rect 25096 16096 25102 16108
rect 25406 16096 25412 16108
rect 25096 16068 25412 16096
rect 25096 16056 25102 16068
rect 25406 16056 25412 16068
rect 25464 16096 25470 16108
rect 25608 16105 25636 16204
rect 25958 16192 25964 16204
rect 26016 16232 26022 16244
rect 26016 16204 26648 16232
rect 26016 16192 26022 16204
rect 25593 16099 25651 16105
rect 25593 16096 25605 16099
rect 25464 16068 25605 16096
rect 25464 16056 25470 16068
rect 25593 16065 25605 16068
rect 25639 16065 25651 16099
rect 26620 16096 26648 16204
rect 26786 16192 26792 16244
rect 26844 16232 26850 16244
rect 29549 16235 29607 16241
rect 26844 16204 28488 16232
rect 26844 16192 26850 16204
rect 28460 16164 28488 16204
rect 29549 16201 29561 16235
rect 29595 16232 29607 16235
rect 29638 16232 29644 16244
rect 29595 16204 29644 16232
rect 29595 16201 29607 16204
rect 29549 16195 29607 16201
rect 29638 16192 29644 16204
rect 29696 16192 29702 16244
rect 29914 16192 29920 16244
rect 29972 16232 29978 16244
rect 32217 16235 32275 16241
rect 32217 16232 32229 16235
rect 29972 16204 32229 16232
rect 29972 16192 29978 16204
rect 32217 16201 32229 16204
rect 32263 16201 32275 16235
rect 32217 16195 32275 16201
rect 33042 16192 33048 16244
rect 33100 16232 33106 16244
rect 33229 16235 33287 16241
rect 33229 16232 33241 16235
rect 33100 16204 33241 16232
rect 33100 16192 33106 16204
rect 33229 16201 33241 16204
rect 33275 16201 33287 16235
rect 33229 16195 33287 16201
rect 33778 16192 33784 16244
rect 33836 16192 33842 16244
rect 37461 16235 37519 16241
rect 37461 16201 37473 16235
rect 37507 16232 37519 16235
rect 38102 16232 38108 16244
rect 37507 16204 38108 16232
rect 37507 16201 37519 16204
rect 37461 16195 37519 16201
rect 38102 16192 38108 16204
rect 38160 16192 38166 16244
rect 28460 16136 28994 16164
rect 27522 16096 27528 16108
rect 26620 16068 27528 16096
rect 25593 16059 25651 16065
rect 27522 16056 27528 16068
rect 27580 16056 27586 16108
rect 28966 16096 28994 16136
rect 30190 16124 30196 16176
rect 30248 16164 30254 16176
rect 31202 16164 31208 16176
rect 30248 16136 31208 16164
rect 30248 16124 30254 16136
rect 30929 16099 30987 16105
rect 30929 16096 30941 16099
rect 28966 16068 30941 16096
rect 30929 16065 30941 16068
rect 30975 16065 30987 16099
rect 30929 16059 30987 16065
rect 1854 16028 1860 16040
rect 1815 16000 1860 16028
rect 1854 15988 1860 16000
rect 1912 15988 1918 16040
rect 22557 16031 22615 16037
rect 22557 15997 22569 16031
rect 22603 16028 22615 16031
rect 22646 16028 22652 16040
rect 22603 16000 22652 16028
rect 22603 15997 22615 16000
rect 22557 15991 22615 15997
rect 22646 15988 22652 16000
rect 22704 16028 22710 16040
rect 23934 16028 23940 16040
rect 22704 16000 23940 16028
rect 22704 15988 22710 16000
rect 23934 15988 23940 16000
rect 23992 16028 23998 16040
rect 24302 16028 24308 16040
rect 23992 16000 24308 16028
rect 23992 15988 23998 16000
rect 24302 15988 24308 16000
rect 24360 15988 24366 16040
rect 25860 16031 25918 16037
rect 25860 15997 25872 16031
rect 25906 16028 25918 16031
rect 27430 16028 27436 16040
rect 25906 16000 27436 16028
rect 25906 15997 25918 16000
rect 25860 15991 25918 15997
rect 27430 15988 27436 16000
rect 27488 15988 27494 16040
rect 27792 16031 27850 16037
rect 27540 16000 27752 16028
rect 22824 15963 22882 15969
rect 22824 15929 22836 15963
rect 22870 15960 22882 15963
rect 23014 15960 23020 15972
rect 22870 15932 23020 15960
rect 22870 15929 22882 15932
rect 22824 15923 22882 15929
rect 23014 15920 23020 15932
rect 23072 15920 23078 15972
rect 23842 15920 23848 15972
rect 23900 15960 23906 15972
rect 27540 15960 27568 16000
rect 23900 15932 27568 15960
rect 27724 15960 27752 16000
rect 27792 15997 27804 16031
rect 27838 16028 27850 16031
rect 28534 16028 28540 16040
rect 27838 16000 28540 16028
rect 27838 15997 27850 16000
rect 27792 15991 27850 15997
rect 28534 15988 28540 16000
rect 28592 15988 28598 16040
rect 28718 15988 28724 16040
rect 28776 16028 28782 16040
rect 29365 16031 29423 16037
rect 29365 16028 29377 16031
rect 28776 16000 29377 16028
rect 28776 15988 28782 16000
rect 29365 15997 29377 16000
rect 29411 15997 29423 16031
rect 30650 16028 30656 16040
rect 30611 16000 30656 16028
rect 29365 15991 29423 15997
rect 30650 15988 30656 16000
rect 30708 15988 30714 16040
rect 31036 16037 31064 16136
rect 31202 16124 31208 16136
rect 31260 16124 31266 16176
rect 32306 16056 32312 16108
rect 32364 16096 32370 16108
rect 32364 16068 32536 16096
rect 32364 16056 32370 16068
rect 30745 16031 30803 16037
rect 30745 15997 30757 16031
rect 30791 15997 30803 16031
rect 30745 15991 30803 15997
rect 31021 16031 31079 16037
rect 31021 15997 31033 16031
rect 31067 15997 31079 16031
rect 31021 15991 31079 15997
rect 29914 15960 29920 15972
rect 27724 15932 29920 15960
rect 23900 15920 23906 15932
rect 29914 15920 29920 15932
rect 29972 15920 29978 15972
rect 1949 15895 2007 15901
rect 1949 15861 1961 15895
rect 1995 15892 2007 15895
rect 16390 15892 16396 15904
rect 1995 15864 16396 15892
rect 1995 15861 2007 15864
rect 1949 15855 2007 15861
rect 16390 15852 16396 15864
rect 16448 15852 16454 15904
rect 26234 15852 26240 15904
rect 26292 15892 26298 15904
rect 26973 15895 27031 15901
rect 26973 15892 26985 15895
rect 26292 15864 26985 15892
rect 26292 15852 26298 15864
rect 26973 15861 26985 15864
rect 27019 15892 27031 15895
rect 27338 15892 27344 15904
rect 27019 15864 27344 15892
rect 27019 15861 27031 15864
rect 26973 15855 27031 15861
rect 27338 15852 27344 15864
rect 27396 15852 27402 15904
rect 27430 15852 27436 15904
rect 27488 15892 27494 15904
rect 28534 15892 28540 15904
rect 27488 15864 28540 15892
rect 27488 15852 27494 15864
rect 28534 15852 28540 15864
rect 28592 15852 28598 15904
rect 28626 15852 28632 15904
rect 28684 15892 28690 15904
rect 28905 15895 28963 15901
rect 28905 15892 28917 15895
rect 28684 15864 28917 15892
rect 28684 15852 28690 15864
rect 28905 15861 28917 15864
rect 28951 15861 28963 15895
rect 30466 15892 30472 15904
rect 30427 15864 30472 15892
rect 28905 15855 28963 15861
rect 30466 15852 30472 15864
rect 30524 15852 30530 15904
rect 30760 15892 30788 15991
rect 31202 15988 31208 16040
rect 31260 16028 31266 16040
rect 31662 16028 31668 16040
rect 31260 16000 31668 16028
rect 31260 15988 31266 16000
rect 31662 15988 31668 16000
rect 31720 15988 31726 16040
rect 32398 16028 32404 16040
rect 32359 16000 32404 16028
rect 32398 15988 32404 16000
rect 32456 15988 32462 16040
rect 32508 16037 32536 16068
rect 33318 16056 33324 16108
rect 33376 16096 33382 16108
rect 33376 16068 33548 16096
rect 33376 16056 33382 16068
rect 32493 16031 32551 16037
rect 32493 15997 32505 16031
rect 32539 15997 32551 16031
rect 32493 15991 32551 15997
rect 32636 16031 32694 16037
rect 32636 15997 32648 16031
rect 32682 15997 32694 16031
rect 32766 16028 32772 16040
rect 32727 16000 32772 16028
rect 32636 15991 32694 15997
rect 31570 15960 31576 15972
rect 31531 15932 31576 15960
rect 31570 15920 31576 15932
rect 31628 15920 31634 15972
rect 31757 15963 31815 15969
rect 31757 15929 31769 15963
rect 31803 15960 31815 15963
rect 32651 15960 32679 15991
rect 32766 15988 32772 16000
rect 32824 15988 32830 16040
rect 33042 15988 33048 16040
rect 33100 16028 33106 16040
rect 33520 16037 33548 16068
rect 33796 16037 33824 16192
rect 34517 16167 34575 16173
rect 34517 16133 34529 16167
rect 34563 16164 34575 16167
rect 34698 16164 34704 16176
rect 34563 16136 34704 16164
rect 34563 16133 34575 16136
rect 34517 16127 34575 16133
rect 34698 16124 34704 16136
rect 34756 16124 34762 16176
rect 33413 16031 33471 16037
rect 33413 16028 33425 16031
rect 33100 16000 33425 16028
rect 33100 15988 33106 16000
rect 33413 15997 33425 16000
rect 33459 15997 33471 16031
rect 33413 15991 33471 15997
rect 33505 16031 33563 16037
rect 33505 15997 33517 16031
rect 33551 15997 33563 16031
rect 33505 15991 33563 15997
rect 33689 16031 33747 16037
rect 33689 15997 33701 16031
rect 33735 15997 33747 16031
rect 33689 15991 33747 15997
rect 33781 16031 33839 16037
rect 33781 15997 33793 16031
rect 33827 15997 33839 16031
rect 37274 16028 37280 16040
rect 37235 16000 37280 16028
rect 33781 15991 33839 15997
rect 33134 15960 33140 15972
rect 31803 15932 33140 15960
rect 31803 15929 31815 15932
rect 31757 15923 31815 15929
rect 33134 15920 33140 15932
rect 33192 15920 33198 15972
rect 33704 15960 33732 15991
rect 37274 15988 37280 16000
rect 37332 15988 37338 16040
rect 37918 16028 37924 16040
rect 37879 16000 37924 16028
rect 37918 15988 37924 16000
rect 37976 15988 37982 16040
rect 33704 15932 33824 15960
rect 33796 15904 33824 15932
rect 33962 15920 33968 15972
rect 34020 15960 34026 15972
rect 34333 15963 34391 15969
rect 34333 15960 34345 15963
rect 34020 15932 34345 15960
rect 34020 15920 34026 15932
rect 34333 15929 34345 15932
rect 34379 15929 34391 15963
rect 34333 15923 34391 15929
rect 32582 15892 32588 15904
rect 30760 15864 32588 15892
rect 32582 15852 32588 15864
rect 32640 15852 32646 15904
rect 33778 15852 33784 15904
rect 33836 15892 33842 15904
rect 34606 15892 34612 15904
rect 33836 15864 34612 15892
rect 33836 15852 33842 15864
rect 34606 15852 34612 15864
rect 34664 15852 34670 15904
rect 1104 15802 38824 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 38824 15802
rect 1104 15728 38824 15750
rect 22646 15648 22652 15700
rect 22704 15688 22710 15700
rect 22741 15691 22799 15697
rect 22741 15688 22753 15691
rect 22704 15660 22753 15688
rect 22704 15648 22710 15660
rect 22741 15657 22753 15660
rect 22787 15657 22799 15691
rect 22741 15651 22799 15657
rect 23658 15648 23664 15700
rect 23716 15688 23722 15700
rect 32766 15688 32772 15700
rect 23716 15660 24624 15688
rect 23716 15648 23722 15660
rect 1854 15552 1860 15564
rect 1815 15524 1860 15552
rect 1854 15512 1860 15524
rect 1912 15512 1918 15564
rect 22922 15552 22928 15564
rect 22883 15524 22928 15552
rect 22922 15512 22928 15524
rect 22980 15512 22986 15564
rect 23566 15552 23572 15564
rect 23527 15524 23572 15552
rect 23566 15512 23572 15524
rect 23624 15512 23630 15564
rect 23661 15555 23719 15561
rect 23661 15521 23673 15555
rect 23707 15552 23719 15555
rect 23842 15552 23848 15564
rect 23707 15524 23848 15552
rect 23707 15521 23719 15524
rect 23661 15515 23719 15521
rect 23842 15512 23848 15524
rect 23900 15512 23906 15564
rect 24596 15561 24624 15660
rect 24688 15660 32772 15688
rect 24688 15561 24716 15660
rect 32766 15648 32772 15660
rect 32824 15648 32830 15700
rect 33318 15648 33324 15700
rect 33376 15648 33382 15700
rect 24762 15580 24768 15632
rect 24820 15620 24826 15632
rect 27890 15620 27896 15632
rect 24820 15592 27896 15620
rect 24820 15580 24826 15592
rect 27890 15580 27896 15592
rect 27948 15580 27954 15632
rect 28068 15623 28126 15629
rect 28068 15589 28080 15623
rect 28114 15620 28126 15623
rect 28994 15620 29000 15632
rect 28114 15592 29000 15620
rect 28114 15589 28126 15592
rect 28068 15583 28126 15589
rect 28994 15580 29000 15592
rect 29052 15580 29058 15632
rect 31386 15620 31392 15632
rect 29932 15592 31392 15620
rect 23937 15555 23995 15561
rect 23937 15521 23949 15555
rect 23983 15521 23995 15555
rect 23937 15515 23995 15521
rect 24581 15555 24639 15561
rect 24581 15521 24593 15555
rect 24627 15521 24639 15555
rect 24581 15515 24639 15521
rect 24673 15555 24731 15561
rect 24673 15521 24685 15555
rect 24719 15521 24731 15555
rect 24673 15515 24731 15521
rect 24949 15555 25007 15561
rect 24949 15521 24961 15555
rect 24995 15552 25007 15555
rect 25406 15552 25412 15564
rect 24995 15524 25268 15552
rect 25367 15524 25412 15552
rect 24995 15521 25007 15524
rect 24949 15515 25007 15521
rect 23952 15484 23980 15515
rect 24210 15484 24216 15496
rect 23952 15456 24216 15484
rect 24210 15444 24216 15456
rect 24268 15484 24274 15496
rect 24964 15484 24992 15515
rect 24268 15456 24992 15484
rect 24268 15444 24274 15456
rect 1949 15351 2007 15357
rect 1949 15317 1961 15351
rect 1995 15348 2007 15351
rect 16114 15348 16120 15360
rect 1995 15320 16120 15348
rect 1995 15317 2007 15320
rect 1949 15311 2007 15317
rect 16114 15308 16120 15320
rect 16172 15308 16178 15360
rect 23198 15308 23204 15360
rect 23256 15348 23262 15360
rect 23385 15351 23443 15357
rect 23385 15348 23397 15351
rect 23256 15320 23397 15348
rect 23256 15308 23262 15320
rect 23385 15317 23397 15320
rect 23431 15317 23443 15351
rect 23842 15348 23848 15360
rect 23803 15320 23848 15348
rect 23385 15311 23443 15317
rect 23842 15308 23848 15320
rect 23900 15308 23906 15360
rect 24394 15348 24400 15360
rect 24355 15320 24400 15348
rect 24394 15308 24400 15320
rect 24452 15308 24458 15360
rect 24854 15348 24860 15360
rect 24815 15320 24860 15348
rect 24854 15308 24860 15320
rect 24912 15308 24918 15360
rect 25240 15348 25268 15524
rect 25406 15512 25412 15524
rect 25464 15512 25470 15564
rect 25676 15555 25734 15561
rect 25676 15521 25688 15555
rect 25722 15552 25734 15555
rect 28350 15552 28356 15564
rect 25722 15524 28356 15552
rect 25722 15521 25734 15524
rect 25676 15515 25734 15521
rect 28350 15512 28356 15524
rect 28408 15512 28414 15564
rect 29822 15552 29828 15564
rect 29783 15524 29828 15552
rect 29822 15512 29828 15524
rect 29880 15512 29886 15564
rect 29932 15561 29960 15592
rect 31386 15580 31392 15592
rect 31444 15580 31450 15632
rect 33336 15620 33364 15648
rect 34054 15620 34060 15632
rect 33336 15592 34060 15620
rect 29917 15555 29975 15561
rect 29917 15521 29929 15555
rect 29963 15521 29975 15555
rect 30190 15552 30196 15564
rect 30151 15524 30196 15552
rect 29917 15515 29975 15521
rect 30190 15512 30196 15524
rect 30248 15512 30254 15564
rect 30834 15552 30840 15564
rect 30795 15524 30840 15552
rect 30834 15512 30840 15524
rect 30892 15512 30898 15564
rect 30975 15555 31033 15561
rect 30975 15521 30987 15555
rect 31021 15552 31033 15555
rect 31205 15555 31263 15561
rect 31021 15524 31156 15552
rect 31021 15521 31033 15524
rect 30975 15515 31033 15521
rect 27522 15444 27528 15496
rect 27580 15484 27586 15496
rect 27801 15487 27859 15493
rect 27801 15484 27813 15487
rect 27580 15456 27813 15484
rect 27580 15444 27586 15456
rect 27801 15453 27813 15456
rect 27847 15453 27859 15487
rect 30101 15487 30159 15493
rect 30101 15484 30113 15487
rect 27801 15447 27859 15453
rect 28828 15456 30113 15484
rect 27154 15416 27160 15428
rect 26344 15388 27160 15416
rect 26344 15348 26372 15388
rect 27154 15376 27160 15388
rect 27212 15376 27218 15428
rect 25240 15320 26372 15348
rect 26602 15308 26608 15360
rect 26660 15348 26666 15360
rect 26789 15351 26847 15357
rect 26789 15348 26801 15351
rect 26660 15320 26801 15348
rect 26660 15308 26666 15320
rect 26789 15317 26801 15320
rect 26835 15317 26847 15351
rect 26789 15311 26847 15317
rect 28442 15308 28448 15360
rect 28500 15348 28506 15360
rect 28828 15348 28856 15456
rect 30101 15453 30113 15456
rect 30147 15453 30159 15487
rect 31128 15484 31156 15524
rect 31205 15521 31217 15555
rect 31251 15552 31263 15555
rect 31846 15552 31852 15564
rect 31251 15524 31852 15552
rect 31251 15521 31263 15524
rect 31205 15515 31263 15521
rect 31846 15512 31852 15524
rect 31904 15512 31910 15564
rect 32950 15512 32956 15564
rect 33008 15552 33014 15564
rect 33428 15561 33456 15592
rect 34054 15580 34060 15592
rect 34112 15580 34118 15632
rect 34238 15620 34244 15632
rect 34164 15592 34244 15620
rect 33321 15555 33379 15561
rect 33321 15552 33333 15555
rect 33008 15524 33333 15552
rect 33008 15512 33014 15524
rect 33321 15521 33333 15524
rect 33367 15521 33379 15555
rect 33321 15515 33379 15521
rect 33413 15555 33471 15561
rect 33413 15521 33425 15555
rect 33459 15521 33471 15555
rect 33413 15515 33471 15521
rect 33597 15555 33655 15561
rect 33597 15521 33609 15555
rect 33643 15521 33655 15555
rect 33597 15515 33655 15521
rect 33689 15555 33747 15561
rect 33689 15521 33701 15555
rect 33735 15552 33747 15555
rect 34164 15552 34192 15592
rect 34238 15580 34244 15592
rect 34296 15580 34302 15632
rect 34330 15552 34336 15564
rect 33735 15524 34192 15552
rect 34243 15524 34336 15552
rect 33735 15521 33747 15524
rect 33689 15515 33747 15521
rect 32582 15484 32588 15496
rect 31128 15456 32588 15484
rect 30101 15447 30159 15453
rect 32582 15444 32588 15456
rect 32640 15444 32646 15496
rect 28902 15376 28908 15428
rect 28960 15416 28966 15428
rect 29641 15419 29699 15425
rect 29641 15416 29653 15419
rect 28960 15388 29653 15416
rect 28960 15376 28966 15388
rect 29641 15385 29653 15388
rect 29687 15385 29699 15419
rect 29641 15379 29699 15385
rect 31113 15419 31171 15425
rect 31113 15385 31125 15419
rect 31159 15416 31171 15419
rect 31386 15416 31392 15428
rect 31159 15388 31392 15416
rect 31159 15385 31171 15388
rect 31113 15379 31171 15385
rect 31386 15376 31392 15388
rect 31444 15376 31450 15428
rect 28500 15320 28856 15348
rect 28500 15308 28506 15320
rect 28994 15308 29000 15360
rect 29052 15348 29058 15360
rect 29181 15351 29239 15357
rect 29181 15348 29193 15351
rect 29052 15320 29193 15348
rect 29052 15308 29058 15320
rect 29181 15317 29193 15320
rect 29227 15348 29239 15351
rect 29454 15348 29460 15360
rect 29227 15320 29460 15348
rect 29227 15317 29239 15320
rect 29181 15311 29239 15317
rect 29454 15308 29460 15320
rect 29512 15308 29518 15360
rect 29730 15308 29736 15360
rect 29788 15348 29794 15360
rect 30653 15351 30711 15357
rect 30653 15348 30665 15351
rect 29788 15320 30665 15348
rect 29788 15308 29794 15320
rect 30653 15317 30665 15320
rect 30699 15317 30711 15351
rect 33134 15348 33140 15360
rect 33095 15320 33140 15348
rect 30653 15311 30711 15317
rect 33134 15308 33140 15320
rect 33192 15308 33198 15360
rect 33612 15348 33640 15515
rect 34330 15512 34336 15524
rect 34388 15512 34394 15564
rect 34425 15555 34483 15561
rect 34425 15521 34437 15555
rect 34471 15521 34483 15555
rect 34606 15552 34612 15564
rect 34567 15524 34612 15552
rect 34425 15515 34483 15521
rect 34238 15376 34244 15428
rect 34296 15416 34302 15428
rect 34348 15416 34376 15512
rect 34440 15484 34468 15515
rect 34606 15512 34612 15524
rect 34664 15512 34670 15564
rect 34701 15555 34759 15561
rect 34701 15521 34713 15555
rect 34747 15552 34759 15555
rect 35618 15552 35624 15564
rect 34747 15524 35624 15552
rect 34747 15521 34759 15524
rect 34701 15515 34759 15521
rect 35618 15512 35624 15524
rect 35676 15512 35682 15564
rect 37182 15552 37188 15564
rect 37143 15524 37188 15552
rect 37182 15512 37188 15524
rect 37240 15512 37246 15564
rect 35434 15484 35440 15496
rect 34440 15456 35440 15484
rect 35434 15444 35440 15456
rect 35492 15444 35498 15496
rect 35894 15416 35900 15428
rect 34296 15388 35900 15416
rect 34296 15376 34302 15388
rect 35894 15376 35900 15388
rect 35952 15376 35958 15428
rect 33778 15348 33784 15360
rect 33612 15320 33784 15348
rect 33778 15308 33784 15320
rect 33836 15308 33842 15360
rect 33962 15308 33968 15360
rect 34020 15348 34026 15360
rect 34149 15351 34207 15357
rect 34149 15348 34161 15351
rect 34020 15320 34161 15348
rect 34020 15308 34026 15320
rect 34149 15317 34161 15320
rect 34195 15317 34207 15351
rect 34149 15311 34207 15317
rect 1104 15258 38824 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 38824 15258
rect 1104 15184 38824 15206
rect 23032 15116 26740 15144
rect 22830 14900 22836 14952
rect 22888 14940 22894 14952
rect 23032 14949 23060 15116
rect 23201 15079 23259 15085
rect 23201 15045 23213 15079
rect 23247 15076 23259 15079
rect 23290 15076 23296 15088
rect 23247 15048 23296 15076
rect 23247 15045 23259 15048
rect 23201 15039 23259 15045
rect 23290 15036 23296 15048
rect 23348 15036 23354 15088
rect 23934 15036 23940 15088
rect 23992 15076 23998 15088
rect 24213 15079 24271 15085
rect 24213 15076 24225 15079
rect 23992 15048 24225 15076
rect 23992 15036 23998 15048
rect 24213 15045 24225 15048
rect 24259 15045 24271 15079
rect 24213 15039 24271 15045
rect 24302 15036 24308 15088
rect 24360 15076 24366 15088
rect 26712 15076 26740 15116
rect 27890 15104 27896 15156
rect 27948 15144 27954 15156
rect 28902 15144 28908 15156
rect 27948 15116 28908 15144
rect 27948 15104 27954 15116
rect 28902 15104 28908 15116
rect 28960 15104 28966 15156
rect 31662 15144 31668 15156
rect 29104 15116 31668 15144
rect 29104 15076 29132 15116
rect 31662 15104 31668 15116
rect 31720 15104 31726 15156
rect 32582 15104 32588 15156
rect 32640 15144 32646 15156
rect 33965 15147 34023 15153
rect 33965 15144 33977 15147
rect 32640 15116 33977 15144
rect 32640 15104 32646 15116
rect 33965 15113 33977 15116
rect 34011 15113 34023 15147
rect 35894 15144 35900 15156
rect 35855 15116 35900 15144
rect 33965 15107 34023 15113
rect 35894 15104 35900 15116
rect 35952 15104 35958 15156
rect 29457 15079 29515 15085
rect 29457 15076 29469 15079
rect 24360 15048 25268 15076
rect 26712 15048 29132 15076
rect 29196 15048 29469 15076
rect 24360 15036 24366 15048
rect 24486 15008 24492 15020
rect 24044 14980 24492 15008
rect 22925 14943 22983 14949
rect 22925 14940 22937 14943
rect 22888 14912 22937 14940
rect 22888 14900 22894 14912
rect 22925 14909 22937 14912
rect 22971 14909 22983 14943
rect 22925 14903 22983 14909
rect 23017 14943 23075 14949
rect 23017 14909 23029 14943
rect 23063 14909 23075 14943
rect 23017 14903 23075 14909
rect 23293 14943 23351 14949
rect 23293 14909 23305 14943
rect 23339 14940 23351 14943
rect 23566 14940 23572 14952
rect 23339 14912 23572 14940
rect 23339 14909 23351 14912
rect 23293 14903 23351 14909
rect 23566 14900 23572 14912
rect 23624 14900 23630 14952
rect 23750 14900 23756 14952
rect 23808 14940 23814 14952
rect 24044 14949 24072 14980
rect 24486 14968 24492 14980
rect 24544 14968 24550 15020
rect 25240 15017 25268 15048
rect 25225 15011 25283 15017
rect 25225 14977 25237 15011
rect 25271 14977 25283 15011
rect 25225 14971 25283 14977
rect 26602 14968 26608 15020
rect 26660 15008 26666 15020
rect 29196 15008 29224 15048
rect 29457 15045 29469 15048
rect 29503 15045 29515 15079
rect 29457 15039 29515 15045
rect 32122 15036 32128 15088
rect 32180 15036 32186 15088
rect 36078 15076 36084 15088
rect 34072 15048 36084 15076
rect 32140 15008 32168 15036
rect 26660 14980 29224 15008
rect 29288 14980 32168 15008
rect 26660 14968 26666 14980
rect 23937 14943 23995 14949
rect 23937 14940 23949 14943
rect 23808 14912 23949 14940
rect 23808 14900 23814 14912
rect 23937 14909 23949 14912
rect 23983 14909 23995 14943
rect 23937 14903 23995 14909
rect 24029 14943 24087 14949
rect 24029 14909 24041 14943
rect 24075 14909 24087 14943
rect 24029 14903 24087 14909
rect 24210 14900 24216 14952
rect 24268 14940 24274 14952
rect 24305 14943 24363 14949
rect 24305 14940 24317 14943
rect 24268 14912 24317 14940
rect 24268 14900 24274 14912
rect 24305 14909 24317 14912
rect 24351 14909 24363 14943
rect 24305 14903 24363 14909
rect 26970 14900 26976 14952
rect 27028 14940 27034 14952
rect 27249 14943 27307 14949
rect 27249 14940 27261 14943
rect 27028 14912 27261 14940
rect 27028 14900 27034 14912
rect 27249 14909 27261 14912
rect 27295 14940 27307 14943
rect 27338 14940 27344 14952
rect 27295 14912 27344 14940
rect 27295 14909 27307 14912
rect 27249 14903 27307 14909
rect 27338 14900 27344 14912
rect 27396 14900 27402 14952
rect 27430 14900 27436 14952
rect 27488 14940 27494 14952
rect 28077 14943 28135 14949
rect 28077 14940 28089 14943
rect 27488 14912 28089 14940
rect 27488 14900 27494 14912
rect 28077 14909 28089 14912
rect 28123 14909 28135 14943
rect 28077 14903 28135 14909
rect 28445 14943 28503 14949
rect 28445 14909 28457 14943
rect 28491 14940 28503 14943
rect 28902 14940 28908 14952
rect 28491 14912 28908 14940
rect 28491 14909 28503 14912
rect 28445 14903 28503 14909
rect 28902 14900 28908 14912
rect 28960 14900 28966 14952
rect 29178 14940 29184 14952
rect 29139 14912 29184 14940
rect 29178 14900 29184 14912
rect 29236 14900 29242 14952
rect 29288 14949 29316 14980
rect 32766 14968 32772 15020
rect 32824 15008 32830 15020
rect 32953 15011 33011 15017
rect 32953 15008 32965 15011
rect 32824 14980 32965 15008
rect 32824 14968 32830 14980
rect 32953 14977 32965 14980
rect 32999 14977 33011 15011
rect 34072 15008 34100 15048
rect 36078 15036 36084 15048
rect 36136 15036 36142 15088
rect 35894 15008 35900 15020
rect 32953 14971 33011 14977
rect 33152 14980 34100 15008
rect 34164 14980 35900 15008
rect 29273 14943 29331 14949
rect 29273 14909 29285 14943
rect 29319 14909 29331 14943
rect 29273 14903 29331 14909
rect 29549 14943 29607 14949
rect 29549 14909 29561 14943
rect 29595 14940 29607 14943
rect 30190 14940 30196 14952
rect 29595 14912 30196 14940
rect 29595 14909 29607 14912
rect 29549 14903 29607 14909
rect 30190 14900 30196 14912
rect 30248 14900 30254 14952
rect 32125 14943 32183 14949
rect 32125 14909 32137 14943
rect 32171 14909 32183 14943
rect 32125 14903 32183 14909
rect 32217 14943 32275 14949
rect 32217 14909 32229 14943
rect 32263 14909 32275 14943
rect 32217 14903 32275 14909
rect 14090 14832 14096 14884
rect 14148 14872 14154 14884
rect 25314 14872 25320 14884
rect 14148 14844 25320 14872
rect 14148 14832 14154 14844
rect 25314 14832 25320 14844
rect 25372 14832 25378 14884
rect 25492 14875 25550 14881
rect 25492 14841 25504 14875
rect 25538 14872 25550 14875
rect 30466 14872 30472 14884
rect 25538 14844 30472 14872
rect 25538 14841 25550 14844
rect 25492 14835 25550 14841
rect 30466 14832 30472 14844
rect 30524 14832 30530 14884
rect 22738 14804 22744 14816
rect 22699 14776 22744 14804
rect 22738 14764 22744 14776
rect 22796 14764 22802 14816
rect 23750 14804 23756 14816
rect 23711 14776 23756 14804
rect 23750 14764 23756 14776
rect 23808 14764 23814 14816
rect 25682 14764 25688 14816
rect 25740 14804 25746 14816
rect 26605 14807 26663 14813
rect 26605 14804 26617 14807
rect 25740 14776 26617 14804
rect 25740 14764 25746 14776
rect 26605 14773 26617 14776
rect 26651 14804 26663 14807
rect 26786 14804 26792 14816
rect 26651 14776 26792 14804
rect 26651 14773 26663 14776
rect 26605 14767 26663 14773
rect 26786 14764 26792 14776
rect 26844 14764 26850 14816
rect 28350 14764 28356 14816
rect 28408 14804 28414 14816
rect 28997 14807 29055 14813
rect 28997 14804 29009 14807
rect 28408 14776 29009 14804
rect 28408 14764 28414 14776
rect 28997 14773 29009 14776
rect 29043 14773 29055 14807
rect 31938 14804 31944 14816
rect 31899 14776 31944 14804
rect 28997 14767 29055 14773
rect 31938 14764 31944 14776
rect 31996 14764 32002 14816
rect 32140 14804 32168 14903
rect 32232 14872 32260 14903
rect 32306 14900 32312 14952
rect 32364 14940 32370 14952
rect 32401 14943 32459 14949
rect 32401 14940 32413 14943
rect 32364 14912 32413 14940
rect 32364 14900 32370 14912
rect 32401 14909 32413 14912
rect 32447 14909 32459 14943
rect 32401 14903 32459 14909
rect 32493 14943 32551 14949
rect 32493 14909 32505 14943
rect 32539 14940 32551 14943
rect 32858 14940 32864 14952
rect 32539 14912 32864 14940
rect 32539 14909 32551 14912
rect 32493 14903 32551 14909
rect 32858 14900 32864 14912
rect 32916 14900 32922 14952
rect 33152 14949 33180 14980
rect 33137 14943 33195 14949
rect 33137 14909 33149 14943
rect 33183 14909 33195 14943
rect 33137 14903 33195 14909
rect 33229 14943 33287 14949
rect 33229 14909 33241 14943
rect 33275 14940 33287 14943
rect 33318 14940 33324 14952
rect 33275 14912 33324 14940
rect 33275 14909 33287 14912
rect 33229 14903 33287 14909
rect 33244 14872 33272 14903
rect 33318 14900 33324 14912
rect 33376 14900 33382 14952
rect 33413 14943 33471 14949
rect 33413 14909 33425 14943
rect 33459 14909 33471 14943
rect 33413 14903 33471 14909
rect 32232 14844 33272 14872
rect 33428 14872 33456 14903
rect 33502 14900 33508 14952
rect 33560 14940 33566 14952
rect 34164 14949 34192 14980
rect 35894 14968 35900 14980
rect 35952 14968 35958 15020
rect 34149 14943 34207 14949
rect 33560 14912 33605 14940
rect 33560 14900 33566 14912
rect 34149 14909 34161 14943
rect 34195 14909 34207 14943
rect 34149 14903 34207 14909
rect 34238 14900 34244 14952
rect 34296 14940 34302 14952
rect 34425 14943 34483 14949
rect 34296 14912 34341 14940
rect 34296 14900 34302 14912
rect 34425 14909 34437 14943
rect 34471 14909 34483 14943
rect 34425 14903 34483 14909
rect 34517 14943 34575 14949
rect 34517 14909 34529 14943
rect 34563 14940 34575 14943
rect 35526 14940 35532 14952
rect 34563 14912 35532 14940
rect 34563 14909 34575 14912
rect 34517 14903 34575 14909
rect 33778 14872 33784 14884
rect 33428 14844 33784 14872
rect 33778 14832 33784 14844
rect 33836 14832 33842 14884
rect 34440 14872 34468 14903
rect 35526 14900 35532 14912
rect 35584 14900 35590 14952
rect 37918 14940 37924 14952
rect 37879 14912 37924 14940
rect 37918 14900 37924 14912
rect 37976 14900 37982 14952
rect 34606 14872 34612 14884
rect 34440 14844 34612 14872
rect 34606 14832 34612 14844
rect 34664 14832 34670 14884
rect 35805 14875 35863 14881
rect 35805 14841 35817 14875
rect 35851 14841 35863 14875
rect 35805 14835 35863 14841
rect 33502 14804 33508 14816
rect 32140 14776 33508 14804
rect 33502 14764 33508 14776
rect 33560 14764 33566 14816
rect 34330 14764 34336 14816
rect 34388 14804 34394 14816
rect 35820 14804 35848 14835
rect 34388 14776 35848 14804
rect 34388 14764 34394 14776
rect 1104 14714 38824 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 38824 14714
rect 1104 14640 38824 14662
rect 23474 14600 23480 14612
rect 23435 14572 23480 14600
rect 23474 14560 23480 14572
rect 23532 14560 23538 14612
rect 23566 14560 23572 14612
rect 23624 14600 23630 14612
rect 24302 14600 24308 14612
rect 23624 14572 24308 14600
rect 23624 14560 23630 14572
rect 1854 14532 1860 14544
rect 1815 14504 1860 14532
rect 1854 14492 1860 14504
rect 1912 14492 1918 14544
rect 14918 14492 14924 14544
rect 14976 14532 14982 14544
rect 14976 14504 23980 14532
rect 14976 14492 14982 14504
rect 3050 14424 3056 14476
rect 3108 14464 3114 14476
rect 23014 14464 23020 14476
rect 3108 14436 23020 14464
rect 3108 14424 3114 14436
rect 23014 14424 23020 14436
rect 23072 14464 23078 14476
rect 23385 14467 23443 14473
rect 23385 14464 23397 14467
rect 23072 14436 23397 14464
rect 23072 14424 23078 14436
rect 23385 14433 23397 14436
rect 23431 14464 23443 14467
rect 23474 14464 23480 14476
rect 23431 14436 23480 14464
rect 23431 14433 23443 14436
rect 23385 14427 23443 14433
rect 23474 14424 23480 14436
rect 23532 14424 23538 14476
rect 18690 14356 18696 14408
rect 18748 14396 18754 14408
rect 23658 14396 23664 14408
rect 18748 14368 23664 14396
rect 18748 14356 18754 14368
rect 23658 14356 23664 14368
rect 23716 14356 23722 14408
rect 1949 14263 2007 14269
rect 1949 14229 1961 14263
rect 1995 14260 2007 14263
rect 15470 14260 15476 14272
rect 1995 14232 15476 14260
rect 1995 14229 2007 14232
rect 1949 14223 2007 14229
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 23952 14260 23980 14504
rect 24044 14473 24072 14572
rect 24302 14560 24308 14572
rect 24360 14560 24366 14612
rect 33134 14600 33140 14612
rect 24596 14572 26372 14600
rect 24029 14467 24087 14473
rect 24029 14433 24041 14467
rect 24075 14433 24087 14467
rect 24029 14427 24087 14433
rect 24296 14467 24354 14473
rect 24296 14433 24308 14467
rect 24342 14464 24354 14467
rect 24596 14464 24624 14572
rect 24342 14436 24624 14464
rect 24342 14433 24354 14436
rect 24296 14427 24354 14433
rect 24670 14424 24676 14476
rect 24728 14464 24734 14476
rect 26234 14464 26240 14476
rect 24728 14436 26240 14464
rect 24728 14424 24734 14436
rect 26234 14424 26240 14436
rect 26292 14424 26298 14476
rect 26344 14396 26372 14572
rect 26620 14572 33140 14600
rect 26510 14464 26516 14476
rect 26471 14436 26516 14464
rect 26510 14424 26516 14436
rect 26568 14424 26574 14476
rect 26620 14473 26648 14572
rect 33134 14560 33140 14572
rect 33192 14560 33198 14612
rect 33778 14600 33784 14612
rect 33520 14572 33784 14600
rect 27154 14532 27160 14544
rect 26896 14504 27160 14532
rect 26896 14473 26924 14504
rect 27154 14492 27160 14504
rect 27212 14492 27218 14544
rect 28068 14535 28126 14541
rect 28068 14501 28080 14535
rect 28114 14532 28126 14535
rect 29362 14532 29368 14544
rect 28114 14504 29368 14532
rect 28114 14501 28126 14504
rect 28068 14495 28126 14501
rect 29362 14492 29368 14504
rect 29420 14492 29426 14544
rect 29730 14532 29736 14544
rect 29643 14504 29736 14532
rect 29730 14492 29736 14504
rect 29788 14532 29794 14544
rect 31570 14532 31576 14544
rect 29788 14504 31576 14532
rect 29788 14492 29794 14504
rect 31570 14492 31576 14504
rect 31628 14492 31634 14544
rect 26605 14467 26663 14473
rect 26605 14433 26617 14467
rect 26651 14433 26663 14467
rect 26605 14427 26663 14433
rect 26881 14467 26939 14473
rect 26881 14433 26893 14467
rect 26927 14433 26939 14467
rect 29270 14464 29276 14476
rect 26881 14427 26939 14433
rect 26988 14436 29276 14464
rect 26988 14396 27016 14436
rect 29270 14424 29276 14436
rect 29328 14424 29334 14476
rect 29914 14424 29920 14476
rect 29972 14464 29978 14476
rect 33045 14467 33103 14473
rect 33045 14464 33057 14467
rect 29972 14436 33057 14464
rect 29972 14424 29978 14436
rect 33045 14433 33057 14436
rect 33091 14433 33103 14467
rect 33045 14427 33103 14433
rect 33229 14467 33287 14473
rect 33229 14433 33241 14467
rect 33275 14433 33287 14467
rect 33229 14427 33287 14433
rect 26344 14368 27016 14396
rect 27522 14356 27528 14408
rect 27580 14396 27586 14408
rect 27801 14399 27859 14405
rect 27801 14396 27813 14399
rect 27580 14368 27813 14396
rect 27580 14356 27586 14368
rect 27801 14365 27813 14368
rect 27847 14365 27859 14399
rect 27801 14359 27859 14365
rect 29178 14356 29184 14408
rect 29236 14396 29242 14408
rect 30282 14396 30288 14408
rect 29236 14368 30288 14396
rect 29236 14356 29242 14368
rect 30282 14356 30288 14368
rect 30340 14356 30346 14408
rect 33244 14396 33272 14427
rect 33318 14424 33324 14476
rect 33376 14464 33382 14476
rect 33520 14473 33548 14572
rect 33778 14560 33784 14572
rect 33836 14560 33842 14612
rect 34606 14560 34612 14612
rect 34664 14560 34670 14612
rect 37369 14603 37427 14609
rect 37369 14569 37381 14603
rect 37415 14600 37427 14603
rect 38010 14600 38016 14612
rect 37415 14572 38016 14600
rect 37415 14569 37427 14572
rect 37369 14563 37427 14569
rect 38010 14560 38016 14572
rect 38068 14560 38074 14612
rect 34624 14532 34652 14560
rect 34532 14504 34652 14532
rect 33505 14467 33563 14473
rect 33376 14436 33421 14464
rect 33376 14424 33382 14436
rect 33505 14433 33517 14467
rect 33551 14433 33563 14467
rect 33505 14427 33563 14433
rect 33244 14368 33364 14396
rect 33336 14340 33364 14368
rect 25314 14288 25320 14340
rect 25372 14328 25378 14340
rect 25409 14331 25467 14337
rect 25409 14328 25421 14331
rect 25372 14300 25421 14328
rect 25372 14288 25378 14300
rect 25409 14297 25421 14300
rect 25455 14328 25467 14331
rect 31846 14328 31852 14340
rect 25455 14300 26924 14328
rect 25455 14297 25467 14300
rect 25409 14291 25467 14297
rect 24670 14260 24676 14272
rect 23952 14232 24676 14260
rect 24670 14220 24676 14232
rect 24728 14220 24734 14272
rect 26326 14260 26332 14272
rect 26287 14232 26332 14260
rect 26326 14220 26332 14232
rect 26384 14220 26390 14272
rect 26786 14260 26792 14272
rect 26747 14232 26792 14260
rect 26786 14220 26792 14232
rect 26844 14220 26850 14272
rect 26896 14260 26924 14300
rect 28736 14300 31852 14328
rect 28736 14260 28764 14300
rect 31846 14288 31852 14300
rect 31904 14288 31910 14340
rect 32674 14288 32680 14340
rect 32732 14328 32738 14340
rect 33226 14328 33232 14340
rect 32732 14300 33232 14328
rect 32732 14288 32738 14300
rect 33226 14288 33232 14300
rect 33284 14288 33290 14340
rect 33318 14288 33324 14340
rect 33376 14288 33382 14340
rect 29178 14260 29184 14272
rect 26896 14232 28764 14260
rect 29139 14232 29184 14260
rect 29178 14220 29184 14232
rect 29236 14220 29242 14272
rect 29825 14263 29883 14269
rect 29825 14229 29837 14263
rect 29871 14260 29883 14263
rect 33520 14260 33548 14427
rect 33594 14424 33600 14476
rect 33652 14464 33658 14476
rect 33652 14436 33697 14464
rect 33652 14424 33658 14436
rect 33778 14424 33784 14476
rect 33836 14464 33842 14476
rect 34241 14467 34299 14473
rect 34241 14464 34253 14467
rect 33836 14436 34253 14464
rect 33836 14424 33842 14436
rect 34241 14433 34253 14436
rect 34287 14433 34299 14467
rect 34241 14427 34299 14433
rect 34330 14424 34336 14476
rect 34388 14464 34394 14476
rect 34532 14473 34560 14504
rect 34517 14467 34575 14473
rect 34388 14436 34433 14464
rect 34388 14424 34394 14436
rect 34517 14433 34529 14467
rect 34563 14433 34575 14467
rect 34517 14427 34575 14433
rect 34609 14467 34667 14473
rect 34609 14433 34621 14467
rect 34655 14464 34667 14467
rect 35710 14464 35716 14476
rect 34655 14436 35716 14464
rect 34655 14433 34667 14436
rect 34609 14427 34667 14433
rect 35710 14424 35716 14436
rect 35768 14424 35774 14476
rect 37182 14464 37188 14476
rect 37143 14436 37188 14464
rect 37182 14424 37188 14436
rect 37240 14424 37246 14476
rect 34054 14260 34060 14272
rect 29871 14232 33548 14260
rect 34015 14232 34060 14260
rect 29871 14229 29883 14232
rect 29825 14223 29883 14229
rect 34054 14220 34060 14232
rect 34112 14220 34118 14272
rect 1104 14170 38824 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 38824 14170
rect 1104 14096 38824 14118
rect 2133 14059 2191 14065
rect 2133 14025 2145 14059
rect 2179 14056 2191 14059
rect 2222 14056 2228 14068
rect 2179 14028 2228 14056
rect 2179 14025 2191 14028
rect 2133 14019 2191 14025
rect 2222 14016 2228 14028
rect 2280 14016 2286 14068
rect 23566 14056 23572 14068
rect 22940 14028 23572 14056
rect 22554 13880 22560 13932
rect 22612 13920 22618 13932
rect 22940 13929 22968 14028
rect 23566 14016 23572 14028
rect 23624 14016 23630 14068
rect 23842 14016 23848 14068
rect 23900 14056 23906 14068
rect 24302 14056 24308 14068
rect 23900 14028 24308 14056
rect 23900 14016 23906 14028
rect 24302 14016 24308 14028
rect 24360 14016 24366 14068
rect 24486 14016 24492 14068
rect 24544 14056 24550 14068
rect 28442 14056 28448 14068
rect 24544 14028 28028 14056
rect 28403 14028 28448 14056
rect 24544 14016 24550 14028
rect 26234 13948 26240 14000
rect 26292 13988 26298 14000
rect 26605 13991 26663 13997
rect 26605 13988 26617 13991
rect 26292 13960 26617 13988
rect 26292 13948 26298 13960
rect 26605 13957 26617 13960
rect 26651 13957 26663 13991
rect 28000 13988 28028 14028
rect 28442 14016 28448 14028
rect 28500 14016 28506 14068
rect 28534 14016 28540 14068
rect 28592 14056 28598 14068
rect 29273 14059 29331 14065
rect 29273 14056 29285 14059
rect 28592 14028 29285 14056
rect 28592 14016 28598 14028
rect 29273 14025 29285 14028
rect 29319 14025 29331 14059
rect 32861 14059 32919 14065
rect 32861 14056 32873 14059
rect 29273 14019 29331 14025
rect 31726 14028 32873 14056
rect 31726 13988 31754 14028
rect 32861 14025 32873 14028
rect 32907 14025 32919 14059
rect 32861 14019 32919 14025
rect 33962 14016 33968 14068
rect 34020 14056 34026 14068
rect 34149 14059 34207 14065
rect 34149 14056 34161 14059
rect 34020 14028 34161 14056
rect 34020 14016 34026 14028
rect 34149 14025 34161 14028
rect 34195 14025 34207 14059
rect 34149 14019 34207 14025
rect 34330 14016 34336 14068
rect 34388 14056 34394 14068
rect 34793 14059 34851 14065
rect 34793 14056 34805 14059
rect 34388 14028 34805 14056
rect 34388 14016 34394 14028
rect 34793 14025 34805 14028
rect 34839 14025 34851 14059
rect 34793 14019 34851 14025
rect 38105 14059 38163 14065
rect 38105 14025 38117 14059
rect 38151 14056 38163 14059
rect 38746 14056 38752 14068
rect 38151 14028 38752 14056
rect 38151 14025 38163 14028
rect 38105 14019 38163 14025
rect 38746 14016 38752 14028
rect 38804 14016 38810 14068
rect 34606 13988 34612 14000
rect 28000 13960 31754 13988
rect 32876 13960 34612 13988
rect 26605 13951 26663 13957
rect 22925 13923 22983 13929
rect 22925 13920 22937 13923
rect 22612 13892 22937 13920
rect 22612 13880 22618 13892
rect 22925 13889 22937 13892
rect 22971 13889 22983 13923
rect 22925 13883 22983 13889
rect 24026 13880 24032 13932
rect 24084 13920 24090 13932
rect 24084 13892 25360 13920
rect 24084 13880 24090 13892
rect 1854 13852 1860 13864
rect 1815 13824 1860 13852
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 23198 13861 23204 13864
rect 23192 13852 23204 13861
rect 23159 13824 23204 13852
rect 23192 13815 23204 13824
rect 23198 13812 23204 13815
rect 23256 13812 23262 13864
rect 25222 13852 25228 13864
rect 25183 13824 25228 13852
rect 25222 13812 25228 13824
rect 25280 13812 25286 13864
rect 25332 13852 25360 13892
rect 28810 13880 28816 13932
rect 28868 13920 28874 13932
rect 28905 13923 28963 13929
rect 28905 13920 28917 13923
rect 28868 13892 28917 13920
rect 28868 13880 28874 13892
rect 28905 13889 28917 13892
rect 28951 13889 28963 13923
rect 28905 13883 28963 13889
rect 25481 13855 25539 13861
rect 25481 13852 25493 13855
rect 25332 13824 25493 13852
rect 25481 13821 25493 13824
rect 25527 13821 25539 13855
rect 25481 13815 25539 13821
rect 26234 13812 26240 13864
rect 26292 13852 26298 13864
rect 27065 13855 27123 13861
rect 27065 13852 27077 13855
rect 26292 13824 27077 13852
rect 26292 13812 26298 13824
rect 26896 13796 26924 13824
rect 27065 13821 27077 13824
rect 27111 13821 27123 13855
rect 27065 13815 27123 13821
rect 27332 13855 27390 13861
rect 27332 13821 27344 13855
rect 27378 13852 27390 13855
rect 27890 13852 27896 13864
rect 27378 13824 27896 13852
rect 27378 13821 27390 13824
rect 27332 13815 27390 13821
rect 27890 13812 27896 13824
rect 27948 13812 27954 13864
rect 29089 13855 29147 13861
rect 29089 13852 29101 13855
rect 28000 13824 29101 13852
rect 20898 13744 20904 13796
rect 20956 13784 20962 13796
rect 20956 13756 26648 13784
rect 20956 13744 20962 13756
rect 21082 13676 21088 13728
rect 21140 13716 21146 13728
rect 22278 13716 22284 13728
rect 21140 13688 22284 13716
rect 21140 13676 21146 13688
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 22370 13676 22376 13728
rect 22428 13716 22434 13728
rect 26510 13716 26516 13728
rect 22428 13688 26516 13716
rect 22428 13676 22434 13688
rect 26510 13676 26516 13688
rect 26568 13676 26574 13728
rect 26620 13716 26648 13756
rect 26878 13744 26884 13796
rect 26936 13744 26942 13796
rect 28000 13716 28028 13824
rect 29089 13821 29101 13824
rect 29135 13821 29147 13855
rect 29730 13852 29736 13864
rect 29089 13815 29147 13821
rect 29196 13824 29736 13852
rect 26620 13688 28028 13716
rect 28258 13676 28264 13728
rect 28316 13716 28322 13728
rect 28442 13716 28448 13728
rect 28316 13688 28448 13716
rect 28316 13676 28322 13688
rect 28442 13676 28448 13688
rect 28500 13676 28506 13728
rect 28718 13676 28724 13728
rect 28776 13716 28782 13728
rect 29196 13716 29224 13824
rect 29730 13812 29736 13824
rect 29788 13812 29794 13864
rect 30282 13812 30288 13864
rect 30340 13852 30346 13864
rect 32306 13852 32312 13864
rect 30340 13824 32312 13852
rect 30340 13812 30346 13824
rect 32306 13812 32312 13824
rect 32364 13852 32370 13864
rect 32876 13852 32904 13960
rect 34606 13948 34612 13960
rect 34664 13948 34670 14000
rect 37461 13991 37519 13997
rect 37461 13957 37473 13991
rect 37507 13988 37519 13991
rect 38378 13988 38384 14000
rect 37507 13960 38384 13988
rect 37507 13957 37519 13960
rect 37461 13951 37519 13957
rect 38378 13948 38384 13960
rect 38436 13948 38442 14000
rect 34330 13920 34336 13932
rect 33152 13892 34336 13920
rect 33042 13852 33048 13864
rect 32364 13824 32904 13852
rect 33003 13824 33048 13852
rect 32364 13812 32370 13824
rect 32876 13784 32904 13824
rect 33042 13812 33048 13824
rect 33100 13812 33106 13864
rect 33152 13861 33180 13892
rect 34330 13880 34336 13892
rect 34388 13880 34394 13932
rect 33137 13855 33195 13861
rect 33137 13821 33149 13855
rect 33183 13821 33195 13855
rect 33321 13855 33379 13861
rect 33321 13852 33333 13855
rect 33137 13815 33195 13821
rect 33244 13824 33333 13852
rect 33244 13784 33272 13824
rect 33321 13821 33333 13824
rect 33367 13821 33379 13855
rect 33321 13815 33379 13821
rect 33410 13812 33416 13864
rect 33468 13852 33474 13864
rect 33962 13852 33968 13864
rect 33468 13824 33513 13852
rect 33875 13824 33968 13852
rect 33468 13812 33474 13824
rect 33962 13812 33968 13824
rect 34020 13852 34026 13864
rect 34238 13852 34244 13864
rect 34020 13824 34244 13852
rect 34020 13812 34026 13824
rect 34238 13812 34244 13824
rect 34296 13852 34302 13864
rect 34609 13855 34667 13861
rect 34609 13852 34621 13855
rect 34296 13824 34621 13852
rect 34296 13812 34302 13824
rect 34609 13821 34621 13824
rect 34655 13821 34667 13855
rect 37274 13852 37280 13864
rect 37235 13824 37280 13852
rect 34609 13815 34667 13821
rect 37274 13812 37280 13824
rect 37332 13812 37338 13864
rect 37918 13852 37924 13864
rect 37879 13824 37924 13852
rect 37918 13812 37924 13824
rect 37976 13812 37982 13864
rect 32876 13756 33272 13784
rect 28776 13688 29224 13716
rect 28776 13676 28782 13688
rect 32306 13676 32312 13728
rect 32364 13716 32370 13728
rect 32490 13716 32496 13728
rect 32364 13688 32496 13716
rect 32364 13676 32370 13688
rect 32490 13676 32496 13688
rect 32548 13676 32554 13728
rect 1104 13626 38824 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 38824 13626
rect 1104 13552 38824 13574
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 24854 13512 24860 13524
rect 11940 13484 24860 13512
rect 11940 13472 11946 13484
rect 24854 13472 24860 13484
rect 24912 13512 24918 13524
rect 25869 13515 25927 13521
rect 25869 13512 25881 13515
rect 24912 13484 25881 13512
rect 24912 13472 24918 13484
rect 25869 13481 25881 13484
rect 25915 13481 25927 13515
rect 26694 13512 26700 13524
rect 25869 13475 25927 13481
rect 26528 13484 26700 13512
rect 22278 13404 22284 13456
rect 22336 13444 22342 13456
rect 24210 13444 24216 13456
rect 22336 13416 24216 13444
rect 22336 13404 22342 13416
rect 24210 13404 24216 13416
rect 24268 13404 24274 13456
rect 24394 13404 24400 13456
rect 24452 13444 24458 13456
rect 24734 13447 24792 13453
rect 24734 13444 24746 13447
rect 24452 13416 24746 13444
rect 24452 13404 24458 13416
rect 24734 13413 24746 13416
rect 24780 13413 24792 13447
rect 24734 13407 24792 13413
rect 25148 13416 26464 13444
rect 1854 13376 1860 13388
rect 1815 13348 1860 13376
rect 1854 13336 1860 13348
rect 1912 13336 1918 13388
rect 21542 13336 21548 13388
rect 21600 13376 21606 13388
rect 22370 13376 22376 13388
rect 21600 13348 22376 13376
rect 21600 13336 21606 13348
rect 22370 13336 22376 13348
rect 22428 13336 22434 13388
rect 22554 13376 22560 13388
rect 22515 13348 22560 13376
rect 22554 13336 22560 13348
rect 22612 13336 22618 13388
rect 22824 13379 22882 13385
rect 22824 13345 22836 13379
rect 22870 13376 22882 13379
rect 25148 13376 25176 13416
rect 22870 13348 25176 13376
rect 22870 13345 22882 13348
rect 22824 13339 22882 13345
rect 25222 13336 25228 13388
rect 25280 13376 25286 13388
rect 26234 13376 26240 13388
rect 25280 13348 26240 13376
rect 25280 13336 25286 13348
rect 26234 13336 26240 13348
rect 26292 13336 26298 13388
rect 23566 13268 23572 13320
rect 23624 13308 23630 13320
rect 24486 13308 24492 13320
rect 23624 13280 24492 13308
rect 23624 13268 23630 13280
rect 24486 13268 24492 13280
rect 24544 13268 24550 13320
rect 26142 13308 26148 13320
rect 25884 13280 26148 13308
rect 2133 13175 2191 13181
rect 2133 13141 2145 13175
rect 2179 13172 2191 13175
rect 17034 13172 17040 13184
rect 2179 13144 17040 13172
rect 2179 13141 2191 13144
rect 2133 13135 2191 13141
rect 17034 13132 17040 13144
rect 17092 13132 17098 13184
rect 23842 13132 23848 13184
rect 23900 13172 23906 13184
rect 23937 13175 23995 13181
rect 23937 13172 23949 13175
rect 23900 13144 23949 13172
rect 23900 13132 23906 13144
rect 23937 13141 23949 13144
rect 23983 13172 23995 13175
rect 24762 13172 24768 13184
rect 23983 13144 24768 13172
rect 23983 13141 23995 13144
rect 23937 13135 23995 13141
rect 24762 13132 24768 13144
rect 24820 13132 24826 13184
rect 24854 13132 24860 13184
rect 24912 13172 24918 13184
rect 25884 13172 25912 13280
rect 26142 13268 26148 13280
rect 26200 13268 26206 13320
rect 26436 13308 26464 13416
rect 26528 13385 26556 13484
rect 26694 13472 26700 13484
rect 26752 13472 26758 13524
rect 27798 13472 27804 13524
rect 27856 13512 27862 13524
rect 28718 13512 28724 13524
rect 27856 13484 28724 13512
rect 27856 13472 27862 13484
rect 28718 13472 28724 13484
rect 28776 13472 28782 13524
rect 29178 13512 29184 13524
rect 29091 13484 29184 13512
rect 29178 13472 29184 13484
rect 29236 13512 29242 13524
rect 29546 13512 29552 13524
rect 29236 13484 29552 13512
rect 29236 13472 29242 13484
rect 29546 13472 29552 13484
rect 29604 13472 29610 13524
rect 36722 13472 36728 13524
rect 36780 13512 36786 13524
rect 37369 13515 37427 13521
rect 37369 13512 37381 13515
rect 36780 13484 37381 13512
rect 36780 13472 36786 13484
rect 37369 13481 37381 13484
rect 37415 13481 37427 13515
rect 37369 13475 37427 13481
rect 31938 13444 31944 13456
rect 26620 13416 31944 13444
rect 26620 13385 26648 13416
rect 31938 13404 31944 13416
rect 31996 13404 32002 13456
rect 26513 13379 26571 13385
rect 26513 13345 26525 13379
rect 26559 13345 26571 13379
rect 26513 13339 26571 13345
rect 26605 13379 26663 13385
rect 26605 13345 26617 13379
rect 26651 13345 26663 13379
rect 26605 13339 26663 13345
rect 26881 13379 26939 13385
rect 26881 13345 26893 13379
rect 26927 13376 26939 13379
rect 27154 13376 27160 13388
rect 26927 13348 27160 13376
rect 26927 13345 26939 13348
rect 26881 13339 26939 13345
rect 27154 13336 27160 13348
rect 27212 13336 27218 13388
rect 28068 13379 28126 13385
rect 28068 13345 28080 13379
rect 28114 13376 28126 13379
rect 29086 13376 29092 13388
rect 28114 13348 29092 13376
rect 28114 13345 28126 13348
rect 28068 13339 28126 13345
rect 29086 13336 29092 13348
rect 29144 13336 29150 13388
rect 37182 13376 37188 13388
rect 37143 13348 37188 13376
rect 37182 13336 37188 13348
rect 37240 13336 37246 13388
rect 27614 13308 27620 13320
rect 26436 13280 27620 13308
rect 27614 13268 27620 13280
rect 27672 13268 27678 13320
rect 27801 13311 27859 13317
rect 27801 13277 27813 13311
rect 27847 13277 27859 13311
rect 27801 13271 27859 13277
rect 26050 13200 26056 13252
rect 26108 13240 26114 13252
rect 26789 13243 26847 13249
rect 26789 13240 26801 13243
rect 26108 13212 26801 13240
rect 26108 13200 26114 13212
rect 26789 13209 26801 13212
rect 26835 13209 26847 13243
rect 26789 13203 26847 13209
rect 26878 13200 26884 13252
rect 26936 13240 26942 13252
rect 27522 13240 27528 13252
rect 26936 13212 27528 13240
rect 26936 13200 26942 13212
rect 27522 13200 27528 13212
rect 27580 13240 27586 13252
rect 27816 13240 27844 13271
rect 27580 13212 27844 13240
rect 27580 13200 27586 13212
rect 24912 13144 25912 13172
rect 24912 13132 24918 13144
rect 25958 13132 25964 13184
rect 26016 13172 26022 13184
rect 26329 13175 26387 13181
rect 26329 13172 26341 13175
rect 26016 13144 26341 13172
rect 26016 13132 26022 13144
rect 26329 13141 26341 13144
rect 26375 13141 26387 13175
rect 26329 13135 26387 13141
rect 27614 13132 27620 13184
rect 27672 13172 27678 13184
rect 28902 13172 28908 13184
rect 27672 13144 28908 13172
rect 27672 13132 27678 13144
rect 28902 13132 28908 13144
rect 28960 13132 28966 13184
rect 1104 13082 38824 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 38824 13082
rect 1104 13008 38824 13030
rect 20898 12968 20904 12980
rect 20859 12940 20904 12968
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 21928 12940 23152 12968
rect 19886 12792 19892 12844
rect 19944 12832 19950 12844
rect 21542 12832 21548 12844
rect 19944 12804 21312 12832
rect 21503 12804 21548 12832
rect 19944 12792 19950 12804
rect 21082 12764 21088 12776
rect 21043 12736 21088 12764
rect 21082 12724 21088 12736
rect 21140 12724 21146 12776
rect 21284 12773 21312 12804
rect 21542 12792 21548 12804
rect 21600 12792 21606 12844
rect 21269 12767 21327 12773
rect 21269 12733 21281 12767
rect 21315 12733 21327 12767
rect 21269 12727 21327 12733
rect 21407 12767 21465 12773
rect 21407 12733 21419 12767
rect 21453 12764 21465 12767
rect 21928 12764 21956 12940
rect 23124 12832 23152 12940
rect 24210 12928 24216 12980
rect 24268 12968 24274 12980
rect 26602 12968 26608 12980
rect 24268 12940 26188 12968
rect 26515 12940 26608 12968
rect 24268 12928 24274 12940
rect 23382 12900 23388 12912
rect 23343 12872 23388 12900
rect 23382 12860 23388 12872
rect 23440 12860 23446 12912
rect 26160 12900 26188 12940
rect 26602 12928 26608 12940
rect 26660 12968 26666 12980
rect 26786 12968 26792 12980
rect 26660 12940 26792 12968
rect 26660 12928 26666 12940
rect 26786 12928 26792 12940
rect 26844 12928 26850 12980
rect 28534 12968 28540 12980
rect 26896 12940 28540 12968
rect 26896 12900 26924 12940
rect 28534 12928 28540 12940
rect 28592 12928 28598 12980
rect 28813 12971 28871 12977
rect 28813 12937 28825 12971
rect 28859 12968 28871 12971
rect 30282 12968 30288 12980
rect 28859 12940 30288 12968
rect 28859 12937 28871 12940
rect 28813 12931 28871 12937
rect 30282 12928 30288 12940
rect 30340 12928 30346 12980
rect 36354 12928 36360 12980
rect 36412 12968 36418 12980
rect 37461 12971 37519 12977
rect 37461 12968 37473 12971
rect 36412 12940 37473 12968
rect 36412 12928 36418 12940
rect 37461 12937 37473 12940
rect 37507 12937 37519 12971
rect 37461 12931 37519 12937
rect 38105 12971 38163 12977
rect 38105 12937 38117 12971
rect 38151 12968 38163 12971
rect 38286 12968 38292 12980
rect 38151 12940 38292 12968
rect 38151 12937 38163 12940
rect 38105 12931 38163 12937
rect 38286 12928 38292 12940
rect 38344 12928 38350 12980
rect 34054 12900 34060 12912
rect 26160 12872 26924 12900
rect 27356 12872 34060 12900
rect 24854 12832 24860 12844
rect 23124 12804 24860 12832
rect 24854 12792 24860 12804
rect 24912 12792 24918 12844
rect 25222 12832 25228 12844
rect 25183 12804 25228 12832
rect 25222 12792 25228 12804
rect 25280 12792 25286 12844
rect 26510 12792 26516 12844
rect 26568 12832 26574 12844
rect 27062 12832 27068 12844
rect 26568 12804 27068 12832
rect 26568 12792 26574 12804
rect 27062 12792 27068 12804
rect 27120 12792 27126 12844
rect 21453 12736 21956 12764
rect 22005 12767 22063 12773
rect 21453 12733 21465 12736
rect 21407 12727 21465 12733
rect 22005 12733 22017 12767
rect 22051 12733 22063 12767
rect 22005 12727 22063 12733
rect 22272 12767 22330 12773
rect 22272 12733 22284 12767
rect 22318 12764 22330 12767
rect 24946 12764 24952 12776
rect 22318 12736 24952 12764
rect 22318 12733 22330 12736
rect 22272 12727 22330 12733
rect 21177 12699 21235 12705
rect 21177 12665 21189 12699
rect 21223 12665 21235 12699
rect 22020 12696 22048 12727
rect 24946 12724 24952 12736
rect 25004 12724 25010 12776
rect 25492 12767 25550 12773
rect 25492 12733 25504 12767
rect 25538 12764 25550 12767
rect 26326 12764 26332 12776
rect 25538 12736 26332 12764
rect 25538 12733 25550 12736
rect 25492 12727 25550 12733
rect 26326 12724 26332 12736
rect 26384 12724 26390 12776
rect 26418 12724 26424 12776
rect 26476 12764 26482 12776
rect 27356 12773 27384 12872
rect 34054 12860 34060 12872
rect 34112 12860 34118 12912
rect 27525 12835 27583 12841
rect 27525 12801 27537 12835
rect 27571 12801 27583 12835
rect 27525 12795 27583 12801
rect 27249 12767 27307 12773
rect 27249 12764 27261 12767
rect 26476 12736 27261 12764
rect 26476 12724 26482 12736
rect 27249 12733 27261 12736
rect 27295 12733 27307 12767
rect 27249 12727 27307 12733
rect 27341 12767 27399 12773
rect 27341 12733 27353 12767
rect 27387 12733 27399 12767
rect 27341 12727 27399 12733
rect 22554 12696 22560 12708
rect 22020 12668 22560 12696
rect 21177 12659 21235 12665
rect 21192 12628 21220 12659
rect 22554 12656 22560 12668
rect 22612 12656 22618 12708
rect 23658 12656 23664 12708
rect 23716 12696 23722 12708
rect 27540 12696 27568 12795
rect 37826 12792 37832 12844
rect 37884 12832 37890 12844
rect 38286 12832 38292 12844
rect 37884 12804 38292 12832
rect 37884 12792 37890 12804
rect 38286 12792 38292 12804
rect 38344 12792 38350 12844
rect 27614 12724 27620 12776
rect 27672 12764 27678 12776
rect 28718 12764 28724 12776
rect 27672 12736 27717 12764
rect 28679 12736 28724 12764
rect 27672 12724 27678 12736
rect 28718 12724 28724 12736
rect 28776 12724 28782 12776
rect 37274 12764 37280 12776
rect 37235 12736 37280 12764
rect 37274 12724 37280 12736
rect 37332 12724 37338 12776
rect 37918 12764 37924 12776
rect 37879 12736 37924 12764
rect 37918 12724 37924 12736
rect 37976 12724 37982 12776
rect 23716 12668 27568 12696
rect 23716 12656 23722 12668
rect 24210 12628 24216 12640
rect 21192 12600 24216 12628
rect 24210 12588 24216 12600
rect 24268 12588 24274 12640
rect 24394 12588 24400 12640
rect 24452 12628 24458 12640
rect 27065 12631 27123 12637
rect 27065 12628 27077 12631
rect 24452 12600 27077 12628
rect 24452 12588 24458 12600
rect 27065 12597 27077 12600
rect 27111 12597 27123 12631
rect 27065 12591 27123 12597
rect 1104 12538 38824 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 38824 12538
rect 1104 12464 38824 12486
rect 10318 12384 10324 12436
rect 10376 12424 10382 12436
rect 10376 12396 22094 12424
rect 10376 12384 10382 12396
rect 1854 12288 1860 12300
rect 1815 12260 1860 12288
rect 1854 12248 1860 12260
rect 1912 12248 1918 12300
rect 2133 12155 2191 12161
rect 2133 12121 2145 12155
rect 2179 12152 2191 12155
rect 16942 12152 16948 12164
rect 2179 12124 16948 12152
rect 2179 12121 2191 12124
rect 2133 12115 2191 12121
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 22066 12084 22094 12396
rect 22186 12384 22192 12436
rect 22244 12424 22250 12436
rect 23290 12424 23296 12436
rect 22244 12396 23296 12424
rect 22244 12384 22250 12396
rect 23290 12384 23296 12396
rect 23348 12424 23354 12436
rect 23937 12427 23995 12433
rect 23937 12424 23949 12427
rect 23348 12396 23949 12424
rect 23348 12384 23354 12396
rect 23937 12393 23949 12396
rect 23983 12393 23995 12427
rect 23937 12387 23995 12393
rect 26234 12384 26240 12436
rect 26292 12424 26298 12436
rect 26329 12427 26387 12433
rect 26329 12424 26341 12427
rect 26292 12396 26341 12424
rect 26292 12384 26298 12396
rect 26329 12393 26341 12396
rect 26375 12393 26387 12427
rect 26329 12387 26387 12393
rect 22738 12316 22744 12368
rect 22796 12365 22802 12368
rect 22796 12359 22860 12365
rect 22796 12325 22814 12359
rect 22848 12325 22860 12359
rect 22796 12319 22860 12325
rect 22796 12316 22802 12319
rect 22922 12316 22928 12368
rect 22980 12356 22986 12368
rect 24756 12359 24814 12365
rect 22980 12328 24624 12356
rect 22980 12316 22986 12328
rect 22554 12288 22560 12300
rect 22515 12260 22560 12288
rect 22554 12248 22560 12260
rect 22612 12248 22618 12300
rect 24486 12288 24492 12300
rect 24447 12260 24492 12288
rect 24486 12248 24492 12260
rect 24544 12248 24550 12300
rect 24596 12288 24624 12328
rect 24756 12325 24768 12359
rect 24802 12356 24814 12359
rect 25958 12356 25964 12368
rect 24802 12328 25964 12356
rect 24802 12325 24814 12328
rect 24756 12319 24814 12325
rect 25958 12316 25964 12328
rect 26016 12316 26022 12368
rect 34698 12316 34704 12368
rect 34756 12356 34762 12368
rect 35342 12356 35348 12368
rect 34756 12328 35348 12356
rect 34756 12316 34762 12328
rect 35342 12316 35348 12328
rect 35400 12316 35406 12368
rect 26513 12291 26571 12297
rect 26513 12288 26525 12291
rect 24596 12260 26525 12288
rect 26513 12257 26525 12260
rect 26559 12257 26571 12291
rect 26513 12251 26571 12257
rect 32950 12248 32956 12300
rect 33008 12288 33014 12300
rect 35618 12288 35624 12300
rect 33008 12260 35624 12288
rect 33008 12248 33014 12260
rect 35618 12248 35624 12260
rect 35676 12248 35682 12300
rect 25869 12087 25927 12093
rect 25869 12084 25881 12087
rect 22066 12056 25881 12084
rect 25869 12053 25881 12056
rect 25915 12084 25927 12087
rect 26050 12084 26056 12096
rect 25915 12056 26056 12084
rect 25915 12053 25927 12056
rect 25869 12047 25927 12053
rect 26050 12044 26056 12056
rect 26108 12044 26114 12096
rect 33318 12044 33324 12096
rect 33376 12084 33382 12096
rect 36814 12084 36820 12096
rect 33376 12056 36820 12084
rect 33376 12044 33382 12056
rect 36814 12044 36820 12056
rect 36872 12044 36878 12096
rect 1104 11994 38824 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 38824 11994
rect 1104 11920 38824 11942
rect 4982 11840 4988 11892
rect 5040 11880 5046 11892
rect 22186 11880 22192 11892
rect 5040 11852 22192 11880
rect 5040 11840 5046 11852
rect 22186 11840 22192 11852
rect 22244 11840 22250 11892
rect 22554 11880 22560 11892
rect 22296 11852 22560 11880
rect 22296 11753 22324 11852
rect 22554 11840 22560 11852
rect 22612 11840 22618 11892
rect 36538 11840 36544 11892
rect 36596 11880 36602 11892
rect 37461 11883 37519 11889
rect 37461 11880 37473 11883
rect 36596 11852 37473 11880
rect 36596 11840 36602 11852
rect 37461 11849 37473 11852
rect 37507 11849 37519 11883
rect 37461 11843 37519 11849
rect 36630 11772 36636 11824
rect 36688 11812 36694 11824
rect 38105 11815 38163 11821
rect 38105 11812 38117 11815
rect 36688 11784 38117 11812
rect 36688 11772 36694 11784
rect 38105 11781 38117 11784
rect 38151 11781 38163 11815
rect 38105 11775 38163 11781
rect 22281 11747 22339 11753
rect 22281 11713 22293 11747
rect 22327 11713 22339 11747
rect 22281 11707 22339 11713
rect 33318 11704 33324 11756
rect 33376 11744 33382 11756
rect 33870 11744 33876 11756
rect 33376 11716 33876 11744
rect 33376 11704 33382 11716
rect 33870 11704 33876 11716
rect 33928 11704 33934 11756
rect 22548 11679 22606 11685
rect 22548 11645 22560 11679
rect 22594 11676 22606 11679
rect 24394 11676 24400 11688
rect 22594 11648 24400 11676
rect 22594 11645 22606 11648
rect 22548 11639 22606 11645
rect 24394 11636 24400 11648
rect 24452 11636 24458 11688
rect 34514 11636 34520 11688
rect 34572 11676 34578 11688
rect 34790 11676 34796 11688
rect 34572 11648 34796 11676
rect 34572 11636 34578 11648
rect 34790 11636 34796 11648
rect 34848 11636 34854 11688
rect 37274 11676 37280 11688
rect 37235 11648 37280 11676
rect 37274 11636 37280 11648
rect 37332 11636 37338 11688
rect 37921 11679 37979 11685
rect 37921 11645 37933 11679
rect 37967 11676 37979 11679
rect 38933 11679 38991 11685
rect 38933 11676 38945 11679
rect 37967 11648 38945 11676
rect 37967 11645 37979 11648
rect 37921 11639 37979 11645
rect 38933 11645 38945 11648
rect 38979 11645 38991 11679
rect 38933 11639 38991 11645
rect 1854 11608 1860 11620
rect 1815 11580 1860 11608
rect 1854 11568 1860 11580
rect 1912 11568 1918 11620
rect 2133 11543 2191 11549
rect 2133 11509 2145 11543
rect 2179 11540 2191 11543
rect 17862 11540 17868 11552
rect 2179 11512 17868 11540
rect 2179 11509 2191 11512
rect 2133 11503 2191 11509
rect 17862 11500 17868 11512
rect 17920 11500 17926 11552
rect 23658 11540 23664 11552
rect 23619 11512 23664 11540
rect 23658 11500 23664 11512
rect 23716 11500 23722 11552
rect 1104 11450 38824 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 38824 11450
rect 1104 11376 38824 11398
rect 31294 11296 31300 11348
rect 31352 11296 31358 11348
rect 37090 11296 37096 11348
rect 37148 11336 37154 11348
rect 37369 11339 37427 11345
rect 37369 11336 37381 11339
rect 37148 11308 37381 11336
rect 37148 11296 37154 11308
rect 37369 11305 37381 11308
rect 37415 11305 37427 11339
rect 37369 11299 37427 11305
rect 22824 11271 22882 11277
rect 22824 11237 22836 11271
rect 22870 11268 22882 11271
rect 23750 11268 23756 11280
rect 22870 11240 23756 11268
rect 22870 11237 22882 11240
rect 22824 11231 22882 11237
rect 23750 11228 23756 11240
rect 23808 11228 23814 11280
rect 31312 11268 31340 11296
rect 31220 11240 31340 11268
rect 22554 11200 22560 11212
rect 22515 11172 22560 11200
rect 22554 11160 22560 11172
rect 22612 11160 22618 11212
rect 30374 11160 30380 11212
rect 30432 11200 30438 11212
rect 30745 11203 30803 11209
rect 30745 11200 30757 11203
rect 30432 11172 30757 11200
rect 30432 11160 30438 11172
rect 30745 11169 30757 11172
rect 30791 11169 30803 11203
rect 30745 11163 30803 11169
rect 30926 11160 30932 11212
rect 30984 11200 30990 11212
rect 31220 11209 31248 11240
rect 31220 11203 31288 11209
rect 31220 11200 31242 11203
rect 30984 11172 31242 11200
rect 30984 11160 30990 11172
rect 31230 11169 31242 11172
rect 31276 11169 31288 11203
rect 37182 11200 37188 11212
rect 37143 11172 37188 11200
rect 31230 11163 31288 11169
rect 37182 11160 37188 11172
rect 37240 11160 37246 11212
rect 30006 11092 30012 11144
rect 30064 11132 30070 11144
rect 30282 11132 30288 11144
rect 30064 11104 30288 11132
rect 30064 11092 30070 11104
rect 30282 11092 30288 11104
rect 30340 11132 30346 11144
rect 31021 11135 31079 11141
rect 31021 11132 31033 11135
rect 30340 11104 31033 11132
rect 30340 11092 30346 11104
rect 31021 11101 31033 11104
rect 31067 11101 31079 11135
rect 31021 11095 31079 11101
rect 31110 11092 31116 11144
rect 31168 11132 31174 11144
rect 31168 11104 31213 11132
rect 31168 11092 31174 11104
rect 23934 11064 23940 11076
rect 23895 11036 23940 11064
rect 23934 11024 23940 11036
rect 23992 11024 23998 11076
rect 31389 11067 31447 11073
rect 31389 11033 31401 11067
rect 31435 11064 31447 11067
rect 32950 11064 32956 11076
rect 31435 11036 32956 11064
rect 31435 11033 31447 11036
rect 31389 11027 31447 11033
rect 32950 11024 32956 11036
rect 33008 11024 33014 11076
rect 38930 11064 38936 11076
rect 38891 11036 38936 11064
rect 38930 11024 38936 11036
rect 38988 11024 38994 11076
rect 1104 10906 38824 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 38824 10906
rect 1104 10832 38824 10854
rect 2133 10795 2191 10801
rect 2133 10761 2145 10795
rect 2179 10792 2191 10795
rect 8938 10792 8944 10804
rect 2179 10764 8944 10792
rect 2179 10761 2191 10764
rect 2133 10755 2191 10761
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 36446 10752 36452 10804
rect 36504 10792 36510 10804
rect 37461 10795 37519 10801
rect 37461 10792 37473 10795
rect 36504 10764 37473 10792
rect 36504 10752 36510 10764
rect 37461 10761 37473 10764
rect 37507 10761 37519 10795
rect 37461 10755 37519 10761
rect 35802 10684 35808 10736
rect 35860 10724 35866 10736
rect 38105 10727 38163 10733
rect 38105 10724 38117 10727
rect 35860 10696 38117 10724
rect 35860 10684 35866 10696
rect 38105 10693 38117 10696
rect 38151 10693 38163 10727
rect 38105 10687 38163 10693
rect 1854 10588 1860 10600
rect 1815 10560 1860 10588
rect 1854 10548 1860 10560
rect 1912 10548 1918 10600
rect 37274 10588 37280 10600
rect 37235 10560 37280 10588
rect 37274 10548 37280 10560
rect 37332 10548 37338 10600
rect 37918 10588 37924 10600
rect 37879 10560 37924 10588
rect 37918 10548 37924 10560
rect 37976 10548 37982 10600
rect 1104 10362 38824 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 38824 10362
rect 1104 10288 38824 10310
rect 1854 10112 1860 10124
rect 1815 10084 1860 10112
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 25774 10072 25780 10124
rect 25832 10112 25838 10124
rect 30377 10115 30435 10121
rect 30377 10112 30389 10115
rect 25832 10084 30389 10112
rect 25832 10072 25838 10084
rect 30377 10081 30389 10084
rect 30423 10081 30435 10115
rect 30377 10075 30435 10081
rect 2133 9911 2191 9917
rect 2133 9877 2145 9911
rect 2179 9908 2191 9911
rect 15930 9908 15936 9920
rect 2179 9880 15936 9908
rect 2179 9877 2191 9880
rect 2133 9871 2191 9877
rect 15930 9868 15936 9880
rect 15988 9868 15994 9920
rect 30561 9911 30619 9917
rect 30561 9877 30573 9911
rect 30607 9908 30619 9911
rect 32490 9908 32496 9920
rect 30607 9880 32496 9908
rect 30607 9877 30619 9880
rect 30561 9871 30619 9877
rect 32490 9868 32496 9880
rect 32548 9868 32554 9920
rect 1104 9818 38824 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 38824 9818
rect 1104 9744 38824 9766
rect 38105 9639 38163 9645
rect 38105 9605 38117 9639
rect 38151 9636 38163 9639
rect 38470 9636 38476 9648
rect 38151 9608 38476 9636
rect 38151 9605 38163 9608
rect 38105 9599 38163 9605
rect 38470 9596 38476 9608
rect 38528 9596 38534 9648
rect 37274 9500 37280 9512
rect 37235 9472 37280 9500
rect 37274 9460 37280 9472
rect 37332 9460 37338 9512
rect 37918 9500 37924 9512
rect 37879 9472 37924 9500
rect 37918 9460 37924 9472
rect 37976 9460 37982 9512
rect 37461 9367 37519 9373
rect 37461 9333 37473 9367
rect 37507 9364 37519 9367
rect 38562 9364 38568 9376
rect 37507 9336 38568 9364
rect 37507 9333 37519 9336
rect 37461 9327 37519 9333
rect 38562 9324 38568 9336
rect 38620 9324 38626 9376
rect 1104 9274 38824 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 38824 9274
rect 1104 9200 38824 9222
rect 37366 9160 37372 9172
rect 37327 9132 37372 9160
rect 37366 9120 37372 9132
rect 37424 9120 37430 9172
rect 1854 9024 1860 9036
rect 1815 8996 1860 9024
rect 1854 8984 1860 8996
rect 1912 8984 1918 9036
rect 37182 9024 37188 9036
rect 37143 8996 37188 9024
rect 37182 8984 37188 8996
rect 37240 8984 37246 9036
rect 30190 8916 30196 8968
rect 30248 8956 30254 8968
rect 33686 8956 33692 8968
rect 30248 8928 33692 8956
rect 30248 8916 30254 8928
rect 33686 8916 33692 8928
rect 33744 8916 33750 8968
rect 2133 8823 2191 8829
rect 2133 8789 2145 8823
rect 2179 8820 2191 8823
rect 15286 8820 15292 8832
rect 2179 8792 15292 8820
rect 2179 8789 2191 8792
rect 2133 8783 2191 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 1104 8730 38824 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 38824 8730
rect 1104 8656 38824 8678
rect 34606 8576 34612 8628
rect 34664 8616 34670 8628
rect 37461 8619 37519 8625
rect 37461 8616 37473 8619
rect 34664 8588 37473 8616
rect 34664 8576 34670 8588
rect 37461 8585 37473 8588
rect 37507 8585 37519 8619
rect 37461 8579 37519 8585
rect 35710 8508 35716 8560
rect 35768 8548 35774 8560
rect 38105 8551 38163 8557
rect 38105 8548 38117 8551
rect 35768 8520 38117 8548
rect 35768 8508 35774 8520
rect 38105 8517 38117 8520
rect 38151 8517 38163 8551
rect 38105 8511 38163 8517
rect 37182 8372 37188 8424
rect 37240 8412 37246 8424
rect 37277 8415 37335 8421
rect 37277 8412 37289 8415
rect 37240 8384 37289 8412
rect 37240 8372 37246 8384
rect 37277 8381 37289 8384
rect 37323 8381 37335 8415
rect 37918 8412 37924 8424
rect 37879 8384 37924 8412
rect 37277 8375 37335 8381
rect 37918 8372 37924 8384
rect 37976 8372 37982 8424
rect 1854 8344 1860 8356
rect 1815 8316 1860 8344
rect 1854 8304 1860 8316
rect 1912 8304 1918 8356
rect 2225 8347 2283 8353
rect 2225 8313 2237 8347
rect 2271 8344 2283 8347
rect 17402 8344 17408 8356
rect 2271 8316 17408 8344
rect 2271 8313 2283 8316
rect 2225 8307 2283 8313
rect 17402 8304 17408 8316
rect 17460 8304 17466 8356
rect 1104 8186 38824 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 38824 8186
rect 1104 8112 38824 8134
rect 28534 8032 28540 8084
rect 28592 8072 28598 8084
rect 29457 8075 29515 8081
rect 29457 8072 29469 8075
rect 28592 8044 29469 8072
rect 28592 8032 28598 8044
rect 29457 8041 29469 8044
rect 29503 8041 29515 8075
rect 29457 8035 29515 8041
rect 26510 7964 26516 8016
rect 26568 8004 26574 8016
rect 26568 7976 29868 8004
rect 26568 7964 26574 7976
rect 22738 7896 22744 7948
rect 22796 7936 22802 7948
rect 28442 7936 28448 7948
rect 22796 7908 28448 7936
rect 22796 7896 22802 7908
rect 28442 7896 28448 7908
rect 28500 7896 28506 7948
rect 29457 7939 29515 7945
rect 29457 7905 29469 7939
rect 29503 7936 29515 7939
rect 29546 7936 29552 7948
rect 29503 7908 29552 7936
rect 29503 7905 29515 7908
rect 29457 7899 29515 7905
rect 29546 7896 29552 7908
rect 29604 7896 29610 7948
rect 29840 7945 29868 7976
rect 29641 7939 29699 7945
rect 29641 7905 29653 7939
rect 29687 7905 29699 7939
rect 29641 7899 29699 7905
rect 29825 7939 29883 7945
rect 29825 7905 29837 7939
rect 29871 7905 29883 7939
rect 29825 7899 29883 7905
rect 30101 7939 30159 7945
rect 30101 7905 30113 7939
rect 30147 7936 30159 7939
rect 31294 7936 31300 7948
rect 30147 7908 31300 7936
rect 30147 7905 30159 7908
rect 30101 7899 30159 7905
rect 27614 7828 27620 7880
rect 27672 7868 27678 7880
rect 29656 7868 29684 7899
rect 31294 7896 31300 7908
rect 31352 7896 31358 7948
rect 27672 7840 29684 7868
rect 27672 7828 27678 7840
rect 10870 7760 10876 7812
rect 10928 7800 10934 7812
rect 24302 7800 24308 7812
rect 10928 7772 24308 7800
rect 10928 7760 10934 7772
rect 24302 7760 24308 7772
rect 24360 7760 24366 7812
rect 5166 7692 5172 7744
rect 5224 7732 5230 7744
rect 5350 7732 5356 7744
rect 5224 7704 5356 7732
rect 5224 7692 5230 7704
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 26602 7732 26608 7744
rect 12860 7704 26608 7732
rect 12860 7692 12866 7704
rect 26602 7692 26608 7704
rect 26660 7692 26666 7744
rect 1104 7642 38824 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 38824 7642
rect 1104 7568 38824 7590
rect 2133 7531 2191 7537
rect 2133 7497 2145 7531
rect 2179 7528 2191 7531
rect 3418 7528 3424 7540
rect 2179 7500 3424 7528
rect 2179 7497 2191 7500
rect 2133 7491 2191 7497
rect 3418 7488 3424 7500
rect 3476 7488 3482 7540
rect 37461 7531 37519 7537
rect 37461 7497 37473 7531
rect 37507 7528 37519 7531
rect 38286 7528 38292 7540
rect 37507 7500 38292 7528
rect 37507 7497 37519 7500
rect 37461 7491 37519 7497
rect 38286 7488 38292 7500
rect 38344 7488 38350 7540
rect 36906 7420 36912 7472
rect 36964 7460 36970 7472
rect 38105 7463 38163 7469
rect 38105 7460 38117 7463
rect 36964 7432 38117 7460
rect 36964 7420 36970 7432
rect 38105 7429 38117 7432
rect 38151 7429 38163 7463
rect 38105 7423 38163 7429
rect 1854 7324 1860 7336
rect 1815 7296 1860 7324
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 37274 7324 37280 7336
rect 37235 7296 37280 7324
rect 37274 7284 37280 7296
rect 37332 7284 37338 7336
rect 37918 7324 37924 7336
rect 37879 7296 37924 7324
rect 37918 7284 37924 7296
rect 37976 7284 37982 7336
rect 1104 7098 38824 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 38824 7098
rect 1104 7024 38824 7046
rect 1854 6848 1860 6860
rect 1815 6820 1860 6848
rect 1854 6808 1860 6820
rect 1912 6808 1918 6860
rect 19334 6808 19340 6860
rect 19392 6848 19398 6860
rect 23661 6851 23719 6857
rect 23661 6848 23673 6851
rect 19392 6820 23673 6848
rect 19392 6808 19398 6820
rect 23661 6817 23673 6820
rect 23707 6817 23719 6851
rect 23661 6811 23719 6817
rect 24581 6851 24639 6857
rect 24581 6817 24593 6851
rect 24627 6848 24639 6851
rect 31110 6848 31116 6860
rect 24627 6820 31116 6848
rect 24627 6817 24639 6820
rect 24581 6811 24639 6817
rect 31110 6808 31116 6820
rect 31168 6808 31174 6860
rect 37182 6848 37188 6860
rect 37143 6820 37188 6848
rect 37182 6808 37188 6820
rect 37240 6808 37246 6860
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 33318 6672 33324 6724
rect 33376 6712 33382 6724
rect 37369 6715 37427 6721
rect 37369 6712 37381 6715
rect 33376 6684 37381 6712
rect 33376 6672 33382 6684
rect 37369 6681 37381 6684
rect 37415 6681 37427 6715
rect 37369 6675 37427 6681
rect 1104 6554 38824 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 38824 6554
rect 1104 6480 38824 6502
rect 20622 6400 20628 6452
rect 20680 6440 20686 6452
rect 28994 6440 29000 6452
rect 20680 6412 29000 6440
rect 20680 6400 20686 6412
rect 28994 6400 29000 6412
rect 29052 6400 29058 6452
rect 36814 6440 36820 6452
rect 36775 6412 36820 6440
rect 36814 6400 36820 6412
rect 36872 6400 36878 6452
rect 37458 6440 37464 6452
rect 37419 6412 37464 6440
rect 37458 6400 37464 6412
rect 37516 6400 37522 6452
rect 17678 6332 17684 6384
rect 17736 6372 17742 6384
rect 26694 6372 26700 6384
rect 17736 6344 26700 6372
rect 17736 6332 17742 6344
rect 26694 6332 26700 6344
rect 26752 6332 26758 6384
rect 36170 6332 36176 6384
rect 36228 6372 36234 6384
rect 38105 6375 38163 6381
rect 38105 6372 38117 6375
rect 36228 6344 38117 6372
rect 36228 6332 36234 6344
rect 38105 6341 38117 6344
rect 38151 6341 38163 6375
rect 38105 6335 38163 6341
rect 15746 6264 15752 6316
rect 15804 6304 15810 6316
rect 25682 6304 25688 6316
rect 15804 6276 25688 6304
rect 15804 6264 15810 6276
rect 25682 6264 25688 6276
rect 25740 6264 25746 6316
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 23934 6236 23940 6248
rect 8996 6208 23940 6236
rect 8996 6196 9002 6208
rect 23934 6196 23940 6208
rect 23992 6196 23998 6248
rect 36633 6239 36691 6245
rect 36633 6205 36645 6239
rect 36679 6236 36691 6239
rect 36906 6236 36912 6248
rect 36679 6208 36912 6236
rect 36679 6205 36691 6208
rect 36633 6199 36691 6205
rect 36906 6196 36912 6208
rect 36964 6196 36970 6248
rect 37274 6236 37280 6248
rect 37235 6208 37280 6236
rect 37274 6196 37280 6208
rect 37332 6196 37338 6248
rect 37921 6239 37979 6245
rect 37921 6205 37933 6239
rect 37967 6236 37979 6239
rect 38933 6239 38991 6245
rect 38933 6236 38945 6239
rect 37967 6208 38945 6236
rect 37967 6205 37979 6208
rect 37921 6199 37979 6205
rect 38933 6205 38945 6208
rect 38979 6205 38991 6239
rect 38933 6199 38991 6205
rect 8018 6128 8024 6180
rect 8076 6168 8082 6180
rect 23658 6168 23664 6180
rect 8076 6140 23664 6168
rect 8076 6128 8082 6140
rect 23658 6128 23664 6140
rect 23716 6128 23722 6180
rect 21266 6060 21272 6112
rect 21324 6100 21330 6112
rect 28626 6100 28632 6112
rect 21324 6072 28632 6100
rect 21324 6060 21330 6072
rect 28626 6060 28632 6072
rect 28684 6060 28690 6112
rect 1104 6010 38824 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 38824 6010
rect 1104 5936 38824 5958
rect 35434 5896 35440 5908
rect 35395 5868 35440 5896
rect 35434 5856 35440 5868
rect 35492 5856 35498 5908
rect 35894 5856 35900 5908
rect 35952 5856 35958 5908
rect 36078 5896 36084 5908
rect 36039 5868 36084 5896
rect 36078 5856 36084 5868
rect 36136 5856 36142 5908
rect 36725 5899 36783 5905
rect 36725 5865 36737 5899
rect 36771 5865 36783 5899
rect 36725 5859 36783 5865
rect 1854 5828 1860 5840
rect 1815 5800 1860 5828
rect 1854 5788 1860 5800
rect 1912 5788 1918 5840
rect 2130 5788 2136 5840
rect 2188 5828 2194 5840
rect 6270 5828 6276 5840
rect 2188 5800 6276 5828
rect 2188 5788 2194 5800
rect 6270 5788 6276 5800
rect 6328 5788 6334 5840
rect 35912 5828 35940 5856
rect 36740 5828 36768 5859
rect 35912 5800 36768 5828
rect 2406 5720 2412 5772
rect 2464 5760 2470 5772
rect 3881 5763 3939 5769
rect 3881 5760 3893 5763
rect 2464 5732 3893 5760
rect 2464 5720 2470 5732
rect 3881 5729 3893 5732
rect 3927 5729 3939 5763
rect 3881 5723 3939 5729
rect 34514 5720 34520 5772
rect 34572 5760 34578 5772
rect 34701 5763 34759 5769
rect 34701 5760 34713 5763
rect 34572 5732 34713 5760
rect 34572 5720 34578 5732
rect 34701 5729 34713 5732
rect 34747 5729 34759 5763
rect 34701 5723 34759 5729
rect 35253 5763 35311 5769
rect 35253 5729 35265 5763
rect 35299 5760 35311 5763
rect 35526 5760 35532 5772
rect 35299 5732 35532 5760
rect 35299 5729 35311 5732
rect 35253 5723 35311 5729
rect 35526 5720 35532 5732
rect 35584 5720 35590 5772
rect 35894 5720 35900 5772
rect 35952 5760 35958 5772
rect 36541 5763 36599 5769
rect 35952 5732 35997 5760
rect 35952 5720 35958 5732
rect 36541 5729 36553 5763
rect 36587 5729 36599 5763
rect 37182 5760 37188 5772
rect 37143 5732 37188 5760
rect 36541 5723 36599 5729
rect 2222 5652 2228 5704
rect 2280 5692 2286 5704
rect 6362 5692 6368 5704
rect 2280 5664 6368 5692
rect 2280 5652 2286 5664
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 35802 5652 35808 5704
rect 35860 5692 35866 5704
rect 36556 5692 36584 5723
rect 37182 5720 37188 5732
rect 37240 5720 37246 5772
rect 35860 5664 36584 5692
rect 35860 5652 35866 5664
rect 2133 5627 2191 5633
rect 2133 5593 2145 5627
rect 2179 5624 2191 5627
rect 3697 5627 3755 5633
rect 2179 5596 3648 5624
rect 2179 5593 2191 5596
rect 2133 5587 2191 5593
rect 3234 5556 3240 5568
rect 3195 5528 3240 5556
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 3620 5556 3648 5596
rect 3697 5593 3709 5627
rect 3743 5624 3755 5627
rect 12618 5624 12624 5636
rect 3743 5596 12624 5624
rect 3743 5593 3755 5596
rect 3697 5587 3755 5593
rect 12618 5584 12624 5596
rect 12676 5584 12682 5636
rect 34698 5584 34704 5636
rect 34756 5624 34762 5636
rect 37369 5627 37427 5633
rect 37369 5624 37381 5627
rect 34756 5596 37381 5624
rect 34756 5584 34762 5596
rect 37369 5593 37381 5596
rect 37415 5593 37427 5627
rect 37369 5587 37427 5593
rect 14458 5556 14464 5568
rect 3620 5528 14464 5556
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 31754 5516 31760 5568
rect 31812 5556 31818 5568
rect 34517 5559 34575 5565
rect 34517 5556 34529 5559
rect 31812 5528 34529 5556
rect 31812 5516 31818 5528
rect 34517 5525 34529 5528
rect 34563 5525 34575 5559
rect 38930 5556 38936 5568
rect 38891 5528 38936 5556
rect 34517 5519 34575 5525
rect 38930 5516 38936 5528
rect 38988 5516 38994 5568
rect 1104 5466 38824 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 38824 5466
rect 1104 5392 38824 5414
rect 2130 5352 2136 5364
rect 2091 5324 2136 5352
rect 2130 5312 2136 5324
rect 2188 5312 2194 5364
rect 24670 5312 24676 5364
rect 24728 5352 24734 5364
rect 30742 5352 30748 5364
rect 24728 5324 30748 5352
rect 24728 5312 24734 5324
rect 30742 5312 30748 5324
rect 30800 5312 30806 5364
rect 34790 5352 34796 5364
rect 34751 5324 34796 5352
rect 34790 5312 34796 5324
rect 34848 5312 34854 5364
rect 35342 5312 35348 5364
rect 35400 5352 35406 5364
rect 36725 5355 36783 5361
rect 36725 5352 36737 5355
rect 35400 5324 36737 5352
rect 35400 5312 35406 5324
rect 36725 5321 36737 5324
rect 36771 5321 36783 5355
rect 36725 5315 36783 5321
rect 23566 5244 23572 5296
rect 23624 5284 23630 5296
rect 31018 5284 31024 5296
rect 23624 5256 31024 5284
rect 23624 5244 23630 5256
rect 31018 5244 31024 5256
rect 31076 5244 31082 5296
rect 33778 5244 33784 5296
rect 33836 5284 33842 5296
rect 36081 5287 36139 5293
rect 36081 5284 36093 5287
rect 33836 5256 36093 5284
rect 33836 5244 33842 5256
rect 36081 5253 36093 5256
rect 36127 5253 36139 5287
rect 36081 5247 36139 5253
rect 2774 5176 2780 5228
rect 2832 5216 2838 5228
rect 2961 5219 3019 5225
rect 2961 5216 2973 5219
rect 2832 5188 2973 5216
rect 2832 5176 2838 5188
rect 2961 5185 2973 5188
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 18230 5176 18236 5228
rect 18288 5216 18294 5228
rect 30282 5216 30288 5228
rect 18288 5188 30288 5216
rect 18288 5176 18294 5188
rect 30282 5176 30288 5188
rect 30340 5176 30346 5228
rect 35912 5188 36124 5216
rect 16758 5108 16764 5160
rect 16816 5148 16822 5160
rect 28350 5148 28356 5160
rect 16816 5120 28356 5148
rect 16816 5108 16822 5120
rect 28350 5108 28356 5120
rect 28408 5108 28414 5160
rect 34606 5148 34612 5160
rect 34567 5120 34612 5148
rect 34606 5108 34612 5120
rect 34664 5108 34670 5160
rect 35912 5157 35940 5188
rect 36096 5160 36124 5188
rect 35897 5151 35955 5157
rect 35897 5117 35909 5151
rect 35943 5117 35955 5151
rect 35897 5111 35955 5117
rect 36078 5108 36084 5160
rect 36136 5108 36142 5160
rect 36541 5151 36599 5157
rect 36541 5117 36553 5151
rect 36587 5148 36599 5151
rect 36722 5148 36728 5160
rect 36587 5120 36728 5148
rect 36587 5117 36599 5120
rect 36541 5111 36599 5117
rect 36722 5108 36728 5120
rect 36780 5108 36786 5160
rect 37090 5108 37096 5160
rect 37148 5148 37154 5160
rect 37185 5151 37243 5157
rect 37185 5148 37197 5151
rect 37148 5120 37197 5148
rect 37148 5108 37154 5120
rect 37185 5117 37197 5120
rect 37231 5117 37243 5151
rect 37185 5111 37243 5117
rect 1854 5080 1860 5092
rect 1815 5052 1860 5080
rect 1854 5040 1860 5052
rect 1912 5040 1918 5092
rect 2777 5083 2835 5089
rect 2777 5049 2789 5083
rect 2823 5080 2835 5083
rect 4338 5080 4344 5092
rect 2823 5052 4344 5080
rect 2823 5049 2835 5052
rect 2777 5043 2835 5049
rect 4338 5040 4344 5052
rect 4396 5040 4402 5092
rect 16390 5040 16396 5092
rect 16448 5080 16454 5092
rect 30926 5080 30932 5092
rect 16448 5052 30932 5080
rect 16448 5040 16454 5052
rect 30926 5040 30932 5052
rect 30984 5040 30990 5092
rect 34698 5040 34704 5092
rect 34756 5080 34762 5092
rect 37921 5083 37979 5089
rect 37921 5080 37933 5083
rect 34756 5052 37933 5080
rect 34756 5040 34762 5052
rect 37921 5049 37933 5052
rect 37967 5049 37979 5083
rect 37921 5043 37979 5049
rect 38105 5083 38163 5089
rect 38105 5049 38117 5083
rect 38151 5080 38163 5083
rect 39390 5080 39396 5092
rect 38151 5052 39396 5080
rect 38151 5049 38163 5052
rect 38105 5043 38163 5049
rect 39390 5040 39396 5052
rect 39448 5040 39454 5092
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 23842 5012 23848 5024
rect 6972 4984 23848 5012
rect 6972 4972 6978 4984
rect 23842 4972 23848 4984
rect 23900 4972 23906 5024
rect 32398 4972 32404 5024
rect 32456 5012 32462 5024
rect 37369 5015 37427 5021
rect 37369 5012 37381 5015
rect 32456 4984 37381 5012
rect 32456 4972 32462 4984
rect 37369 4981 37381 4984
rect 37415 4981 37427 5015
rect 37369 4975 37427 4981
rect 1104 4922 38824 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 38824 4922
rect 1104 4848 38824 4870
rect 4614 4768 4620 4820
rect 4672 4808 4678 4820
rect 23382 4808 23388 4820
rect 4672 4780 23388 4808
rect 4672 4768 4678 4780
rect 23382 4768 23388 4780
rect 23440 4768 23446 4820
rect 33042 4768 33048 4820
rect 33100 4808 33106 4820
rect 34701 4811 34759 4817
rect 34701 4808 34713 4811
rect 33100 4780 34713 4808
rect 33100 4768 33106 4780
rect 34701 4777 34713 4780
rect 34747 4777 34759 4811
rect 34701 4771 34759 4777
rect 35710 4768 35716 4820
rect 35768 4808 35774 4820
rect 36633 4811 36691 4817
rect 36633 4808 36645 4811
rect 35768 4780 36645 4808
rect 35768 4768 35774 4780
rect 36633 4777 36645 4780
rect 36679 4777 36691 4811
rect 36633 4771 36691 4777
rect 2222 4740 2228 4752
rect 2183 4712 2228 4740
rect 2222 4700 2228 4712
rect 2280 4700 2286 4752
rect 2777 4743 2835 4749
rect 2777 4709 2789 4743
rect 2823 4740 2835 4743
rect 3142 4740 3148 4752
rect 2823 4712 3148 4740
rect 2823 4709 2835 4712
rect 2777 4703 2835 4709
rect 3142 4700 3148 4712
rect 3200 4700 3206 4752
rect 3234 4700 3240 4752
rect 3292 4740 3298 4752
rect 3513 4743 3571 4749
rect 3513 4740 3525 4743
rect 3292 4712 3525 4740
rect 3292 4700 3298 4712
rect 3513 4709 3525 4712
rect 3559 4709 3571 4743
rect 3513 4703 3571 4709
rect 34422 4700 34428 4752
rect 34480 4740 34486 4752
rect 35253 4743 35311 4749
rect 35253 4740 35265 4743
rect 34480 4712 35265 4740
rect 34480 4700 34486 4712
rect 35253 4709 35265 4712
rect 35299 4709 35311 4743
rect 35253 4703 35311 4709
rect 36354 4700 36360 4752
rect 36412 4740 36418 4752
rect 37185 4743 37243 4749
rect 37185 4740 37197 4743
rect 36412 4712 37197 4740
rect 36412 4700 36418 4712
rect 37185 4709 37197 4712
rect 37231 4709 37243 4743
rect 37185 4703 37243 4709
rect 1854 4672 1860 4684
rect 1815 4644 1860 4672
rect 1854 4632 1860 4644
rect 1912 4632 1918 4684
rect 4338 4672 4344 4684
rect 4299 4644 4344 4672
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 4985 4675 5043 4681
rect 4985 4641 4997 4675
rect 5031 4672 5043 4675
rect 5166 4672 5172 4684
rect 5031 4644 5172 4672
rect 5031 4641 5043 4644
rect 4985 4635 5043 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 31938 4632 31944 4684
rect 31996 4672 32002 4684
rect 32125 4675 32183 4681
rect 32125 4672 32137 4675
rect 31996 4644 32137 4672
rect 31996 4632 32002 4644
rect 32125 4641 32137 4644
rect 32171 4641 32183 4675
rect 32125 4635 32183 4641
rect 33594 4632 33600 4684
rect 33652 4672 33658 4684
rect 33781 4675 33839 4681
rect 33781 4672 33793 4675
rect 33652 4644 33793 4672
rect 33652 4632 33658 4644
rect 33781 4641 33793 4644
rect 33827 4641 33839 4675
rect 33781 4635 33839 4641
rect 34517 4675 34575 4681
rect 34517 4641 34529 4675
rect 34563 4672 34575 4675
rect 35618 4672 35624 4684
rect 34563 4644 35624 4672
rect 34563 4641 34575 4644
rect 34517 4635 34575 4641
rect 35618 4632 35624 4644
rect 35676 4632 35682 4684
rect 36446 4672 36452 4684
rect 36407 4644 36452 4672
rect 36446 4632 36452 4644
rect 36504 4632 36510 4684
rect 2961 4539 3019 4545
rect 2961 4505 2973 4539
rect 3007 4536 3019 4539
rect 3142 4536 3148 4548
rect 3007 4508 3148 4536
rect 3007 4505 3019 4508
rect 2961 4499 3019 4505
rect 3142 4496 3148 4508
rect 3200 4496 3206 4548
rect 31941 4539 31999 4545
rect 31941 4505 31953 4539
rect 31987 4536 31999 4539
rect 34790 4536 34796 4548
rect 31987 4508 34796 4536
rect 31987 4505 31999 4508
rect 31941 4499 31999 4505
rect 34790 4496 34796 4508
rect 34848 4496 34854 4548
rect 37369 4539 37427 4545
rect 37369 4505 37381 4539
rect 37415 4536 37427 4539
rect 39758 4536 39764 4548
rect 37415 4508 39764 4536
rect 37415 4505 37427 4508
rect 37369 4499 37427 4505
rect 39758 4496 39764 4508
rect 39816 4496 39822 4548
rect 3602 4468 3608 4480
rect 3563 4440 3608 4468
rect 3602 4428 3608 4440
rect 3660 4428 3666 4480
rect 4801 4471 4859 4477
rect 4801 4437 4813 4471
rect 4847 4468 4859 4471
rect 12434 4468 12440 4480
rect 4847 4440 12440 4468
rect 4847 4437 4859 4440
rect 4801 4431 4859 4437
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 29270 4428 29276 4480
rect 29328 4468 29334 4480
rect 31846 4468 31852 4480
rect 29328 4440 31852 4468
rect 29328 4428 29334 4440
rect 31846 4428 31852 4440
rect 31904 4428 31910 4480
rect 32030 4428 32036 4480
rect 32088 4468 32094 4480
rect 33597 4471 33655 4477
rect 33597 4468 33609 4471
rect 32088 4440 33609 4468
rect 32088 4428 32094 4440
rect 33597 4437 33609 4440
rect 33643 4437 33655 4471
rect 33597 4431 33655 4437
rect 35250 4428 35256 4480
rect 35308 4468 35314 4480
rect 35345 4471 35403 4477
rect 35345 4468 35357 4471
rect 35308 4440 35357 4468
rect 35308 4428 35314 4440
rect 35345 4437 35357 4440
rect 35391 4437 35403 4471
rect 35345 4431 35403 4437
rect 1104 4378 38824 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 38824 4378
rect 1104 4304 38824 4326
rect 2866 4264 2872 4276
rect 2827 4236 2872 4264
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 23477 4267 23535 4273
rect 23477 4233 23489 4267
rect 23523 4264 23535 4267
rect 27982 4264 27988 4276
rect 23523 4236 27988 4264
rect 23523 4233 23535 4236
rect 23477 4227 23535 4233
rect 27982 4224 27988 4236
rect 28040 4224 28046 4276
rect 28552 4236 28764 4264
rect 5169 4199 5227 4205
rect 5169 4165 5181 4199
rect 5215 4165 5227 4199
rect 5169 4159 5227 4165
rect 26145 4199 26203 4205
rect 26145 4165 26157 4199
rect 26191 4196 26203 4199
rect 27890 4196 27896 4208
rect 26191 4168 27896 4196
rect 26191 4165 26203 4168
rect 26145 4159 26203 4165
rect 2038 4088 2044 4140
rect 2096 4128 2102 4140
rect 2133 4131 2191 4137
rect 2133 4128 2145 4131
rect 2096 4100 2145 4128
rect 2096 4088 2102 4100
rect 2133 4097 2145 4100
rect 2179 4097 2191 4131
rect 5184 4128 5212 4159
rect 27890 4156 27896 4168
rect 27948 4156 27954 4208
rect 20714 4128 20720 4140
rect 5184 4100 20720 4128
rect 2133 4091 2191 4097
rect 20714 4088 20720 4100
rect 20772 4088 20778 4140
rect 28552 4128 28580 4236
rect 25700 4100 28580 4128
rect 28736 4128 28764 4236
rect 31588 4236 31892 4264
rect 31588 4128 31616 4236
rect 28736 4100 31616 4128
rect 1486 4020 1492 4072
rect 1544 4060 1550 4072
rect 3602 4060 3608 4072
rect 1544 4032 3608 4060
rect 1544 4020 1550 4032
rect 3602 4020 3608 4032
rect 3660 4020 3666 4072
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4060 4399 4063
rect 4614 4060 4620 4072
rect 4387 4032 4620 4060
rect 4387 4029 4399 4032
rect 4341 4023 4399 4029
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 4706 4020 4712 4072
rect 4764 4060 4770 4072
rect 4985 4063 5043 4069
rect 4985 4060 4997 4063
rect 4764 4032 4997 4060
rect 4764 4020 4770 4032
rect 4985 4029 4997 4032
rect 5031 4029 5043 4063
rect 4985 4023 5043 4029
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 5629 4063 5687 4069
rect 5629 4060 5641 4063
rect 5316 4032 5641 4060
rect 5316 4020 5322 4032
rect 5629 4029 5641 4032
rect 5675 4029 5687 4063
rect 6546 4060 6552 4072
rect 6507 4032 6552 4060
rect 5629 4023 5687 4029
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 11882 4060 11888 4072
rect 11843 4032 11888 4060
rect 11882 4020 11888 4032
rect 11940 4020 11946 4072
rect 12802 4060 12808 4072
rect 12763 4032 12808 4060
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 14366 4020 14372 4072
rect 14424 4060 14430 4072
rect 14737 4063 14795 4069
rect 14737 4060 14749 4063
rect 14424 4032 14749 4060
rect 14424 4020 14430 4032
rect 14737 4029 14749 4032
rect 14783 4029 14795 4063
rect 18690 4060 18696 4072
rect 14737 4023 14795 4029
rect 14936 4032 18552 4060
rect 18651 4032 18696 4060
rect 1854 3992 1860 4004
rect 1815 3964 1860 3992
rect 1854 3952 1860 3964
rect 1912 3952 1918 4004
rect 2682 3952 2688 4004
rect 2740 3992 2746 4004
rect 2777 3995 2835 4001
rect 2777 3992 2789 3995
rect 2740 3964 2789 3992
rect 2740 3952 2746 3964
rect 2777 3961 2789 3964
rect 2823 3961 2835 3995
rect 2777 3955 2835 3961
rect 3602 3884 3608 3936
rect 3660 3924 3666 3936
rect 4433 3927 4491 3933
rect 4433 3924 4445 3927
rect 3660 3896 4445 3924
rect 3660 3884 3666 3896
rect 4433 3893 4445 3896
rect 4479 3893 4491 3927
rect 4433 3887 4491 3893
rect 11790 3884 11796 3936
rect 11848 3924 11854 3936
rect 11977 3927 12035 3933
rect 11977 3924 11989 3927
rect 11848 3896 11989 3924
rect 11848 3884 11854 3896
rect 11977 3893 11989 3896
rect 12023 3893 12035 3927
rect 11977 3887 12035 3893
rect 12710 3884 12716 3936
rect 12768 3924 12774 3936
rect 14936 3933 14964 4032
rect 16758 3992 16764 4004
rect 16719 3964 16764 3992
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 17678 3992 17684 4004
rect 17639 3964 17684 3992
rect 17678 3952 17684 3964
rect 17736 3952 17742 4004
rect 18524 3992 18552 4032
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 19978 4020 19984 4072
rect 20036 4060 20042 4072
rect 20165 4063 20223 4069
rect 20165 4060 20177 4063
rect 20036 4032 20177 4060
rect 20036 4020 20042 4032
rect 20165 4029 20177 4032
rect 20211 4029 20223 4063
rect 20165 4023 20223 4029
rect 21818 4020 21824 4072
rect 21876 4060 21882 4072
rect 22005 4063 22063 4069
rect 22005 4060 22017 4063
rect 21876 4032 22017 4060
rect 21876 4020 21882 4032
rect 22005 4029 22017 4032
rect 22051 4029 22063 4063
rect 22005 4023 22063 4029
rect 22830 4020 22836 4072
rect 22888 4060 22894 4072
rect 23017 4063 23075 4069
rect 23017 4060 23029 4063
rect 22888 4032 23029 4060
rect 22888 4020 22894 4032
rect 23017 4029 23029 4032
rect 23063 4029 23075 4063
rect 23017 4023 23075 4029
rect 23198 4020 23204 4072
rect 23256 4060 23262 4072
rect 23661 4063 23719 4069
rect 23661 4060 23673 4063
rect 23256 4032 23673 4060
rect 23256 4020 23262 4032
rect 23661 4029 23673 4032
rect 23707 4029 23719 4063
rect 23661 4023 23719 4029
rect 24118 4020 24124 4072
rect 24176 4060 24182 4072
rect 24305 4063 24363 4069
rect 24305 4060 24317 4063
rect 24176 4032 24317 4060
rect 24176 4020 24182 4032
rect 24305 4029 24317 4032
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 24762 4020 24768 4072
rect 24820 4060 24826 4072
rect 25409 4063 25467 4069
rect 25409 4060 25421 4063
rect 24820 4032 25421 4060
rect 24820 4020 24826 4032
rect 25409 4029 25421 4032
rect 25455 4029 25467 4063
rect 25409 4023 25467 4029
rect 20070 3992 20076 4004
rect 18524 3964 20076 3992
rect 20070 3952 20076 3964
rect 20128 3952 20134 4004
rect 20990 3952 20996 4004
rect 21048 3992 21054 4004
rect 25700 3992 25728 4100
rect 31662 4088 31668 4140
rect 31720 4128 31726 4140
rect 31754 4128 31760 4140
rect 31720 4100 31760 4128
rect 31720 4088 31726 4100
rect 31754 4088 31760 4100
rect 31812 4088 31818 4140
rect 31864 4128 31892 4236
rect 32950 4156 32956 4208
rect 33008 4196 33014 4208
rect 33008 4168 34468 4196
rect 33008 4156 33014 4168
rect 32122 4128 32128 4140
rect 31864 4100 32128 4128
rect 32122 4088 32128 4100
rect 32180 4088 32186 4140
rect 33134 4088 33140 4140
rect 33192 4128 33198 4140
rect 34330 4128 34336 4140
rect 33192 4100 34336 4128
rect 33192 4088 33198 4100
rect 34330 4088 34336 4100
rect 34388 4088 34394 4140
rect 34440 4128 34468 4168
rect 34440 4100 37964 4128
rect 25958 4060 25964 4072
rect 25919 4032 25964 4060
rect 25958 4020 25964 4032
rect 26016 4020 26022 4072
rect 26789 4063 26847 4069
rect 26789 4029 26801 4063
rect 26835 4029 26847 4063
rect 26789 4023 26847 4029
rect 21048 3964 25728 3992
rect 21048 3952 21054 3964
rect 25774 3952 25780 4004
rect 25832 3992 25838 4004
rect 26804 3992 26832 4023
rect 26878 4020 26884 4072
rect 26936 4060 26942 4072
rect 27433 4063 27491 4069
rect 27433 4060 27445 4063
rect 26936 4032 27445 4060
rect 26936 4020 26942 4032
rect 27433 4029 27445 4032
rect 27479 4029 27491 4063
rect 28902 4060 28908 4072
rect 28863 4032 28908 4060
rect 27433 4023 27491 4029
rect 28902 4020 28908 4032
rect 28960 4020 28966 4072
rect 29546 4060 29552 4072
rect 29507 4032 29552 4060
rect 29546 4020 29552 4032
rect 29604 4020 29610 4072
rect 29638 4020 29644 4072
rect 29696 4060 29702 4072
rect 30653 4063 30711 4069
rect 30653 4060 30665 4063
rect 29696 4032 30665 4060
rect 29696 4020 29702 4032
rect 30653 4029 30665 4032
rect 30699 4029 30711 4063
rect 30653 4023 30711 4029
rect 30742 4020 30748 4072
rect 30800 4060 30806 4072
rect 31297 4063 31355 4069
rect 31297 4060 31309 4063
rect 30800 4032 31309 4060
rect 30800 4020 30806 4032
rect 31297 4029 31309 4032
rect 31343 4029 31355 4063
rect 31297 4023 31355 4029
rect 31496 4032 31800 4060
rect 25832 3964 26832 3992
rect 25832 3952 25838 3964
rect 27522 3952 27528 4004
rect 27580 3992 27586 4004
rect 29270 3992 29276 4004
rect 27580 3964 29276 3992
rect 27580 3952 27586 3964
rect 29270 3952 29276 3964
rect 29328 3952 29334 4004
rect 31496 3992 31524 4032
rect 29380 3964 31524 3992
rect 31772 3992 31800 4032
rect 31846 4020 31852 4072
rect 31904 4060 31910 4072
rect 31941 4063 31999 4069
rect 31941 4060 31953 4063
rect 31904 4032 31953 4060
rect 31904 4020 31910 4032
rect 31941 4029 31953 4032
rect 31987 4029 31999 4063
rect 31941 4023 31999 4029
rect 32582 4020 32588 4072
rect 32640 4060 32646 4072
rect 32769 4063 32827 4069
rect 32769 4060 32781 4063
rect 32640 4032 32781 4060
rect 32640 4020 32646 4032
rect 32769 4029 32781 4032
rect 32815 4029 32827 4063
rect 33410 4060 33416 4072
rect 33371 4032 33416 4060
rect 32769 4023 32827 4029
rect 33410 4020 33416 4032
rect 33468 4020 33474 4072
rect 34241 4063 34299 4069
rect 34241 4029 34253 4063
rect 34287 4029 34299 4063
rect 34241 4023 34299 4029
rect 34256 3992 34284 4023
rect 34790 4020 34796 4072
rect 34848 4060 34854 4072
rect 37936 4069 37964 4100
rect 35897 4063 35955 4069
rect 35897 4060 35909 4063
rect 34848 4032 35909 4060
rect 34848 4020 34854 4032
rect 35897 4029 35909 4032
rect 35943 4029 35955 4063
rect 37921 4063 37979 4069
rect 35897 4023 35955 4029
rect 36556 4032 37872 4060
rect 31772 3964 34284 3992
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 12768 3896 12909 3924
rect 12768 3884 12774 3896
rect 12897 3893 12909 3896
rect 12943 3893 12955 3927
rect 12897 3887 12955 3893
rect 14921 3927 14979 3933
rect 14921 3893 14933 3927
rect 14967 3893 14979 3927
rect 14921 3887 14979 3893
rect 16666 3884 16672 3936
rect 16724 3924 16730 3936
rect 16853 3927 16911 3933
rect 16853 3924 16865 3927
rect 16724 3896 16865 3924
rect 16724 3884 16730 3896
rect 16853 3893 16865 3896
rect 16899 3893 16911 3927
rect 17770 3924 17776 3936
rect 17731 3896 17776 3924
rect 16853 3887 16911 3893
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 18690 3884 18696 3936
rect 18748 3924 18754 3936
rect 18785 3927 18843 3933
rect 18785 3924 18797 3927
rect 18748 3896 18797 3924
rect 18748 3884 18754 3896
rect 18785 3893 18797 3896
rect 18831 3893 18843 3927
rect 18785 3887 18843 3893
rect 19981 3927 20039 3933
rect 19981 3893 19993 3927
rect 20027 3924 20039 3927
rect 20254 3924 20260 3936
rect 20027 3896 20260 3924
rect 20027 3893 20039 3896
rect 19981 3887 20039 3893
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 20438 3884 20444 3936
rect 20496 3924 20502 3936
rect 21821 3927 21879 3933
rect 21821 3924 21833 3927
rect 20496 3896 21833 3924
rect 20496 3884 20502 3896
rect 21821 3893 21833 3896
rect 21867 3893 21879 3927
rect 21821 3887 21879 3893
rect 21910 3884 21916 3936
rect 21968 3924 21974 3936
rect 22833 3927 22891 3933
rect 22833 3924 22845 3927
rect 21968 3896 22845 3924
rect 21968 3884 21974 3896
rect 22833 3893 22845 3896
rect 22879 3893 22891 3927
rect 22833 3887 22891 3893
rect 24121 3927 24179 3933
rect 24121 3893 24133 3927
rect 24167 3924 24179 3927
rect 25130 3924 25136 3936
rect 24167 3896 25136 3924
rect 24167 3893 24179 3896
rect 24121 3887 24179 3893
rect 25130 3884 25136 3896
rect 25188 3884 25194 3936
rect 25225 3927 25283 3933
rect 25225 3893 25237 3927
rect 25271 3924 25283 3927
rect 25590 3924 25596 3936
rect 25271 3896 25596 3924
rect 25271 3893 25283 3896
rect 25225 3887 25283 3893
rect 25590 3884 25596 3896
rect 25648 3884 25654 3936
rect 26234 3884 26240 3936
rect 26292 3924 26298 3936
rect 26605 3927 26663 3933
rect 26605 3924 26617 3927
rect 26292 3896 26617 3924
rect 26292 3884 26298 3896
rect 26605 3893 26617 3896
rect 26651 3893 26663 3927
rect 26605 3887 26663 3893
rect 26694 3884 26700 3936
rect 26752 3924 26758 3936
rect 27249 3927 27307 3933
rect 27249 3924 27261 3927
rect 26752 3896 27261 3924
rect 26752 3884 26758 3896
rect 27249 3893 27261 3896
rect 27295 3893 27307 3927
rect 27249 3887 27307 3893
rect 28074 3884 28080 3936
rect 28132 3924 28138 3936
rect 29380 3933 29408 3964
rect 34606 3952 34612 4004
rect 34664 3992 34670 4004
rect 36449 3995 36507 4001
rect 36449 3992 36461 3995
rect 34664 3964 36461 3992
rect 34664 3952 34670 3964
rect 36449 3961 36461 3964
rect 36495 3961 36507 3995
rect 36449 3955 36507 3961
rect 28721 3927 28779 3933
rect 28721 3924 28733 3927
rect 28132 3896 28733 3924
rect 28132 3884 28138 3896
rect 28721 3893 28733 3896
rect 28767 3893 28779 3927
rect 28721 3887 28779 3893
rect 29365 3927 29423 3933
rect 29365 3893 29377 3927
rect 29411 3893 29423 3927
rect 29365 3887 29423 3893
rect 29454 3884 29460 3936
rect 29512 3924 29518 3936
rect 30469 3927 30527 3933
rect 30469 3924 30481 3927
rect 29512 3896 30481 3924
rect 29512 3884 29518 3896
rect 30469 3893 30481 3896
rect 30515 3893 30527 3927
rect 30469 3887 30527 3893
rect 30558 3884 30564 3936
rect 30616 3924 30622 3936
rect 31113 3927 31171 3933
rect 31113 3924 31125 3927
rect 30616 3896 31125 3924
rect 30616 3884 30622 3896
rect 31113 3893 31125 3896
rect 31159 3893 31171 3927
rect 31754 3924 31760 3936
rect 31715 3896 31760 3924
rect 31113 3887 31171 3893
rect 31754 3884 31760 3896
rect 31812 3884 31818 3936
rect 31846 3884 31852 3936
rect 31904 3924 31910 3936
rect 32585 3927 32643 3933
rect 32585 3924 32597 3927
rect 31904 3896 32597 3924
rect 31904 3884 31910 3896
rect 32585 3893 32597 3896
rect 32631 3893 32643 3927
rect 32585 3887 32643 3893
rect 33502 3884 33508 3936
rect 33560 3924 33566 3936
rect 33597 3927 33655 3933
rect 33597 3924 33609 3927
rect 33560 3896 33609 3924
rect 33560 3884 33566 3896
rect 33597 3893 33609 3896
rect 33643 3893 33655 3927
rect 33597 3887 33655 3893
rect 34057 3927 34115 3933
rect 34057 3893 34069 3927
rect 34103 3924 34115 3927
rect 34698 3924 34704 3936
rect 34103 3896 34704 3924
rect 34103 3893 34115 3896
rect 34057 3887 34115 3893
rect 34698 3884 34704 3896
rect 34756 3884 34762 3936
rect 35713 3927 35771 3933
rect 35713 3893 35725 3927
rect 35759 3924 35771 3927
rect 36354 3924 36360 3936
rect 35759 3896 36360 3924
rect 35759 3893 35771 3896
rect 35713 3887 35771 3893
rect 36354 3884 36360 3896
rect 36412 3884 36418 3936
rect 36556 3933 36584 4032
rect 36630 3952 36636 4004
rect 36688 3992 36694 4004
rect 37185 3995 37243 4001
rect 37185 3992 37197 3995
rect 36688 3964 37197 3992
rect 36688 3952 36694 3964
rect 37185 3961 37197 3964
rect 37231 3961 37243 3995
rect 37844 3992 37872 4032
rect 37921 4029 37933 4063
rect 37967 4029 37979 4063
rect 39114 4060 39120 4072
rect 37921 4023 37979 4029
rect 38028 4032 39120 4060
rect 38028 3992 38056 4032
rect 39114 4020 39120 4032
rect 39172 4020 39178 4072
rect 37844 3964 38056 3992
rect 38105 3995 38163 4001
rect 37185 3955 37243 3961
rect 38105 3961 38117 3995
rect 38151 3992 38163 3995
rect 38470 3992 38476 4004
rect 38151 3964 38476 3992
rect 38151 3961 38163 3964
rect 38105 3955 38163 3961
rect 38470 3952 38476 3964
rect 38528 3952 38534 4004
rect 36541 3927 36599 3933
rect 36541 3893 36553 3927
rect 36587 3893 36599 3927
rect 36541 3887 36599 3893
rect 37277 3927 37335 3933
rect 37277 3893 37289 3927
rect 37323 3924 37335 3927
rect 38746 3924 38752 3936
rect 37323 3896 38752 3924
rect 37323 3893 37335 3896
rect 37277 3887 37335 3893
rect 38746 3884 38752 3896
rect 38804 3884 38810 3936
rect 1104 3834 38824 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 38824 3834
rect 1104 3760 38824 3782
rect 1026 3680 1032 3732
rect 1084 3720 1090 3732
rect 2774 3720 2780 3732
rect 1084 3692 2780 3720
rect 1084 3680 1090 3692
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 3510 3720 3516 3732
rect 3471 3692 3516 3720
rect 3510 3680 3516 3692
rect 3568 3680 3574 3732
rect 8389 3723 8447 3729
rect 8389 3689 8401 3723
rect 8435 3720 8447 3723
rect 18141 3723 18199 3729
rect 8435 3692 14228 3720
rect 8435 3689 8447 3692
rect 8389 3683 8447 3689
rect 2225 3655 2283 3661
rect 2225 3621 2237 3655
rect 2271 3652 2283 3655
rect 2498 3652 2504 3664
rect 2271 3624 2504 3652
rect 2271 3621 2283 3624
rect 2225 3615 2283 3621
rect 2498 3612 2504 3624
rect 2556 3612 2562 3664
rect 4341 3655 4399 3661
rect 4341 3621 4353 3655
rect 4387 3652 4399 3655
rect 6638 3652 6644 3664
rect 4387 3624 6644 3652
rect 4387 3621 4399 3624
rect 4341 3615 4399 3621
rect 6638 3612 6644 3624
rect 6696 3612 6702 3664
rect 6914 3652 6920 3664
rect 6875 3624 6920 3652
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 8938 3652 8944 3664
rect 8899 3624 8944 3652
rect 8938 3612 8944 3624
rect 8996 3612 9002 3664
rect 10870 3652 10876 3664
rect 10831 3624 10876 3652
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 12483 3655 12541 3661
rect 12483 3621 12495 3655
rect 12529 3652 12541 3655
rect 12618 3652 12624 3664
rect 12529 3624 12624 3652
rect 12529 3621 12541 3624
rect 12483 3615 12541 3621
rect 12618 3612 12624 3624
rect 12676 3612 12682 3664
rect 13262 3612 13268 3664
rect 13320 3652 13326 3664
rect 13357 3655 13415 3661
rect 13357 3652 13369 3655
rect 13320 3624 13369 3652
rect 13320 3612 13326 3624
rect 13357 3621 13369 3624
rect 13403 3621 13415 3655
rect 14090 3652 14096 3664
rect 14051 3624 14096 3652
rect 13357 3615 13415 3621
rect 14090 3612 14096 3624
rect 14148 3612 14154 3664
rect 14200 3652 14228 3692
rect 18141 3689 18153 3723
rect 18187 3720 18199 3723
rect 19242 3720 19248 3732
rect 18187 3692 19248 3720
rect 18187 3689 18199 3692
rect 18141 3683 18199 3689
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 19426 3720 19432 3732
rect 19387 3692 19432 3720
rect 19426 3680 19432 3692
rect 19484 3680 19490 3732
rect 20070 3680 20076 3732
rect 20128 3720 20134 3732
rect 25958 3720 25964 3732
rect 20128 3692 25964 3720
rect 20128 3680 20134 3692
rect 25958 3680 25964 3692
rect 26016 3680 26022 3732
rect 27890 3680 27896 3732
rect 27948 3720 27954 3732
rect 27948 3692 37228 3720
rect 27948 3680 27954 3692
rect 14200 3624 22094 3652
rect 1394 3544 1400 3596
rect 1452 3584 1458 3596
rect 1857 3587 1915 3593
rect 1857 3584 1869 3587
rect 1452 3556 1869 3584
rect 1452 3544 1458 3556
rect 1857 3553 1869 3556
rect 1903 3553 1915 3587
rect 1857 3547 1915 3553
rect 3326 3544 3332 3596
rect 3384 3584 3390 3596
rect 3421 3587 3479 3593
rect 3421 3584 3433 3587
rect 3384 3556 3433 3584
rect 3384 3544 3390 3556
rect 3421 3553 3433 3556
rect 3467 3553 3479 3587
rect 3421 3547 3479 3553
rect 4982 3544 4988 3596
rect 5040 3584 5046 3596
rect 5077 3587 5135 3593
rect 5077 3584 5089 3587
rect 5040 3556 5089 3584
rect 5040 3544 5046 3556
rect 5077 3553 5089 3556
rect 5123 3553 5135 3587
rect 5077 3547 5135 3553
rect 5721 3587 5779 3593
rect 5721 3553 5733 3587
rect 5767 3553 5779 3587
rect 5721 3547 5779 3553
rect 7561 3587 7619 3593
rect 7561 3553 7573 3587
rect 7607 3584 7619 3587
rect 7834 3584 7840 3596
rect 7607 3556 7840 3584
rect 7607 3553 7619 3556
rect 7561 3547 7619 3553
rect 106 3476 112 3528
rect 164 3516 170 3528
rect 1302 3516 1308 3528
rect 164 3488 1308 3516
rect 164 3476 170 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 3970 3476 3976 3528
rect 4028 3516 4034 3528
rect 5736 3516 5764 3547
rect 7834 3544 7840 3556
rect 7892 3544 7898 3596
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3584 8263 3587
rect 8478 3584 8484 3596
rect 8251 3556 8484 3584
rect 8251 3553 8263 3556
rect 8205 3547 8263 3553
rect 8478 3544 8484 3556
rect 8536 3544 8542 3596
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 9585 3587 9643 3593
rect 9585 3584 9597 3587
rect 9548 3556 9597 3584
rect 9548 3544 9554 3556
rect 9585 3553 9597 3556
rect 9631 3553 9643 3587
rect 9585 3547 9643 3553
rect 12802 3544 12808 3596
rect 12860 3584 12866 3596
rect 13081 3587 13139 3593
rect 13081 3584 13093 3587
rect 12860 3556 13093 3584
rect 12860 3544 12866 3556
rect 13081 3553 13093 3556
rect 13127 3553 13139 3587
rect 13081 3547 13139 3553
rect 14829 3587 14887 3593
rect 14829 3553 14841 3587
rect 14875 3584 14887 3587
rect 14918 3584 14924 3596
rect 14875 3556 14924 3584
rect 14875 3553 14887 3556
rect 14829 3547 14887 3553
rect 14918 3544 14924 3556
rect 14976 3544 14982 3596
rect 15746 3584 15752 3596
rect 15707 3556 15752 3584
rect 15746 3544 15752 3556
rect 15804 3544 15810 3596
rect 17954 3584 17960 3596
rect 17915 3556 17960 3584
rect 17954 3544 17960 3556
rect 18012 3544 18018 3596
rect 19242 3584 19248 3596
rect 19203 3556 19248 3584
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 20073 3587 20131 3593
rect 20073 3553 20085 3587
rect 20119 3584 20131 3587
rect 20622 3584 20628 3596
rect 20119 3556 20628 3584
rect 20119 3553 20131 3556
rect 20073 3547 20131 3553
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 20772 3556 20817 3584
rect 20772 3544 20778 3556
rect 20898 3544 20904 3596
rect 20956 3584 20962 3596
rect 21545 3587 21603 3593
rect 21545 3584 21557 3587
rect 20956 3556 21557 3584
rect 20956 3544 20962 3556
rect 21545 3553 21557 3556
rect 21591 3553 21603 3587
rect 22066 3584 22094 3624
rect 25314 3612 25320 3664
rect 25372 3652 25378 3664
rect 26694 3652 26700 3664
rect 25372 3624 26700 3652
rect 25372 3612 25378 3624
rect 26694 3612 26700 3624
rect 26752 3612 26758 3664
rect 27982 3612 27988 3664
rect 28040 3652 28046 3664
rect 29362 3652 29368 3664
rect 28040 3624 29368 3652
rect 28040 3612 28046 3624
rect 29362 3612 29368 3624
rect 29420 3612 29426 3664
rect 29457 3655 29515 3661
rect 29457 3621 29469 3655
rect 29503 3652 29515 3655
rect 30190 3652 30196 3664
rect 29503 3624 30196 3652
rect 29503 3621 29515 3624
rect 29457 3615 29515 3621
rect 30190 3612 30196 3624
rect 30248 3612 30254 3664
rect 30377 3655 30435 3661
rect 30377 3621 30389 3655
rect 30423 3652 30435 3655
rect 30423 3624 30512 3652
rect 30423 3621 30435 3624
rect 30377 3615 30435 3621
rect 22557 3587 22615 3593
rect 22557 3584 22569 3587
rect 22066 3556 22569 3584
rect 21545 3547 21603 3553
rect 22557 3553 22569 3556
rect 22603 3553 22615 3587
rect 22557 3547 22615 3553
rect 23201 3587 23259 3593
rect 23201 3553 23213 3587
rect 23247 3553 23259 3587
rect 23201 3547 23259 3553
rect 4028 3488 5764 3516
rect 12069 3519 12127 3525
rect 4028 3476 4034 3488
rect 12069 3485 12081 3519
rect 12115 3516 12127 3519
rect 16574 3516 16580 3528
rect 12115 3488 16580 3516
rect 12115 3485 12127 3488
rect 12069 3479 12127 3485
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 4525 3451 4583 3457
rect 4525 3448 4537 3451
rect 2746 3420 4537 3448
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 2746 3380 2774 3420
rect 4525 3417 4537 3420
rect 4571 3417 4583 3451
rect 4525 3411 4583 3417
rect 9769 3451 9827 3457
rect 9769 3417 9781 3451
rect 9815 3448 9827 3451
rect 23216 3448 23244 3547
rect 23842 3544 23848 3596
rect 23900 3584 23906 3596
rect 24029 3587 24087 3593
rect 24029 3584 24041 3587
rect 23900 3556 24041 3584
rect 23900 3544 23906 3556
rect 24029 3553 24041 3556
rect 24075 3553 24087 3587
rect 24029 3547 24087 3553
rect 24581 3587 24639 3593
rect 24581 3553 24593 3587
rect 24627 3584 24639 3587
rect 24670 3584 24676 3596
rect 24627 3556 24676 3584
rect 24627 3553 24639 3556
rect 24581 3547 24639 3553
rect 24670 3544 24676 3556
rect 24728 3544 24734 3596
rect 25501 3587 25559 3593
rect 25501 3553 25513 3587
rect 25547 3584 25559 3587
rect 26326 3584 26332 3596
rect 25547 3556 26332 3584
rect 25547 3553 25559 3556
rect 25501 3547 25559 3553
rect 26326 3544 26332 3556
rect 26384 3544 26390 3596
rect 26421 3587 26479 3593
rect 26421 3553 26433 3587
rect 26467 3553 26479 3587
rect 27893 3587 27951 3593
rect 27893 3584 27905 3587
rect 26421 3547 26479 3553
rect 27724 3556 27905 3584
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 26436 3516 26464 3547
rect 24268 3488 26464 3516
rect 24268 3476 24274 3488
rect 27522 3476 27528 3528
rect 27580 3516 27586 3528
rect 27724 3516 27752 3556
rect 27893 3553 27905 3556
rect 27939 3553 27951 3587
rect 27893 3547 27951 3553
rect 28721 3587 28779 3593
rect 28721 3553 28733 3587
rect 28767 3553 28779 3587
rect 28721 3547 28779 3553
rect 27580 3488 27752 3516
rect 27580 3476 27586 3488
rect 27798 3476 27804 3528
rect 27856 3516 27862 3528
rect 28736 3516 28764 3547
rect 27856 3488 28764 3516
rect 27856 3476 27862 3488
rect 28810 3476 28816 3528
rect 28868 3516 28874 3528
rect 29454 3516 29460 3528
rect 28868 3488 29460 3516
rect 28868 3476 28874 3488
rect 29454 3476 29460 3488
rect 29512 3476 29518 3528
rect 30484 3516 30512 3624
rect 31570 3612 31576 3664
rect 31628 3652 31634 3664
rect 35529 3655 35587 3661
rect 35529 3652 35541 3655
rect 31628 3624 35541 3652
rect 31628 3612 31634 3624
rect 35529 3621 35541 3624
rect 35575 3621 35587 3655
rect 36262 3652 36268 3664
rect 36223 3624 36268 3652
rect 35529 3615 35587 3621
rect 36262 3612 36268 3624
rect 36320 3612 36326 3664
rect 37200 3661 37228 3692
rect 37185 3655 37243 3661
rect 37185 3621 37197 3655
rect 37231 3621 37243 3655
rect 37185 3615 37243 3621
rect 31018 3584 31024 3596
rect 30979 3556 31024 3584
rect 31018 3544 31024 3556
rect 31076 3544 31082 3596
rect 31110 3544 31116 3596
rect 31168 3584 31174 3596
rect 31665 3587 31723 3593
rect 31665 3584 31677 3587
rect 31168 3556 31677 3584
rect 31168 3544 31174 3556
rect 31665 3553 31677 3556
rect 31711 3553 31723 3587
rect 31665 3547 31723 3553
rect 31754 3544 31760 3596
rect 31812 3584 31818 3596
rect 33597 3587 33655 3593
rect 33597 3584 33609 3587
rect 31812 3556 33609 3584
rect 31812 3544 31818 3556
rect 33597 3553 33609 3556
rect 33643 3553 33655 3587
rect 34330 3584 34336 3596
rect 34291 3556 34336 3584
rect 33597 3547 33655 3553
rect 34330 3544 34336 3556
rect 34388 3544 34394 3596
rect 36630 3584 36636 3596
rect 35866 3556 36636 3584
rect 30484 3488 30788 3516
rect 25038 3448 25044 3460
rect 9815 3420 23244 3448
rect 23308 3420 25044 3448
rect 9815 3417 9827 3420
rect 9769 3411 9827 3417
rect 1728 3352 2774 3380
rect 1728 3340 1734 3352
rect 4982 3340 4988 3392
rect 5040 3380 5046 3392
rect 5169 3383 5227 3389
rect 5169 3380 5181 3383
rect 5040 3352 5181 3380
rect 5040 3340 5046 3352
rect 5169 3349 5181 3352
rect 5215 3349 5227 3383
rect 5169 3343 5227 3349
rect 6270 3340 6276 3392
rect 6328 3380 6334 3392
rect 7009 3383 7067 3389
rect 7009 3380 7021 3383
rect 6328 3352 7021 3380
rect 6328 3340 6334 3352
rect 7009 3349 7021 3352
rect 7055 3349 7067 3383
rect 7009 3343 7067 3349
rect 8846 3340 8852 3392
rect 8904 3380 8910 3392
rect 9033 3383 9091 3389
rect 9033 3380 9045 3383
rect 8904 3352 9045 3380
rect 8904 3340 8910 3352
rect 9033 3349 9045 3352
rect 9079 3349 9091 3383
rect 9033 3343 9091 3349
rect 10778 3340 10784 3392
rect 10836 3380 10842 3392
rect 10965 3383 11023 3389
rect 10965 3380 10977 3383
rect 10836 3352 10977 3380
rect 10836 3340 10842 3352
rect 10965 3349 10977 3352
rect 11011 3349 11023 3383
rect 10965 3343 11023 3349
rect 12434 3340 12440 3392
rect 12492 3380 12498 3392
rect 12621 3383 12679 3389
rect 12492 3352 12537 3380
rect 12492 3340 12498 3352
rect 12621 3349 12633 3383
rect 12667 3380 12679 3383
rect 13354 3380 13360 3392
rect 12667 3352 13360 3380
rect 12667 3349 12679 3352
rect 12621 3343 12679 3349
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 13630 3340 13636 3392
rect 13688 3380 13694 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 13688 3352 14197 3380
rect 13688 3340 13694 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 14185 3343 14243 3349
rect 14734 3340 14740 3392
rect 14792 3380 14798 3392
rect 14921 3383 14979 3389
rect 14921 3380 14933 3383
rect 14792 3352 14933 3380
rect 14792 3340 14798 3352
rect 14921 3349 14933 3352
rect 14967 3349 14979 3383
rect 14921 3343 14979 3349
rect 15654 3340 15660 3392
rect 15712 3380 15718 3392
rect 15841 3383 15899 3389
rect 15841 3380 15853 3383
rect 15712 3352 15853 3380
rect 15712 3340 15718 3352
rect 15841 3349 15853 3352
rect 15887 3349 15899 3383
rect 15841 3343 15899 3349
rect 19886 3340 19892 3392
rect 19944 3380 19950 3392
rect 20165 3383 20223 3389
rect 20165 3380 20177 3383
rect 19944 3352 20177 3380
rect 19944 3340 19950 3352
rect 20165 3349 20177 3352
rect 20211 3349 20223 3383
rect 20165 3343 20223 3349
rect 20901 3383 20959 3389
rect 20901 3349 20913 3383
rect 20947 3380 20959 3383
rect 20990 3380 20996 3392
rect 20947 3352 20996 3380
rect 20947 3349 20959 3352
rect 20901 3343 20959 3349
rect 20990 3340 20996 3352
rect 21048 3340 21054 3392
rect 21358 3380 21364 3392
rect 21319 3352 21364 3380
rect 21358 3340 21364 3352
rect 21416 3340 21422 3392
rect 22741 3383 22799 3389
rect 22741 3349 22753 3383
rect 22787 3380 22799 3383
rect 23308 3380 23336 3420
rect 25038 3408 25044 3420
rect 25096 3408 25102 3460
rect 25130 3408 25136 3460
rect 25188 3448 25194 3460
rect 30006 3448 30012 3460
rect 25188 3420 30012 3448
rect 25188 3408 25194 3420
rect 30006 3408 30012 3420
rect 30064 3408 30070 3460
rect 30374 3408 30380 3460
rect 30432 3448 30438 3460
rect 30561 3451 30619 3457
rect 30561 3448 30573 3451
rect 30432 3420 30573 3448
rect 30432 3408 30438 3420
rect 30561 3417 30573 3420
rect 30607 3417 30619 3451
rect 30561 3411 30619 3417
rect 22787 3352 23336 3380
rect 23385 3383 23443 3389
rect 22787 3349 22799 3352
rect 22741 3343 22799 3349
rect 23385 3349 23397 3383
rect 23431 3380 23443 3383
rect 23750 3380 23756 3392
rect 23431 3352 23756 3380
rect 23431 3349 23443 3352
rect 23385 3343 23443 3349
rect 23750 3340 23756 3352
rect 23808 3340 23814 3392
rect 23845 3383 23903 3389
rect 23845 3349 23857 3383
rect 23891 3380 23903 3383
rect 24394 3380 24400 3392
rect 23891 3352 24400 3380
rect 23891 3349 23903 3352
rect 23845 3343 23903 3349
rect 24394 3340 24400 3352
rect 24452 3340 24458 3392
rect 24486 3340 24492 3392
rect 24544 3380 24550 3392
rect 24673 3383 24731 3389
rect 24673 3380 24685 3383
rect 24544 3352 24685 3380
rect 24544 3340 24550 3352
rect 24673 3349 24685 3352
rect 24719 3349 24731 3383
rect 24673 3343 24731 3349
rect 25406 3340 25412 3392
rect 25464 3380 25470 3392
rect 25593 3383 25651 3389
rect 25593 3380 25605 3383
rect 25464 3352 25605 3380
rect 25464 3340 25470 3352
rect 25593 3349 25605 3352
rect 25639 3349 25651 3383
rect 26602 3380 26608 3392
rect 26563 3352 26608 3380
rect 25593 3343 25651 3349
rect 26602 3340 26608 3352
rect 26660 3340 26666 3392
rect 27430 3340 27436 3392
rect 27488 3380 27494 3392
rect 27985 3383 28043 3389
rect 27985 3380 27997 3383
rect 27488 3352 27997 3380
rect 27488 3340 27494 3352
rect 27985 3349 27997 3352
rect 28031 3349 28043 3383
rect 28534 3380 28540 3392
rect 28495 3352 28540 3380
rect 27985 3343 28043 3349
rect 28534 3340 28540 3352
rect 28592 3340 28598 3392
rect 29362 3340 29368 3392
rect 29420 3380 29426 3392
rect 29549 3383 29607 3389
rect 29549 3380 29561 3383
rect 29420 3352 29561 3380
rect 29420 3340 29426 3352
rect 29549 3349 29561 3352
rect 29595 3349 29607 3383
rect 30760 3380 30788 3488
rect 30834 3476 30840 3528
rect 30892 3516 30898 3528
rect 31478 3516 31484 3528
rect 30892 3488 31484 3516
rect 30892 3476 30898 3488
rect 31478 3476 31484 3488
rect 31536 3476 31542 3528
rect 35866 3516 35894 3556
rect 36630 3544 36636 3556
rect 36688 3544 36694 3596
rect 31726 3488 35894 3516
rect 31205 3451 31263 3457
rect 31205 3417 31217 3451
rect 31251 3448 31263 3451
rect 31726 3448 31754 3488
rect 31251 3420 31754 3448
rect 31849 3451 31907 3457
rect 31251 3417 31263 3420
rect 31205 3411 31263 3417
rect 31849 3417 31861 3451
rect 31895 3448 31907 3451
rect 34606 3448 34612 3460
rect 31895 3420 34612 3448
rect 31895 3417 31907 3420
rect 31849 3411 31907 3417
rect 34606 3408 34612 3420
rect 34664 3408 34670 3460
rect 35713 3451 35771 3457
rect 35713 3417 35725 3451
rect 35759 3448 35771 3451
rect 36814 3448 36820 3460
rect 35759 3420 36820 3448
rect 35759 3417 35771 3420
rect 35713 3411 35771 3417
rect 36814 3408 36820 3420
rect 36872 3408 36878 3460
rect 37369 3451 37427 3457
rect 37369 3417 37381 3451
rect 37415 3448 37427 3451
rect 37826 3448 37832 3460
rect 37415 3420 37832 3448
rect 37415 3417 37427 3420
rect 37369 3411 37427 3417
rect 37826 3408 37832 3420
rect 37884 3408 37890 3460
rect 32306 3380 32312 3392
rect 30760 3352 32312 3380
rect 29549 3343 29607 3349
rect 32306 3340 32312 3352
rect 32364 3340 32370 3392
rect 33686 3380 33692 3392
rect 33647 3352 33692 3380
rect 33686 3340 33692 3352
rect 33744 3340 33750 3392
rect 34238 3340 34244 3392
rect 34296 3380 34302 3392
rect 34425 3383 34483 3389
rect 34425 3380 34437 3383
rect 34296 3352 34437 3380
rect 34296 3340 34302 3352
rect 34425 3349 34437 3352
rect 34471 3349 34483 3383
rect 34425 3343 34483 3349
rect 36170 3340 36176 3392
rect 36228 3380 36234 3392
rect 36357 3383 36415 3389
rect 36357 3380 36369 3383
rect 36228 3352 36369 3380
rect 36228 3340 36234 3352
rect 36357 3349 36369 3352
rect 36403 3349 36415 3383
rect 36357 3343 36415 3349
rect 1104 3290 38824 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 38824 3290
rect 1104 3216 38824 3238
rect 2133 3179 2191 3185
rect 2133 3145 2145 3179
rect 2179 3176 2191 3179
rect 2314 3176 2320 3188
rect 2179 3148 2320 3176
rect 2179 3145 2191 3148
rect 2133 3139 2191 3145
rect 2314 3136 2320 3148
rect 2372 3136 2378 3188
rect 3050 3176 3056 3188
rect 3011 3148 3056 3176
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 7374 3176 7380 3188
rect 7335 3148 7380 3176
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 9674 3176 9680 3188
rect 9635 3148 9680 3176
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 16482 3176 16488 3188
rect 9784 3148 15608 3176
rect 16443 3148 16488 3176
rect 2038 3068 2044 3120
rect 2096 3108 2102 3120
rect 5166 3108 5172 3120
rect 2096 3080 5172 3108
rect 2096 3068 2102 3080
rect 5166 3068 5172 3080
rect 5224 3068 5230 3120
rect 7558 3068 7564 3120
rect 7616 3108 7622 3120
rect 9784 3108 9812 3148
rect 7616 3080 9812 3108
rect 7616 3068 7622 3080
rect 10502 3068 10508 3120
rect 10560 3108 10566 3120
rect 10560 3080 13308 3108
rect 10560 3068 10566 3080
rect 4798 3040 4804 3052
rect 4759 3012 4804 3040
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 6178 3040 6184 3052
rect 6139 3012 6184 3040
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 11422 3040 11428 3052
rect 11383 3012 11428 3040
rect 11422 3000 11428 3012
rect 11480 3000 11486 3052
rect 12342 3040 12348 3052
rect 12303 3012 12348 3040
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 12526 3000 12532 3052
rect 12584 3040 12590 3052
rect 12802 3040 12808 3052
rect 12584 3012 12808 3040
rect 12584 3000 12590 3012
rect 12802 3000 12808 3012
rect 12860 3000 12866 3052
rect 13280 3049 13308 3080
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3009 13323 3043
rect 13265 3003 13323 3009
rect 13354 3000 13360 3052
rect 13412 3040 13418 3052
rect 15580 3049 15608 3148
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 20254 3176 20260 3188
rect 20215 3148 20260 3176
rect 20254 3136 20260 3148
rect 20312 3136 20318 3188
rect 20346 3136 20352 3188
rect 20404 3176 20410 3188
rect 24210 3176 24216 3188
rect 20404 3148 24216 3176
rect 20404 3136 20410 3148
rect 24210 3136 24216 3148
rect 24268 3136 24274 3188
rect 24394 3136 24400 3188
rect 24452 3176 24458 3188
rect 25501 3179 25559 3185
rect 25501 3176 25513 3179
rect 24452 3148 25513 3176
rect 24452 3136 24458 3148
rect 25501 3145 25513 3148
rect 25547 3145 25559 3179
rect 25501 3139 25559 3145
rect 25869 3179 25927 3185
rect 25869 3145 25881 3179
rect 25915 3176 25927 3179
rect 27522 3176 27528 3188
rect 25915 3148 27528 3176
rect 25915 3145 25927 3148
rect 25869 3139 25927 3145
rect 27522 3136 27528 3148
rect 27580 3136 27586 3188
rect 27801 3179 27859 3185
rect 27801 3145 27813 3179
rect 27847 3176 27859 3179
rect 28534 3176 28540 3188
rect 27847 3148 28540 3176
rect 27847 3145 27859 3148
rect 27801 3139 27859 3145
rect 28534 3136 28540 3148
rect 28592 3136 28598 3188
rect 28626 3136 28632 3188
rect 28684 3176 28690 3188
rect 30650 3176 30656 3188
rect 28684 3148 30656 3176
rect 28684 3136 28690 3148
rect 30650 3136 30656 3148
rect 30708 3136 30714 3188
rect 30834 3176 30840 3188
rect 30795 3148 30840 3176
rect 30834 3136 30840 3148
rect 30892 3136 30898 3188
rect 30929 3179 30987 3185
rect 30929 3145 30941 3179
rect 30975 3176 30987 3179
rect 33686 3176 33692 3188
rect 30975 3148 33692 3176
rect 30975 3145 30987 3148
rect 30929 3139 30987 3145
rect 33686 3136 33692 3148
rect 33744 3136 33750 3188
rect 35897 3179 35955 3185
rect 35897 3145 35909 3179
rect 35943 3176 35955 3179
rect 38194 3176 38200 3188
rect 35943 3148 38200 3176
rect 35943 3145 35955 3148
rect 35897 3139 35955 3145
rect 38194 3136 38200 3148
rect 38252 3136 38258 3188
rect 19794 3108 19800 3120
rect 15672 3080 19800 3108
rect 15565 3043 15623 3049
rect 13412 3012 15516 3040
rect 13412 3000 13418 3012
rect 382 2932 388 2984
rect 440 2972 446 2984
rect 2777 2975 2835 2981
rect 2777 2972 2789 2975
rect 440 2944 2789 2972
rect 440 2932 446 2944
rect 2777 2941 2789 2944
rect 2823 2941 2835 2975
rect 4614 2972 4620 2984
rect 4575 2944 4620 2972
rect 2777 2935 2835 2941
rect 4614 2932 4620 2944
rect 4672 2932 4678 2984
rect 5902 2972 5908 2984
rect 5863 2944 5908 2972
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 7190 2972 7196 2984
rect 7151 2944 7196 2972
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 8018 2972 8024 2984
rect 7979 2944 8024 2972
rect 8018 2932 8024 2944
rect 8076 2932 8082 2984
rect 9214 2932 9220 2984
rect 9272 2972 9278 2984
rect 9493 2975 9551 2981
rect 9493 2972 9505 2975
rect 9272 2944 9505 2972
rect 9272 2932 9278 2944
rect 9493 2941 9505 2944
rect 9539 2941 9551 2975
rect 10318 2972 10324 2984
rect 10279 2944 10324 2972
rect 9493 2935 9551 2941
rect 10318 2932 10324 2944
rect 10376 2932 10382 2984
rect 11146 2972 11152 2984
rect 11107 2944 11152 2972
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 11440 2944 12081 2972
rect 11440 2916 11468 2944
rect 12069 2941 12081 2944
rect 12115 2941 12127 2975
rect 13078 2972 13084 2984
rect 13039 2944 13084 2972
rect 12069 2935 12127 2941
rect 13078 2932 13084 2944
rect 13136 2932 13142 2984
rect 14737 2975 14795 2981
rect 14737 2941 14749 2975
rect 14783 2972 14795 2975
rect 15010 2972 15016 2984
rect 14783 2944 15016 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 15010 2932 15016 2944
rect 15068 2932 15074 2984
rect 15378 2972 15384 2984
rect 15339 2944 15384 2972
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 15488 2972 15516 3012
rect 15565 3009 15577 3043
rect 15611 3009 15623 3043
rect 15565 3003 15623 3009
rect 15672 2972 15700 3080
rect 19794 3068 19800 3080
rect 19852 3068 19858 3120
rect 20146 3111 20204 3117
rect 20146 3077 20158 3111
rect 20192 3108 20204 3111
rect 21910 3108 21916 3120
rect 20192 3080 21916 3108
rect 20192 3077 20204 3080
rect 20146 3071 20204 3077
rect 21910 3068 21916 3080
rect 21968 3068 21974 3120
rect 25314 3068 25320 3120
rect 25372 3117 25378 3120
rect 25372 3111 25421 3117
rect 25372 3077 25375 3111
rect 25409 3077 25421 3111
rect 25372 3071 25421 3077
rect 27690 3111 27748 3117
rect 27690 3077 27702 3111
rect 27736 3108 27748 3111
rect 28994 3108 29000 3120
rect 27736 3080 29000 3108
rect 27736 3077 27748 3080
rect 27690 3071 27748 3077
rect 25372 3068 25378 3071
rect 28994 3068 29000 3080
rect 29052 3068 29058 3120
rect 31754 3108 31760 3120
rect 30576 3080 31760 3108
rect 17586 3040 17592 3052
rect 17547 3012 17592 3040
rect 17586 3000 17592 3012
rect 17644 3000 17650 3052
rect 18598 3040 18604 3052
rect 18559 3012 18604 3040
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 20349 3043 20407 3049
rect 20349 3009 20361 3043
rect 20395 3040 20407 3043
rect 21358 3040 21364 3052
rect 20395 3012 21364 3040
rect 20395 3009 20407 3012
rect 20349 3003 20407 3009
rect 21358 3000 21364 3012
rect 21416 3000 21422 3052
rect 25590 3000 25596 3052
rect 25648 3040 25654 3052
rect 27893 3043 27951 3049
rect 25648 3012 25690 3040
rect 25648 3000 25654 3012
rect 27893 3009 27905 3043
rect 27939 3040 27951 3043
rect 28074 3040 28080 3052
rect 27939 3012 28080 3040
rect 27939 3009 27951 3012
rect 27893 3003 27951 3009
rect 28074 3000 28080 3012
rect 28132 3000 28138 3052
rect 28261 3043 28319 3049
rect 28261 3009 28273 3043
rect 28307 3040 28319 3043
rect 29730 3040 29736 3052
rect 28307 3012 29736 3040
rect 28307 3009 28319 3012
rect 28261 3003 28319 3009
rect 29730 3000 29736 3012
rect 29788 3000 29794 3052
rect 30469 3043 30527 3049
rect 30469 3009 30481 3043
rect 30515 3040 30527 3043
rect 30576 3040 30604 3080
rect 31754 3068 31760 3080
rect 31812 3068 31818 3120
rect 32122 3068 32128 3120
rect 32180 3108 32186 3120
rect 34425 3111 34483 3117
rect 34425 3108 34437 3111
rect 32180 3080 34437 3108
rect 32180 3068 32186 3080
rect 34425 3077 34437 3080
rect 34471 3077 34483 3111
rect 34425 3071 34483 3077
rect 34793 3111 34851 3117
rect 34793 3077 34805 3111
rect 34839 3108 34851 3111
rect 37182 3108 37188 3120
rect 34839 3080 37188 3108
rect 34839 3077 34851 3080
rect 34793 3071 34851 3077
rect 37182 3068 37188 3080
rect 37240 3068 37246 3120
rect 30515 3012 30604 3040
rect 31021 3043 31079 3049
rect 30515 3009 30527 3012
rect 30469 3003 30527 3009
rect 31021 3009 31033 3043
rect 31067 3040 31079 3043
rect 32030 3040 32036 3052
rect 31067 3012 32036 3040
rect 31067 3009 31079 3012
rect 31021 3003 31079 3009
rect 32030 3000 32036 3012
rect 32088 3000 32094 3052
rect 16298 2972 16304 2984
rect 15488 2944 15700 2972
rect 16259 2944 16304 2972
rect 16298 2932 16304 2944
rect 16356 2932 16362 2984
rect 17310 2972 17316 2984
rect 17271 2944 17316 2972
rect 17310 2932 17316 2944
rect 17368 2932 17374 2984
rect 18322 2972 18328 2984
rect 18283 2944 18328 2972
rect 18322 2932 18328 2944
rect 18380 2932 18386 2984
rect 19981 2975 20039 2981
rect 19981 2941 19993 2975
rect 20027 2972 20039 2975
rect 20438 2972 20444 2984
rect 20027 2944 20444 2972
rect 20027 2941 20039 2944
rect 19981 2935 20039 2941
rect 20438 2932 20444 2944
rect 20496 2932 20502 2984
rect 20530 2932 20536 2984
rect 20588 2972 20594 2984
rect 21453 2975 21511 2981
rect 21453 2972 21465 2975
rect 20588 2944 21465 2972
rect 20588 2932 20594 2944
rect 21453 2941 21465 2944
rect 21499 2941 21511 2975
rect 22738 2972 22744 2984
rect 22699 2944 22744 2972
rect 21453 2935 21511 2941
rect 22738 2932 22744 2944
rect 22796 2932 22802 2984
rect 23566 2972 23572 2984
rect 23527 2944 23572 2972
rect 23566 2932 23572 2944
rect 23624 2932 23630 2984
rect 23750 2932 23756 2984
rect 23808 2972 23814 2984
rect 25225 2975 25283 2981
rect 23808 2944 25176 2972
rect 23808 2932 23814 2944
rect 1854 2904 1860 2916
rect 1815 2876 1860 2904
rect 1854 2864 1860 2876
rect 1912 2864 1918 2916
rect 11422 2864 11428 2916
rect 11480 2864 11486 2916
rect 16574 2864 16580 2916
rect 16632 2904 16638 2916
rect 21266 2904 21272 2916
rect 16632 2876 20668 2904
rect 21227 2876 21272 2904
rect 16632 2864 16638 2876
rect 750 2796 756 2848
rect 808 2836 814 2848
rect 3142 2836 3148 2848
rect 808 2808 3148 2836
rect 808 2796 814 2808
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 7558 2796 7564 2848
rect 7616 2836 7622 2848
rect 8113 2839 8171 2845
rect 8113 2836 8125 2839
rect 7616 2808 8125 2836
rect 7616 2796 7622 2808
rect 8113 2805 8125 2808
rect 8159 2805 8171 2839
rect 8113 2799 8171 2805
rect 9858 2796 9864 2848
rect 9916 2836 9922 2848
rect 10413 2839 10471 2845
rect 10413 2836 10425 2839
rect 9916 2808 10425 2836
rect 9916 2796 9922 2808
rect 10413 2805 10425 2808
rect 10459 2805 10471 2839
rect 10413 2799 10471 2805
rect 14921 2839 14979 2845
rect 14921 2805 14933 2839
rect 14967 2836 14979 2839
rect 20346 2836 20352 2848
rect 14967 2808 20352 2836
rect 14967 2805 14979 2808
rect 14921 2799 14979 2805
rect 20346 2796 20352 2808
rect 20404 2796 20410 2848
rect 20640 2845 20668 2876
rect 21266 2864 21272 2876
rect 21324 2864 21330 2916
rect 22005 2907 22063 2913
rect 22005 2873 22017 2907
rect 22051 2904 22063 2907
rect 25148 2904 25176 2944
rect 25225 2941 25237 2975
rect 25271 2972 25283 2975
rect 26234 2972 26240 2984
rect 25271 2944 26240 2972
rect 25271 2941 25283 2944
rect 25225 2935 25283 2941
rect 26234 2932 26240 2944
rect 26292 2932 26298 2984
rect 26513 2975 26571 2981
rect 26513 2941 26525 2975
rect 26559 2972 26571 2975
rect 26786 2972 26792 2984
rect 26559 2944 26792 2972
rect 26559 2941 26571 2944
rect 26513 2935 26571 2941
rect 26786 2932 26792 2944
rect 26844 2932 26850 2984
rect 27525 2975 27583 2981
rect 27525 2941 27537 2975
rect 27571 2972 27583 2975
rect 28534 2972 28540 2984
rect 27571 2944 28540 2972
rect 27571 2941 27583 2944
rect 27525 2935 27583 2941
rect 28534 2932 28540 2944
rect 28592 2932 28598 2984
rect 28813 2975 28871 2981
rect 28813 2941 28825 2975
rect 28859 2972 28871 2975
rect 31202 2972 31208 2984
rect 28859 2944 31208 2972
rect 28859 2941 28871 2944
rect 28813 2935 28871 2941
rect 31202 2932 31208 2944
rect 31260 2932 31266 2984
rect 31294 2932 31300 2984
rect 31352 2972 31358 2984
rect 31389 2975 31447 2981
rect 31389 2972 31401 2975
rect 31352 2944 31401 2972
rect 31352 2932 31358 2944
rect 31389 2941 31401 2944
rect 31435 2941 31447 2975
rect 31389 2935 31447 2941
rect 31941 2975 31999 2981
rect 31941 2941 31953 2975
rect 31987 2972 31999 2975
rect 32214 2972 32220 2984
rect 31987 2944 32220 2972
rect 31987 2941 31999 2944
rect 31941 2935 31999 2941
rect 32214 2932 32220 2944
rect 32272 2932 32278 2984
rect 32677 2975 32735 2981
rect 32677 2941 32689 2975
rect 32723 2972 32735 2975
rect 33226 2972 33232 2984
rect 32723 2944 33232 2972
rect 32723 2941 32735 2944
rect 32677 2935 32735 2941
rect 33226 2932 33232 2944
rect 33284 2932 33290 2984
rect 33413 2975 33471 2981
rect 33413 2941 33425 2975
rect 33459 2972 33471 2975
rect 34146 2972 34152 2984
rect 33459 2944 34152 2972
rect 33459 2941 33471 2944
rect 33413 2935 33471 2941
rect 34146 2932 34152 2944
rect 34204 2932 34210 2984
rect 34425 2975 34483 2981
rect 34425 2941 34437 2975
rect 34471 2972 34483 2975
rect 34471 2944 34744 2972
rect 34471 2941 34483 2944
rect 34425 2935 34483 2941
rect 34609 2907 34667 2913
rect 34609 2904 34621 2907
rect 22051 2876 23796 2904
rect 25148 2876 34621 2904
rect 22051 2873 22063 2876
rect 22005 2867 22063 2873
rect 20625 2839 20683 2845
rect 20625 2805 20637 2839
rect 20671 2805 20683 2839
rect 20625 2799 20683 2805
rect 21542 2796 21548 2848
rect 21600 2836 21606 2848
rect 22097 2839 22155 2845
rect 22097 2836 22109 2839
rect 21600 2808 22109 2836
rect 21600 2796 21606 2808
rect 22097 2805 22109 2808
rect 22143 2805 22155 2839
rect 22097 2799 22155 2805
rect 22554 2796 22560 2848
rect 22612 2836 22618 2848
rect 22833 2839 22891 2845
rect 22833 2836 22845 2839
rect 22612 2808 22845 2836
rect 22612 2796 22618 2808
rect 22833 2805 22845 2808
rect 22879 2805 22891 2839
rect 22833 2799 22891 2805
rect 23474 2796 23480 2848
rect 23532 2836 23538 2848
rect 23661 2839 23719 2845
rect 23661 2836 23673 2839
rect 23532 2808 23673 2836
rect 23532 2796 23538 2808
rect 23661 2805 23673 2808
rect 23707 2805 23719 2839
rect 23768 2836 23796 2876
rect 34609 2873 34621 2876
rect 34655 2873 34667 2907
rect 34716 2904 34744 2944
rect 34790 2932 34796 2984
rect 34848 2972 34854 2984
rect 35713 2975 35771 2981
rect 35713 2972 35725 2975
rect 34848 2944 35725 2972
rect 34848 2932 34854 2944
rect 35713 2941 35725 2944
rect 35759 2941 35771 2975
rect 37918 2972 37924 2984
rect 37879 2944 37924 2972
rect 35713 2935 35771 2941
rect 37918 2932 37924 2944
rect 37976 2932 37982 2984
rect 36633 2907 36691 2913
rect 36633 2904 36645 2907
rect 34716 2876 36645 2904
rect 34609 2867 34667 2873
rect 36633 2873 36645 2876
rect 36679 2873 36691 2907
rect 38102 2904 38108 2916
rect 38063 2876 38108 2904
rect 36633 2867 36691 2873
rect 38102 2864 38108 2876
rect 38160 2864 38166 2916
rect 26326 2836 26332 2848
rect 23768 2808 26332 2836
rect 23661 2799 23719 2805
rect 26326 2796 26332 2808
rect 26384 2796 26390 2848
rect 26418 2796 26424 2848
rect 26476 2836 26482 2848
rect 26605 2839 26663 2845
rect 26605 2836 26617 2839
rect 26476 2808 26617 2836
rect 26476 2796 26482 2808
rect 26605 2805 26617 2808
rect 26651 2805 26663 2839
rect 26605 2799 26663 2805
rect 28350 2796 28356 2848
rect 28408 2836 28414 2848
rect 28905 2839 28963 2845
rect 28905 2836 28917 2839
rect 28408 2808 28917 2836
rect 28408 2796 28414 2808
rect 28905 2805 28917 2808
rect 28951 2805 28963 2839
rect 28905 2799 28963 2805
rect 31294 2796 31300 2848
rect 31352 2836 31358 2848
rect 32033 2839 32091 2845
rect 32033 2836 32045 2839
rect 31352 2808 32045 2836
rect 31352 2796 31358 2808
rect 32033 2805 32045 2808
rect 32079 2805 32091 2839
rect 32033 2799 32091 2805
rect 32306 2796 32312 2848
rect 32364 2836 32370 2848
rect 32769 2839 32827 2845
rect 32769 2836 32781 2839
rect 32364 2808 32781 2836
rect 32364 2796 32370 2808
rect 32769 2805 32781 2808
rect 32815 2805 32827 2839
rect 32769 2799 32827 2805
rect 33226 2796 33232 2848
rect 33284 2836 33290 2848
rect 33505 2839 33563 2845
rect 33505 2836 33517 2839
rect 33284 2808 33517 2836
rect 33284 2796 33290 2808
rect 33505 2805 33517 2808
rect 33551 2805 33563 2839
rect 33505 2799 33563 2805
rect 36538 2796 36544 2848
rect 36596 2836 36602 2848
rect 36725 2839 36783 2845
rect 36725 2836 36737 2839
rect 36596 2808 36737 2836
rect 36596 2796 36602 2808
rect 36725 2805 36737 2808
rect 36771 2805 36783 2839
rect 36725 2799 36783 2805
rect 1104 2746 38824 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 38824 2746
rect 1104 2672 38824 2694
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3053 2635 3111 2641
rect 3053 2632 3065 2635
rect 3016 2604 3065 2632
rect 3016 2592 3022 2604
rect 3053 2601 3065 2604
rect 3099 2601 3111 2635
rect 3053 2595 3111 2601
rect 4890 2592 4896 2644
rect 4948 2632 4954 2644
rect 11238 2632 11244 2644
rect 4948 2604 10456 2632
rect 11199 2604 11244 2632
rect 4948 2592 4954 2604
rect 1857 2567 1915 2573
rect 1857 2533 1869 2567
rect 1903 2564 1915 2567
rect 2866 2564 2872 2576
rect 1903 2536 2872 2564
rect 1903 2533 1915 2536
rect 1857 2527 1915 2533
rect 2866 2524 2872 2536
rect 2924 2524 2930 2576
rect 5350 2524 5356 2576
rect 5408 2564 5414 2576
rect 5813 2567 5871 2573
rect 5813 2564 5825 2567
rect 5408 2536 5825 2564
rect 5408 2524 5414 2536
rect 5813 2533 5825 2536
rect 5859 2533 5871 2567
rect 5813 2527 5871 2533
rect 8386 2524 8392 2576
rect 8444 2564 8450 2576
rect 8481 2567 8539 2573
rect 8481 2564 8493 2567
rect 8444 2536 8493 2564
rect 8444 2524 8450 2536
rect 8481 2533 8493 2536
rect 8527 2533 8539 2567
rect 8481 2527 8539 2533
rect 9950 2524 9956 2576
rect 10008 2564 10014 2576
rect 10428 2573 10456 2604
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 12894 2592 12900 2644
rect 12952 2632 12958 2644
rect 23106 2632 23112 2644
rect 12952 2604 16574 2632
rect 23067 2604 23112 2632
rect 12952 2592 12958 2604
rect 10413 2567 10471 2573
rect 10008 2536 10272 2564
rect 10008 2524 10014 2536
rect 2774 2496 2780 2508
rect 2735 2468 2780 2496
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 2958 2456 2964 2508
rect 3016 2496 3022 2508
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 3016 2468 4261 2496
rect 3016 2456 3022 2468
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 4249 2459 4307 2465
rect 5537 2499 5595 2505
rect 5537 2465 5549 2499
rect 5583 2496 5595 2499
rect 5626 2496 5632 2508
rect 5583 2468 5632 2496
rect 5583 2465 5595 2468
rect 5537 2459 5595 2465
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 8202 2496 8208 2508
rect 6972 2468 7017 2496
rect 8163 2468 8208 2496
rect 6972 2456 6978 2468
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 10134 2496 10140 2508
rect 10095 2468 10140 2496
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 10244 2496 10272 2536
rect 10413 2533 10425 2567
rect 10459 2533 10471 2567
rect 13722 2564 13728 2576
rect 10413 2527 10471 2533
rect 10520 2536 12572 2564
rect 13683 2536 13728 2564
rect 10520 2496 10548 2536
rect 10244 2468 10548 2496
rect 11057 2499 11115 2505
rect 11057 2465 11069 2499
rect 11103 2496 11115 2499
rect 12066 2496 12072 2508
rect 11103 2468 12072 2496
rect 11103 2465 11115 2468
rect 11057 2459 11115 2465
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 12253 2499 12311 2505
rect 12253 2465 12265 2499
rect 12299 2465 12311 2499
rect 12253 2459 12311 2465
rect 1578 2388 1584 2440
rect 1636 2428 1642 2440
rect 4433 2431 4491 2437
rect 4433 2428 4445 2431
rect 1636 2400 4445 2428
rect 1636 2388 1642 2400
rect 4433 2397 4445 2400
rect 4479 2397 4491 2431
rect 4433 2391 4491 2397
rect 5442 2388 5448 2440
rect 5500 2428 5506 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 5500 2400 7113 2428
rect 5500 2388 5506 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 10502 2388 10508 2440
rect 10560 2428 10566 2440
rect 12268 2428 12296 2459
rect 10560 2400 12296 2428
rect 12437 2431 12495 2437
rect 10560 2388 10566 2400
rect 12437 2397 12449 2431
rect 12483 2397 12495 2431
rect 12544 2428 12572 2536
rect 13722 2524 13728 2536
rect 13780 2524 13786 2576
rect 16390 2564 16396 2576
rect 16351 2536 16396 2564
rect 16390 2524 16396 2536
rect 16448 2524 16454 2576
rect 16546 2564 16574 2604
rect 23106 2592 23112 2604
rect 23164 2592 23170 2644
rect 24578 2632 24584 2644
rect 24539 2604 24584 2632
rect 24578 2592 24584 2604
rect 24636 2592 24642 2644
rect 27706 2592 27712 2644
rect 27764 2632 27770 2644
rect 28445 2635 28503 2641
rect 28445 2632 28457 2635
rect 27764 2604 28457 2632
rect 27764 2592 27770 2604
rect 28445 2601 28457 2604
rect 28491 2601 28503 2635
rect 28445 2595 28503 2601
rect 33410 2592 33416 2644
rect 33468 2632 33474 2644
rect 34606 2632 34612 2644
rect 33468 2604 34612 2632
rect 33468 2592 33474 2604
rect 34606 2592 34612 2604
rect 34664 2592 34670 2644
rect 35621 2635 35679 2641
rect 35621 2601 35633 2635
rect 35667 2632 35679 2635
rect 36449 2635 36507 2641
rect 36449 2632 36461 2635
rect 35667 2604 36461 2632
rect 35667 2601 35679 2604
rect 35621 2595 35679 2601
rect 36449 2601 36461 2604
rect 36495 2601 36507 2635
rect 36449 2595 36507 2601
rect 26329 2567 26387 2573
rect 26329 2564 26341 2567
rect 16546 2536 26341 2564
rect 26329 2533 26341 2536
rect 26375 2533 26387 2567
rect 32490 2564 32496 2576
rect 32451 2536 32496 2564
rect 26329 2527 26387 2533
rect 32490 2524 32496 2536
rect 32548 2524 32554 2576
rect 34057 2567 34115 2573
rect 34057 2533 34069 2567
rect 34103 2564 34115 2567
rect 35986 2564 35992 2576
rect 34103 2536 35992 2564
rect 34103 2533 34115 2536
rect 34057 2527 34115 2533
rect 35986 2524 35992 2536
rect 36044 2524 36050 2576
rect 37642 2524 37648 2576
rect 37700 2564 37706 2576
rect 37737 2567 37795 2573
rect 37737 2564 37749 2567
rect 37700 2536 37749 2564
rect 37700 2524 37706 2536
rect 37737 2533 37749 2536
rect 37783 2533 37795 2567
rect 37737 2527 37795 2533
rect 13357 2499 13415 2505
rect 13357 2465 13369 2499
rect 13403 2496 13415 2499
rect 13446 2496 13452 2508
rect 13403 2468 13452 2496
rect 13403 2465 13415 2468
rect 13357 2459 13415 2465
rect 13446 2456 13452 2468
rect 13504 2456 13510 2508
rect 14090 2456 14096 2508
rect 14148 2496 14154 2508
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14148 2468 14933 2496
rect 14148 2456 14154 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 16022 2496 16028 2508
rect 14921 2459 14979 2465
rect 15028 2468 15240 2496
rect 15983 2468 16028 2496
rect 15028 2428 15056 2468
rect 12544 2400 15056 2428
rect 15105 2431 15163 2437
rect 12437 2391 12495 2397
rect 15105 2397 15117 2431
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 5074 2320 5080 2372
rect 5132 2360 5138 2372
rect 12452 2360 12480 2391
rect 5132 2332 12480 2360
rect 5132 2320 5138 2332
rect 2133 2295 2191 2301
rect 2133 2261 2145 2295
rect 2179 2292 2191 2295
rect 6454 2292 6460 2304
rect 2179 2264 6460 2292
rect 2179 2261 2191 2264
rect 2133 2255 2191 2261
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 7006 2252 7012 2304
rect 7064 2292 7070 2304
rect 15120 2292 15148 2391
rect 15212 2360 15240 2468
rect 16022 2456 16028 2468
rect 16080 2456 16086 2508
rect 16942 2456 16948 2508
rect 17000 2496 17006 2508
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17000 2468 17693 2496
rect 17000 2456 17006 2468
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 18230 2496 18236 2508
rect 18191 2468 18236 2496
rect 17681 2459 17739 2465
rect 18230 2456 18236 2468
rect 18288 2456 18294 2508
rect 18966 2496 18972 2508
rect 18927 2468 18972 2496
rect 18966 2456 18972 2468
rect 19024 2456 19030 2508
rect 20254 2496 20260 2508
rect 20215 2468 20260 2496
rect 20254 2456 20260 2468
rect 20312 2456 20318 2508
rect 21174 2496 21180 2508
rect 21135 2468 21180 2496
rect 21174 2456 21180 2468
rect 21232 2456 21238 2508
rect 21450 2496 21456 2508
rect 21411 2468 21456 2496
rect 21450 2456 21456 2468
rect 21508 2456 21514 2508
rect 22186 2456 22192 2508
rect 22244 2496 22250 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22244 2468 23029 2496
rect 22244 2456 22250 2468
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 23017 2459 23075 2465
rect 24397 2499 24455 2505
rect 24397 2465 24409 2499
rect 24443 2496 24455 2499
rect 25130 2496 25136 2508
rect 24443 2468 25136 2496
rect 24443 2465 24455 2468
rect 24397 2459 24455 2465
rect 25130 2456 25136 2468
rect 25188 2456 25194 2508
rect 26050 2496 26056 2508
rect 26011 2468 26056 2496
rect 26050 2456 26056 2468
rect 26108 2456 26114 2508
rect 27062 2496 27068 2508
rect 27023 2468 27068 2496
rect 27062 2456 27068 2468
rect 27120 2456 27126 2508
rect 28074 2456 28080 2508
rect 28132 2496 28138 2508
rect 28261 2499 28319 2505
rect 28261 2496 28273 2499
rect 28132 2468 28273 2496
rect 28132 2456 28138 2468
rect 28261 2465 28273 2468
rect 28307 2465 28319 2499
rect 28261 2459 28319 2465
rect 29549 2499 29607 2505
rect 29549 2465 29561 2499
rect 29595 2496 29607 2499
rect 30006 2496 30012 2508
rect 29595 2468 30012 2496
rect 29595 2465 29607 2468
rect 29549 2459 29607 2465
rect 30006 2456 30012 2468
rect 30064 2456 30070 2508
rect 30926 2456 30932 2508
rect 30984 2496 30990 2508
rect 31021 2499 31079 2505
rect 31021 2496 31033 2499
rect 30984 2468 31033 2496
rect 30984 2456 30990 2468
rect 31021 2465 31033 2468
rect 31067 2465 31079 2499
rect 31021 2459 31079 2465
rect 32950 2456 32956 2508
rect 33008 2496 33014 2508
rect 33689 2499 33747 2505
rect 33689 2496 33701 2499
rect 33008 2468 33701 2496
rect 33008 2456 33014 2468
rect 33689 2465 33701 2468
rect 33735 2465 33747 2499
rect 33689 2459 33747 2465
rect 33870 2456 33876 2508
rect 33928 2496 33934 2508
rect 34517 2499 34575 2505
rect 34517 2496 34529 2499
rect 33928 2468 34529 2496
rect 33928 2456 33934 2468
rect 34517 2465 34529 2468
rect 34563 2465 34575 2499
rect 34517 2459 34575 2465
rect 35894 2456 35900 2508
rect 35952 2496 35958 2508
rect 36357 2499 36415 2505
rect 36357 2496 36369 2499
rect 35952 2468 36369 2496
rect 35952 2456 35958 2468
rect 36357 2465 36369 2468
rect 36403 2465 36415 2499
rect 37458 2496 37464 2508
rect 37419 2468 37464 2496
rect 36357 2459 36415 2465
rect 37458 2456 37464 2468
rect 37516 2456 37522 2508
rect 20441 2431 20499 2437
rect 20441 2397 20453 2431
rect 20487 2397 20499 2431
rect 29730 2428 29736 2440
rect 29691 2400 29736 2428
rect 20441 2391 20499 2397
rect 20456 2360 20484 2391
rect 29730 2388 29736 2400
rect 29788 2388 29794 2440
rect 33962 2388 33968 2440
rect 34020 2428 34026 2440
rect 35621 2431 35679 2437
rect 35621 2428 35633 2431
rect 34020 2400 35633 2428
rect 34020 2388 34026 2400
rect 35621 2397 35633 2400
rect 35667 2397 35679 2431
rect 35621 2391 35679 2397
rect 15212 2332 20484 2360
rect 27249 2363 27307 2369
rect 27249 2329 27261 2363
rect 27295 2360 27307 2363
rect 28166 2360 28172 2372
rect 27295 2332 28172 2360
rect 27295 2329 27307 2332
rect 27249 2323 27307 2329
rect 28166 2320 28172 2332
rect 28224 2320 28230 2372
rect 32677 2363 32735 2369
rect 32677 2329 32689 2363
rect 32723 2360 32735 2363
rect 35526 2360 35532 2372
rect 32723 2332 35532 2360
rect 32723 2329 32735 2332
rect 32677 2323 32735 2329
rect 35526 2320 35532 2332
rect 35584 2320 35590 2372
rect 7064 2264 15148 2292
rect 19245 2295 19303 2301
rect 7064 2252 7070 2264
rect 19245 2261 19257 2295
rect 19291 2292 19303 2295
rect 27338 2292 27344 2304
rect 19291 2264 27344 2292
rect 19291 2261 19303 2264
rect 19245 2255 19303 2261
rect 27338 2252 27344 2264
rect 27396 2252 27402 2304
rect 31110 2292 31116 2304
rect 31071 2264 31116 2292
rect 31110 2252 31116 2264
rect 31168 2252 31174 2304
rect 34701 2295 34759 2301
rect 34701 2261 34713 2295
rect 34747 2292 34759 2295
rect 36998 2292 37004 2304
rect 34747 2264 37004 2292
rect 34747 2261 34759 2264
rect 34701 2255 34759 2261
rect 36998 2252 37004 2264
rect 37056 2252 37062 2304
rect 1104 2202 38824 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 38824 2202
rect 1104 2128 38824 2150
rect 4246 1980 4252 2032
rect 4304 2020 4310 2032
rect 4706 2020 4712 2032
rect 4304 1992 4712 2020
rect 4304 1980 4310 1992
rect 4706 1980 4712 1992
rect 4764 1980 4770 2032
rect 15470 1980 15476 2032
rect 15528 2020 15534 2032
rect 31110 2020 31116 2032
rect 15528 1992 31116 2020
rect 15528 1980 15534 1992
rect 31110 1980 31116 1992
rect 31168 1980 31174 2032
rect 14826 1912 14832 1964
rect 14884 1952 14890 1964
rect 29730 1952 29736 1964
rect 14884 1924 29736 1952
rect 14884 1912 14890 1924
rect 29730 1912 29736 1924
rect 29788 1912 29794 1964
rect 28994 1504 29000 1556
rect 29052 1544 29058 1556
rect 29546 1544 29552 1556
rect 29052 1516 29552 1544
rect 29052 1504 29058 1516
rect 29546 1504 29552 1516
rect 29604 1504 29610 1556
<< via1 >>
rect 4712 118192 4764 118244
rect 34796 118192 34848 118244
rect 34796 117988 34848 118040
rect 4712 117920 4764 117972
rect 25044 117648 25096 117700
rect 29276 117648 29328 117700
rect 34704 117648 34756 117700
rect 34980 117648 35032 117700
rect 24400 117580 24452 117632
rect 28816 117580 28868 117632
rect 4246 117478 4298 117530
rect 4310 117478 4362 117530
rect 4374 117478 4426 117530
rect 4438 117478 4490 117530
rect 34966 117478 35018 117530
rect 35030 117478 35082 117530
rect 35094 117478 35146 117530
rect 35158 117478 35210 117530
rect 296 117376 348 117428
rect 2964 117376 3016 117428
rect 1216 117308 1268 117360
rect 112 117240 164 117292
rect 756 117172 808 117224
rect 6184 117240 6236 117292
rect 11152 117376 11204 117428
rect 17408 117376 17460 117428
rect 17960 117376 18012 117428
rect 18144 117376 18196 117428
rect 16304 117308 16356 117360
rect 16488 117308 16540 117360
rect 16764 117308 16816 117360
rect 20904 117376 20956 117428
rect 9128 117240 9180 117292
rect 10508 117240 10560 117292
rect 11888 117240 11940 117292
rect 13360 117240 13412 117292
rect 17592 117240 17644 117292
rect 19524 117308 19576 117360
rect 22928 117376 22980 117428
rect 27344 117376 27396 117428
rect 22284 117308 22336 117360
rect 1860 117147 1912 117156
rect 1860 117113 1869 117147
rect 1869 117113 1903 117147
rect 1903 117113 1912 117147
rect 1860 117104 1912 117113
rect 4068 117104 4120 117156
rect 1032 117036 1084 117088
rect 5448 117172 5500 117224
rect 9772 117172 9824 117224
rect 13912 117172 13964 117224
rect 17316 117172 17368 117224
rect 4528 117104 4580 117156
rect 6828 117104 6880 117156
rect 7564 117104 7616 117156
rect 7748 117147 7800 117156
rect 7748 117113 7757 117147
rect 7757 117113 7791 117147
rect 7791 117113 7800 117147
rect 7748 117104 7800 117113
rect 9680 117147 9732 117156
rect 9680 117113 9689 117147
rect 9689 117113 9723 117147
rect 9723 117113 9732 117147
rect 9680 117104 9732 117113
rect 10416 117147 10468 117156
rect 10416 117113 10425 117147
rect 10425 117113 10459 117147
rect 10459 117113 10468 117147
rect 10416 117104 10468 117113
rect 11152 117147 11204 117156
rect 11152 117113 11161 117147
rect 11161 117113 11195 117147
rect 11195 117113 11204 117147
rect 11152 117104 11204 117113
rect 11612 117104 11664 117156
rect 13084 117147 13136 117156
rect 13084 117113 13093 117147
rect 13093 117113 13127 117147
rect 13127 117113 13136 117147
rect 13084 117104 13136 117113
rect 13820 117147 13872 117156
rect 13820 117113 13829 117147
rect 13829 117113 13863 117147
rect 13863 117113 13872 117147
rect 13820 117104 13872 117113
rect 14004 117104 14056 117156
rect 15200 117104 15252 117156
rect 16212 117104 16264 117156
rect 17684 117147 17736 117156
rect 17684 117113 17693 117147
rect 17693 117113 17727 117147
rect 17727 117113 17736 117147
rect 17684 117104 17736 117113
rect 19156 117147 19208 117156
rect 19156 117113 19165 117147
rect 19165 117113 19199 117147
rect 19199 117113 19208 117147
rect 19156 117104 19208 117113
rect 19340 117104 19392 117156
rect 20536 117104 20588 117156
rect 21272 117104 21324 117156
rect 26424 117308 26476 117360
rect 28908 117308 28960 117360
rect 27160 117240 27212 117292
rect 34796 117376 34848 117428
rect 22928 117172 22980 117224
rect 27712 117172 27764 117224
rect 35440 117172 35492 117224
rect 37096 117172 37148 117224
rect 23020 117147 23072 117156
rect 7380 117036 7432 117088
rect 7840 117036 7892 117088
rect 12532 117036 12584 117088
rect 14648 117036 14700 117088
rect 17040 117036 17092 117088
rect 17960 117036 18012 117088
rect 21916 117079 21968 117088
rect 21916 117045 21925 117079
rect 21925 117045 21959 117079
rect 21959 117045 21968 117079
rect 21916 117036 21968 117045
rect 23020 117113 23029 117147
rect 23029 117113 23063 117147
rect 23063 117113 23072 117147
rect 23020 117104 23072 117113
rect 23296 117104 23348 117156
rect 24492 117147 24544 117156
rect 24492 117113 24501 117147
rect 24501 117113 24535 117147
rect 24535 117113 24544 117147
rect 24492 117104 24544 117113
rect 24676 117104 24728 117156
rect 26424 117147 26476 117156
rect 26424 117113 26433 117147
rect 26433 117113 26467 117147
rect 26467 117113 26476 117147
rect 26424 117104 26476 117113
rect 27160 117147 27212 117156
rect 27160 117113 27169 117147
rect 27169 117113 27203 117147
rect 27203 117113 27212 117147
rect 27160 117104 27212 117113
rect 28356 117147 28408 117156
rect 28356 117113 28365 117147
rect 28365 117113 28399 117147
rect 28399 117113 28408 117147
rect 28356 117104 28408 117113
rect 28632 117104 28684 117156
rect 29828 117147 29880 117156
rect 29828 117113 29837 117147
rect 29837 117113 29871 117147
rect 29871 117113 29880 117147
rect 29828 117104 29880 117113
rect 30012 117104 30064 117156
rect 31392 117104 31444 117156
rect 33324 117104 33376 117156
rect 34152 117104 34204 117156
rect 34612 117104 34664 117156
rect 23204 117036 23256 117088
rect 28172 117036 28224 117088
rect 28816 117036 28868 117088
rect 29276 117036 29328 117088
rect 30932 117036 30984 117088
rect 31208 117036 31260 117088
rect 33048 117036 33100 117088
rect 38568 117104 38620 117156
rect 36452 117079 36504 117088
rect 36452 117045 36461 117079
rect 36461 117045 36495 117079
rect 36495 117045 36504 117079
rect 36452 117036 36504 117045
rect 36544 117036 36596 117088
rect 37740 117036 37792 117088
rect 19606 116934 19658 116986
rect 19670 116934 19722 116986
rect 19734 116934 19786 116986
rect 19798 116934 19850 116986
rect 1676 116832 1728 116884
rect 4068 116832 4120 116884
rect 2136 116764 2188 116816
rect 4620 116764 4672 116816
rect 4896 116832 4948 116884
rect 6276 116832 6328 116884
rect 7104 116832 7156 116884
rect 8392 116832 8444 116884
rect 9312 116832 9364 116884
rect 10048 116832 10100 116884
rect 11428 116832 11480 116884
rect 12808 116832 12860 116884
rect 14188 116832 14240 116884
rect 15568 116832 15620 116884
rect 16948 116832 17000 116884
rect 17776 116832 17828 116884
rect 18328 116832 18380 116884
rect 19064 116832 19116 116884
rect 20444 116832 20496 116884
rect 21824 116832 21876 116884
rect 23112 116832 23164 116884
rect 24584 116832 24636 116884
rect 25320 116832 25372 116884
rect 25964 116832 26016 116884
rect 27804 116832 27856 116884
rect 28080 116832 28132 116884
rect 28908 116832 28960 116884
rect 31208 116832 31260 116884
rect 31760 116832 31812 116884
rect 32312 116832 32364 116884
rect 36544 116832 36596 116884
rect 36636 116832 36688 116884
rect 6000 116764 6052 116816
rect 12072 116764 12124 116816
rect 13452 116764 13504 116816
rect 19892 116764 19944 116816
rect 3240 116696 3292 116748
rect 3884 116696 3936 116748
rect 5080 116739 5132 116748
rect 5080 116705 5089 116739
rect 5089 116705 5123 116739
rect 5123 116705 5132 116739
rect 5080 116696 5132 116705
rect 6920 116739 6972 116748
rect 6920 116705 6929 116739
rect 6929 116705 6963 116739
rect 6963 116705 6972 116739
rect 6920 116696 6972 116705
rect 7104 116696 7156 116748
rect 8392 116739 8444 116748
rect 8392 116705 8401 116739
rect 8401 116705 8435 116739
rect 8435 116705 8444 116739
rect 8392 116696 8444 116705
rect 9128 116739 9180 116748
rect 9128 116705 9137 116739
rect 9137 116705 9171 116739
rect 9171 116705 9180 116739
rect 9128 116696 9180 116705
rect 9864 116739 9916 116748
rect 9864 116705 9873 116739
rect 9873 116705 9907 116739
rect 9907 116705 9916 116739
rect 9864 116696 9916 116705
rect 10600 116739 10652 116748
rect 10600 116705 10609 116739
rect 10609 116705 10643 116739
rect 10643 116705 10652 116739
rect 10600 116696 10652 116705
rect 12164 116739 12216 116748
rect 12164 116705 12173 116739
rect 12173 116705 12207 116739
rect 12207 116705 12216 116739
rect 12164 116696 12216 116705
rect 12900 116739 12952 116748
rect 12900 116705 12909 116739
rect 12909 116705 12943 116739
rect 12943 116705 12952 116739
rect 12900 116696 12952 116705
rect 12992 116696 13044 116748
rect 14372 116739 14424 116748
rect 14372 116705 14381 116739
rect 14381 116705 14415 116739
rect 14415 116705 14424 116739
rect 14372 116696 14424 116705
rect 15108 116739 15160 116748
rect 15108 116705 15117 116739
rect 15117 116705 15151 116739
rect 15151 116705 15160 116739
rect 15108 116696 15160 116705
rect 15844 116739 15896 116748
rect 15844 116705 15853 116739
rect 15853 116705 15887 116739
rect 15887 116705 15896 116739
rect 15844 116696 15896 116705
rect 17408 116739 17460 116748
rect 17408 116705 17417 116739
rect 17417 116705 17451 116739
rect 17451 116705 17460 116739
rect 17408 116696 17460 116705
rect 18144 116739 18196 116748
rect 18144 116705 18153 116739
rect 18153 116705 18187 116739
rect 18187 116705 18196 116739
rect 18144 116696 18196 116705
rect 18880 116739 18932 116748
rect 18880 116705 18889 116739
rect 18889 116705 18923 116739
rect 18923 116705 18932 116739
rect 18880 116696 18932 116705
rect 19432 116696 19484 116748
rect 20352 116739 20404 116748
rect 20352 116705 20361 116739
rect 20361 116705 20395 116739
rect 20395 116705 20404 116739
rect 20352 116696 20404 116705
rect 20444 116696 20496 116748
rect 21272 116764 21324 116816
rect 22468 116764 22520 116816
rect 21088 116739 21140 116748
rect 21088 116705 21097 116739
rect 21097 116705 21131 116739
rect 21131 116705 21140 116739
rect 21088 116696 21140 116705
rect 22652 116739 22704 116748
rect 22652 116705 22661 116739
rect 22661 116705 22695 116739
rect 22695 116705 22704 116739
rect 22652 116696 22704 116705
rect 4988 116628 5040 116680
rect 5540 116628 5592 116680
rect 7748 116628 7800 116680
rect 18788 116628 18840 116680
rect 21916 116628 21968 116680
rect 22376 116628 22428 116680
rect 24768 116696 24820 116748
rect 28448 116764 28500 116816
rect 28540 116764 28592 116816
rect 34152 116764 34204 116816
rect 35256 116764 35308 116816
rect 38200 116764 38252 116816
rect 6276 116560 6328 116612
rect 20260 116560 20312 116612
rect 23204 116560 23256 116612
rect 25688 116628 25740 116680
rect 24492 116560 24544 116612
rect 27896 116739 27948 116748
rect 27896 116705 27905 116739
rect 27905 116705 27939 116739
rect 27939 116705 27948 116739
rect 27896 116696 27948 116705
rect 28632 116739 28684 116748
rect 28632 116705 28641 116739
rect 28641 116705 28675 116739
rect 28675 116705 28684 116739
rect 28632 116696 28684 116705
rect 28816 116696 28868 116748
rect 29368 116739 29420 116748
rect 28540 116628 28592 116680
rect 29368 116705 29377 116739
rect 29377 116705 29411 116739
rect 29411 116705 29420 116739
rect 29368 116696 29420 116705
rect 30472 116739 30524 116748
rect 30472 116705 30481 116739
rect 30481 116705 30515 116739
rect 30515 116705 30524 116739
rect 30472 116696 30524 116705
rect 31024 116696 31076 116748
rect 31852 116696 31904 116748
rect 33968 116696 34020 116748
rect 31392 116628 31444 116680
rect 34704 116696 34756 116748
rect 35440 116696 35492 116748
rect 36360 116739 36412 116748
rect 36360 116705 36369 116739
rect 36369 116705 36403 116739
rect 36403 116705 36412 116739
rect 36360 116696 36412 116705
rect 36544 116696 36596 116748
rect 36268 116628 36320 116680
rect 28908 116560 28960 116612
rect 34244 116560 34296 116612
rect 36820 116560 36872 116612
rect 2964 116492 3016 116544
rect 5724 116492 5776 116544
rect 7656 116492 7708 116544
rect 20720 116492 20772 116544
rect 23296 116492 23348 116544
rect 25872 116492 25924 116544
rect 30012 116492 30064 116544
rect 32772 116492 32824 116544
rect 33876 116492 33928 116544
rect 34152 116492 34204 116544
rect 36728 116492 36780 116544
rect 4246 116390 4298 116442
rect 4310 116390 4362 116442
rect 4374 116390 4426 116442
rect 4438 116390 4490 116442
rect 34966 116390 35018 116442
rect 35030 116390 35082 116442
rect 35094 116390 35146 116442
rect 35158 116390 35210 116442
rect 2412 116288 2464 116340
rect 3792 116288 3844 116340
rect 5448 116288 5500 116340
rect 5632 116288 5684 116340
rect 5908 116288 5960 116340
rect 6644 116288 6696 116340
rect 8668 116288 8720 116340
rect 10692 116288 10744 116340
rect 11612 116331 11664 116340
rect 11612 116297 11621 116331
rect 11621 116297 11655 116331
rect 11655 116297 11664 116331
rect 11612 116288 11664 116297
rect 13084 116288 13136 116340
rect 14004 116288 14056 116340
rect 14832 116288 14884 116340
rect 17684 116288 17736 116340
rect 19340 116288 19392 116340
rect 21180 116288 21232 116340
rect 1860 116220 1912 116272
rect 7196 116220 7248 116272
rect 13820 116220 13872 116272
rect 16580 116263 16632 116272
rect 16580 116229 16589 116263
rect 16589 116229 16623 116263
rect 16623 116229 16632 116263
rect 16580 116220 16632 116229
rect 19156 116220 19208 116272
rect 23020 116288 23072 116340
rect 23848 116288 23900 116340
rect 24768 116288 24820 116340
rect 26608 116288 26660 116340
rect 26700 116288 26752 116340
rect 26976 116288 27028 116340
rect 21548 116220 21600 116272
rect 22928 116220 22980 116272
rect 2044 116195 2096 116204
rect 2044 116161 2053 116195
rect 2053 116161 2087 116195
rect 2087 116161 2096 116195
rect 2044 116152 2096 116161
rect 5448 116152 5500 116204
rect 20536 116152 20588 116204
rect 22468 116195 22520 116204
rect 5724 116127 5776 116136
rect 5724 116093 5733 116127
rect 5733 116093 5767 116127
rect 5767 116093 5776 116127
rect 5724 116084 5776 116093
rect 15292 116084 15344 116136
rect 17040 116084 17092 116136
rect 1768 116016 1820 116068
rect 3148 116059 3200 116068
rect 3148 116025 3157 116059
rect 3157 116025 3191 116059
rect 3191 116025 3200 116059
rect 3148 116016 3200 116025
rect 4896 116016 4948 116068
rect 6460 116059 6512 116068
rect 6460 116025 6469 116059
rect 6469 116025 6503 116059
rect 6503 116025 6512 116059
rect 6460 116016 6512 116025
rect 7012 116016 7064 116068
rect 7932 116059 7984 116068
rect 7932 116025 7941 116059
rect 7941 116025 7975 116059
rect 7975 116025 7984 116059
rect 7932 116016 7984 116025
rect 9588 116059 9640 116068
rect 9588 116025 9597 116059
rect 9597 116025 9631 116059
rect 9631 116025 9640 116059
rect 9588 116016 9640 116025
rect 10784 116059 10836 116068
rect 10784 116025 10793 116059
rect 10793 116025 10827 116059
rect 10827 116025 10836 116059
rect 10784 116016 10836 116025
rect 14924 116059 14976 116068
rect 14924 116025 14933 116059
rect 14933 116025 14967 116059
rect 14967 116025 14976 116059
rect 14924 116016 14976 116025
rect 16396 116059 16448 116068
rect 16396 116025 16405 116059
rect 16405 116025 16439 116059
rect 16439 116025 16448 116059
rect 16396 116016 16448 116025
rect 21180 116059 21232 116068
rect 21180 116025 21189 116059
rect 21189 116025 21223 116059
rect 21223 116025 21232 116059
rect 21180 116016 21232 116025
rect 22468 116161 22477 116195
rect 22477 116161 22511 116195
rect 22511 116161 22520 116195
rect 22468 116152 22520 116161
rect 27160 116220 27212 116272
rect 27712 116288 27764 116340
rect 28264 116288 28316 116340
rect 28724 116288 28776 116340
rect 29276 116288 29328 116340
rect 30932 116220 30984 116272
rect 31484 116220 31536 116272
rect 32404 116288 32456 116340
rect 32772 116288 32824 116340
rect 35716 116288 35768 116340
rect 35900 116331 35952 116340
rect 35900 116297 35909 116331
rect 35909 116297 35943 116331
rect 35943 116297 35952 116331
rect 35900 116288 35952 116297
rect 29828 116152 29880 116204
rect 31392 116195 31444 116204
rect 31392 116161 31401 116195
rect 31401 116161 31435 116195
rect 31435 116161 31444 116195
rect 31392 116152 31444 116161
rect 31576 116152 31628 116204
rect 32220 116220 32272 116272
rect 32864 116220 32916 116272
rect 33692 116263 33744 116272
rect 33692 116229 33701 116263
rect 33701 116229 33735 116263
rect 33735 116229 33744 116263
rect 33692 116220 33744 116229
rect 34244 116220 34296 116272
rect 36360 116220 36412 116272
rect 38016 116220 38068 116272
rect 32036 116152 32088 116204
rect 32588 116195 32640 116204
rect 32588 116161 32597 116195
rect 32597 116161 32631 116195
rect 32631 116161 32640 116195
rect 32588 116152 32640 116161
rect 33508 116152 33560 116204
rect 33784 116195 33836 116204
rect 33784 116161 33793 116195
rect 33793 116161 33827 116195
rect 33827 116161 33836 116195
rect 33784 116152 33836 116161
rect 23480 116084 23532 116136
rect 26700 116016 26752 116068
rect 26976 116084 27028 116136
rect 31668 116084 31720 116136
rect 31760 116084 31812 116136
rect 34520 116084 34572 116136
rect 34888 116084 34940 116136
rect 36084 116084 36136 116136
rect 37556 116127 37608 116136
rect 37556 116093 37565 116127
rect 37565 116093 37599 116127
rect 37599 116093 37608 116127
rect 37556 116084 37608 116093
rect 24676 115948 24728 116000
rect 25872 115991 25924 116000
rect 25872 115957 25881 115991
rect 25881 115957 25915 115991
rect 25915 115957 25924 115991
rect 25872 115948 25924 115957
rect 28724 116016 28776 116068
rect 30932 116016 30984 116068
rect 30288 115948 30340 116000
rect 33232 116016 33284 116068
rect 35808 116059 35860 116068
rect 31208 115948 31260 116000
rect 32772 115948 32824 116000
rect 33048 115948 33100 116000
rect 34336 115948 34388 116000
rect 35808 116025 35817 116059
rect 35817 116025 35851 116059
rect 35851 116025 35860 116059
rect 35808 116016 35860 116025
rect 37004 116016 37056 116068
rect 19606 115846 19658 115898
rect 19670 115846 19722 115898
rect 19734 115846 19786 115898
rect 19798 115846 19850 115898
rect 572 115744 624 115796
rect 2964 115744 3016 115796
rect 3056 115744 3108 115796
rect 3516 115744 3568 115796
rect 4804 115676 4856 115728
rect 5172 115744 5224 115796
rect 7840 115744 7892 115796
rect 8024 115744 8076 115796
rect 9128 115744 9180 115796
rect 23480 115744 23532 115796
rect 24768 115744 24820 115796
rect 8392 115676 8444 115728
rect 21364 115676 21416 115728
rect 21916 115676 21968 115728
rect 4068 115608 4120 115660
rect 4620 115608 4672 115660
rect 5264 115651 5316 115660
rect 5264 115617 5273 115651
rect 5273 115617 5307 115651
rect 5307 115617 5316 115651
rect 5264 115608 5316 115617
rect 8300 115608 8352 115660
rect 9680 115608 9732 115660
rect 10416 115608 10468 115660
rect 11152 115608 11204 115660
rect 12164 115608 12216 115660
rect 12900 115651 12952 115660
rect 12900 115617 12909 115651
rect 12909 115617 12943 115651
rect 12943 115617 12952 115651
rect 12900 115608 12952 115617
rect 15108 115608 15160 115660
rect 17316 115608 17368 115660
rect 17408 115608 17460 115660
rect 18144 115651 18196 115660
rect 18144 115617 18153 115651
rect 18153 115617 18187 115651
rect 18187 115617 18196 115651
rect 18144 115608 18196 115617
rect 19432 115651 19484 115660
rect 19432 115617 19441 115651
rect 19441 115617 19475 115651
rect 19475 115617 19484 115651
rect 19432 115608 19484 115617
rect 20720 115608 20772 115660
rect 21180 115608 21232 115660
rect 3240 115540 3292 115592
rect 4436 115540 4488 115592
rect 4804 115540 4856 115592
rect 5172 115540 5224 115592
rect 8484 115540 8536 115592
rect 15200 115540 15252 115592
rect 16120 115540 16172 115592
rect 17592 115540 17644 115592
rect 20444 115540 20496 115592
rect 22376 115540 22428 115592
rect 1492 115472 1544 115524
rect 6184 115472 6236 115524
rect 16212 115472 16264 115524
rect 17776 115472 17828 115524
rect 1952 115447 2004 115456
rect 1952 115413 1961 115447
rect 1961 115413 1995 115447
rect 1995 115413 2004 115447
rect 1952 115404 2004 115413
rect 7748 115404 7800 115456
rect 20996 115404 21048 115456
rect 23664 115608 23716 115660
rect 25228 115676 25280 115728
rect 26976 115676 27028 115728
rect 27068 115676 27120 115728
rect 29552 115744 29604 115796
rect 30288 115744 30340 115796
rect 35348 115744 35400 115796
rect 35716 115744 35768 115796
rect 38660 115744 38712 115796
rect 24952 115540 25004 115592
rect 23480 115472 23532 115524
rect 25228 115472 25280 115524
rect 25688 115515 25740 115524
rect 25688 115481 25697 115515
rect 25697 115481 25731 115515
rect 25731 115481 25740 115515
rect 25688 115472 25740 115481
rect 27712 115540 27764 115592
rect 27896 115608 27948 115660
rect 28080 115608 28132 115660
rect 28816 115608 28868 115660
rect 29460 115676 29512 115728
rect 34520 115676 34572 115728
rect 28172 115472 28224 115524
rect 29552 115540 29604 115592
rect 29184 115472 29236 115524
rect 24216 115404 24268 115456
rect 30932 115608 30984 115660
rect 31760 115608 31812 115660
rect 33600 115608 33652 115660
rect 34796 115540 34848 115592
rect 31576 115404 31628 115456
rect 33324 115404 33376 115456
rect 36176 115676 36228 115728
rect 36360 115676 36412 115728
rect 39580 115676 39632 115728
rect 35716 115651 35768 115660
rect 35716 115617 35725 115651
rect 35725 115617 35759 115651
rect 35759 115617 35768 115651
rect 35716 115608 35768 115617
rect 35992 115608 36044 115660
rect 36820 115608 36872 115660
rect 37280 115540 37332 115592
rect 36360 115472 36412 115524
rect 37372 115515 37424 115524
rect 37372 115481 37381 115515
rect 37381 115481 37415 115515
rect 37415 115481 37424 115515
rect 37372 115472 37424 115481
rect 35256 115404 35308 115456
rect 36544 115447 36596 115456
rect 36544 115413 36553 115447
rect 36553 115413 36587 115447
rect 36587 115413 36596 115447
rect 36544 115404 36596 115413
rect 4246 115302 4298 115354
rect 4310 115302 4362 115354
rect 4374 115302 4426 115354
rect 4438 115302 4490 115354
rect 34966 115302 35018 115354
rect 35030 115302 35082 115354
rect 35094 115302 35146 115354
rect 35158 115302 35210 115354
rect 1400 115200 1452 115252
rect 5080 115200 5132 115252
rect 6920 115200 6972 115252
rect 7104 115200 7156 115252
rect 7932 115200 7984 115252
rect 8300 115243 8352 115252
rect 8300 115209 8309 115243
rect 8309 115209 8343 115243
rect 8343 115209 8352 115243
rect 8300 115200 8352 115209
rect 9864 115200 9916 115252
rect 10600 115200 10652 115252
rect 10784 115200 10836 115252
rect 12992 115200 13044 115252
rect 14372 115200 14424 115252
rect 14924 115243 14976 115252
rect 14924 115209 14933 115243
rect 14933 115209 14967 115243
rect 14967 115209 14976 115243
rect 14924 115200 14976 115209
rect 15844 115200 15896 115252
rect 16396 115200 16448 115252
rect 18880 115200 18932 115252
rect 20352 115200 20404 115252
rect 21088 115200 21140 115252
rect 25412 115200 25464 115252
rect 28632 115200 28684 115252
rect 28908 115200 28960 115252
rect 29644 115200 29696 115252
rect 31392 115200 31444 115252
rect 31484 115200 31536 115252
rect 35348 115200 35400 115252
rect 2780 115175 2832 115184
rect 2780 115141 2789 115175
rect 2789 115141 2823 115175
rect 2823 115141 2832 115175
rect 2780 115132 2832 115141
rect 5540 115132 5592 115184
rect 21456 115132 21508 115184
rect 24032 115132 24084 115184
rect 24216 115132 24268 115184
rect 30012 115132 30064 115184
rect 4988 115064 5040 115116
rect 6920 115064 6972 115116
rect 8760 115064 8812 115116
rect 15292 115064 15344 115116
rect 21824 115064 21876 115116
rect 8668 114996 8720 115048
rect 10968 114996 11020 115048
rect 16488 114996 16540 115048
rect 17224 114996 17276 115048
rect 18604 114996 18656 115048
rect 20628 114996 20680 115048
rect 21916 115039 21968 115048
rect 21916 115005 21925 115039
rect 21925 115005 21959 115039
rect 21959 115005 21968 115039
rect 21916 114996 21968 115005
rect 22468 114996 22520 115048
rect 23020 114996 23072 115048
rect 24400 115064 24452 115116
rect 27068 115064 27120 115116
rect 31576 115064 31628 115116
rect 26424 115039 26476 115048
rect 7656 114928 7708 114980
rect 13360 114928 13412 114980
rect 5172 114860 5224 114912
rect 5540 114860 5592 114912
rect 10692 114860 10744 114912
rect 22836 114928 22888 114980
rect 26424 115005 26433 115039
rect 26433 115005 26467 115039
rect 26467 115005 26476 115039
rect 26424 114996 26476 115005
rect 28816 114996 28868 115048
rect 29184 114996 29236 115048
rect 29368 115039 29420 115048
rect 29368 115005 29377 115039
rect 29377 115005 29411 115039
rect 29411 115005 29420 115039
rect 29368 114996 29420 115005
rect 32128 115132 32180 115184
rect 31944 114996 31996 115048
rect 21088 114860 21140 114912
rect 23480 114903 23532 114912
rect 23480 114869 23489 114903
rect 23489 114869 23523 114903
rect 23523 114869 23532 114903
rect 23480 114860 23532 114869
rect 23572 114860 23624 114912
rect 24308 114860 24360 114912
rect 24400 114860 24452 114912
rect 26700 114860 26752 114912
rect 30380 114928 30432 114980
rect 30656 114860 30708 114912
rect 31392 114860 31444 114912
rect 31484 114860 31536 114912
rect 34152 115064 34204 115116
rect 35532 115132 35584 115184
rect 39856 115064 39908 115116
rect 32404 114996 32456 115048
rect 34796 114996 34848 115048
rect 36084 114996 36136 115048
rect 34244 114928 34296 114980
rect 34520 114928 34572 114980
rect 35532 114928 35584 114980
rect 37924 114971 37976 114980
rect 37924 114937 37933 114971
rect 37933 114937 37967 114971
rect 37967 114937 37976 114971
rect 37924 114928 37976 114937
rect 35256 114860 35308 114912
rect 37740 114860 37792 114912
rect 19606 114758 19658 114810
rect 19670 114758 19722 114810
rect 19734 114758 19786 114810
rect 19798 114758 19850 114810
rect 3424 114699 3476 114708
rect 3424 114665 3433 114699
rect 3433 114665 3467 114699
rect 3467 114665 3476 114699
rect 3424 114656 3476 114665
rect 6828 114656 6880 114708
rect 8300 114656 8352 114708
rect 13360 114699 13412 114708
rect 13360 114665 13369 114699
rect 13369 114665 13403 114699
rect 13403 114665 13412 114699
rect 13360 114656 13412 114665
rect 15292 114699 15344 114708
rect 7196 114588 7248 114640
rect 15292 114665 15301 114699
rect 15301 114665 15335 114699
rect 15335 114665 15344 114699
rect 15292 114656 15344 114665
rect 17776 114656 17828 114708
rect 21824 114656 21876 114708
rect 23572 114656 23624 114708
rect 24124 114656 24176 114708
rect 2596 114563 2648 114572
rect 2596 114529 2605 114563
rect 2605 114529 2639 114563
rect 2639 114529 2648 114563
rect 2596 114520 2648 114529
rect 3700 114520 3752 114572
rect 5264 114520 5316 114572
rect 6276 114520 6328 114572
rect 7380 114520 7432 114572
rect 7656 114563 7708 114572
rect 2044 114495 2096 114504
rect 2044 114461 2053 114495
rect 2053 114461 2087 114495
rect 2087 114461 2096 114495
rect 2044 114452 2096 114461
rect 2872 114452 2924 114504
rect 4068 114452 4120 114504
rect 4896 114452 4948 114504
rect 7012 114495 7064 114504
rect 7012 114461 7021 114495
rect 7021 114461 7055 114495
rect 7055 114461 7064 114495
rect 7012 114452 7064 114461
rect 7656 114529 7665 114563
rect 7665 114529 7699 114563
rect 7699 114529 7708 114563
rect 7656 114520 7708 114529
rect 8760 114563 8812 114572
rect 8760 114529 8769 114563
rect 8769 114529 8803 114563
rect 8803 114529 8812 114563
rect 8760 114520 8812 114529
rect 8852 114520 8904 114572
rect 9496 114520 9548 114572
rect 10232 114520 10284 114572
rect 11704 114520 11756 114572
rect 12348 114520 12400 114572
rect 13176 114520 13228 114572
rect 13728 114520 13780 114572
rect 14464 114520 14516 114572
rect 15016 114520 15068 114572
rect 15752 114520 15804 114572
rect 17868 114520 17920 114572
rect 19248 114520 19300 114572
rect 19984 114520 20036 114572
rect 10692 114427 10744 114436
rect 10692 114393 10701 114427
rect 10701 114393 10735 114427
rect 10735 114393 10744 114427
rect 10692 114384 10744 114393
rect 20996 114520 21048 114572
rect 21088 114520 21140 114572
rect 22468 114520 22520 114572
rect 22836 114563 22888 114572
rect 22836 114529 22845 114563
rect 22845 114529 22879 114563
rect 22879 114529 22888 114563
rect 22836 114520 22888 114529
rect 22928 114520 22980 114572
rect 24400 114520 24452 114572
rect 25504 114656 25556 114708
rect 24860 114588 24912 114640
rect 26608 114656 26660 114708
rect 28448 114699 28500 114708
rect 28448 114665 28457 114699
rect 28457 114665 28491 114699
rect 28491 114665 28500 114699
rect 28448 114656 28500 114665
rect 28540 114656 28592 114708
rect 29920 114656 29972 114708
rect 30288 114656 30340 114708
rect 31668 114656 31720 114708
rect 30012 114563 30064 114572
rect 30012 114529 30021 114563
rect 30021 114529 30055 114563
rect 30055 114529 30064 114563
rect 30012 114520 30064 114529
rect 30104 114520 30156 114572
rect 33692 114588 33744 114640
rect 31484 114563 31536 114572
rect 30656 114452 30708 114504
rect 30748 114384 30800 114436
rect 31484 114529 31493 114563
rect 31493 114529 31527 114563
rect 31527 114529 31536 114563
rect 31484 114520 31536 114529
rect 32680 114520 32732 114572
rect 33048 114520 33100 114572
rect 33324 114520 33376 114572
rect 35900 114656 35952 114708
rect 36268 114699 36320 114708
rect 36268 114665 36277 114699
rect 36277 114665 36311 114699
rect 36311 114665 36320 114699
rect 36268 114656 36320 114665
rect 34796 114563 34848 114572
rect 34796 114529 34805 114563
rect 34805 114529 34839 114563
rect 34839 114529 34848 114563
rect 34796 114520 34848 114529
rect 32128 114384 32180 114436
rect 34152 114384 34204 114436
rect 35532 114520 35584 114572
rect 35716 114563 35768 114572
rect 35716 114529 35725 114563
rect 35725 114529 35759 114563
rect 35759 114529 35768 114563
rect 35716 114520 35768 114529
rect 36176 114563 36228 114572
rect 36176 114529 36185 114563
rect 36185 114529 36219 114563
rect 36219 114529 36228 114563
rect 36176 114520 36228 114529
rect 36084 114384 36136 114436
rect 36268 114384 36320 114436
rect 12716 114359 12768 114368
rect 12716 114325 12725 114359
rect 12725 114325 12759 114359
rect 12759 114325 12768 114359
rect 12716 114316 12768 114325
rect 14648 114359 14700 114368
rect 14648 114325 14657 114359
rect 14657 114325 14691 114359
rect 14691 114325 14700 114359
rect 14648 114316 14700 114325
rect 34428 114316 34480 114368
rect 4246 114214 4298 114266
rect 4310 114214 4362 114266
rect 4374 114214 4426 114266
rect 4438 114214 4490 114266
rect 34966 114214 35018 114266
rect 35030 114214 35082 114266
rect 35094 114214 35146 114266
rect 35158 114214 35210 114266
rect 3148 114112 3200 114164
rect 4620 114112 4672 114164
rect 5448 114112 5500 114164
rect 6460 114112 6512 114164
rect 7564 114112 7616 114164
rect 30380 114112 30432 114164
rect 32036 114112 32088 114164
rect 32864 114112 32916 114164
rect 33508 114112 33560 114164
rect 35532 114112 35584 114164
rect 3884 114044 3936 114096
rect 29368 114044 29420 114096
rect 31208 114044 31260 114096
rect 34428 114044 34480 114096
rect 5540 113908 5592 113960
rect 6920 113908 6972 113960
rect 12716 113976 12768 114028
rect 1860 113883 1912 113892
rect 1860 113849 1869 113883
rect 1869 113849 1903 113883
rect 1903 113849 1912 113883
rect 1860 113840 1912 113849
rect 2688 113840 2740 113892
rect 4804 113840 4856 113892
rect 14648 113908 14700 113960
rect 22008 113951 22060 113960
rect 22008 113917 22017 113951
rect 22017 113917 22051 113951
rect 22051 113917 22060 113951
rect 22008 113908 22060 113917
rect 23388 113951 23440 113960
rect 23388 113917 23397 113951
rect 23397 113917 23431 113951
rect 23431 113917 23440 113951
rect 23388 113908 23440 113917
rect 26240 113951 26292 113960
rect 26240 113917 26249 113951
rect 26249 113917 26283 113951
rect 26283 113917 26292 113951
rect 26240 113908 26292 113917
rect 26884 113951 26936 113960
rect 26884 113917 26893 113951
rect 26893 113917 26927 113951
rect 26927 113917 26936 113951
rect 26884 113908 26936 113917
rect 27620 113951 27672 113960
rect 27620 113917 27629 113951
rect 27629 113917 27663 113951
rect 27663 113917 27672 113951
rect 27620 113908 27672 113917
rect 30564 113908 30616 113960
rect 31392 113908 31444 113960
rect 33876 113976 33928 114028
rect 34612 113976 34664 114028
rect 32496 113908 32548 113960
rect 32956 113908 33008 113960
rect 6000 113772 6052 113824
rect 8300 113840 8352 113892
rect 25780 113840 25832 113892
rect 31760 113840 31812 113892
rect 34612 113883 34664 113892
rect 34612 113849 34621 113883
rect 34621 113849 34655 113883
rect 34655 113849 34664 113883
rect 34612 113840 34664 113849
rect 35256 114044 35308 114096
rect 36084 113908 36136 113960
rect 36268 113951 36320 113960
rect 36268 113917 36277 113951
rect 36277 113917 36311 113951
rect 36311 113917 36320 113951
rect 36268 113908 36320 113917
rect 39396 113908 39448 113960
rect 37924 113883 37976 113892
rect 37924 113849 37933 113883
rect 37933 113849 37967 113883
rect 37967 113849 37976 113883
rect 37924 113840 37976 113849
rect 33968 113772 34020 113824
rect 37372 113772 37424 113824
rect 19606 113670 19658 113722
rect 19670 113670 19722 113722
rect 19734 113670 19786 113722
rect 19798 113670 19850 113722
rect 30932 113568 30984 113620
rect 6736 113500 6788 113552
rect 2136 113475 2188 113484
rect 2136 113441 2145 113475
rect 2145 113441 2179 113475
rect 2179 113441 2188 113475
rect 2136 113432 2188 113441
rect 2780 113475 2832 113484
rect 2780 113441 2789 113475
rect 2789 113441 2823 113475
rect 2823 113441 2832 113475
rect 2780 113432 2832 113441
rect 3332 113432 3384 113484
rect 3976 113432 4028 113484
rect 4712 113432 4764 113484
rect 5356 113432 5408 113484
rect 6092 113432 6144 113484
rect 8208 113500 8260 113552
rect 7564 113432 7616 113484
rect 25044 113500 25096 113552
rect 30840 113432 30892 113484
rect 31116 113432 31168 113484
rect 29184 113296 29236 113348
rect 32588 113568 32640 113620
rect 34152 113568 34204 113620
rect 33140 113432 33192 113484
rect 34152 113364 34204 113416
rect 35808 113568 35860 113620
rect 34888 113500 34940 113552
rect 35256 113500 35308 113552
rect 37188 113568 37240 113620
rect 36912 113500 36964 113552
rect 34796 113432 34848 113484
rect 35716 113475 35768 113484
rect 35716 113441 35725 113475
rect 35725 113441 35759 113475
rect 35759 113441 35768 113475
rect 35716 113432 35768 113441
rect 36544 113432 36596 113484
rect 37188 113475 37240 113484
rect 37188 113441 37197 113475
rect 37197 113441 37231 113475
rect 37231 113441 37240 113475
rect 37188 113432 37240 113441
rect 34428 113364 34480 113416
rect 35532 113364 35584 113416
rect 35808 113364 35860 113416
rect 37004 113296 37056 113348
rect 37280 113271 37332 113280
rect 37280 113237 37289 113271
rect 37289 113237 37323 113271
rect 37323 113237 37332 113271
rect 37280 113228 37332 113237
rect 4246 113126 4298 113178
rect 4310 113126 4362 113178
rect 4374 113126 4426 113178
rect 4438 113126 4490 113178
rect 34966 113126 35018 113178
rect 35030 113126 35082 113178
rect 35094 113126 35146 113178
rect 35158 113126 35210 113178
rect 1952 113067 2004 113076
rect 1952 113033 1961 113067
rect 1961 113033 1995 113067
rect 1995 113033 2004 113067
rect 1952 113024 2004 113033
rect 30656 113024 30708 113076
rect 32128 113024 32180 113076
rect 33232 113024 33284 113076
rect 34704 113067 34756 113076
rect 34704 113033 34713 113067
rect 34713 113033 34747 113067
rect 34747 113033 34756 113067
rect 34704 113024 34756 113033
rect 36268 113024 36320 113076
rect 39120 113024 39172 113076
rect 29276 112956 29328 113008
rect 30748 112956 30800 113008
rect 38936 112956 38988 113008
rect 35256 112888 35308 112940
rect 2228 112752 2280 112804
rect 30380 112820 30432 112872
rect 31300 112820 31352 112872
rect 32220 112820 32272 112872
rect 32312 112820 32364 112872
rect 33416 112820 33468 112872
rect 34152 112820 34204 112872
rect 34336 112820 34388 112872
rect 34796 112820 34848 112872
rect 35624 112820 35676 112872
rect 38476 112888 38528 112940
rect 37924 112863 37976 112872
rect 37924 112829 37933 112863
rect 37933 112829 37967 112863
rect 37967 112829 37976 112863
rect 37924 112820 37976 112829
rect 29000 112684 29052 112736
rect 31852 112684 31904 112736
rect 32772 112684 32824 112736
rect 34336 112727 34388 112736
rect 34336 112693 34345 112727
rect 34345 112693 34379 112727
rect 34379 112693 34388 112727
rect 36268 112752 36320 112804
rect 37188 112795 37240 112804
rect 37188 112761 37197 112795
rect 37197 112761 37231 112795
rect 37231 112761 37240 112795
rect 37188 112752 37240 112761
rect 34336 112684 34388 112693
rect 34704 112684 34756 112736
rect 37648 112684 37700 112736
rect 19606 112582 19658 112634
rect 19670 112582 19722 112634
rect 19734 112582 19786 112634
rect 19798 112582 19850 112634
rect 33784 112480 33836 112532
rect 35532 112480 35584 112532
rect 29460 112412 29512 112464
rect 37188 112412 37240 112464
rect 6276 112344 6328 112396
rect 34060 112344 34112 112396
rect 35348 112344 35400 112396
rect 36084 112344 36136 112396
rect 37096 112387 37148 112396
rect 37096 112353 37105 112387
rect 37105 112353 37139 112387
rect 37139 112353 37148 112387
rect 37096 112344 37148 112353
rect 2044 112319 2096 112328
rect 2044 112285 2053 112319
rect 2053 112285 2087 112319
rect 2087 112285 2096 112319
rect 2044 112276 2096 112285
rect 35348 112208 35400 112260
rect 35900 112183 35952 112192
rect 35900 112149 35909 112183
rect 35909 112149 35943 112183
rect 35943 112149 35952 112183
rect 35900 112140 35952 112149
rect 4246 112038 4298 112090
rect 4310 112038 4362 112090
rect 4374 112038 4426 112090
rect 4438 112038 4490 112090
rect 34966 112038 35018 112090
rect 35030 112038 35082 112090
rect 35094 112038 35146 112090
rect 35158 112038 35210 112090
rect 34796 111800 34848 111852
rect 35624 111732 35676 111784
rect 37096 111775 37148 111784
rect 37096 111741 37105 111775
rect 37105 111741 37139 111775
rect 37139 111741 37148 111775
rect 37096 111732 37148 111741
rect 37832 111775 37884 111784
rect 37832 111741 37841 111775
rect 37841 111741 37875 111775
rect 37875 111741 37884 111775
rect 37832 111732 37884 111741
rect 35532 111664 35584 111716
rect 36176 111707 36228 111716
rect 36176 111673 36210 111707
rect 36210 111673 36228 111707
rect 36176 111664 36228 111673
rect 33784 111596 33836 111648
rect 34336 111596 34388 111648
rect 36360 111639 36412 111648
rect 36360 111605 36369 111639
rect 36369 111605 36403 111639
rect 36403 111605 36412 111639
rect 36360 111596 36412 111605
rect 38476 111664 38528 111716
rect 39120 111596 39172 111648
rect 19606 111494 19658 111546
rect 19670 111494 19722 111546
rect 19734 111494 19786 111546
rect 19798 111494 19850 111546
rect 1952 111435 2004 111444
rect 1952 111401 1961 111435
rect 1961 111401 1995 111435
rect 1995 111401 2004 111435
rect 1952 111392 2004 111401
rect 35992 111435 36044 111444
rect 35992 111401 36001 111435
rect 36001 111401 36035 111435
rect 36035 111401 36044 111435
rect 35992 111392 36044 111401
rect 35624 111324 35676 111376
rect 2504 111256 2556 111308
rect 34060 111256 34112 111308
rect 34428 111256 34480 111308
rect 33508 111188 33560 111240
rect 34152 111188 34204 111240
rect 35532 111256 35584 111308
rect 37096 111299 37148 111308
rect 37096 111265 37105 111299
rect 37105 111265 37139 111299
rect 37139 111265 37148 111299
rect 37096 111256 37148 111265
rect 34428 111052 34480 111104
rect 4246 110950 4298 111002
rect 4310 110950 4362 111002
rect 4374 110950 4426 111002
rect 4438 110950 4490 111002
rect 34966 110950 35018 111002
rect 35030 110950 35082 111002
rect 35094 110950 35146 111002
rect 35158 110950 35210 111002
rect 2136 110644 2188 110696
rect 13728 110644 13780 110696
rect 37832 110687 37884 110696
rect 37832 110653 37841 110687
rect 37841 110653 37875 110687
rect 37875 110653 37884 110687
rect 37832 110644 37884 110653
rect 2044 110619 2096 110628
rect 2044 110585 2053 110619
rect 2053 110585 2087 110619
rect 2087 110585 2096 110619
rect 2044 110576 2096 110585
rect 36084 110576 36136 110628
rect 32588 110508 32640 110560
rect 19606 110406 19658 110458
rect 19670 110406 19722 110458
rect 19734 110406 19786 110458
rect 19798 110406 19850 110458
rect 37096 110211 37148 110220
rect 37096 110177 37105 110211
rect 37105 110177 37139 110211
rect 37139 110177 37148 110211
rect 37096 110168 37148 110177
rect 33232 110032 33284 110084
rect 34704 110032 34756 110084
rect 31944 109964 31996 110016
rect 35808 109964 35860 110016
rect 38660 109964 38712 110016
rect 4246 109862 4298 109914
rect 4310 109862 4362 109914
rect 4374 109862 4426 109914
rect 4438 109862 4490 109914
rect 34966 109862 35018 109914
rect 35030 109862 35082 109914
rect 35094 109862 35146 109914
rect 35158 109862 35210 109914
rect 1952 109803 2004 109812
rect 1952 109769 1961 109803
rect 1961 109769 1995 109803
rect 1995 109769 2004 109803
rect 1952 109760 2004 109769
rect 2688 109556 2740 109608
rect 32680 109599 32732 109608
rect 1952 109488 2004 109540
rect 32680 109565 32689 109599
rect 32689 109565 32723 109599
rect 32723 109565 32732 109599
rect 32680 109556 32732 109565
rect 35440 109760 35492 109812
rect 35808 109760 35860 109812
rect 35900 109624 35952 109676
rect 33232 109599 33284 109608
rect 33232 109565 33241 109599
rect 33241 109565 33275 109599
rect 33275 109565 33284 109599
rect 33232 109556 33284 109565
rect 34796 109556 34848 109608
rect 37096 109599 37148 109608
rect 37096 109565 37105 109599
rect 37105 109565 37139 109599
rect 37139 109565 37148 109599
rect 37096 109556 37148 109565
rect 37832 109599 37884 109608
rect 37832 109565 37841 109599
rect 37841 109565 37875 109599
rect 37875 109565 37884 109599
rect 37832 109556 37884 109565
rect 34152 109488 34204 109540
rect 33140 109420 33192 109472
rect 34060 109420 34112 109472
rect 34336 109463 34388 109472
rect 34336 109429 34345 109463
rect 34345 109429 34379 109463
rect 34379 109429 34388 109463
rect 34336 109420 34388 109429
rect 38844 109420 38896 109472
rect 19606 109318 19658 109370
rect 19670 109318 19722 109370
rect 19734 109318 19786 109370
rect 19798 109318 19850 109370
rect 34520 109216 34572 109268
rect 36912 109216 36964 109268
rect 33416 109148 33468 109200
rect 34336 109148 34388 109200
rect 1860 109123 1912 109132
rect 1860 109089 1869 109123
rect 1869 109089 1903 109123
rect 1903 109089 1912 109123
rect 1860 109080 1912 109089
rect 33232 109080 33284 109132
rect 27160 109012 27212 109064
rect 30564 109012 30616 109064
rect 34796 109080 34848 109132
rect 37096 109123 37148 109132
rect 37096 109089 37105 109123
rect 37105 109089 37139 109123
rect 37139 109089 37148 109123
rect 37096 109080 37148 109089
rect 34888 109012 34940 109064
rect 4246 108774 4298 108826
rect 4310 108774 4362 108826
rect 4374 108774 4426 108826
rect 4438 108774 4490 108826
rect 34966 108774 35018 108826
rect 35030 108774 35082 108826
rect 35094 108774 35146 108826
rect 35158 108774 35210 108826
rect 8484 108672 8536 108724
rect 36544 108672 36596 108724
rect 32864 108604 32916 108656
rect 35440 108536 35492 108588
rect 12900 108511 12952 108520
rect 12900 108477 12909 108511
rect 12909 108477 12943 108511
rect 12943 108477 12952 108511
rect 12900 108468 12952 108477
rect 17592 108468 17644 108520
rect 33416 108468 33468 108520
rect 34152 108511 34204 108520
rect 34152 108477 34161 108511
rect 34161 108477 34195 108511
rect 34195 108477 34204 108511
rect 34152 108468 34204 108477
rect 37832 108511 37884 108520
rect 37832 108477 37841 108511
rect 37841 108477 37875 108511
rect 37875 108477 37884 108511
rect 37832 108468 37884 108477
rect 33508 108400 33560 108452
rect 34520 108332 34572 108384
rect 35532 108332 35584 108384
rect 19606 108230 19658 108282
rect 19670 108230 19722 108282
rect 19734 108230 19786 108282
rect 19798 108230 19850 108282
rect 1952 108171 2004 108180
rect 1952 108137 1961 108171
rect 1961 108137 1995 108171
rect 1995 108137 2004 108171
rect 1952 108128 2004 108137
rect 34244 108060 34296 108112
rect 34428 108060 34480 108112
rect 3516 107992 3568 108044
rect 33232 107992 33284 108044
rect 37188 108035 37240 108044
rect 37188 108001 37197 108035
rect 37197 108001 37231 108035
rect 37231 108001 37240 108035
rect 37188 107992 37240 108001
rect 32496 107856 32548 107908
rect 33784 107788 33836 107840
rect 35256 107788 35308 107840
rect 4246 107686 4298 107738
rect 4310 107686 4362 107738
rect 4374 107686 4426 107738
rect 4438 107686 4490 107738
rect 34966 107686 35018 107738
rect 35030 107686 35082 107738
rect 35094 107686 35146 107738
rect 35158 107686 35210 107738
rect 35440 107516 35492 107568
rect 2412 107380 2464 107432
rect 31116 107380 31168 107432
rect 33416 107380 33468 107432
rect 37188 107423 37240 107432
rect 37188 107389 37197 107423
rect 37197 107389 37231 107423
rect 37231 107389 37240 107423
rect 37188 107380 37240 107389
rect 2044 107355 2096 107364
rect 2044 107321 2053 107355
rect 2053 107321 2087 107355
rect 2087 107321 2096 107355
rect 2044 107312 2096 107321
rect 35624 107312 35676 107364
rect 37924 107355 37976 107364
rect 34336 107244 34388 107296
rect 37924 107321 37933 107355
rect 37933 107321 37967 107355
rect 37967 107321 37976 107355
rect 37924 107312 37976 107321
rect 19606 107142 19658 107194
rect 19670 107142 19722 107194
rect 19734 107142 19786 107194
rect 19798 107142 19850 107194
rect 2872 106904 2924 106956
rect 37188 106947 37240 106956
rect 37188 106913 37197 106947
rect 37197 106913 37231 106947
rect 37231 106913 37240 106947
rect 37188 106904 37240 106913
rect 1952 106743 2004 106752
rect 1952 106709 1961 106743
rect 1961 106709 1995 106743
rect 1995 106709 2004 106743
rect 1952 106700 2004 106709
rect 35532 106700 35584 106752
rect 4246 106598 4298 106650
rect 4310 106598 4362 106650
rect 4374 106598 4426 106650
rect 4438 106598 4490 106650
rect 34966 106598 35018 106650
rect 35030 106598 35082 106650
rect 35094 106598 35146 106650
rect 35158 106598 35210 106650
rect 34060 106360 34112 106412
rect 37924 106335 37976 106344
rect 37924 106301 37933 106335
rect 37933 106301 37967 106335
rect 37967 106301 37976 106335
rect 37924 106292 37976 106301
rect 19606 106054 19658 106106
rect 19670 106054 19722 106106
rect 19734 106054 19786 106106
rect 19798 106054 19850 106106
rect 8668 105952 8720 106004
rect 33140 105927 33192 105936
rect 33140 105893 33149 105927
rect 33149 105893 33183 105927
rect 33183 105893 33192 105927
rect 33140 105884 33192 105893
rect 35256 105927 35308 105936
rect 35256 105893 35265 105927
rect 35265 105893 35299 105927
rect 35299 105893 35308 105927
rect 35256 105884 35308 105893
rect 1400 105859 1452 105868
rect 1400 105825 1409 105859
rect 1409 105825 1443 105859
rect 1443 105825 1452 105859
rect 1400 105816 1452 105825
rect 9956 105859 10008 105868
rect 9956 105825 9965 105859
rect 9965 105825 9999 105859
rect 9999 105825 10008 105859
rect 9956 105816 10008 105825
rect 34520 105816 34572 105868
rect 35440 105816 35492 105868
rect 37188 105859 37240 105868
rect 37188 105825 37197 105859
rect 37197 105825 37231 105859
rect 37231 105825 37240 105859
rect 37188 105816 37240 105825
rect 1584 105791 1636 105800
rect 1584 105757 1593 105791
rect 1593 105757 1627 105791
rect 1627 105757 1636 105791
rect 1584 105748 1636 105757
rect 27068 105748 27120 105800
rect 33508 105748 33560 105800
rect 34704 105791 34756 105800
rect 34704 105757 34713 105791
rect 34713 105757 34747 105791
rect 34747 105757 34756 105791
rect 34704 105748 34756 105757
rect 27620 105612 27672 105664
rect 35440 105612 35492 105664
rect 4246 105510 4298 105562
rect 4310 105510 4362 105562
rect 4374 105510 4426 105562
rect 4438 105510 4490 105562
rect 34966 105510 35018 105562
rect 35030 105510 35082 105562
rect 35094 105510 35146 105562
rect 35158 105510 35210 105562
rect 37924 105247 37976 105256
rect 37924 105213 37933 105247
rect 37933 105213 37967 105247
rect 37967 105213 37976 105247
rect 37924 105204 37976 105213
rect 2320 105136 2372 105188
rect 1952 105111 2004 105120
rect 1952 105077 1961 105111
rect 1961 105077 1995 105111
rect 1995 105077 2004 105111
rect 1952 105068 2004 105077
rect 33968 105068 34020 105120
rect 19606 104966 19658 105018
rect 19670 104966 19722 105018
rect 19734 104966 19786 105018
rect 19798 104966 19850 105018
rect 37188 104839 37240 104848
rect 37188 104805 37197 104839
rect 37197 104805 37231 104839
rect 37231 104805 37240 104839
rect 37188 104796 37240 104805
rect 35992 104524 36044 104576
rect 4246 104422 4298 104474
rect 4310 104422 4362 104474
rect 4374 104422 4426 104474
rect 4438 104422 4490 104474
rect 34966 104422 35018 104474
rect 35030 104422 35082 104474
rect 35094 104422 35146 104474
rect 35158 104422 35210 104474
rect 34796 104320 34848 104372
rect 1492 104159 1544 104168
rect 1492 104125 1501 104159
rect 1501 104125 1535 104159
rect 1535 104125 1544 104159
rect 1492 104116 1544 104125
rect 30656 104116 30708 104168
rect 37188 104159 37240 104168
rect 37188 104125 37197 104159
rect 37197 104125 37231 104159
rect 37231 104125 37240 104159
rect 37188 104116 37240 104125
rect 3608 104048 3660 104100
rect 31208 104048 31260 104100
rect 37924 104091 37976 104100
rect 36176 103980 36228 104032
rect 37924 104057 37933 104091
rect 37933 104057 37967 104091
rect 37967 104057 37976 104091
rect 37924 104048 37976 104057
rect 19606 103878 19658 103930
rect 19670 103878 19722 103930
rect 19734 103878 19786 103930
rect 19798 103878 19850 103930
rect 33232 103776 33284 103828
rect 33876 103708 33928 103760
rect 1676 103640 1728 103692
rect 30012 103683 30064 103692
rect 30012 103649 30021 103683
rect 30021 103649 30055 103683
rect 30055 103649 30064 103683
rect 30012 103640 30064 103649
rect 37188 103683 37240 103692
rect 37188 103649 37197 103683
rect 37197 103649 37231 103683
rect 37231 103649 37240 103683
rect 37188 103640 37240 103649
rect 2044 103547 2096 103556
rect 2044 103513 2053 103547
rect 2053 103513 2087 103547
rect 2087 103513 2096 103547
rect 2044 103504 2096 103513
rect 38200 103504 38252 103556
rect 4246 103334 4298 103386
rect 4310 103334 4362 103386
rect 4374 103334 4426 103386
rect 4438 103334 4490 103386
rect 34966 103334 35018 103386
rect 35030 103334 35082 103386
rect 35094 103334 35146 103386
rect 35158 103334 35210 103386
rect 7104 103275 7156 103284
rect 7104 103241 7113 103275
rect 7113 103241 7147 103275
rect 7147 103241 7156 103275
rect 7104 103232 7156 103241
rect 34152 103232 34204 103284
rect 36820 103096 36872 103148
rect 7012 103028 7064 103080
rect 30656 103028 30708 103080
rect 11428 102960 11480 103012
rect 37924 103003 37976 103012
rect 37924 102969 37933 103003
rect 37933 102969 37967 103003
rect 37967 102969 37976 103003
rect 37924 102960 37976 102969
rect 31576 102892 31628 102944
rect 19606 102790 19658 102842
rect 19670 102790 19722 102842
rect 19734 102790 19786 102842
rect 19798 102790 19850 102842
rect 7748 102731 7800 102740
rect 7748 102697 7757 102731
rect 7757 102697 7791 102731
rect 7791 102697 7800 102731
rect 7748 102688 7800 102697
rect 1492 102552 1544 102604
rect 2044 102595 2096 102604
rect 2044 102561 2053 102595
rect 2053 102561 2087 102595
rect 2087 102561 2096 102595
rect 2044 102552 2096 102561
rect 7564 102595 7616 102604
rect 7564 102561 7573 102595
rect 7573 102561 7607 102595
rect 7607 102561 7616 102595
rect 7564 102552 7616 102561
rect 37188 102595 37240 102604
rect 37188 102561 37197 102595
rect 37197 102561 37231 102595
rect 37231 102561 37240 102595
rect 37188 102552 37240 102561
rect 37004 102348 37056 102400
rect 4246 102246 4298 102298
rect 4310 102246 4362 102298
rect 4374 102246 4426 102298
rect 4438 102246 4490 102298
rect 34966 102246 35018 102298
rect 35030 102246 35082 102298
rect 35094 102246 35146 102298
rect 35158 102246 35210 102298
rect 30656 102144 30708 102196
rect 31300 102144 31352 102196
rect 32772 102144 32824 102196
rect 36728 102144 36780 102196
rect 25780 102076 25832 102128
rect 1400 101983 1452 101992
rect 1400 101949 1409 101983
rect 1409 101949 1443 101983
rect 1443 101949 1452 101983
rect 1400 101940 1452 101949
rect 18604 101940 18656 101992
rect 37188 101983 37240 101992
rect 37188 101949 37197 101983
rect 37197 101949 37231 101983
rect 37231 101949 37240 101983
rect 37188 101940 37240 101949
rect 38752 101940 38804 101992
rect 12348 101872 12400 101924
rect 37924 101915 37976 101924
rect 37924 101881 37933 101915
rect 37933 101881 37967 101915
rect 37967 101881 37976 101915
rect 37924 101872 37976 101881
rect 1860 101804 1912 101856
rect 36728 101804 36780 101856
rect 19606 101702 19658 101754
rect 19670 101702 19722 101754
rect 19734 101702 19786 101754
rect 19798 101702 19850 101754
rect 37188 101507 37240 101516
rect 37188 101473 37197 101507
rect 37197 101473 37231 101507
rect 37231 101473 37240 101507
rect 37188 101464 37240 101473
rect 35808 101396 35860 101448
rect 37740 101396 37792 101448
rect 31392 101260 31444 101312
rect 4246 101158 4298 101210
rect 4310 101158 4362 101210
rect 4374 101158 4426 101210
rect 4438 101158 4490 101210
rect 34966 101158 35018 101210
rect 35030 101158 35082 101210
rect 35094 101158 35146 101210
rect 35158 101158 35210 101210
rect 2228 101056 2280 101108
rect 1400 100895 1452 100904
rect 1400 100861 1409 100895
rect 1409 100861 1443 100895
rect 1443 100861 1452 100895
rect 1400 100852 1452 100861
rect 10508 100852 10560 100904
rect 37924 100827 37976 100836
rect 37924 100793 37933 100827
rect 37933 100793 37967 100827
rect 37967 100793 37976 100827
rect 37924 100784 37976 100793
rect 36268 100716 36320 100768
rect 19606 100614 19658 100666
rect 19670 100614 19722 100666
rect 19734 100614 19786 100666
rect 19798 100614 19850 100666
rect 34152 100444 34204 100496
rect 37648 100444 37700 100496
rect 1400 100419 1452 100428
rect 1400 100385 1409 100419
rect 1409 100385 1443 100419
rect 1443 100385 1452 100419
rect 1400 100376 1452 100385
rect 37188 100419 37240 100428
rect 37188 100385 37197 100419
rect 37197 100385 37231 100419
rect 37231 100385 37240 100419
rect 37188 100376 37240 100385
rect 33048 100172 33100 100224
rect 4246 100070 4298 100122
rect 4310 100070 4362 100122
rect 4374 100070 4426 100122
rect 4438 100070 4490 100122
rect 34966 100070 35018 100122
rect 35030 100070 35082 100122
rect 35094 100070 35146 100122
rect 35158 100070 35210 100122
rect 6276 100011 6328 100020
rect 6276 99977 6285 100011
rect 6285 99977 6319 100011
rect 6319 99977 6328 100011
rect 6276 99968 6328 99977
rect 36544 99968 36596 100020
rect 37280 99968 37332 100020
rect 34520 99900 34572 99952
rect 13268 99764 13320 99816
rect 37280 99807 37332 99816
rect 37280 99773 37289 99807
rect 37289 99773 37323 99807
rect 37323 99773 37332 99807
rect 37280 99764 37332 99773
rect 37924 99807 37976 99816
rect 37924 99773 37933 99807
rect 37933 99773 37967 99807
rect 37967 99773 37976 99807
rect 37924 99764 37976 99773
rect 36820 99628 36872 99680
rect 19606 99526 19658 99578
rect 19670 99526 19722 99578
rect 19734 99526 19786 99578
rect 19798 99526 19850 99578
rect 1400 99331 1452 99340
rect 1400 99297 1409 99331
rect 1409 99297 1443 99331
rect 1443 99297 1452 99331
rect 1400 99288 1452 99297
rect 5080 99331 5132 99340
rect 5080 99297 5089 99331
rect 5089 99297 5123 99331
rect 5123 99297 5132 99331
rect 5080 99288 5132 99297
rect 37188 99331 37240 99340
rect 37188 99297 37197 99331
rect 37197 99297 37231 99331
rect 37231 99297 37240 99331
rect 37188 99288 37240 99297
rect 2504 99152 2556 99204
rect 34796 99084 34848 99136
rect 4246 98982 4298 99034
rect 4310 98982 4362 99034
rect 4374 98982 4426 99034
rect 4438 98982 4490 99034
rect 34966 98982 35018 99034
rect 35030 98982 35082 99034
rect 35094 98982 35146 99034
rect 35158 98982 35210 99034
rect 35348 98880 35400 98932
rect 1400 98719 1452 98728
rect 1400 98685 1409 98719
rect 1409 98685 1443 98719
rect 1443 98685 1452 98719
rect 1400 98676 1452 98685
rect 37924 98719 37976 98728
rect 37924 98685 37933 98719
rect 37933 98685 37967 98719
rect 37967 98685 37976 98719
rect 37924 98676 37976 98685
rect 35348 98608 35400 98660
rect 35440 98540 35492 98592
rect 19606 98438 19658 98490
rect 19670 98438 19722 98490
rect 19734 98438 19786 98490
rect 19798 98438 19850 98490
rect 2136 98336 2188 98388
rect 4896 98243 4948 98252
rect 4896 98209 4905 98243
rect 4905 98209 4939 98243
rect 4939 98209 4948 98243
rect 4896 98200 4948 98209
rect 37096 98243 37148 98252
rect 37096 98209 37105 98243
rect 37105 98209 37139 98243
rect 37139 98209 37148 98243
rect 37096 98200 37148 98209
rect 33416 97996 33468 98048
rect 4246 97894 4298 97946
rect 4310 97894 4362 97946
rect 4374 97894 4426 97946
rect 4438 97894 4490 97946
rect 34966 97894 35018 97946
rect 35030 97894 35082 97946
rect 35094 97894 35146 97946
rect 35158 97894 35210 97946
rect 1952 97792 2004 97844
rect 1400 97631 1452 97640
rect 1400 97597 1409 97631
rect 1409 97597 1443 97631
rect 1443 97597 1452 97631
rect 1400 97588 1452 97597
rect 8392 97588 8444 97640
rect 37832 97631 37884 97640
rect 37832 97597 37841 97631
rect 37841 97597 37875 97631
rect 37875 97597 37884 97631
rect 37832 97588 37884 97597
rect 33508 97452 33560 97504
rect 19606 97350 19658 97402
rect 19670 97350 19722 97402
rect 19734 97350 19786 97402
rect 19798 97350 19850 97402
rect 1400 97155 1452 97164
rect 1400 97121 1409 97155
rect 1409 97121 1443 97155
rect 1443 97121 1452 97155
rect 1400 97112 1452 97121
rect 37096 97155 37148 97164
rect 37096 97121 37105 97155
rect 37105 97121 37139 97155
rect 37139 97121 37148 97155
rect 37096 97112 37148 97121
rect 33140 96908 33192 96960
rect 4246 96806 4298 96858
rect 4310 96806 4362 96858
rect 4374 96806 4426 96858
rect 4438 96806 4490 96858
rect 34966 96806 35018 96858
rect 35030 96806 35082 96858
rect 35094 96806 35146 96858
rect 35158 96806 35210 96858
rect 37096 96543 37148 96552
rect 37096 96509 37105 96543
rect 37105 96509 37139 96543
rect 37139 96509 37148 96543
rect 37096 96500 37148 96509
rect 32220 96432 32272 96484
rect 37924 96475 37976 96484
rect 33692 96364 33744 96416
rect 37924 96441 37933 96475
rect 37933 96441 37967 96475
rect 37967 96441 37976 96475
rect 37924 96432 37976 96441
rect 19606 96262 19658 96314
rect 19670 96262 19722 96314
rect 19734 96262 19786 96314
rect 19798 96262 19850 96314
rect 3516 96203 3568 96212
rect 3516 96169 3525 96203
rect 3525 96169 3559 96203
rect 3559 96169 3568 96203
rect 3516 96160 3568 96169
rect 1400 96067 1452 96076
rect 1400 96033 1409 96067
rect 1409 96033 1443 96067
rect 1443 96033 1452 96067
rect 1400 96024 1452 96033
rect 5264 96024 5316 96076
rect 37188 96067 37240 96076
rect 37188 96033 37197 96067
rect 37197 96033 37231 96067
rect 37231 96033 37240 96067
rect 37188 96024 37240 96033
rect 23480 95888 23532 95940
rect 38568 95956 38620 96008
rect 38384 95888 38436 95940
rect 4246 95718 4298 95770
rect 4310 95718 4362 95770
rect 4374 95718 4426 95770
rect 4438 95718 4490 95770
rect 34966 95718 35018 95770
rect 35030 95718 35082 95770
rect 35094 95718 35146 95770
rect 35158 95718 35210 95770
rect 2412 95616 2464 95668
rect 30748 95616 30800 95668
rect 32404 95616 32456 95668
rect 1400 95455 1452 95464
rect 1400 95421 1409 95455
rect 1409 95421 1443 95455
rect 1443 95421 1452 95455
rect 1400 95412 1452 95421
rect 6184 95412 6236 95464
rect 31484 95412 31536 95464
rect 37924 95387 37976 95396
rect 37924 95353 37933 95387
rect 37933 95353 37967 95387
rect 37967 95353 37976 95387
rect 37924 95344 37976 95353
rect 19606 95174 19658 95226
rect 19670 95174 19722 95226
rect 19734 95174 19786 95226
rect 19798 95174 19850 95226
rect 37188 94979 37240 94988
rect 37188 94945 37197 94979
rect 37197 94945 37231 94979
rect 37231 94945 37240 94979
rect 37188 94936 37240 94945
rect 32036 94800 32088 94852
rect 35256 94800 35308 94852
rect 33876 94732 33928 94784
rect 34060 94732 34112 94784
rect 35440 94732 35492 94784
rect 35900 94732 35952 94784
rect 37004 94732 37056 94784
rect 4246 94630 4298 94682
rect 4310 94630 4362 94682
rect 4374 94630 4426 94682
rect 4438 94630 4490 94682
rect 34966 94630 35018 94682
rect 35030 94630 35082 94682
rect 35094 94630 35146 94682
rect 35158 94630 35210 94682
rect 2872 94571 2924 94580
rect 2872 94537 2881 94571
rect 2881 94537 2915 94571
rect 2915 94537 2924 94571
rect 2872 94528 2924 94537
rect 32404 94460 32456 94512
rect 34336 94460 34388 94512
rect 35256 94460 35308 94512
rect 35624 94460 35676 94512
rect 1400 94367 1452 94376
rect 1400 94333 1409 94367
rect 1409 94333 1443 94367
rect 1443 94333 1452 94367
rect 1400 94324 1452 94333
rect 5356 94324 5408 94376
rect 35440 94324 35492 94376
rect 35808 94324 35860 94376
rect 37188 94367 37240 94376
rect 37188 94333 37197 94367
rect 37197 94333 37231 94367
rect 37231 94333 37240 94367
rect 37188 94324 37240 94333
rect 37924 94299 37976 94308
rect 37924 94265 37933 94299
rect 37933 94265 37967 94299
rect 37967 94265 37976 94299
rect 37924 94256 37976 94265
rect 35808 94188 35860 94240
rect 37556 94188 37608 94240
rect 19606 94086 19658 94138
rect 19670 94086 19722 94138
rect 19734 94086 19786 94138
rect 19798 94086 19850 94138
rect 33968 93984 34020 94036
rect 1400 93891 1452 93900
rect 1400 93857 1409 93891
rect 1409 93857 1443 93891
rect 1443 93857 1452 93891
rect 1400 93848 1452 93857
rect 37188 93891 37240 93900
rect 37188 93857 37197 93891
rect 37197 93857 37231 93891
rect 37231 93857 37240 93891
rect 37188 93848 37240 93857
rect 36636 93780 36688 93832
rect 37372 93780 37424 93832
rect 4246 93542 4298 93594
rect 4310 93542 4362 93594
rect 4374 93542 4426 93594
rect 4438 93542 4490 93594
rect 34966 93542 35018 93594
rect 35030 93542 35082 93594
rect 35094 93542 35146 93594
rect 35158 93542 35210 93594
rect 30840 93304 30892 93356
rect 33876 93304 33928 93356
rect 1400 93279 1452 93288
rect 1400 93245 1409 93279
rect 1409 93245 1443 93279
rect 1443 93245 1452 93279
rect 1400 93236 1452 93245
rect 37280 93279 37332 93288
rect 37280 93245 37289 93279
rect 37289 93245 37323 93279
rect 37323 93245 37332 93279
rect 37280 93236 37332 93245
rect 37924 93279 37976 93288
rect 37924 93245 37933 93279
rect 37933 93245 37967 93279
rect 37967 93245 37976 93279
rect 37924 93236 37976 93245
rect 35624 93100 35676 93152
rect 38108 93143 38160 93152
rect 38108 93109 38117 93143
rect 38117 93109 38151 93143
rect 38151 93109 38160 93143
rect 38108 93100 38160 93109
rect 19606 92998 19658 93050
rect 19670 92998 19722 93050
rect 19734 92998 19786 93050
rect 19798 92998 19850 93050
rect 2320 92939 2372 92948
rect 2320 92905 2329 92939
rect 2329 92905 2363 92939
rect 2363 92905 2372 92939
rect 2320 92896 2372 92905
rect 30748 92871 30800 92880
rect 30748 92837 30757 92871
rect 30757 92837 30791 92871
rect 30791 92837 30800 92871
rect 30748 92828 30800 92837
rect 4804 92760 4856 92812
rect 21364 92760 21416 92812
rect 4246 92454 4298 92506
rect 4310 92454 4362 92506
rect 4374 92454 4426 92506
rect 4438 92454 4490 92506
rect 34966 92454 35018 92506
rect 35030 92454 35082 92506
rect 35094 92454 35146 92506
rect 35158 92454 35210 92506
rect 1400 92191 1452 92200
rect 1400 92157 1409 92191
rect 1409 92157 1443 92191
rect 1443 92157 1452 92191
rect 1400 92148 1452 92157
rect 37280 92191 37332 92200
rect 37280 92157 37289 92191
rect 37289 92157 37323 92191
rect 37323 92157 37332 92191
rect 37280 92148 37332 92157
rect 37924 92191 37976 92200
rect 37924 92157 37933 92191
rect 37933 92157 37967 92191
rect 37967 92157 37976 92191
rect 37924 92148 37976 92157
rect 37372 92012 37424 92064
rect 37832 92012 37884 92064
rect 19606 91910 19658 91962
rect 19670 91910 19722 91962
rect 19734 91910 19786 91962
rect 19798 91910 19850 91962
rect 21548 91808 21600 91860
rect 32956 91808 33008 91860
rect 19340 91740 19392 91792
rect 33600 91740 33652 91792
rect 1400 91715 1452 91724
rect 1400 91681 1409 91715
rect 1409 91681 1443 91715
rect 1443 91681 1452 91715
rect 1400 91672 1452 91681
rect 37188 91715 37240 91724
rect 37188 91681 37197 91715
rect 37197 91681 37231 91715
rect 37231 91681 37240 91715
rect 37188 91672 37240 91681
rect 33968 91536 34020 91588
rect 35624 91536 35676 91588
rect 37280 91468 37332 91520
rect 4246 91366 4298 91418
rect 4310 91366 4362 91418
rect 4374 91366 4426 91418
rect 4438 91366 4490 91418
rect 34966 91366 35018 91418
rect 35030 91366 35082 91418
rect 35094 91366 35146 91418
rect 35158 91366 35210 91418
rect 1676 91264 1728 91316
rect 37740 91196 37792 91248
rect 27988 91128 28040 91180
rect 31760 91128 31812 91180
rect 1400 91103 1452 91112
rect 1400 91069 1409 91103
rect 1409 91069 1443 91103
rect 1443 91069 1452 91103
rect 1400 91060 1452 91069
rect 31668 91060 31720 91112
rect 33048 91060 33100 91112
rect 37188 91060 37240 91112
rect 37924 91103 37976 91112
rect 37924 91069 37933 91103
rect 37933 91069 37967 91103
rect 37967 91069 37976 91103
rect 37924 91060 37976 91069
rect 37464 90967 37516 90976
rect 37464 90933 37473 90967
rect 37473 90933 37507 90967
rect 37507 90933 37516 90967
rect 37464 90924 37516 90933
rect 19606 90822 19658 90874
rect 19670 90822 19722 90874
rect 19734 90822 19786 90874
rect 19798 90822 19850 90874
rect 1492 90720 1544 90772
rect 2044 90627 2096 90636
rect 2044 90593 2053 90627
rect 2053 90593 2087 90627
rect 2087 90593 2096 90627
rect 2044 90584 2096 90593
rect 2872 90516 2924 90568
rect 4246 90278 4298 90330
rect 4310 90278 4362 90330
rect 4374 90278 4426 90330
rect 4438 90278 4490 90330
rect 34966 90278 35018 90330
rect 35030 90278 35082 90330
rect 35094 90278 35146 90330
rect 35158 90278 35210 90330
rect 35164 90108 35216 90160
rect 35900 90108 35952 90160
rect 36084 90108 36136 90160
rect 34888 90040 34940 90092
rect 35440 90040 35492 90092
rect 1400 90015 1452 90024
rect 1400 89981 1409 90015
rect 1409 89981 1443 90015
rect 1443 89981 1452 90015
rect 1400 89972 1452 89981
rect 37280 90015 37332 90024
rect 37280 89981 37289 90015
rect 37289 89981 37323 90015
rect 37323 89981 37332 90015
rect 37280 89972 37332 89981
rect 37464 89972 37516 90024
rect 37924 90015 37976 90024
rect 37924 89981 37933 90015
rect 37933 89981 37967 90015
rect 37967 89981 37976 90015
rect 37924 89972 37976 89981
rect 33600 89904 33652 89956
rect 35256 89904 35308 89956
rect 35900 89904 35952 89956
rect 34796 89836 34848 89888
rect 35440 89836 35492 89888
rect 37464 89879 37516 89888
rect 37464 89845 37473 89879
rect 37473 89845 37507 89879
rect 37507 89845 37516 89879
rect 37464 89836 37516 89845
rect 19606 89734 19658 89786
rect 19670 89734 19722 89786
rect 19734 89734 19786 89786
rect 19798 89734 19850 89786
rect 37188 89539 37240 89548
rect 37188 89505 37197 89539
rect 37197 89505 37231 89539
rect 37231 89505 37240 89539
rect 37188 89496 37240 89505
rect 37648 89292 37700 89344
rect 4246 89190 4298 89242
rect 4310 89190 4362 89242
rect 4374 89190 4426 89242
rect 4438 89190 4490 89242
rect 34966 89190 35018 89242
rect 35030 89190 35082 89242
rect 35094 89190 35146 89242
rect 35158 89190 35210 89242
rect 1400 88927 1452 88936
rect 1400 88893 1409 88927
rect 1409 88893 1443 88927
rect 1443 88893 1452 88927
rect 1400 88884 1452 88893
rect 37280 88927 37332 88936
rect 37280 88893 37289 88927
rect 37289 88893 37323 88927
rect 37323 88893 37332 88927
rect 37280 88884 37332 88893
rect 37924 88927 37976 88936
rect 37924 88893 37933 88927
rect 37933 88893 37967 88927
rect 37967 88893 37976 88927
rect 37924 88884 37976 88893
rect 37832 88748 37884 88800
rect 38292 88748 38344 88800
rect 19606 88646 19658 88698
rect 19670 88646 19722 88698
rect 19734 88646 19786 88698
rect 19798 88646 19850 88698
rect 1400 88451 1452 88460
rect 1400 88417 1409 88451
rect 1409 88417 1443 88451
rect 1443 88417 1452 88451
rect 1400 88408 1452 88417
rect 35624 88340 35676 88392
rect 37556 88340 37608 88392
rect 30748 88272 30800 88324
rect 34060 88272 34112 88324
rect 4246 88102 4298 88154
rect 4310 88102 4362 88154
rect 4374 88102 4426 88154
rect 4438 88102 4490 88154
rect 34966 88102 35018 88154
rect 35030 88102 35082 88154
rect 35094 88102 35146 88154
rect 35158 88102 35210 88154
rect 34152 87864 34204 87916
rect 33784 87839 33836 87848
rect 33784 87805 33793 87839
rect 33793 87805 33827 87839
rect 33827 87805 33836 87839
rect 34060 87839 34112 87848
rect 33784 87796 33836 87805
rect 34060 87805 34069 87839
rect 34069 87805 34103 87839
rect 34103 87805 34112 87839
rect 34060 87796 34112 87805
rect 34336 87839 34388 87848
rect 34336 87805 34345 87839
rect 34345 87805 34379 87839
rect 34379 87805 34388 87839
rect 34336 87796 34388 87805
rect 35256 87796 35308 87848
rect 37280 87839 37332 87848
rect 37280 87805 37289 87839
rect 37289 87805 37323 87839
rect 37323 87805 37332 87839
rect 37280 87796 37332 87805
rect 37924 87839 37976 87848
rect 37924 87805 37933 87839
rect 37933 87805 37967 87839
rect 37967 87805 37976 87839
rect 37924 87796 37976 87805
rect 27896 87728 27948 87780
rect 35256 87660 35308 87712
rect 37464 87703 37516 87712
rect 37464 87669 37473 87703
rect 37473 87669 37507 87703
rect 37507 87669 37516 87703
rect 37464 87660 37516 87669
rect 19606 87558 19658 87610
rect 19670 87558 19722 87610
rect 19734 87558 19786 87610
rect 19798 87558 19850 87610
rect 1400 87363 1452 87372
rect 1400 87329 1409 87363
rect 1409 87329 1443 87363
rect 1443 87329 1452 87363
rect 1400 87320 1452 87329
rect 21180 87320 21232 87372
rect 36636 87456 36688 87508
rect 37188 87456 37240 87508
rect 34152 87388 34204 87440
rect 35900 87388 35952 87440
rect 33784 87363 33836 87372
rect 33784 87329 33793 87363
rect 33793 87329 33827 87363
rect 33827 87329 33836 87363
rect 33784 87320 33836 87329
rect 34336 87363 34388 87372
rect 34336 87329 34345 87363
rect 34345 87329 34379 87363
rect 34379 87329 34388 87363
rect 34336 87320 34388 87329
rect 35440 87320 35492 87372
rect 37188 87363 37240 87372
rect 37188 87329 37197 87363
rect 37197 87329 37231 87363
rect 37231 87329 37240 87363
rect 37188 87320 37240 87329
rect 34704 87252 34756 87304
rect 20352 87184 20404 87236
rect 34060 87184 34112 87236
rect 36636 87184 36688 87236
rect 36912 87184 36964 87236
rect 37188 87184 37240 87236
rect 28632 87116 28684 87168
rect 34704 87116 34756 87168
rect 35900 87116 35952 87168
rect 4246 87014 4298 87066
rect 4310 87014 4362 87066
rect 4374 87014 4426 87066
rect 4438 87014 4490 87066
rect 34966 87014 35018 87066
rect 35030 87014 35082 87066
rect 35094 87014 35146 87066
rect 35158 87014 35210 87066
rect 30932 86844 30984 86896
rect 33784 86844 33836 86896
rect 36728 86844 36780 86896
rect 33324 86776 33376 86828
rect 1400 86751 1452 86760
rect 1400 86717 1409 86751
rect 1409 86717 1443 86751
rect 1443 86717 1452 86751
rect 1400 86708 1452 86717
rect 27160 86708 27212 86760
rect 32128 86708 32180 86760
rect 32772 86708 32824 86760
rect 34796 86776 34848 86828
rect 35440 86776 35492 86828
rect 35624 86776 35676 86828
rect 33784 86751 33836 86760
rect 33784 86717 33793 86751
rect 33793 86717 33827 86751
rect 33827 86717 33836 86751
rect 33784 86708 33836 86717
rect 34336 86751 34388 86760
rect 28356 86640 28408 86692
rect 29644 86572 29696 86624
rect 32312 86572 32364 86624
rect 32772 86572 32824 86624
rect 34336 86717 34345 86751
rect 34345 86717 34379 86751
rect 34379 86717 34388 86751
rect 34336 86708 34388 86717
rect 36820 86708 36872 86760
rect 37280 86751 37332 86760
rect 37280 86717 37289 86751
rect 37289 86717 37323 86751
rect 37323 86717 37332 86751
rect 37280 86708 37332 86717
rect 37924 86751 37976 86760
rect 37924 86717 37933 86751
rect 37933 86717 37967 86751
rect 37967 86717 37976 86751
rect 37924 86708 37976 86717
rect 34796 86640 34848 86692
rect 37188 86640 37240 86692
rect 35624 86572 35676 86624
rect 19606 86470 19658 86522
rect 19670 86470 19722 86522
rect 19734 86470 19786 86522
rect 19798 86470 19850 86522
rect 20536 86232 20588 86284
rect 20444 86096 20496 86148
rect 32772 86096 32824 86148
rect 33784 86275 33836 86284
rect 33784 86241 33793 86275
rect 33793 86241 33827 86275
rect 33827 86241 33836 86275
rect 33784 86232 33836 86241
rect 34336 86275 34388 86284
rect 34336 86241 34345 86275
rect 34345 86241 34379 86275
rect 34379 86241 34388 86275
rect 34336 86232 34388 86241
rect 34520 86275 34572 86284
rect 34520 86241 34529 86275
rect 34529 86241 34563 86275
rect 34563 86241 34572 86275
rect 34520 86232 34572 86241
rect 36544 86164 36596 86216
rect 36176 86096 36228 86148
rect 37096 86096 37148 86148
rect 32956 86028 33008 86080
rect 34152 86028 34204 86080
rect 34336 86028 34388 86080
rect 4246 85926 4298 85978
rect 4310 85926 4362 85978
rect 4374 85926 4426 85978
rect 4438 85926 4490 85978
rect 34966 85926 35018 85978
rect 35030 85926 35082 85978
rect 35094 85926 35146 85978
rect 35158 85926 35210 85978
rect 31760 85824 31812 85876
rect 32312 85824 32364 85876
rect 32772 85824 32824 85876
rect 36176 85824 36228 85876
rect 16948 85756 17000 85808
rect 32312 85688 32364 85740
rect 1400 85663 1452 85672
rect 1400 85629 1409 85663
rect 1409 85629 1443 85663
rect 1443 85629 1452 85663
rect 1400 85620 1452 85629
rect 27160 85663 27212 85672
rect 27160 85629 27169 85663
rect 27169 85629 27203 85663
rect 27203 85629 27212 85663
rect 27160 85620 27212 85629
rect 32404 85663 32456 85672
rect 32404 85629 32413 85663
rect 32413 85629 32447 85663
rect 32447 85629 32456 85663
rect 32404 85620 32456 85629
rect 33324 85756 33376 85808
rect 36636 85756 36688 85808
rect 33968 85620 34020 85672
rect 37280 85663 37332 85672
rect 37280 85629 37289 85663
rect 37289 85629 37323 85663
rect 37323 85629 37332 85663
rect 37280 85620 37332 85629
rect 37924 85663 37976 85672
rect 37924 85629 37933 85663
rect 37933 85629 37967 85663
rect 37967 85629 37976 85663
rect 37924 85620 37976 85629
rect 28264 85552 28316 85604
rect 34520 85552 34572 85604
rect 35624 85552 35676 85604
rect 32404 85484 32456 85536
rect 33600 85484 33652 85536
rect 19606 85382 19658 85434
rect 19670 85382 19722 85434
rect 19734 85382 19786 85434
rect 19798 85382 19850 85434
rect 1400 85187 1452 85196
rect 1400 85153 1409 85187
rect 1409 85153 1443 85187
rect 1443 85153 1452 85187
rect 1400 85144 1452 85153
rect 32128 85144 32180 85196
rect 33600 84940 33652 84992
rect 4246 84838 4298 84890
rect 4310 84838 4362 84890
rect 4374 84838 4426 84890
rect 4438 84838 4490 84890
rect 34966 84838 35018 84890
rect 35030 84838 35082 84890
rect 35094 84838 35146 84890
rect 35158 84838 35210 84890
rect 33048 84736 33100 84788
rect 36544 84736 36596 84788
rect 34152 84668 34204 84720
rect 17684 84600 17736 84652
rect 26976 84575 27028 84584
rect 26976 84541 26985 84575
rect 26985 84541 27019 84575
rect 27019 84541 27028 84575
rect 26976 84532 27028 84541
rect 27160 84532 27212 84584
rect 32128 84532 32180 84584
rect 32496 84575 32548 84584
rect 32496 84541 32505 84575
rect 32505 84541 32539 84575
rect 32539 84541 32548 84575
rect 32496 84532 32548 84541
rect 32772 84575 32824 84584
rect 32772 84541 32781 84575
rect 32781 84541 32815 84575
rect 32815 84541 32824 84575
rect 32772 84532 32824 84541
rect 33324 84532 33376 84584
rect 33876 84532 33928 84584
rect 37280 84575 37332 84584
rect 37280 84541 37289 84575
rect 37289 84541 37323 84575
rect 37323 84541 37332 84575
rect 37280 84532 37332 84541
rect 37924 84575 37976 84584
rect 37924 84541 37933 84575
rect 37933 84541 37967 84575
rect 37967 84541 37976 84575
rect 37924 84532 37976 84541
rect 29368 84464 29420 84516
rect 34060 84464 34112 84516
rect 33784 84396 33836 84448
rect 36820 84396 36872 84448
rect 39396 84396 39448 84448
rect 19606 84294 19658 84346
rect 19670 84294 19722 84346
rect 19734 84294 19786 84346
rect 19798 84294 19850 84346
rect 32128 84192 32180 84244
rect 32496 84192 32548 84244
rect 33324 84192 33376 84244
rect 1400 84099 1452 84108
rect 1400 84065 1409 84099
rect 1409 84065 1443 84099
rect 1443 84065 1452 84099
rect 1400 84056 1452 84065
rect 30840 84056 30892 84108
rect 32404 84124 32456 84176
rect 32772 84124 32824 84176
rect 34060 84124 34112 84176
rect 16488 83988 16540 84040
rect 30380 83920 30432 83972
rect 29184 83852 29236 83904
rect 33968 84056 34020 84108
rect 37372 84124 37424 84176
rect 37188 84099 37240 84108
rect 37188 84065 37197 84099
rect 37197 84065 37231 84099
rect 37231 84065 37240 84099
rect 37188 84056 37240 84065
rect 33324 83852 33376 83904
rect 35532 83920 35584 83972
rect 34796 83852 34848 83904
rect 37372 83895 37424 83904
rect 37372 83861 37381 83895
rect 37381 83861 37415 83895
rect 37415 83861 37424 83895
rect 37372 83852 37424 83861
rect 4246 83750 4298 83802
rect 4310 83750 4362 83802
rect 4374 83750 4426 83802
rect 4438 83750 4490 83802
rect 34966 83750 35018 83802
rect 35030 83750 35082 83802
rect 35094 83750 35146 83802
rect 35158 83750 35210 83802
rect 32772 83648 32824 83700
rect 34336 83648 34388 83700
rect 17776 83512 17828 83564
rect 29276 83512 29328 83564
rect 1400 83487 1452 83496
rect 1400 83453 1409 83487
rect 1409 83453 1443 83487
rect 1443 83453 1452 83487
rect 1400 83444 1452 83453
rect 17868 83444 17920 83496
rect 32312 83487 32364 83496
rect 32312 83453 32321 83487
rect 32321 83453 32355 83487
rect 32355 83453 32364 83487
rect 32312 83444 32364 83453
rect 32404 83487 32456 83496
rect 32404 83453 32413 83487
rect 32413 83453 32447 83487
rect 32447 83453 32456 83487
rect 33324 83512 33376 83564
rect 32404 83444 32456 83453
rect 38108 83512 38160 83564
rect 37280 83487 37332 83496
rect 37280 83453 37289 83487
rect 37289 83453 37323 83487
rect 37323 83453 37332 83487
rect 37280 83444 37332 83453
rect 37924 83487 37976 83496
rect 37924 83453 37933 83487
rect 37933 83453 37967 83487
rect 37967 83453 37976 83487
rect 37924 83444 37976 83453
rect 29552 83376 29604 83428
rect 32128 83308 32180 83360
rect 33600 83376 33652 83428
rect 36544 83308 36596 83360
rect 39028 83308 39080 83360
rect 19606 83206 19658 83258
rect 19670 83206 19722 83258
rect 19734 83206 19786 83258
rect 19798 83206 19850 83258
rect 29276 83104 29328 83156
rect 29276 82968 29328 83020
rect 29552 82968 29604 83020
rect 30656 83011 30708 83020
rect 30656 82977 30665 83011
rect 30665 82977 30699 83011
rect 30699 82977 30708 83011
rect 30656 82968 30708 82977
rect 30748 82968 30800 83020
rect 32128 83036 32180 83088
rect 16028 82900 16080 82952
rect 31760 83011 31812 83020
rect 31760 82977 31769 83011
rect 31769 82977 31803 83011
rect 31803 82977 31812 83011
rect 31760 82968 31812 82977
rect 32772 82968 32824 83020
rect 33600 83011 33652 83020
rect 33600 82977 33609 83011
rect 33609 82977 33643 83011
rect 33643 82977 33652 83011
rect 33600 82968 33652 82977
rect 35992 83036 36044 83088
rect 24216 82832 24268 82884
rect 37740 82968 37792 83020
rect 37556 82832 37608 82884
rect 37740 82832 37792 82884
rect 32772 82764 32824 82816
rect 37096 82764 37148 82816
rect 4246 82662 4298 82714
rect 4310 82662 4362 82714
rect 4374 82662 4426 82714
rect 4438 82662 4490 82714
rect 34966 82662 35018 82714
rect 35030 82662 35082 82714
rect 35094 82662 35146 82714
rect 35158 82662 35210 82714
rect 1400 82399 1452 82408
rect 1400 82365 1409 82399
rect 1409 82365 1443 82399
rect 1443 82365 1452 82399
rect 1400 82356 1452 82365
rect 32036 82492 32088 82544
rect 32128 82424 32180 82476
rect 32312 82399 32364 82408
rect 32312 82365 32321 82399
rect 32321 82365 32355 82399
rect 32355 82365 32364 82399
rect 32312 82356 32364 82365
rect 38016 82424 38068 82476
rect 37280 82399 37332 82408
rect 29828 82288 29880 82340
rect 31760 82220 31812 82272
rect 32404 82220 32456 82272
rect 37280 82365 37289 82399
rect 37289 82365 37323 82399
rect 37323 82365 37332 82399
rect 37280 82356 37332 82365
rect 37924 82399 37976 82408
rect 37924 82365 37933 82399
rect 37933 82365 37967 82399
rect 37967 82365 37976 82399
rect 37924 82356 37976 82365
rect 35532 82220 35584 82272
rect 35808 82220 35860 82272
rect 37556 82220 37608 82272
rect 39948 82220 40000 82272
rect 19606 82118 19658 82170
rect 19670 82118 19722 82170
rect 19734 82118 19786 82170
rect 19798 82118 19850 82170
rect 1400 81923 1452 81932
rect 1400 81889 1409 81923
rect 1409 81889 1443 81923
rect 1443 81889 1452 81923
rect 1400 81880 1452 81889
rect 31208 82016 31260 82068
rect 32128 81948 32180 82000
rect 16672 81812 16724 81864
rect 31760 81923 31812 81932
rect 31760 81889 31769 81923
rect 31769 81889 31803 81923
rect 31803 81889 31812 81923
rect 31760 81880 31812 81889
rect 37648 82016 37700 82068
rect 33600 81923 33652 81932
rect 33600 81889 33609 81923
rect 33609 81889 33643 81923
rect 33643 81889 33652 81923
rect 33600 81880 33652 81889
rect 38200 81948 38252 82000
rect 34152 81923 34204 81932
rect 15844 81744 15896 81796
rect 34152 81889 34161 81923
rect 34161 81889 34195 81923
rect 34195 81889 34204 81923
rect 34152 81880 34204 81889
rect 36084 81880 36136 81932
rect 37188 81923 37240 81932
rect 37188 81889 37197 81923
rect 37197 81889 37231 81923
rect 37231 81889 37240 81923
rect 37188 81880 37240 81889
rect 36268 81744 36320 81796
rect 37188 81744 37240 81796
rect 26516 81676 26568 81728
rect 31760 81676 31812 81728
rect 32772 81676 32824 81728
rect 33140 81719 33192 81728
rect 33140 81685 33149 81719
rect 33149 81685 33183 81719
rect 33183 81685 33192 81719
rect 33140 81676 33192 81685
rect 33600 81676 33652 81728
rect 33784 81676 33836 81728
rect 39672 81676 39724 81728
rect 4246 81574 4298 81626
rect 4310 81574 4362 81626
rect 4374 81574 4426 81626
rect 4438 81574 4490 81626
rect 34966 81574 35018 81626
rect 35030 81574 35082 81626
rect 35094 81574 35146 81626
rect 35158 81574 35210 81626
rect 23572 81472 23624 81524
rect 33140 81472 33192 81524
rect 36268 81472 36320 81524
rect 36728 81472 36780 81524
rect 25596 81404 25648 81456
rect 32312 81404 32364 81456
rect 15568 81336 15620 81388
rect 33600 81336 33652 81388
rect 30840 81268 30892 81320
rect 31576 81268 31628 81320
rect 31760 81311 31812 81320
rect 31760 81277 31769 81311
rect 31769 81277 31803 81311
rect 31803 81277 31812 81311
rect 32036 81311 32088 81320
rect 31760 81268 31812 81277
rect 32036 81277 32045 81311
rect 32045 81277 32079 81311
rect 32079 81277 32088 81311
rect 32036 81268 32088 81277
rect 32404 81311 32456 81320
rect 31576 81132 31628 81184
rect 31760 81132 31812 81184
rect 32404 81277 32413 81311
rect 32413 81277 32447 81311
rect 32447 81277 32456 81311
rect 32404 81268 32456 81277
rect 33968 81336 34020 81388
rect 33784 81311 33836 81320
rect 33784 81277 33793 81311
rect 33793 81277 33827 81311
rect 33827 81277 33836 81311
rect 34060 81311 34112 81320
rect 33784 81268 33836 81277
rect 34060 81277 34069 81311
rect 34069 81277 34103 81311
rect 34103 81277 34112 81311
rect 34060 81268 34112 81277
rect 34152 81268 34204 81320
rect 37464 81336 37516 81388
rect 37648 81336 37700 81388
rect 37280 81311 37332 81320
rect 37280 81277 37289 81311
rect 37289 81277 37323 81311
rect 37323 81277 37332 81311
rect 37280 81268 37332 81277
rect 37740 81268 37792 81320
rect 37924 81311 37976 81320
rect 37924 81277 37933 81311
rect 37933 81277 37967 81311
rect 37967 81277 37976 81311
rect 37924 81268 37976 81277
rect 33324 81175 33376 81184
rect 33324 81141 33333 81175
rect 33333 81141 33367 81175
rect 33367 81141 33376 81175
rect 33324 81132 33376 81141
rect 38292 81132 38344 81184
rect 19606 81030 19658 81082
rect 19670 81030 19722 81082
rect 19734 81030 19786 81082
rect 19798 81030 19850 81082
rect 26424 80928 26476 80980
rect 33600 80928 33652 80980
rect 1400 80835 1452 80844
rect 1400 80801 1409 80835
rect 1409 80801 1443 80835
rect 1443 80801 1452 80835
rect 1400 80792 1452 80801
rect 30840 80792 30892 80844
rect 31208 80835 31260 80844
rect 31208 80801 31217 80835
rect 31217 80801 31251 80835
rect 31251 80801 31260 80835
rect 31208 80792 31260 80801
rect 33784 80835 33836 80844
rect 17500 80724 17552 80776
rect 32036 80724 32088 80776
rect 33784 80801 33793 80835
rect 33793 80801 33827 80835
rect 33827 80801 33836 80835
rect 33784 80792 33836 80801
rect 33968 80928 34020 80980
rect 38752 80928 38804 80980
rect 34152 80835 34204 80844
rect 34152 80801 34161 80835
rect 34161 80801 34195 80835
rect 34195 80801 34204 80835
rect 34152 80792 34204 80801
rect 35900 80792 35952 80844
rect 23756 80656 23808 80708
rect 33324 80656 33376 80708
rect 36912 80724 36964 80776
rect 34152 80656 34204 80708
rect 25504 80588 25556 80640
rect 37832 80588 37884 80640
rect 4246 80486 4298 80538
rect 4310 80486 4362 80538
rect 4374 80486 4426 80538
rect 4438 80486 4490 80538
rect 34966 80486 35018 80538
rect 35030 80486 35082 80538
rect 35094 80486 35146 80538
rect 35158 80486 35210 80538
rect 31208 80384 31260 80436
rect 1400 80223 1452 80232
rect 1400 80189 1409 80223
rect 1409 80189 1443 80223
rect 1443 80189 1452 80223
rect 1400 80180 1452 80189
rect 16212 80180 16264 80232
rect 26792 80112 26844 80164
rect 33784 80384 33836 80436
rect 39856 80316 39908 80368
rect 32036 80223 32088 80232
rect 32036 80189 32045 80223
rect 32045 80189 32079 80223
rect 32079 80189 32088 80223
rect 32036 80180 32088 80189
rect 38200 80248 38252 80300
rect 37280 80223 37332 80232
rect 37280 80189 37289 80223
rect 37289 80189 37323 80223
rect 37323 80189 37332 80223
rect 37280 80180 37332 80189
rect 37924 80223 37976 80232
rect 37924 80189 37933 80223
rect 37933 80189 37967 80223
rect 37967 80189 37976 80223
rect 37924 80180 37976 80189
rect 37096 80044 37148 80096
rect 39488 80044 39540 80096
rect 19606 79942 19658 79994
rect 19670 79942 19722 79994
rect 19734 79942 19786 79994
rect 19798 79942 19850 79994
rect 30748 79840 30800 79892
rect 37188 79840 37240 79892
rect 1400 79747 1452 79756
rect 1400 79713 1409 79747
rect 1409 79713 1443 79747
rect 1443 79713 1452 79747
rect 1400 79704 1452 79713
rect 14832 79747 14884 79756
rect 14832 79713 14841 79747
rect 14841 79713 14875 79747
rect 14875 79713 14884 79747
rect 14832 79704 14884 79713
rect 37188 79747 37240 79756
rect 37188 79713 37197 79747
rect 37197 79713 37231 79747
rect 37231 79713 37240 79747
rect 37188 79704 37240 79713
rect 2596 79500 2648 79552
rect 17132 79500 17184 79552
rect 33876 79500 33928 79552
rect 38568 79500 38620 79552
rect 4246 79398 4298 79450
rect 4310 79398 4362 79450
rect 4374 79398 4426 79450
rect 4438 79398 4490 79450
rect 34966 79398 35018 79450
rect 35030 79398 35082 79450
rect 35094 79398 35146 79450
rect 35158 79398 35210 79450
rect 16304 79296 16356 79348
rect 34060 79296 34112 79348
rect 38752 79228 38804 79280
rect 37280 79135 37332 79144
rect 37280 79101 37289 79135
rect 37289 79101 37323 79135
rect 37323 79101 37332 79135
rect 37280 79092 37332 79101
rect 37924 79135 37976 79144
rect 37924 79101 37933 79135
rect 37933 79101 37967 79135
rect 37967 79101 37976 79135
rect 37924 79092 37976 79101
rect 39120 78956 39172 79008
rect 19606 78854 19658 78906
rect 19670 78854 19722 78906
rect 19734 78854 19786 78906
rect 19798 78854 19850 78906
rect 1400 78659 1452 78668
rect 1400 78625 1409 78659
rect 1409 78625 1443 78659
rect 1443 78625 1452 78659
rect 1400 78616 1452 78625
rect 26976 78616 27028 78668
rect 30840 78412 30892 78464
rect 4246 78310 4298 78362
rect 4310 78310 4362 78362
rect 4374 78310 4426 78362
rect 4438 78310 4490 78362
rect 34966 78310 35018 78362
rect 35030 78310 35082 78362
rect 35094 78310 35146 78362
rect 35158 78310 35210 78362
rect 39304 78140 39356 78192
rect 1400 78047 1452 78056
rect 1400 78013 1409 78047
rect 1409 78013 1443 78047
rect 1443 78013 1452 78047
rect 1400 78004 1452 78013
rect 32496 78004 32548 78056
rect 37280 78047 37332 78056
rect 37280 78013 37289 78047
rect 37289 78013 37323 78047
rect 37323 78013 37332 78047
rect 37280 78004 37332 78013
rect 37924 78047 37976 78056
rect 37924 78013 37933 78047
rect 37933 78013 37967 78047
rect 37967 78013 37976 78047
rect 37924 78004 37976 78013
rect 16396 77936 16448 77988
rect 31760 77936 31812 77988
rect 32496 77868 32548 77920
rect 38200 77868 38252 77920
rect 19606 77766 19658 77818
rect 19670 77766 19722 77818
rect 19734 77766 19786 77818
rect 19798 77766 19850 77818
rect 33048 77324 33100 77376
rect 36268 77324 36320 77376
rect 4246 77222 4298 77274
rect 4310 77222 4362 77274
rect 4374 77222 4426 77274
rect 4438 77222 4490 77274
rect 34966 77222 35018 77274
rect 35030 77222 35082 77274
rect 35094 77222 35146 77274
rect 35158 77222 35210 77274
rect 1400 76959 1452 76968
rect 1400 76925 1409 76959
rect 1409 76925 1443 76959
rect 1443 76925 1452 76959
rect 1400 76916 1452 76925
rect 37280 76959 37332 76968
rect 37280 76925 37289 76959
rect 37289 76925 37323 76959
rect 37323 76925 37332 76959
rect 37280 76916 37332 76925
rect 38016 76916 38068 76968
rect 29920 76848 29972 76900
rect 30932 76848 30984 76900
rect 37648 76780 37700 76832
rect 37832 76780 37884 76832
rect 19606 76678 19658 76730
rect 19670 76678 19722 76730
rect 19734 76678 19786 76730
rect 19798 76678 19850 76730
rect 31024 76576 31076 76628
rect 23480 76551 23532 76560
rect 23480 76517 23489 76551
rect 23489 76517 23523 76551
rect 23523 76517 23532 76551
rect 23480 76508 23532 76517
rect 1400 76483 1452 76492
rect 1400 76449 1409 76483
rect 1409 76449 1443 76483
rect 1443 76449 1452 76483
rect 1400 76440 1452 76449
rect 23112 76440 23164 76492
rect 23848 76304 23900 76356
rect 4246 76134 4298 76186
rect 4310 76134 4362 76186
rect 4374 76134 4426 76186
rect 4438 76134 4490 76186
rect 34966 76134 35018 76186
rect 35030 76134 35082 76186
rect 35094 76134 35146 76186
rect 35158 76134 35210 76186
rect 33784 75964 33836 76016
rect 38384 75964 38436 76016
rect 35256 75896 35308 75948
rect 39212 75896 39264 75948
rect 20076 75871 20128 75880
rect 20076 75837 20085 75871
rect 20085 75837 20119 75871
rect 20119 75837 20128 75871
rect 20076 75828 20128 75837
rect 9036 75760 9088 75812
rect 20536 75828 20588 75880
rect 37280 75871 37332 75880
rect 37280 75837 37289 75871
rect 37289 75837 37323 75871
rect 37323 75837 37332 75871
rect 37280 75828 37332 75837
rect 37924 75871 37976 75880
rect 37924 75837 37933 75871
rect 37933 75837 37967 75871
rect 37967 75837 37976 75871
rect 37924 75828 37976 75837
rect 39764 75760 39816 75812
rect 38660 75692 38712 75744
rect 19606 75590 19658 75642
rect 19670 75590 19722 75642
rect 19734 75590 19786 75642
rect 19798 75590 19850 75642
rect 20444 75488 20496 75540
rect 21180 75531 21232 75540
rect 21180 75497 21189 75531
rect 21189 75497 21223 75531
rect 21223 75497 21232 75531
rect 21180 75488 21232 75497
rect 29552 75488 29604 75540
rect 1400 75395 1452 75404
rect 1400 75361 1409 75395
rect 1409 75361 1443 75395
rect 1443 75361 1452 75395
rect 1400 75352 1452 75361
rect 10324 75352 10376 75404
rect 23848 75420 23900 75472
rect 20996 75395 21048 75404
rect 20076 75284 20128 75336
rect 20996 75361 21005 75395
rect 21005 75361 21039 75395
rect 21039 75361 21048 75395
rect 20996 75352 21048 75361
rect 29644 75395 29696 75404
rect 29644 75361 29653 75395
rect 29653 75361 29687 75395
rect 29687 75361 29696 75395
rect 29644 75352 29696 75361
rect 29920 75395 29972 75404
rect 29920 75361 29929 75395
rect 29929 75361 29963 75395
rect 29963 75361 29972 75395
rect 29920 75352 29972 75361
rect 32036 75488 32088 75540
rect 34520 75488 34572 75540
rect 37188 75395 37240 75404
rect 37188 75361 37197 75395
rect 37197 75361 37231 75395
rect 37231 75361 37240 75395
rect 37188 75352 37240 75361
rect 35900 75284 35952 75336
rect 32312 75216 32364 75268
rect 32956 75216 33008 75268
rect 33876 75216 33928 75268
rect 38936 75216 38988 75268
rect 39396 75216 39448 75268
rect 39580 75216 39632 75268
rect 36268 75148 36320 75200
rect 4246 75046 4298 75098
rect 4310 75046 4362 75098
rect 4374 75046 4426 75098
rect 4438 75046 4490 75098
rect 34966 75046 35018 75098
rect 35030 75046 35082 75098
rect 35094 75046 35146 75098
rect 35158 75046 35210 75098
rect 39672 75080 39724 75132
rect 39304 75012 39356 75064
rect 20352 74987 20404 74996
rect 20352 74953 20361 74987
rect 20361 74953 20395 74987
rect 20395 74953 20404 74987
rect 20352 74944 20404 74953
rect 32956 74944 33008 74996
rect 36360 74944 36412 74996
rect 38292 74944 38344 74996
rect 39672 74944 39724 74996
rect 20076 74808 20128 74860
rect 1400 74783 1452 74792
rect 1400 74749 1409 74783
rect 1409 74749 1443 74783
rect 1443 74749 1452 74783
rect 1400 74740 1452 74749
rect 37280 74783 37332 74792
rect 14556 74672 14608 74724
rect 37280 74749 37289 74783
rect 37289 74749 37323 74783
rect 37323 74749 37332 74783
rect 37280 74740 37332 74749
rect 37924 74783 37976 74792
rect 37924 74749 37933 74783
rect 37933 74749 37967 74783
rect 37967 74749 37976 74783
rect 37924 74740 37976 74749
rect 35624 74604 35676 74656
rect 19606 74502 19658 74554
rect 19670 74502 19722 74554
rect 19734 74502 19786 74554
rect 19798 74502 19850 74554
rect 34060 74400 34112 74452
rect 38844 74400 38896 74452
rect 37188 74307 37240 74316
rect 37188 74273 37197 74307
rect 37197 74273 37231 74307
rect 37231 74273 37240 74307
rect 37188 74264 37240 74273
rect 38844 74060 38896 74112
rect 4246 73958 4298 74010
rect 4310 73958 4362 74010
rect 4374 73958 4426 74010
rect 4438 73958 4490 74010
rect 34966 73958 35018 74010
rect 35030 73958 35082 74010
rect 35094 73958 35146 74010
rect 35158 73958 35210 74010
rect 16120 73788 16172 73840
rect 25596 73788 25648 73840
rect 37096 73788 37148 73840
rect 1400 73695 1452 73704
rect 1400 73661 1409 73695
rect 1409 73661 1443 73695
rect 1443 73661 1452 73695
rect 1400 73652 1452 73661
rect 20168 73652 20220 73704
rect 23480 73652 23532 73704
rect 37280 73695 37332 73704
rect 37280 73661 37289 73695
rect 37289 73661 37323 73695
rect 37323 73661 37332 73695
rect 37280 73652 37332 73661
rect 37924 73695 37976 73704
rect 37924 73661 37933 73695
rect 37933 73661 37967 73695
rect 37967 73661 37976 73695
rect 37924 73652 37976 73661
rect 17316 73584 17368 73636
rect 17408 73516 17460 73568
rect 36176 73516 36228 73568
rect 19606 73414 19658 73466
rect 19670 73414 19722 73466
rect 19734 73414 19786 73466
rect 19798 73414 19850 73466
rect 1400 73219 1452 73228
rect 1400 73185 1409 73219
rect 1409 73185 1443 73219
rect 1443 73185 1452 73219
rect 1400 73176 1452 73185
rect 32404 73108 32456 73160
rect 34796 73108 34848 73160
rect 34336 73040 34388 73092
rect 37004 73040 37056 73092
rect 37740 72972 37792 73024
rect 37924 72972 37976 73024
rect 4246 72870 4298 72922
rect 4310 72870 4362 72922
rect 4374 72870 4426 72922
rect 4438 72870 4490 72922
rect 34966 72870 35018 72922
rect 35030 72870 35082 72922
rect 35094 72870 35146 72922
rect 35158 72870 35210 72922
rect 16120 72811 16172 72820
rect 16120 72777 16129 72811
rect 16129 72777 16163 72811
rect 16163 72777 16172 72811
rect 16120 72768 16172 72777
rect 16948 72811 17000 72820
rect 16948 72777 16957 72811
rect 16957 72777 16991 72811
rect 16991 72777 17000 72811
rect 16948 72768 17000 72777
rect 17868 72768 17920 72820
rect 17316 72700 17368 72752
rect 17408 72675 17460 72684
rect 17408 72641 17417 72675
rect 17417 72641 17451 72675
rect 17451 72641 17460 72675
rect 17408 72632 17460 72641
rect 15936 72607 15988 72616
rect 15936 72573 15945 72607
rect 15945 72573 15979 72607
rect 15979 72573 15988 72607
rect 15936 72564 15988 72573
rect 17040 72564 17092 72616
rect 16948 72496 17000 72548
rect 20168 72564 20220 72616
rect 37280 72607 37332 72616
rect 37280 72573 37289 72607
rect 37289 72573 37323 72607
rect 37323 72573 37332 72607
rect 37280 72564 37332 72573
rect 17224 72428 17276 72480
rect 36360 72428 36412 72480
rect 38384 72428 38436 72480
rect 19606 72326 19658 72378
rect 19670 72326 19722 72378
rect 19734 72326 19786 72378
rect 19798 72326 19850 72378
rect 16488 72224 16540 72276
rect 17684 72267 17736 72276
rect 17684 72233 17693 72267
rect 17693 72233 17727 72267
rect 17727 72233 17736 72267
rect 17684 72224 17736 72233
rect 1400 72131 1452 72140
rect 1400 72097 1409 72131
rect 1409 72097 1443 72131
rect 1443 72097 1452 72131
rect 1400 72088 1452 72097
rect 2228 72088 2280 72140
rect 8944 72088 8996 72140
rect 17408 72131 17460 72140
rect 17408 72097 17417 72131
rect 17417 72097 17451 72131
rect 17451 72097 17460 72131
rect 17408 72088 17460 72097
rect 37188 72131 37240 72140
rect 37188 72097 37197 72131
rect 37197 72097 37231 72131
rect 37231 72097 37240 72131
rect 37188 72088 37240 72097
rect 16580 72020 16632 72072
rect 36912 71884 36964 71936
rect 4246 71782 4298 71834
rect 4310 71782 4362 71834
rect 4374 71782 4426 71834
rect 4438 71782 4490 71834
rect 34966 71782 35018 71834
rect 35030 71782 35082 71834
rect 35094 71782 35146 71834
rect 35158 71782 35210 71834
rect 38936 71791 38988 71800
rect 38936 71757 38945 71791
rect 38945 71757 38979 71791
rect 38979 71757 38988 71791
rect 38936 71748 38988 71757
rect 16856 71680 16908 71732
rect 17132 71680 17184 71732
rect 17776 71723 17828 71732
rect 17776 71689 17785 71723
rect 17785 71689 17819 71723
rect 17819 71689 17828 71723
rect 17776 71680 17828 71689
rect 35900 71723 35952 71732
rect 35900 71689 35909 71723
rect 35909 71689 35943 71723
rect 35943 71689 35952 71723
rect 35900 71680 35952 71689
rect 16028 71612 16080 71664
rect 16580 71587 16632 71596
rect 16580 71553 16589 71587
rect 16589 71553 16623 71587
rect 16623 71553 16632 71587
rect 16580 71544 16632 71553
rect 1400 71519 1452 71528
rect 1400 71485 1409 71519
rect 1409 71485 1443 71519
rect 1443 71485 1452 71519
rect 1400 71476 1452 71485
rect 15292 71476 15344 71528
rect 17868 71612 17920 71664
rect 30840 71612 30892 71664
rect 31024 71612 31076 71664
rect 32128 71612 32180 71664
rect 16856 71544 16908 71596
rect 17316 71544 17368 71596
rect 15752 71408 15804 71460
rect 26608 71544 26660 71596
rect 31392 71544 31444 71596
rect 31760 71544 31812 71596
rect 32496 71544 32548 71596
rect 37556 71544 37608 71596
rect 32128 71519 32180 71528
rect 17408 71340 17460 71392
rect 30840 71408 30892 71460
rect 31208 71340 31260 71392
rect 32128 71485 32137 71519
rect 32137 71485 32171 71519
rect 32171 71485 32180 71519
rect 32128 71476 32180 71485
rect 32404 71519 32456 71528
rect 32404 71485 32413 71519
rect 32413 71485 32447 71519
rect 32447 71485 32456 71519
rect 32404 71476 32456 71485
rect 35992 71476 36044 71528
rect 36452 71476 36504 71528
rect 37464 71519 37516 71528
rect 37464 71485 37473 71519
rect 37473 71485 37507 71519
rect 37507 71485 37516 71519
rect 37464 71476 37516 71485
rect 38108 71519 38160 71528
rect 38108 71485 38117 71519
rect 38117 71485 38151 71519
rect 38151 71485 38160 71519
rect 38108 71476 38160 71485
rect 38844 71476 38896 71528
rect 37280 71383 37332 71392
rect 37280 71349 37289 71383
rect 37289 71349 37323 71383
rect 37323 71349 37332 71383
rect 37280 71340 37332 71349
rect 37556 71340 37608 71392
rect 19606 71238 19658 71290
rect 19670 71238 19722 71290
rect 19734 71238 19786 71290
rect 19798 71238 19850 71290
rect 15568 71179 15620 71188
rect 15568 71145 15577 71179
rect 15577 71145 15611 71179
rect 15611 71145 15620 71179
rect 15568 71136 15620 71145
rect 16396 71179 16448 71188
rect 16396 71145 16405 71179
rect 16405 71145 16439 71179
rect 16439 71145 16448 71179
rect 16396 71136 16448 71145
rect 16764 71136 16816 71188
rect 31208 71136 31260 71188
rect 3424 71068 3476 71120
rect 2504 71000 2556 71052
rect 30748 71000 30800 71052
rect 31392 71043 31444 71052
rect 31392 71009 31401 71043
rect 31401 71009 31435 71043
rect 31435 71009 31444 71043
rect 31392 71000 31444 71009
rect 32128 71068 32180 71120
rect 32404 71068 32456 71120
rect 32036 71043 32088 71052
rect 15476 70932 15528 70984
rect 16580 70932 16632 70984
rect 16856 70932 16908 70984
rect 17776 70932 17828 70984
rect 32036 71009 32045 71043
rect 32045 71009 32079 71043
rect 32079 71009 32088 71043
rect 32036 71000 32088 71009
rect 37372 71043 37424 71052
rect 37372 71009 37381 71043
rect 37381 71009 37415 71043
rect 37415 71009 37424 71043
rect 37372 71000 37424 71009
rect 32128 70932 32180 70984
rect 32956 70932 33008 70984
rect 32036 70864 32088 70916
rect 33048 70864 33100 70916
rect 15476 70796 15528 70848
rect 17224 70796 17276 70848
rect 22836 70796 22888 70848
rect 37096 70796 37148 70848
rect 4246 70694 4298 70746
rect 4310 70694 4362 70746
rect 4374 70694 4426 70746
rect 4438 70694 4490 70746
rect 34966 70694 35018 70746
rect 35030 70694 35082 70746
rect 35094 70694 35146 70746
rect 35158 70694 35210 70746
rect 2136 70592 2188 70644
rect 15844 70635 15896 70644
rect 15844 70601 15853 70635
rect 15853 70601 15887 70635
rect 15887 70601 15896 70635
rect 15844 70592 15896 70601
rect 16672 70635 16724 70644
rect 16672 70601 16681 70635
rect 16681 70601 16715 70635
rect 16715 70601 16724 70635
rect 16672 70592 16724 70601
rect 17500 70635 17552 70644
rect 17500 70601 17509 70635
rect 17509 70601 17543 70635
rect 17543 70601 17552 70635
rect 17500 70592 17552 70601
rect 6276 70456 6328 70508
rect 1400 70431 1452 70440
rect 1400 70397 1409 70431
rect 1409 70397 1443 70431
rect 1443 70397 1452 70431
rect 1400 70388 1452 70397
rect 14464 70388 14516 70440
rect 15476 70431 15528 70440
rect 15476 70397 15485 70431
rect 15485 70397 15519 70431
rect 15519 70397 15528 70431
rect 15476 70388 15528 70397
rect 16396 70456 16448 70508
rect 31392 70524 31444 70576
rect 31760 70524 31812 70576
rect 37832 70524 37884 70576
rect 38016 70524 38068 70576
rect 17224 70431 17276 70440
rect 17224 70397 17233 70431
rect 17233 70397 17267 70431
rect 17267 70397 17276 70431
rect 17224 70388 17276 70397
rect 26608 70388 26660 70440
rect 31392 70431 31444 70440
rect 26332 70320 26384 70372
rect 31392 70397 31401 70431
rect 31401 70397 31435 70431
rect 31435 70397 31444 70431
rect 31392 70388 31444 70397
rect 31668 70431 31720 70440
rect 31668 70397 31677 70431
rect 31677 70397 31711 70431
rect 31711 70397 31720 70431
rect 31668 70388 31720 70397
rect 32036 70431 32088 70440
rect 32036 70397 32045 70431
rect 32045 70397 32079 70431
rect 32079 70397 32088 70431
rect 32036 70388 32088 70397
rect 32404 70388 32456 70440
rect 37464 70431 37516 70440
rect 37464 70397 37473 70431
rect 37473 70397 37507 70431
rect 37507 70397 37516 70431
rect 37464 70388 37516 70397
rect 38292 70388 38344 70440
rect 37740 70320 37792 70372
rect 38660 70320 38712 70372
rect 37924 70252 37976 70304
rect 19606 70150 19658 70202
rect 19670 70150 19722 70202
rect 19734 70150 19786 70202
rect 19798 70150 19850 70202
rect 39304 70363 39356 70372
rect 39304 70329 39313 70363
rect 39313 70329 39347 70363
rect 39347 70329 39356 70363
rect 39304 70320 39356 70329
rect 39120 70116 39172 70168
rect 16212 70048 16264 70100
rect 37372 70048 37424 70100
rect 37648 70048 37700 70100
rect 1400 69955 1452 69964
rect 1400 69921 1409 69955
rect 1409 69921 1443 69955
rect 1443 69921 1452 69955
rect 1400 69912 1452 69921
rect 6368 69912 6420 69964
rect 36728 69955 36780 69964
rect 36728 69921 36737 69955
rect 36737 69921 36771 69955
rect 36771 69921 36780 69955
rect 36728 69912 36780 69921
rect 37372 69955 37424 69964
rect 37372 69921 37381 69955
rect 37381 69921 37415 69955
rect 37415 69921 37424 69955
rect 37372 69912 37424 69921
rect 15476 69844 15528 69896
rect 16120 69844 16172 69896
rect 37004 69776 37056 69828
rect 36912 69708 36964 69760
rect 39764 69683 39816 69692
rect 4246 69606 4298 69658
rect 4310 69606 4362 69658
rect 4374 69606 4426 69658
rect 4438 69606 4490 69658
rect 34966 69606 35018 69658
rect 35030 69606 35082 69658
rect 35094 69606 35146 69658
rect 35158 69606 35210 69658
rect 39764 69649 39773 69683
rect 39773 69649 39807 69683
rect 39807 69649 39816 69683
rect 39764 69640 39816 69649
rect 16304 69504 16356 69556
rect 38200 69504 38252 69556
rect 39764 69504 39816 69556
rect 32404 69436 32456 69488
rect 38384 69436 38436 69488
rect 16120 69411 16172 69420
rect 16120 69377 16129 69411
rect 16129 69377 16163 69411
rect 16163 69377 16172 69411
rect 16120 69368 16172 69377
rect 38200 69368 38252 69420
rect 2044 69300 2096 69352
rect 36636 69343 36688 69352
rect 36636 69309 36645 69343
rect 36645 69309 36679 69343
rect 36679 69309 36688 69343
rect 36636 69300 36688 69309
rect 37280 69300 37332 69352
rect 38384 69300 38436 69352
rect 35900 69232 35952 69284
rect 36728 69232 36780 69284
rect 33968 69164 34020 69216
rect 35348 69164 35400 69216
rect 37280 69164 37332 69216
rect 38016 69164 38068 69216
rect 39212 69207 39264 69216
rect 39212 69173 39221 69207
rect 39221 69173 39255 69207
rect 39255 69173 39264 69207
rect 39212 69164 39264 69173
rect 19606 69062 19658 69114
rect 19670 69062 19722 69114
rect 19734 69062 19786 69114
rect 19798 69062 19850 69114
rect 36728 68960 36780 69012
rect 36084 68892 36136 68944
rect 1400 68867 1452 68876
rect 1400 68833 1409 68867
rect 1409 68833 1443 68867
rect 1443 68833 1452 68867
rect 1400 68824 1452 68833
rect 35808 68824 35860 68876
rect 37280 68892 37332 68944
rect 37096 68867 37148 68876
rect 37096 68833 37105 68867
rect 37105 68833 37139 68867
rect 37139 68833 37148 68867
rect 37096 68824 37148 68833
rect 37188 68688 37240 68740
rect 34520 68620 34572 68672
rect 4246 68518 4298 68570
rect 4310 68518 4362 68570
rect 4374 68518 4426 68570
rect 4438 68518 4490 68570
rect 34966 68518 35018 68570
rect 35030 68518 35082 68570
rect 35094 68518 35146 68570
rect 35158 68518 35210 68570
rect 36268 68416 36320 68468
rect 36452 68416 36504 68468
rect 37372 68416 37424 68468
rect 30104 68348 30156 68400
rect 34520 68348 34572 68400
rect 36728 68348 36780 68400
rect 36176 68280 36228 68332
rect 36636 68280 36688 68332
rect 1400 68255 1452 68264
rect 1400 68221 1409 68255
rect 1409 68221 1443 68255
rect 1443 68221 1452 68255
rect 1400 68212 1452 68221
rect 36268 68255 36320 68264
rect 1584 68144 1636 68196
rect 36268 68221 36277 68255
rect 36277 68221 36311 68255
rect 36311 68221 36320 68255
rect 36268 68212 36320 68221
rect 36820 68212 36872 68264
rect 37372 68280 37424 68332
rect 37924 68280 37976 68332
rect 37556 68212 37608 68264
rect 38200 68212 38252 68264
rect 33048 68144 33100 68196
rect 32956 68076 33008 68128
rect 37280 68144 37332 68196
rect 36176 68076 36228 68128
rect 37924 68119 37976 68128
rect 37924 68085 37933 68119
rect 37933 68085 37967 68119
rect 37967 68085 37976 68119
rect 37924 68076 37976 68085
rect 19606 67974 19658 68026
rect 19670 67974 19722 68026
rect 19734 67974 19786 68026
rect 19798 67974 19850 68026
rect 27528 67872 27580 67924
rect 35348 67872 35400 67924
rect 36728 67872 36780 67924
rect 36820 67872 36872 67924
rect 37648 67872 37700 67924
rect 29920 67804 29972 67856
rect 35900 67736 35952 67788
rect 37280 67804 37332 67856
rect 36728 67779 36780 67788
rect 36728 67745 36737 67779
rect 36737 67745 36771 67779
rect 36771 67745 36780 67779
rect 36728 67736 36780 67745
rect 37096 67779 37148 67788
rect 37096 67745 37105 67779
rect 37105 67745 37139 67779
rect 37139 67745 37148 67779
rect 37096 67736 37148 67745
rect 35716 67600 35768 67652
rect 30196 67532 30248 67584
rect 36084 67532 36136 67584
rect 36636 67532 36688 67584
rect 39212 67532 39264 67584
rect 4246 67430 4298 67482
rect 4310 67430 4362 67482
rect 4374 67430 4426 67482
rect 4438 67430 4490 67482
rect 34966 67430 35018 67482
rect 35030 67430 35082 67482
rect 35094 67430 35146 67482
rect 35158 67430 35210 67482
rect 36084 67328 36136 67380
rect 31208 67260 31260 67312
rect 1400 67167 1452 67176
rect 1400 67133 1409 67167
rect 1409 67133 1443 67167
rect 1443 67133 1452 67167
rect 1400 67124 1452 67133
rect 33048 67124 33100 67176
rect 35992 67124 36044 67176
rect 36544 67167 36596 67176
rect 36544 67133 36553 67167
rect 36553 67133 36587 67167
rect 36587 67133 36596 67167
rect 36544 67124 36596 67133
rect 36912 67167 36964 67176
rect 36912 67133 36921 67167
rect 36921 67133 36955 67167
rect 36955 67133 36964 67167
rect 36912 67124 36964 67133
rect 34152 67056 34204 67108
rect 36728 67099 36780 67108
rect 36728 67065 36737 67099
rect 36737 67065 36771 67099
rect 36771 67065 36780 67099
rect 36728 67056 36780 67065
rect 37096 67056 37148 67108
rect 36084 67031 36136 67040
rect 36084 66997 36093 67031
rect 36093 66997 36127 67031
rect 36127 66997 36136 67031
rect 36084 66988 36136 66997
rect 39580 67260 39632 67312
rect 37832 67192 37884 67244
rect 38384 67124 38436 67176
rect 39580 67124 39632 67176
rect 37648 67056 37700 67108
rect 19606 66886 19658 66938
rect 19670 66886 19722 66938
rect 19734 66886 19786 66938
rect 19798 66886 19850 66938
rect 1400 66691 1452 66700
rect 1400 66657 1409 66691
rect 1409 66657 1443 66691
rect 1443 66657 1452 66691
rect 1400 66648 1452 66657
rect 34796 66648 34848 66700
rect 35348 66691 35400 66700
rect 35348 66657 35357 66691
rect 35357 66657 35391 66691
rect 35391 66657 35400 66691
rect 35348 66648 35400 66657
rect 36636 66784 36688 66836
rect 36912 66784 36964 66836
rect 38844 66784 38896 66836
rect 36728 66716 36780 66768
rect 37280 66716 37332 66768
rect 37648 66716 37700 66768
rect 36176 66691 36228 66700
rect 36176 66657 36185 66691
rect 36185 66657 36219 66691
rect 36219 66657 36228 66691
rect 36176 66648 36228 66657
rect 36912 66648 36964 66700
rect 37096 66691 37148 66700
rect 37096 66657 37105 66691
rect 37105 66657 37139 66691
rect 37139 66657 37148 66691
rect 37096 66648 37148 66657
rect 37188 66691 37240 66700
rect 37188 66657 37197 66691
rect 37197 66657 37231 66691
rect 37231 66657 37240 66691
rect 37188 66648 37240 66657
rect 36268 66580 36320 66632
rect 31392 66512 31444 66564
rect 34520 66487 34572 66496
rect 34520 66453 34529 66487
rect 34529 66453 34563 66487
rect 34563 66453 34572 66487
rect 34520 66444 34572 66453
rect 36912 66444 36964 66496
rect 37832 66444 37884 66496
rect 4246 66342 4298 66394
rect 4310 66342 4362 66394
rect 4374 66342 4426 66394
rect 4438 66342 4490 66394
rect 34966 66342 35018 66394
rect 35030 66342 35082 66394
rect 35094 66342 35146 66394
rect 35158 66342 35210 66394
rect 1400 66079 1452 66088
rect 1400 66045 1409 66079
rect 1409 66045 1443 66079
rect 1443 66045 1452 66079
rect 1400 66036 1452 66045
rect 30288 65968 30340 66020
rect 33048 66036 33100 66088
rect 35992 66036 36044 66088
rect 39028 66104 39080 66156
rect 38108 66036 38160 66088
rect 33600 65968 33652 66020
rect 35808 65968 35860 66020
rect 37280 65968 37332 66020
rect 36636 65900 36688 65952
rect 37096 65900 37148 65952
rect 19606 65798 19658 65850
rect 19670 65798 19722 65850
rect 19734 65798 19786 65850
rect 19798 65798 19850 65850
rect 34428 65696 34480 65748
rect 38844 65696 38896 65748
rect 34520 65628 34572 65680
rect 31760 65560 31812 65612
rect 32772 65560 32824 65612
rect 32864 65560 32916 65612
rect 33048 65560 33100 65612
rect 35072 65603 35124 65612
rect 35072 65569 35081 65603
rect 35081 65569 35115 65603
rect 35115 65569 35124 65603
rect 35072 65560 35124 65569
rect 35716 65603 35768 65612
rect 35716 65569 35725 65603
rect 35725 65569 35759 65603
rect 35759 65569 35768 65603
rect 35716 65560 35768 65569
rect 36452 65560 36504 65612
rect 32036 65492 32088 65544
rect 32680 65492 32732 65544
rect 33324 65492 33376 65544
rect 35532 65492 35584 65544
rect 33140 65424 33192 65476
rect 34428 65424 34480 65476
rect 36728 65492 36780 65544
rect 37096 65603 37148 65612
rect 37096 65569 37105 65603
rect 37105 65569 37139 65603
rect 37139 65569 37148 65603
rect 37648 65628 37700 65680
rect 39396 65628 39448 65680
rect 37096 65560 37148 65569
rect 38568 65424 38620 65476
rect 32864 65356 32916 65408
rect 34796 65356 34848 65408
rect 35440 65356 35492 65408
rect 35532 65399 35584 65408
rect 35532 65365 35541 65399
rect 35541 65365 35575 65399
rect 35575 65365 35584 65399
rect 36176 65399 36228 65408
rect 35532 65356 35584 65365
rect 36176 65365 36185 65399
rect 36185 65365 36219 65399
rect 36219 65365 36228 65399
rect 36176 65356 36228 65365
rect 39028 65356 39080 65408
rect 4246 65254 4298 65306
rect 4310 65254 4362 65306
rect 4374 65254 4426 65306
rect 4438 65254 4490 65306
rect 34966 65254 35018 65306
rect 35030 65254 35082 65306
rect 35094 65254 35146 65306
rect 35158 65254 35210 65306
rect 34520 65152 34572 65204
rect 37188 65152 37240 65204
rect 26148 65016 26200 65068
rect 34612 65016 34664 65068
rect 35164 65016 35216 65068
rect 39672 65152 39724 65204
rect 39396 65084 39448 65136
rect 1400 64991 1452 65000
rect 1400 64957 1409 64991
rect 1409 64957 1443 64991
rect 1443 64957 1452 64991
rect 1400 64948 1452 64957
rect 33048 64948 33100 65000
rect 34796 64991 34848 65000
rect 34796 64957 34805 64991
rect 34805 64957 34839 64991
rect 34839 64957 34848 64991
rect 34796 64948 34848 64957
rect 35992 64948 36044 65000
rect 36912 64991 36964 65000
rect 36912 64957 36921 64991
rect 36921 64957 36955 64991
rect 36955 64957 36964 64991
rect 39948 65016 40000 65068
rect 36912 64948 36964 64957
rect 38016 64948 38068 65000
rect 32404 64880 32456 64932
rect 32956 64880 33008 64932
rect 36728 64923 36780 64932
rect 36728 64889 36737 64923
rect 36737 64889 36771 64923
rect 36771 64889 36780 64923
rect 36728 64880 36780 64889
rect 37096 64880 37148 64932
rect 34612 64855 34664 64864
rect 34612 64821 34621 64855
rect 34621 64821 34655 64855
rect 34655 64821 34664 64855
rect 34612 64812 34664 64821
rect 34796 64812 34848 64864
rect 35348 64812 35400 64864
rect 37464 64812 37516 64864
rect 19606 64710 19658 64762
rect 19670 64710 19722 64762
rect 19734 64710 19786 64762
rect 19798 64710 19850 64762
rect 36268 64608 36320 64660
rect 20168 64583 20220 64592
rect 20168 64549 20177 64583
rect 20177 64549 20211 64583
rect 20211 64549 20220 64583
rect 20168 64540 20220 64549
rect 32496 64540 32548 64592
rect 35072 64540 35124 64592
rect 1400 64515 1452 64524
rect 1400 64481 1409 64515
rect 1409 64481 1443 64515
rect 1443 64481 1452 64515
rect 1400 64472 1452 64481
rect 31024 64472 31076 64524
rect 31668 64515 31720 64524
rect 31668 64481 31677 64515
rect 31677 64481 31711 64515
rect 31711 64481 31720 64515
rect 31668 64472 31720 64481
rect 34152 64472 34204 64524
rect 3148 64336 3200 64388
rect 29000 64336 29052 64388
rect 34152 64336 34204 64388
rect 34888 64472 34940 64524
rect 35348 64404 35400 64456
rect 35716 64336 35768 64388
rect 36728 64540 36780 64592
rect 37096 64583 37148 64592
rect 37096 64549 37105 64583
rect 37105 64549 37139 64583
rect 37139 64549 37148 64583
rect 37096 64540 37148 64549
rect 37464 64540 37516 64592
rect 35992 64515 36044 64524
rect 35992 64481 36001 64515
rect 36001 64481 36035 64515
rect 36035 64481 36044 64515
rect 35992 64472 36044 64481
rect 17316 64268 17368 64320
rect 33140 64268 33192 64320
rect 36912 64472 36964 64524
rect 37556 64472 37608 64524
rect 36268 64404 36320 64456
rect 37648 64404 37700 64456
rect 36360 64311 36412 64320
rect 36360 64277 36369 64311
rect 36369 64277 36403 64311
rect 36403 64277 36412 64311
rect 36360 64268 36412 64277
rect 38568 64268 38620 64320
rect 4246 64166 4298 64218
rect 4310 64166 4362 64218
rect 4374 64166 4426 64218
rect 4438 64166 4490 64218
rect 34966 64166 35018 64218
rect 35030 64166 35082 64218
rect 35094 64166 35146 64218
rect 35158 64166 35210 64218
rect 37280 64064 37332 64116
rect 37556 64064 37608 64116
rect 39856 64064 39908 64116
rect 34796 63903 34848 63912
rect 34796 63869 34805 63903
rect 34805 63869 34839 63903
rect 34839 63869 34848 63903
rect 34796 63860 34848 63869
rect 34980 63860 35032 63912
rect 35348 63860 35400 63912
rect 35808 63860 35860 63912
rect 39488 63928 39540 63980
rect 36912 63903 36964 63912
rect 36912 63869 36921 63903
rect 36921 63869 36955 63903
rect 36955 63869 36964 63903
rect 36912 63860 36964 63869
rect 37556 63903 37608 63912
rect 37556 63869 37565 63903
rect 37565 63869 37599 63903
rect 37599 63869 37608 63903
rect 37556 63860 37608 63869
rect 37648 63860 37700 63912
rect 37924 63903 37976 63912
rect 37924 63869 37933 63903
rect 37933 63869 37967 63903
rect 37967 63869 37976 63903
rect 37924 63860 37976 63869
rect 35992 63792 36044 63844
rect 34612 63767 34664 63776
rect 34612 63733 34621 63767
rect 34621 63733 34655 63767
rect 34655 63733 34664 63767
rect 34612 63724 34664 63733
rect 35716 63724 35768 63776
rect 37464 63792 37516 63844
rect 38844 63792 38896 63844
rect 37096 63767 37148 63776
rect 37096 63733 37105 63767
rect 37105 63733 37139 63767
rect 37139 63733 37148 63767
rect 37096 63724 37148 63733
rect 38108 63767 38160 63776
rect 38108 63733 38117 63767
rect 38117 63733 38151 63767
rect 38151 63733 38160 63767
rect 38108 63724 38160 63733
rect 19606 63622 19658 63674
rect 19670 63622 19722 63674
rect 19734 63622 19786 63674
rect 19798 63622 19850 63674
rect 38936 63588 38988 63640
rect 35808 63520 35860 63572
rect 35992 63520 36044 63572
rect 36452 63520 36504 63572
rect 1400 63427 1452 63436
rect 1400 63393 1409 63427
rect 1409 63393 1443 63427
rect 1443 63393 1452 63427
rect 1400 63384 1452 63393
rect 34980 63384 35032 63436
rect 35164 63427 35216 63436
rect 35164 63393 35173 63427
rect 35173 63393 35207 63427
rect 35207 63393 35216 63427
rect 35164 63384 35216 63393
rect 35532 63384 35584 63436
rect 35808 63427 35860 63436
rect 35808 63393 35817 63427
rect 35817 63393 35851 63427
rect 35851 63393 35860 63427
rect 35808 63384 35860 63393
rect 36176 63427 36228 63436
rect 36176 63393 36185 63427
rect 36185 63393 36219 63427
rect 36219 63393 36228 63427
rect 36176 63384 36228 63393
rect 35716 63316 35768 63368
rect 36728 63452 36780 63504
rect 37556 63452 37608 63504
rect 38384 63452 38436 63504
rect 37280 63384 37332 63436
rect 38752 63316 38804 63368
rect 37464 63248 37516 63300
rect 35808 63180 35860 63232
rect 38292 63180 38344 63232
rect 4246 63078 4298 63130
rect 4310 63078 4362 63130
rect 4374 63078 4426 63130
rect 4438 63078 4490 63130
rect 34966 63078 35018 63130
rect 35030 63078 35082 63130
rect 35094 63078 35146 63130
rect 35158 63078 35210 63130
rect 36544 62976 36596 63028
rect 36912 62976 36964 63028
rect 37280 62908 37332 62960
rect 32496 62840 32548 62892
rect 1400 62815 1452 62824
rect 1400 62781 1409 62815
rect 1409 62781 1443 62815
rect 1443 62781 1452 62815
rect 1400 62772 1452 62781
rect 31668 62772 31720 62824
rect 34612 62840 34664 62892
rect 36084 62815 36136 62824
rect 36084 62781 36093 62815
rect 36093 62781 36127 62815
rect 36127 62781 36136 62815
rect 36084 62772 36136 62781
rect 36636 62840 36688 62892
rect 37556 62908 37608 62960
rect 38752 62908 38804 62960
rect 32496 62704 32548 62756
rect 33600 62704 33652 62756
rect 36728 62704 36780 62756
rect 36452 62636 36504 62688
rect 36636 62679 36688 62688
rect 36636 62645 36645 62679
rect 36645 62645 36679 62679
rect 36679 62645 36688 62679
rect 36636 62636 36688 62645
rect 37464 62815 37516 62824
rect 37464 62781 37478 62815
rect 37478 62781 37512 62815
rect 37512 62781 37516 62815
rect 37464 62772 37516 62781
rect 37648 62636 37700 62688
rect 19606 62534 19658 62586
rect 19670 62534 19722 62586
rect 19734 62534 19786 62586
rect 19798 62534 19850 62586
rect 37464 62432 37516 62484
rect 36544 62364 36596 62416
rect 37280 62364 37332 62416
rect 15384 62339 15436 62348
rect 15384 62305 15393 62339
rect 15393 62305 15427 62339
rect 15427 62305 15436 62339
rect 15384 62296 15436 62305
rect 35716 62296 35768 62348
rect 36268 62339 36320 62348
rect 36268 62305 36277 62339
rect 36277 62305 36311 62339
rect 36311 62305 36320 62339
rect 36268 62296 36320 62305
rect 36728 62160 36780 62212
rect 37464 62296 37516 62348
rect 37556 62228 37608 62280
rect 39120 62160 39172 62212
rect 3700 62092 3752 62144
rect 36176 62092 36228 62144
rect 4246 61990 4298 62042
rect 4310 61990 4362 62042
rect 4374 61990 4426 62042
rect 4438 61990 4490 62042
rect 34966 61990 35018 62042
rect 35030 61990 35082 62042
rect 35094 61990 35146 62042
rect 35158 61990 35210 62042
rect 37464 61820 37516 61872
rect 37740 61820 37792 61872
rect 37372 61752 37424 61804
rect 1400 61727 1452 61736
rect 1400 61693 1409 61727
rect 1409 61693 1443 61727
rect 1443 61693 1452 61727
rect 1400 61684 1452 61693
rect 35808 61684 35860 61736
rect 36728 61684 36780 61736
rect 35532 61616 35584 61668
rect 36544 61616 36596 61668
rect 37280 61659 37332 61668
rect 37280 61625 37289 61659
rect 37289 61625 37323 61659
rect 37323 61625 37332 61659
rect 37280 61616 37332 61625
rect 37556 61616 37608 61668
rect 19606 61446 19658 61498
rect 19670 61446 19722 61498
rect 19734 61446 19786 61498
rect 19798 61446 19850 61498
rect 35440 61344 35492 61396
rect 1400 61251 1452 61260
rect 1400 61217 1409 61251
rect 1409 61217 1443 61251
rect 1443 61217 1452 61251
rect 1400 61208 1452 61217
rect 34888 61251 34940 61260
rect 34888 61217 34897 61251
rect 34897 61217 34931 61251
rect 34931 61217 34940 61251
rect 34888 61208 34940 61217
rect 35532 61251 35584 61260
rect 35532 61217 35541 61251
rect 35541 61217 35575 61251
rect 35575 61217 35584 61251
rect 35532 61208 35584 61217
rect 36268 61208 36320 61260
rect 36728 61251 36780 61260
rect 36728 61217 36737 61251
rect 36737 61217 36771 61251
rect 36771 61217 36780 61251
rect 36728 61208 36780 61217
rect 37556 61344 37608 61396
rect 37280 61276 37332 61328
rect 33048 61004 33100 61056
rect 35348 61047 35400 61056
rect 35348 61013 35357 61047
rect 35357 61013 35391 61047
rect 35391 61013 35400 61047
rect 35348 61004 35400 61013
rect 36728 61004 36780 61056
rect 39580 61004 39632 61056
rect 4246 60902 4298 60954
rect 4310 60902 4362 60954
rect 4374 60902 4426 60954
rect 4438 60902 4490 60954
rect 34966 60902 35018 60954
rect 35030 60902 35082 60954
rect 35094 60902 35146 60954
rect 35158 60902 35210 60954
rect 28540 60732 28592 60784
rect 34888 60732 34940 60784
rect 35164 60732 35216 60784
rect 35532 60732 35584 60784
rect 32680 60664 32732 60716
rect 35256 60596 35308 60648
rect 35532 60596 35584 60648
rect 35992 60639 36044 60648
rect 35992 60605 36001 60639
rect 36001 60605 36035 60639
rect 36035 60605 36044 60639
rect 35992 60596 36044 60605
rect 36544 60664 36596 60716
rect 36728 60664 36780 60716
rect 36452 60639 36504 60648
rect 36452 60605 36455 60639
rect 36455 60605 36504 60639
rect 36452 60596 36504 60605
rect 36912 60596 36964 60648
rect 37280 60639 37332 60648
rect 37280 60605 37289 60639
rect 37289 60605 37323 60639
rect 37323 60605 37332 60639
rect 37280 60596 37332 60605
rect 37464 60639 37516 60648
rect 37464 60605 37478 60639
rect 37478 60605 37512 60639
rect 37512 60605 37516 60639
rect 37464 60596 37516 60605
rect 35440 60528 35492 60580
rect 37556 60528 37608 60580
rect 36544 60503 36596 60512
rect 36544 60469 36561 60503
rect 36561 60469 36595 60503
rect 36595 60469 36596 60503
rect 36544 60460 36596 60469
rect 19606 60358 19658 60410
rect 19670 60358 19722 60410
rect 19734 60358 19786 60410
rect 19798 60358 19850 60410
rect 33140 60256 33192 60308
rect 35348 60256 35400 60308
rect 34520 60188 34572 60240
rect 37372 60188 37424 60240
rect 1400 60163 1452 60172
rect 1400 60129 1409 60163
rect 1409 60129 1443 60163
rect 1443 60129 1452 60163
rect 1400 60120 1452 60129
rect 16580 60120 16632 60172
rect 34060 60120 34112 60172
rect 35164 60163 35216 60172
rect 35164 60129 35173 60163
rect 35173 60129 35207 60163
rect 35207 60129 35216 60163
rect 35164 60120 35216 60129
rect 35624 60163 35676 60172
rect 35624 60129 35633 60163
rect 35633 60129 35667 60163
rect 35667 60129 35676 60163
rect 35624 60120 35676 60129
rect 34152 60052 34204 60104
rect 35992 60163 36044 60172
rect 35992 60129 36006 60163
rect 36006 60129 36040 60163
rect 36040 60129 36044 60163
rect 35992 60120 36044 60129
rect 33784 59984 33836 60036
rect 34520 59984 34572 60036
rect 34888 59984 34940 60036
rect 35348 59984 35400 60036
rect 31668 59916 31720 59968
rect 35808 59916 35860 59968
rect 37280 60052 37332 60104
rect 39304 59984 39356 60036
rect 37188 59916 37240 59968
rect 38660 59916 38712 59968
rect 4246 59814 4298 59866
rect 4310 59814 4362 59866
rect 4374 59814 4426 59866
rect 4438 59814 4490 59866
rect 34966 59814 35018 59866
rect 35030 59814 35082 59866
rect 35094 59814 35146 59866
rect 35158 59814 35210 59866
rect 25688 59576 25740 59628
rect 33140 59576 33192 59628
rect 33600 59712 33652 59764
rect 33876 59712 33928 59764
rect 35992 59712 36044 59764
rect 33324 59644 33376 59696
rect 1400 59551 1452 59560
rect 1400 59517 1409 59551
rect 1409 59517 1443 59551
rect 1443 59517 1452 59551
rect 1400 59508 1452 59517
rect 31760 59508 31812 59560
rect 35624 59644 35676 59696
rect 38384 59644 38436 59696
rect 35808 59576 35860 59628
rect 34796 59551 34848 59560
rect 30748 59440 30800 59492
rect 34796 59517 34805 59551
rect 34805 59517 34839 59551
rect 34839 59517 34848 59551
rect 34796 59508 34848 59517
rect 36084 59508 36136 59560
rect 36728 59508 36780 59560
rect 34152 59440 34204 59492
rect 35440 59440 35492 59492
rect 36912 59440 36964 59492
rect 33600 59372 33652 59424
rect 37188 59440 37240 59492
rect 37372 59483 37424 59492
rect 37372 59449 37381 59483
rect 37381 59449 37415 59483
rect 37415 59449 37424 59483
rect 37372 59440 37424 59449
rect 38844 59372 38896 59424
rect 19606 59270 19658 59322
rect 19670 59270 19722 59322
rect 19734 59270 19786 59322
rect 19798 59270 19850 59322
rect 29644 59168 29696 59220
rect 30104 59168 30156 59220
rect 34152 59168 34204 59220
rect 33140 59100 33192 59152
rect 36728 59168 36780 59220
rect 37188 59168 37240 59220
rect 37372 59100 37424 59152
rect 25596 58964 25648 59016
rect 31484 59075 31536 59084
rect 31484 59041 31494 59075
rect 31494 59041 31528 59075
rect 31528 59041 31536 59075
rect 31484 59032 31536 59041
rect 31944 59032 31996 59084
rect 33600 59075 33652 59084
rect 33600 59041 33609 59075
rect 33609 59041 33643 59075
rect 33643 59041 33652 59075
rect 33600 59032 33652 59041
rect 34152 59075 34204 59084
rect 33784 58964 33836 59016
rect 30104 58896 30156 58948
rect 34152 59041 34161 59075
rect 34161 59041 34195 59075
rect 34195 59041 34204 59075
rect 34152 59032 34204 59041
rect 34336 59075 34388 59084
rect 34336 59041 34345 59075
rect 34345 59041 34379 59075
rect 34379 59041 34388 59075
rect 34336 59032 34388 59041
rect 35440 59032 35492 59084
rect 35992 59075 36044 59084
rect 35992 59041 36006 59075
rect 36006 59041 36040 59075
rect 36040 59041 36044 59075
rect 35992 59032 36044 59041
rect 36820 59032 36872 59084
rect 37280 59032 37332 59084
rect 37924 58896 37976 58948
rect 31024 58828 31076 58880
rect 32404 58828 32456 58880
rect 36176 58871 36228 58880
rect 36176 58837 36185 58871
rect 36185 58837 36219 58871
rect 36219 58837 36228 58871
rect 36176 58828 36228 58837
rect 36728 58828 36780 58880
rect 4246 58726 4298 58778
rect 4310 58726 4362 58778
rect 4374 58726 4426 58778
rect 4438 58726 4490 58778
rect 34966 58726 35018 58778
rect 35030 58726 35082 58778
rect 35094 58726 35146 58778
rect 35158 58726 35210 58778
rect 31208 58624 31260 58676
rect 33784 58624 33836 58676
rect 36452 58667 36504 58676
rect 36452 58633 36461 58667
rect 36461 58633 36495 58667
rect 36495 58633 36504 58667
rect 36452 58624 36504 58633
rect 31392 58556 31444 58608
rect 34060 58556 34112 58608
rect 37280 58624 37332 58676
rect 36728 58556 36780 58608
rect 37832 58556 37884 58608
rect 1400 58463 1452 58472
rect 1400 58429 1409 58463
rect 1409 58429 1443 58463
rect 1443 58429 1452 58463
rect 1400 58420 1452 58429
rect 15660 58420 15712 58472
rect 32864 58463 32916 58472
rect 32864 58429 32873 58463
rect 32873 58429 32907 58463
rect 32907 58429 32916 58463
rect 32864 58420 32916 58429
rect 33140 58463 33192 58472
rect 33140 58429 33149 58463
rect 33149 58429 33183 58463
rect 33183 58429 33192 58463
rect 33140 58420 33192 58429
rect 34152 58488 34204 58540
rect 34796 58420 34848 58472
rect 35808 58420 35860 58472
rect 36268 58420 36320 58472
rect 36728 58420 36780 58472
rect 37004 58420 37056 58472
rect 37188 58420 37240 58472
rect 29736 58352 29788 58404
rect 37280 58395 37332 58404
rect 37280 58361 37289 58395
rect 37289 58361 37323 58395
rect 37323 58361 37332 58395
rect 37280 58352 37332 58361
rect 37372 58395 37424 58404
rect 37372 58361 37381 58395
rect 37381 58361 37415 58395
rect 37415 58361 37424 58395
rect 37372 58352 37424 58361
rect 29920 58284 29972 58336
rect 33600 58284 33652 58336
rect 19606 58182 19658 58234
rect 19670 58182 19722 58234
rect 19734 58182 19786 58234
rect 19798 58182 19850 58234
rect 18788 58080 18840 58132
rect 30104 58080 30156 58132
rect 30196 58080 30248 58132
rect 34060 58080 34112 58132
rect 37188 58080 37240 58132
rect 30288 58012 30340 58064
rect 34336 58012 34388 58064
rect 35992 58012 36044 58064
rect 37280 58012 37332 58064
rect 1400 57987 1452 57996
rect 1400 57953 1409 57987
rect 1409 57953 1443 57987
rect 1443 57953 1452 57987
rect 1400 57944 1452 57953
rect 29644 57944 29696 57996
rect 33324 57944 33376 57996
rect 36820 57944 36872 57996
rect 36912 57944 36964 57996
rect 30472 57876 30524 57928
rect 32036 57876 32088 57928
rect 37188 57944 37240 57996
rect 4246 57638 4298 57690
rect 4310 57638 4362 57690
rect 4374 57638 4426 57690
rect 4438 57638 4490 57690
rect 34966 57638 35018 57690
rect 35030 57638 35082 57690
rect 35094 57638 35146 57690
rect 35158 57638 35210 57690
rect 37280 57579 37332 57588
rect 37280 57545 37289 57579
rect 37289 57545 37323 57579
rect 37323 57545 37332 57579
rect 37280 57536 37332 57545
rect 37464 57375 37516 57384
rect 37464 57341 37473 57375
rect 37473 57341 37507 57375
rect 37507 57341 37516 57375
rect 37464 57332 37516 57341
rect 37924 57375 37976 57384
rect 37924 57341 37933 57375
rect 37933 57341 37967 57375
rect 37967 57341 37976 57375
rect 37924 57332 37976 57341
rect 19606 57094 19658 57146
rect 19670 57094 19722 57146
rect 19734 57094 19786 57146
rect 19798 57094 19850 57146
rect 1400 56899 1452 56908
rect 1400 56865 1409 56899
rect 1409 56865 1443 56899
rect 1443 56865 1452 56899
rect 1400 56856 1452 56865
rect 31944 56652 31996 56704
rect 37648 56652 37700 56704
rect 4246 56550 4298 56602
rect 4310 56550 4362 56602
rect 4374 56550 4426 56602
rect 4438 56550 4490 56602
rect 34966 56550 35018 56602
rect 35030 56550 35082 56602
rect 35094 56550 35146 56602
rect 35158 56550 35210 56602
rect 15752 56491 15804 56500
rect 15752 56457 15761 56491
rect 15761 56457 15795 56491
rect 15795 56457 15804 56491
rect 15752 56448 15804 56457
rect 16856 56448 16908 56500
rect 17776 56448 17828 56500
rect 1400 56287 1452 56296
rect 1400 56253 1409 56287
rect 1409 56253 1443 56287
rect 1443 56253 1452 56287
rect 1400 56244 1452 56253
rect 2964 56176 3016 56228
rect 17316 56287 17368 56296
rect 6460 56108 6512 56160
rect 16764 56176 16816 56228
rect 17316 56253 17325 56287
rect 17325 56253 17359 56287
rect 17359 56253 17368 56287
rect 17316 56244 17368 56253
rect 33048 56287 33100 56296
rect 33048 56253 33057 56287
rect 33057 56253 33091 56287
rect 33091 56253 33100 56287
rect 33048 56244 33100 56253
rect 33692 56312 33744 56364
rect 34244 56312 34296 56364
rect 37464 56287 37516 56296
rect 37464 56253 37473 56287
rect 37473 56253 37507 56287
rect 37507 56253 37516 56287
rect 37464 56244 37516 56253
rect 37924 56287 37976 56296
rect 37924 56253 37933 56287
rect 37933 56253 37967 56287
rect 37967 56253 37976 56287
rect 37924 56244 37976 56253
rect 16856 56108 16908 56160
rect 32496 56176 32548 56228
rect 33876 56176 33928 56228
rect 34152 56108 34204 56160
rect 37556 56108 37608 56160
rect 19606 56006 19658 56058
rect 19670 56006 19722 56058
rect 19734 56006 19786 56058
rect 19798 56006 19850 56058
rect 2412 55904 2464 55956
rect 16856 55904 16908 55956
rect 16028 55836 16080 55888
rect 33048 55836 33100 55888
rect 17684 55768 17736 55820
rect 33508 55904 33560 55956
rect 36452 55904 36504 55956
rect 37004 55904 37056 55956
rect 33876 55836 33928 55888
rect 35256 55836 35308 55888
rect 35808 55836 35860 55888
rect 36084 55836 36136 55888
rect 36820 55836 36872 55888
rect 38476 55836 38528 55888
rect 37188 55811 37240 55820
rect 32496 55700 32548 55752
rect 32864 55700 32916 55752
rect 37188 55777 37197 55811
rect 37197 55777 37231 55811
rect 37231 55777 37240 55811
rect 37188 55768 37240 55777
rect 35256 55700 35308 55752
rect 35716 55700 35768 55752
rect 31944 55632 31996 55684
rect 32496 55564 32548 55616
rect 32680 55564 32732 55616
rect 33140 55564 33192 55616
rect 33600 55564 33652 55616
rect 4246 55462 4298 55514
rect 4310 55462 4362 55514
rect 4374 55462 4426 55514
rect 4438 55462 4490 55514
rect 34966 55462 35018 55514
rect 35030 55462 35082 55514
rect 35094 55462 35146 55514
rect 35158 55462 35210 55514
rect 1400 55199 1452 55208
rect 1400 55165 1409 55199
rect 1409 55165 1443 55199
rect 1443 55165 1452 55199
rect 1400 55156 1452 55165
rect 18512 55088 18564 55140
rect 32220 55199 32272 55208
rect 32220 55165 32227 55199
rect 32227 55165 32272 55199
rect 32220 55156 32272 55165
rect 32864 55224 32916 55276
rect 33508 55224 33560 55276
rect 32588 55156 32640 55208
rect 32680 55156 32732 55208
rect 33416 55199 33468 55208
rect 33416 55165 33423 55199
rect 33423 55165 33468 55199
rect 33416 55156 33468 55165
rect 33876 55224 33928 55276
rect 31760 55020 31812 55072
rect 32864 55088 32916 55140
rect 33968 55156 34020 55208
rect 37464 55199 37516 55208
rect 37464 55165 37473 55199
rect 37473 55165 37507 55199
rect 37507 55165 37516 55199
rect 37464 55156 37516 55165
rect 37924 55199 37976 55208
rect 37924 55165 37933 55199
rect 37933 55165 37967 55199
rect 37967 55165 37976 55199
rect 37924 55156 37976 55165
rect 33692 55020 33744 55072
rect 37372 55020 37424 55072
rect 19606 54918 19658 54970
rect 19670 54918 19722 54970
rect 19734 54918 19786 54970
rect 19798 54918 19850 54970
rect 33876 54816 33928 54868
rect 34244 54816 34296 54868
rect 18696 54748 18748 54800
rect 32680 54748 32732 54800
rect 1400 54723 1452 54732
rect 1400 54689 1409 54723
rect 1409 54689 1443 54723
rect 1443 54689 1452 54723
rect 1400 54680 1452 54689
rect 29644 54680 29696 54732
rect 34428 54748 34480 54800
rect 32864 54612 32916 54664
rect 33508 54723 33560 54732
rect 33508 54689 33517 54723
rect 33517 54689 33551 54723
rect 33551 54689 33560 54723
rect 33508 54680 33560 54689
rect 35532 54680 35584 54732
rect 37188 54723 37240 54732
rect 37188 54689 37197 54723
rect 37197 54689 37231 54723
rect 37231 54689 37240 54723
rect 37188 54680 37240 54689
rect 33416 54476 33468 54528
rect 4246 54374 4298 54426
rect 4310 54374 4362 54426
rect 4374 54374 4426 54426
rect 4438 54374 4490 54426
rect 34966 54374 35018 54426
rect 35030 54374 35082 54426
rect 35094 54374 35146 54426
rect 35158 54374 35210 54426
rect 21548 54315 21600 54324
rect 21548 54281 21557 54315
rect 21557 54281 21591 54315
rect 21591 54281 21600 54315
rect 21548 54272 21600 54281
rect 32128 54315 32180 54324
rect 32128 54281 32137 54315
rect 32137 54281 32171 54315
rect 32171 54281 32180 54315
rect 32128 54272 32180 54281
rect 33232 54315 33284 54324
rect 33232 54281 33241 54315
rect 33241 54281 33275 54315
rect 33275 54281 33284 54315
rect 33232 54272 33284 54281
rect 38936 54272 38988 54324
rect 32036 54204 32088 54256
rect 28172 54068 28224 54120
rect 7380 54000 7432 54052
rect 24400 54000 24452 54052
rect 27712 53932 27764 53984
rect 38200 54000 38252 54052
rect 19606 53830 19658 53882
rect 19670 53830 19722 53882
rect 19734 53830 19786 53882
rect 19798 53830 19850 53882
rect 19340 53771 19392 53780
rect 19340 53737 19349 53771
rect 19349 53737 19383 53771
rect 19383 53737 19392 53771
rect 19340 53728 19392 53737
rect 22928 53771 22980 53780
rect 22928 53737 22937 53771
rect 22937 53737 22971 53771
rect 22971 53737 22980 53771
rect 22928 53728 22980 53737
rect 25044 53771 25096 53780
rect 25044 53737 25053 53771
rect 25053 53737 25087 53771
rect 25087 53737 25096 53771
rect 25044 53728 25096 53737
rect 27988 53771 28040 53780
rect 27988 53737 27997 53771
rect 27997 53737 28031 53771
rect 28031 53737 28040 53771
rect 27988 53728 28040 53737
rect 1400 53635 1452 53644
rect 1400 53601 1409 53635
rect 1409 53601 1443 53635
rect 1443 53601 1452 53635
rect 1400 53592 1452 53601
rect 3516 53592 3568 53644
rect 11244 53524 11296 53576
rect 29460 53660 29512 53712
rect 9680 53456 9732 53508
rect 25044 53592 25096 53644
rect 36728 53635 36780 53644
rect 19432 53388 19484 53440
rect 36728 53601 36737 53635
rect 36737 53601 36771 53635
rect 36771 53601 36780 53635
rect 36728 53592 36780 53601
rect 37188 53635 37240 53644
rect 37188 53601 37197 53635
rect 37197 53601 37231 53635
rect 37231 53601 37240 53635
rect 37188 53592 37240 53601
rect 34244 53388 34296 53440
rect 4246 53286 4298 53338
rect 4310 53286 4362 53338
rect 4374 53286 4426 53338
rect 4438 53286 4490 53338
rect 34966 53286 35018 53338
rect 35030 53286 35082 53338
rect 35094 53286 35146 53338
rect 35158 53286 35210 53338
rect 16488 53184 16540 53236
rect 25044 53184 25096 53236
rect 38660 53116 38712 53168
rect 38936 53116 38988 53168
rect 1400 53023 1452 53032
rect 1400 52989 1409 53023
rect 1409 52989 1443 53023
rect 1443 52989 1452 53023
rect 1400 52980 1452 52989
rect 37280 53023 37332 53032
rect 37280 52989 37289 53023
rect 37289 52989 37323 53023
rect 37323 52989 37332 53023
rect 37280 52980 37332 52989
rect 37924 53023 37976 53032
rect 37924 52989 37933 53023
rect 37933 52989 37967 53023
rect 37967 52989 37976 53023
rect 37924 52980 37976 52989
rect 19606 52742 19658 52794
rect 19670 52742 19722 52794
rect 19734 52742 19786 52794
rect 19798 52742 19850 52794
rect 1400 52547 1452 52556
rect 1400 52513 1409 52547
rect 1409 52513 1443 52547
rect 1443 52513 1452 52547
rect 1400 52504 1452 52513
rect 32680 52368 32732 52420
rect 36268 52368 36320 52420
rect 4246 52198 4298 52250
rect 4310 52198 4362 52250
rect 4374 52198 4426 52250
rect 4438 52198 4490 52250
rect 34966 52198 35018 52250
rect 35030 52198 35082 52250
rect 35094 52198 35146 52250
rect 35158 52198 35210 52250
rect 35532 52028 35584 52080
rect 32956 51892 33008 51944
rect 37556 51960 37608 52012
rect 37464 51935 37516 51944
rect 37464 51901 37473 51935
rect 37473 51901 37507 51935
rect 37507 51901 37516 51935
rect 37464 51892 37516 51901
rect 37924 51935 37976 51944
rect 37924 51901 37933 51935
rect 37933 51901 37967 51935
rect 37967 51901 37976 51935
rect 37924 51892 37976 51901
rect 32864 51799 32916 51808
rect 32864 51765 32873 51799
rect 32873 51765 32907 51799
rect 32907 51765 32916 51799
rect 32864 51756 32916 51765
rect 38752 51824 38804 51876
rect 33508 51756 33560 51808
rect 33600 51756 33652 51808
rect 35440 51756 35492 51808
rect 19606 51654 19658 51706
rect 19670 51654 19722 51706
rect 19734 51654 19786 51706
rect 19798 51654 19850 51706
rect 33600 51552 33652 51604
rect 38752 51552 38804 51604
rect 1400 51459 1452 51468
rect 1400 51425 1409 51459
rect 1409 51425 1443 51459
rect 1443 51425 1452 51459
rect 1400 51416 1452 51425
rect 33232 51416 33284 51468
rect 33508 51416 33560 51468
rect 37372 51484 37424 51536
rect 37188 51459 37240 51468
rect 37188 51425 37197 51459
rect 37197 51425 37231 51459
rect 37231 51425 37240 51459
rect 37188 51416 37240 51425
rect 2320 51212 2372 51264
rect 34612 51212 34664 51264
rect 4246 51110 4298 51162
rect 4310 51110 4362 51162
rect 4374 51110 4426 51162
rect 4438 51110 4490 51162
rect 34966 51110 35018 51162
rect 35030 51110 35082 51162
rect 35094 51110 35146 51162
rect 35158 51110 35210 51162
rect 32588 50940 32640 50992
rect 35624 50940 35676 50992
rect 33692 50872 33744 50924
rect 34060 50872 34112 50924
rect 27528 50804 27580 50856
rect 1860 50779 1912 50788
rect 1860 50745 1869 50779
rect 1869 50745 1903 50779
rect 1903 50745 1912 50779
rect 1860 50736 1912 50745
rect 33508 50804 33560 50856
rect 34244 50804 34296 50856
rect 37464 50847 37516 50856
rect 37464 50813 37473 50847
rect 37473 50813 37507 50847
rect 37507 50813 37516 50847
rect 37464 50804 37516 50813
rect 37924 50847 37976 50856
rect 37924 50813 37933 50847
rect 37933 50813 37967 50847
rect 37967 50813 37976 50847
rect 37924 50804 37976 50813
rect 32864 50668 32916 50720
rect 33324 50668 33376 50720
rect 33600 50668 33652 50720
rect 35808 50668 35860 50720
rect 37556 50668 37608 50720
rect 19606 50566 19658 50618
rect 19670 50566 19722 50618
rect 19734 50566 19786 50618
rect 19798 50566 19850 50618
rect 33692 50464 33744 50516
rect 3608 50328 3660 50380
rect 28908 50371 28960 50380
rect 28908 50337 28917 50371
rect 28917 50337 28951 50371
rect 28951 50337 28960 50371
rect 28908 50328 28960 50337
rect 33140 50328 33192 50380
rect 35440 50396 35492 50448
rect 24860 50260 24912 50312
rect 28908 50192 28960 50244
rect 32128 50192 32180 50244
rect 33600 50192 33652 50244
rect 34520 50328 34572 50380
rect 33508 50124 33560 50176
rect 33692 50124 33744 50176
rect 35624 50124 35676 50176
rect 4246 50022 4298 50074
rect 4310 50022 4362 50074
rect 4374 50022 4426 50074
rect 4438 50022 4490 50074
rect 34966 50022 35018 50074
rect 35030 50022 35082 50074
rect 35094 50022 35146 50074
rect 35158 50022 35210 50074
rect 2320 49852 2372 49904
rect 1860 49759 1912 49768
rect 1860 49725 1869 49759
rect 1869 49725 1903 49759
rect 1903 49725 1912 49759
rect 1860 49716 1912 49725
rect 33508 49852 33560 49904
rect 32128 49784 32180 49836
rect 32220 49759 32272 49768
rect 32220 49725 32229 49759
rect 32229 49725 32263 49759
rect 32263 49725 32272 49759
rect 32220 49716 32272 49725
rect 32772 49716 32824 49768
rect 34520 49716 34572 49768
rect 34796 49716 34848 49768
rect 37924 49759 37976 49768
rect 37924 49725 37933 49759
rect 37933 49725 37967 49759
rect 37967 49725 37976 49759
rect 37924 49716 37976 49725
rect 32036 49623 32088 49632
rect 32036 49589 32045 49623
rect 32045 49589 32079 49623
rect 32079 49589 32088 49623
rect 32036 49580 32088 49589
rect 19606 49478 19658 49530
rect 19670 49478 19722 49530
rect 19734 49478 19786 49530
rect 19798 49478 19850 49530
rect 1860 49283 1912 49292
rect 1860 49249 1869 49283
rect 1869 49249 1903 49283
rect 1903 49249 1912 49283
rect 1860 49240 1912 49249
rect 37372 49283 37424 49292
rect 37372 49249 37381 49283
rect 37381 49249 37415 49283
rect 37415 49249 37424 49283
rect 37372 49240 37424 49249
rect 2320 49172 2372 49224
rect 24860 49172 24912 49224
rect 33324 49036 33376 49088
rect 34520 49036 34572 49088
rect 4246 48934 4298 48986
rect 4310 48934 4362 48986
rect 4374 48934 4426 48986
rect 4438 48934 4490 48986
rect 34966 48934 35018 48986
rect 35030 48934 35082 48986
rect 35094 48934 35146 48986
rect 35158 48934 35210 48986
rect 16764 48628 16816 48680
rect 27620 48671 27672 48680
rect 27620 48637 27629 48671
rect 27629 48637 27663 48671
rect 27663 48637 27672 48671
rect 27620 48628 27672 48637
rect 29552 48764 29604 48816
rect 32036 48696 32088 48748
rect 28540 48671 28592 48680
rect 28540 48637 28549 48671
rect 28549 48637 28583 48671
rect 28583 48637 28592 48671
rect 28540 48628 28592 48637
rect 37280 48671 37332 48680
rect 37280 48637 37289 48671
rect 37289 48637 37323 48671
rect 37323 48637 37332 48671
rect 37280 48628 37332 48637
rect 37924 48671 37976 48680
rect 37924 48637 37933 48671
rect 37933 48637 37967 48671
rect 37967 48637 37976 48671
rect 37924 48628 37976 48637
rect 6644 48560 6696 48612
rect 16856 48535 16908 48544
rect 16856 48501 16865 48535
rect 16865 48501 16899 48535
rect 16899 48501 16908 48535
rect 16856 48492 16908 48501
rect 19606 48390 19658 48442
rect 19670 48390 19722 48442
rect 19734 48390 19786 48442
rect 19798 48390 19850 48442
rect 2320 48220 2372 48272
rect 1860 48195 1912 48204
rect 1860 48161 1869 48195
rect 1869 48161 1903 48195
rect 1903 48161 1912 48195
rect 1860 48152 1912 48161
rect 37372 48195 37424 48204
rect 37372 48161 37381 48195
rect 37381 48161 37415 48195
rect 37415 48161 37424 48195
rect 37372 48152 37424 48161
rect 34612 48084 34664 48136
rect 35440 48084 35492 48136
rect 34612 47948 34664 48000
rect 4246 47846 4298 47898
rect 4310 47846 4362 47898
rect 4374 47846 4426 47898
rect 4438 47846 4490 47898
rect 34966 47846 35018 47898
rect 35030 47846 35082 47898
rect 35094 47846 35146 47898
rect 35158 47846 35210 47898
rect 16764 47583 16816 47592
rect 16764 47549 16773 47583
rect 16773 47549 16807 47583
rect 16807 47549 16816 47583
rect 16764 47540 16816 47549
rect 37280 47583 37332 47592
rect 37280 47549 37289 47583
rect 37289 47549 37323 47583
rect 37323 47549 37332 47583
rect 37280 47540 37332 47549
rect 37924 47583 37976 47592
rect 37924 47549 37933 47583
rect 37933 47549 37967 47583
rect 37967 47549 37976 47583
rect 37924 47540 37976 47549
rect 1860 47515 1912 47524
rect 1860 47481 1869 47515
rect 1869 47481 1903 47515
rect 1903 47481 1912 47515
rect 1860 47472 1912 47481
rect 1952 47447 2004 47456
rect 1952 47413 1961 47447
rect 1961 47413 1995 47447
rect 1995 47413 2004 47447
rect 1952 47404 2004 47413
rect 17316 47404 17368 47456
rect 19606 47302 19658 47354
rect 19670 47302 19722 47354
rect 19734 47302 19786 47354
rect 19798 47302 19850 47354
rect 1952 47200 2004 47252
rect 33968 47107 34020 47116
rect 33968 47073 33977 47107
rect 33977 47073 34011 47107
rect 34011 47073 34020 47107
rect 33968 47064 34020 47073
rect 34244 47107 34296 47116
rect 34244 47073 34253 47107
rect 34253 47073 34287 47107
rect 34287 47073 34296 47107
rect 34244 47064 34296 47073
rect 37556 47064 37608 47116
rect 34428 46928 34480 46980
rect 36084 46928 36136 46980
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 34966 46758 35018 46810
rect 35030 46758 35082 46810
rect 35094 46758 35146 46810
rect 35158 46758 35210 46810
rect 35348 46588 35400 46640
rect 1860 46495 1912 46504
rect 1860 46461 1869 46495
rect 1869 46461 1903 46495
rect 1903 46461 1912 46495
rect 1860 46452 1912 46461
rect 33784 46452 33836 46504
rect 34520 46452 34572 46504
rect 34244 46427 34296 46436
rect 34244 46393 34253 46427
rect 34253 46393 34287 46427
rect 34287 46393 34296 46427
rect 34244 46384 34296 46393
rect 34428 46316 34480 46368
rect 34520 46316 34572 46368
rect 34796 46452 34848 46504
rect 37464 46495 37516 46504
rect 37464 46461 37473 46495
rect 37473 46461 37507 46495
rect 37507 46461 37516 46495
rect 37464 46452 37516 46461
rect 37924 46495 37976 46504
rect 37924 46461 37933 46495
rect 37933 46461 37967 46495
rect 37967 46461 37976 46495
rect 37924 46452 37976 46461
rect 34796 46316 34848 46368
rect 19606 46214 19658 46266
rect 19670 46214 19722 46266
rect 19734 46214 19786 46266
rect 19798 46214 19850 46266
rect 1860 46019 1912 46028
rect 1860 45985 1869 46019
rect 1869 45985 1903 46019
rect 1903 45985 1912 46019
rect 1860 45976 1912 45985
rect 34336 46112 34388 46164
rect 34244 46019 34296 46028
rect 34244 45985 34253 46019
rect 34253 45985 34287 46019
rect 34287 45985 34296 46019
rect 34244 45976 34296 45985
rect 34336 46019 34388 46028
rect 34336 45985 34345 46019
rect 34345 45985 34379 46019
rect 34379 45985 34388 46019
rect 34336 45976 34388 45985
rect 34612 45976 34664 46028
rect 37188 46019 37240 46028
rect 37188 45985 37197 46019
rect 37197 45985 37231 46019
rect 37231 45985 37240 46019
rect 37188 45976 37240 45985
rect 30288 45840 30340 45892
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 34966 45670 35018 45722
rect 35030 45670 35082 45722
rect 35094 45670 35146 45722
rect 35158 45670 35210 45722
rect 36452 45500 36504 45552
rect 35716 45432 35768 45484
rect 34060 45407 34112 45416
rect 34060 45373 34070 45407
rect 34070 45373 34104 45407
rect 34104 45373 34112 45407
rect 34060 45364 34112 45373
rect 34796 45364 34848 45416
rect 37464 45407 37516 45416
rect 37464 45373 37473 45407
rect 37473 45373 37507 45407
rect 37507 45373 37516 45407
rect 37464 45364 37516 45373
rect 37924 45407 37976 45416
rect 37924 45373 37933 45407
rect 37933 45373 37967 45407
rect 37967 45373 37976 45407
rect 37924 45364 37976 45373
rect 34244 45339 34296 45348
rect 34244 45305 34253 45339
rect 34253 45305 34287 45339
rect 34287 45305 34296 45339
rect 34244 45296 34296 45305
rect 34336 45339 34388 45348
rect 34336 45305 34345 45339
rect 34345 45305 34379 45339
rect 34379 45305 34388 45339
rect 34336 45296 34388 45305
rect 34612 45296 34664 45348
rect 35532 45296 35584 45348
rect 35716 45296 35768 45348
rect 35900 45296 35952 45348
rect 34796 45228 34848 45280
rect 19606 45126 19658 45178
rect 19670 45126 19722 45178
rect 19734 45126 19786 45178
rect 19798 45126 19850 45178
rect 33784 45024 33836 45076
rect 39396 45024 39448 45076
rect 1860 44999 1912 45008
rect 1860 44965 1869 44999
rect 1869 44965 1903 44999
rect 1903 44965 1912 44999
rect 1860 44956 1912 44965
rect 34060 44684 34112 44736
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 34966 44582 35018 44634
rect 35030 44582 35082 44634
rect 35094 44582 35146 44634
rect 35158 44582 35210 44634
rect 33416 44412 33468 44464
rect 34060 44412 34112 44464
rect 34336 44412 34388 44464
rect 33692 44344 33744 44396
rect 33876 44319 33928 44328
rect 33876 44285 33885 44319
rect 33885 44285 33919 44319
rect 33919 44285 33928 44319
rect 33876 44276 33928 44285
rect 34244 44344 34296 44396
rect 1860 44251 1912 44260
rect 1860 44217 1869 44251
rect 1869 44217 1903 44251
rect 1903 44217 1912 44251
rect 1860 44208 1912 44217
rect 34796 44276 34848 44328
rect 37188 44276 37240 44328
rect 37924 44319 37976 44328
rect 37924 44285 37933 44319
rect 37933 44285 37967 44319
rect 37967 44285 37976 44319
rect 37924 44276 37976 44285
rect 34060 44208 34112 44260
rect 36728 44140 36780 44192
rect 37280 44183 37332 44192
rect 37280 44149 37289 44183
rect 37289 44149 37323 44183
rect 37323 44149 37332 44183
rect 37280 44140 37332 44149
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 33968 43936 34020 43988
rect 34244 43936 34296 43988
rect 37188 43843 37240 43852
rect 37188 43809 37197 43843
rect 37197 43809 37231 43843
rect 37231 43809 37240 43843
rect 37188 43800 37240 43809
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 15660 43435 15712 43444
rect 15660 43401 15669 43435
rect 15669 43401 15703 43435
rect 15703 43401 15712 43435
rect 15660 43392 15712 43401
rect 16304 43392 16356 43444
rect 25688 43392 25740 43444
rect 18788 43324 18840 43376
rect 16856 43256 16908 43308
rect 1860 43231 1912 43240
rect 1860 43197 1869 43231
rect 1869 43197 1903 43231
rect 1903 43197 1912 43231
rect 1860 43188 1912 43197
rect 15476 43231 15528 43240
rect 15476 43197 15485 43231
rect 15485 43197 15519 43231
rect 15519 43197 15528 43231
rect 15476 43188 15528 43197
rect 16396 43231 16448 43240
rect 16396 43197 16405 43231
rect 16405 43197 16439 43231
rect 16439 43197 16448 43231
rect 16396 43188 16448 43197
rect 37924 43231 37976 43240
rect 37924 43197 37933 43231
rect 37933 43197 37967 43231
rect 37967 43197 37976 43231
rect 37924 43188 37976 43197
rect 1952 43095 2004 43104
rect 1952 43061 1961 43095
rect 1961 43061 1995 43095
rect 1995 43061 2004 43095
rect 1952 43052 2004 43061
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 1952 42848 2004 42900
rect 24860 42848 24912 42900
rect 1860 42755 1912 42764
rect 1860 42721 1869 42755
rect 1869 42721 1903 42755
rect 1903 42721 1912 42755
rect 1860 42712 1912 42721
rect 16120 42755 16172 42764
rect 16120 42721 16129 42755
rect 16129 42721 16163 42755
rect 16163 42721 16172 42755
rect 16120 42712 16172 42721
rect 16304 42755 16356 42764
rect 16304 42721 16313 42755
rect 16313 42721 16347 42755
rect 16347 42721 16356 42755
rect 16304 42712 16356 42721
rect 17500 42755 17552 42764
rect 17500 42721 17509 42755
rect 17509 42721 17543 42755
rect 17543 42721 17552 42755
rect 17500 42712 17552 42721
rect 25596 42712 25648 42764
rect 33048 42712 33100 42764
rect 36820 42712 36872 42764
rect 37372 42755 37424 42764
rect 37372 42721 37381 42755
rect 37381 42721 37415 42755
rect 37415 42721 37424 42755
rect 37372 42712 37424 42721
rect 16856 42644 16908 42696
rect 33876 42576 33928 42628
rect 34428 42508 34480 42560
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 16580 42347 16632 42356
rect 16580 42313 16589 42347
rect 16589 42313 16623 42347
rect 16623 42313 16632 42347
rect 16580 42304 16632 42313
rect 37280 42304 37332 42356
rect 16856 42168 16908 42220
rect 16304 42100 16356 42152
rect 24860 42100 24912 42152
rect 33784 42143 33836 42152
rect 33784 42109 33793 42143
rect 33793 42109 33827 42143
rect 33827 42109 33836 42143
rect 33784 42100 33836 42109
rect 33968 42100 34020 42152
rect 37280 42143 37332 42152
rect 37280 42109 37289 42143
rect 37289 42109 37323 42143
rect 37323 42109 37332 42143
rect 37280 42100 37332 42109
rect 37924 42143 37976 42152
rect 37924 42109 37933 42143
rect 37933 42109 37967 42143
rect 37967 42109 37976 42143
rect 37924 42100 37976 42109
rect 34060 42075 34112 42084
rect 34060 42041 34069 42075
rect 34069 42041 34103 42075
rect 34103 42041 34112 42075
rect 34060 42032 34112 42041
rect 34336 41964 34388 42016
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 1860 41735 1912 41744
rect 1860 41701 1869 41735
rect 1869 41701 1903 41735
rect 1903 41701 1912 41735
rect 1860 41692 1912 41701
rect 34060 41735 34112 41744
rect 34060 41701 34069 41735
rect 34069 41701 34103 41735
rect 34103 41701 34112 41735
rect 34060 41692 34112 41701
rect 2688 41488 2740 41540
rect 30932 41420 30984 41472
rect 32404 41420 32456 41472
rect 33876 41667 33928 41676
rect 33876 41633 33886 41667
rect 33886 41633 33920 41667
rect 33920 41633 33928 41667
rect 33876 41624 33928 41633
rect 33876 41488 33928 41540
rect 34060 41488 34112 41540
rect 34428 41624 34480 41676
rect 37188 41624 37240 41676
rect 39028 41556 39080 41608
rect 35256 41488 35308 41540
rect 35900 41420 35952 41472
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 26148 41080 26200 41132
rect 2688 41012 2740 41064
rect 1860 40987 1912 40996
rect 1860 40953 1869 40987
rect 1869 40953 1903 40987
rect 1903 40953 1912 40987
rect 1860 40944 1912 40953
rect 2596 40944 2648 40996
rect 33876 41012 33928 41064
rect 35256 41012 35308 41064
rect 37280 41055 37332 41064
rect 37280 41021 37289 41055
rect 37289 41021 37323 41055
rect 37323 41021 37332 41055
rect 37280 41012 37332 41021
rect 37924 41055 37976 41064
rect 37924 41021 37933 41055
rect 37933 41021 37967 41055
rect 37967 41021 37976 41055
rect 37924 41012 37976 41021
rect 34060 40987 34112 40996
rect 34060 40953 34069 40987
rect 34069 40953 34103 40987
rect 34103 40953 34112 40987
rect 34060 40944 34112 40953
rect 35440 40876 35492 40928
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 1860 40579 1912 40588
rect 1860 40545 1869 40579
rect 1869 40545 1903 40579
rect 1903 40545 1912 40579
rect 1860 40536 1912 40545
rect 17224 40536 17276 40588
rect 17316 40511 17368 40520
rect 17316 40477 17325 40511
rect 17325 40477 17359 40511
rect 17359 40477 17368 40511
rect 17316 40468 17368 40477
rect 2688 40400 2740 40452
rect 29644 40332 29696 40384
rect 36176 40332 36228 40384
rect 36820 40332 36872 40384
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 17684 40171 17736 40180
rect 17684 40137 17693 40171
rect 17693 40137 17727 40171
rect 17727 40137 17736 40171
rect 17684 40128 17736 40137
rect 17316 40060 17368 40112
rect 2596 39992 2648 40044
rect 9128 39992 9180 40044
rect 16028 40035 16080 40044
rect 16028 40001 16037 40035
rect 16037 40001 16071 40035
rect 16071 40001 16080 40035
rect 16028 39992 16080 40001
rect 16672 39967 16724 39976
rect 16672 39933 16681 39967
rect 16681 39933 16715 39967
rect 16715 39933 16724 39967
rect 16672 39924 16724 39933
rect 36176 40060 36228 40112
rect 36636 40060 36688 40112
rect 17316 39967 17368 39976
rect 17316 39933 17325 39967
rect 17325 39933 17359 39967
rect 17359 39933 17368 39967
rect 17316 39924 17368 39933
rect 17132 39856 17184 39908
rect 18512 40035 18564 40044
rect 18512 40001 18521 40035
rect 18521 40001 18555 40035
rect 18555 40001 18564 40035
rect 18512 39992 18564 40001
rect 18328 39967 18380 39976
rect 18328 39933 18337 39967
rect 18337 39933 18371 39967
rect 18371 39933 18380 39967
rect 18328 39924 18380 39933
rect 38108 39992 38160 40044
rect 18696 39856 18748 39908
rect 33876 39924 33928 39976
rect 37464 39967 37516 39976
rect 34060 39899 34112 39908
rect 34060 39865 34069 39899
rect 34069 39865 34103 39899
rect 34103 39865 34112 39899
rect 34060 39856 34112 39865
rect 36636 39788 36688 39840
rect 37464 39933 37473 39967
rect 37473 39933 37507 39967
rect 37507 39933 37516 39967
rect 37464 39924 37516 39933
rect 37924 39967 37976 39976
rect 37924 39933 37933 39967
rect 37933 39933 37967 39967
rect 37967 39933 37976 39967
rect 37924 39924 37976 39933
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 1860 39491 1912 39500
rect 1860 39457 1869 39491
rect 1869 39457 1903 39491
rect 1903 39457 1912 39491
rect 1860 39448 1912 39457
rect 2688 39448 2740 39500
rect 33876 39516 33928 39568
rect 34060 39491 34112 39500
rect 34060 39457 34069 39491
rect 34069 39457 34103 39491
rect 34103 39457 34112 39491
rect 34060 39448 34112 39457
rect 37280 39448 37332 39500
rect 38568 39380 38620 39432
rect 2688 39312 2740 39364
rect 34428 39244 34480 39296
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 37280 39083 37332 39092
rect 37280 39049 37289 39083
rect 37289 39049 37323 39083
rect 37323 39049 37332 39083
rect 37280 39040 37332 39049
rect 37464 38879 37516 38888
rect 37464 38845 37473 38879
rect 37473 38845 37507 38879
rect 37507 38845 37516 38879
rect 37464 38836 37516 38845
rect 37924 38879 37976 38888
rect 37924 38845 37933 38879
rect 37933 38845 37967 38879
rect 37967 38845 37976 38879
rect 37924 38836 37976 38845
rect 1860 38811 1912 38820
rect 1860 38777 1869 38811
rect 1869 38777 1903 38811
rect 1903 38777 1912 38811
rect 1860 38768 1912 38777
rect 2596 38768 2648 38820
rect 32772 38700 32824 38752
rect 35808 38700 35860 38752
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 33692 38496 33744 38548
rect 34336 38496 34388 38548
rect 34796 38496 34848 38548
rect 28908 38428 28960 38480
rect 33416 38471 33468 38480
rect 33416 38437 33425 38471
rect 33425 38437 33459 38471
rect 33459 38437 33468 38471
rect 33416 38428 33468 38437
rect 33508 38428 33560 38480
rect 36360 38428 36412 38480
rect 33784 38360 33836 38412
rect 34336 38360 34388 38412
rect 34520 38360 34572 38412
rect 37188 38403 37240 38412
rect 37188 38369 37197 38403
rect 37197 38369 37231 38403
rect 37231 38369 37240 38403
rect 37188 38360 37240 38369
rect 33692 38224 33744 38276
rect 33600 38156 33652 38208
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 1860 37791 1912 37800
rect 1860 37757 1869 37791
rect 1869 37757 1903 37791
rect 1903 37757 1912 37791
rect 1860 37748 1912 37757
rect 37096 37816 37148 37868
rect 33600 37791 33652 37800
rect 4068 37680 4120 37732
rect 33600 37757 33609 37791
rect 33609 37757 33643 37791
rect 33643 37757 33652 37791
rect 33600 37748 33652 37757
rect 33692 37791 33744 37800
rect 33692 37757 33701 37791
rect 33701 37757 33735 37791
rect 33735 37757 33744 37791
rect 33692 37748 33744 37757
rect 37188 37748 37240 37800
rect 37924 37791 37976 37800
rect 37924 37757 37933 37791
rect 37933 37757 37967 37791
rect 37967 37757 37976 37791
rect 37924 37748 37976 37757
rect 2688 37612 2740 37664
rect 34060 37612 34112 37664
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 34520 37408 34572 37460
rect 37188 37451 37240 37460
rect 37188 37417 37197 37451
rect 37197 37417 37231 37451
rect 37231 37417 37240 37451
rect 37188 37408 37240 37417
rect 1860 37315 1912 37324
rect 1860 37281 1869 37315
rect 1869 37281 1903 37315
rect 1903 37281 1912 37315
rect 1860 37272 1912 37281
rect 2688 37272 2740 37324
rect 37372 37315 37424 37324
rect 37372 37281 37381 37315
rect 37381 37281 37415 37315
rect 37415 37281 37424 37315
rect 37372 37272 37424 37281
rect 34428 37204 34480 37256
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 33876 36864 33928 36916
rect 36360 36864 36412 36916
rect 36544 36864 36596 36916
rect 38292 36796 38344 36848
rect 33600 36728 33652 36780
rect 37096 36660 37148 36712
rect 37280 36703 37332 36712
rect 37280 36669 37289 36703
rect 37289 36669 37323 36703
rect 37323 36669 37332 36703
rect 37280 36660 37332 36669
rect 37924 36703 37976 36712
rect 37924 36669 37933 36703
rect 37933 36669 37967 36703
rect 37967 36669 37976 36703
rect 37924 36660 37976 36669
rect 2596 36524 2648 36576
rect 34336 36592 34388 36644
rect 33692 36524 33744 36576
rect 33876 36567 33928 36576
rect 33876 36533 33885 36567
rect 33885 36533 33919 36567
rect 33919 36533 33928 36567
rect 33876 36524 33928 36533
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 32404 36320 32456 36372
rect 4068 36252 4120 36304
rect 28724 36295 28776 36304
rect 1860 36227 1912 36236
rect 1860 36193 1869 36227
rect 1869 36193 1903 36227
rect 1903 36193 1912 36227
rect 1860 36184 1912 36193
rect 28724 36261 28733 36295
rect 28733 36261 28767 36295
rect 28767 36261 28776 36295
rect 28724 36252 28776 36261
rect 28908 36252 28960 36304
rect 33600 36320 33652 36372
rect 33692 36320 33744 36372
rect 33968 36320 34020 36372
rect 37096 36320 37148 36372
rect 33876 36252 33928 36304
rect 34704 36252 34756 36304
rect 33968 36184 34020 36236
rect 34888 36184 34940 36236
rect 37372 36227 37424 36236
rect 37372 36193 37381 36227
rect 37381 36193 37415 36227
rect 37415 36193 37424 36227
rect 37372 36184 37424 36193
rect 33508 36116 33560 36168
rect 35348 36116 35400 36168
rect 36268 36116 36320 36168
rect 2688 36048 2740 36100
rect 35348 35980 35400 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 33140 35776 33192 35828
rect 36176 35776 36228 35828
rect 2596 35572 2648 35624
rect 35256 35708 35308 35760
rect 33600 35640 33652 35692
rect 1860 35547 1912 35556
rect 1860 35513 1869 35547
rect 1869 35513 1903 35547
rect 1903 35513 1912 35547
rect 1860 35504 1912 35513
rect 2412 35504 2464 35556
rect 28724 35504 28776 35556
rect 36176 35572 36228 35624
rect 37280 35615 37332 35624
rect 37280 35581 37289 35615
rect 37289 35581 37323 35615
rect 37323 35581 37332 35615
rect 37280 35572 37332 35581
rect 37924 35615 37976 35624
rect 37924 35581 37933 35615
rect 37933 35581 37967 35615
rect 37967 35581 37976 35615
rect 37924 35572 37976 35581
rect 34428 35547 34480 35556
rect 33416 35436 33468 35488
rect 33508 35436 33560 35488
rect 34428 35513 34437 35547
rect 34437 35513 34471 35547
rect 34471 35513 34480 35547
rect 34428 35504 34480 35513
rect 33692 35436 33744 35488
rect 33876 35479 33928 35488
rect 33876 35445 33885 35479
rect 33885 35445 33919 35479
rect 33919 35445 33928 35479
rect 33876 35436 33928 35445
rect 34336 35436 34388 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 33600 35232 33652 35284
rect 33784 35164 33836 35216
rect 34428 35164 34480 35216
rect 33140 35139 33192 35148
rect 33140 35105 33149 35139
rect 33149 35105 33183 35139
rect 33183 35105 33192 35139
rect 33140 35096 33192 35105
rect 33508 35139 33560 35148
rect 33508 35105 33517 35139
rect 33517 35105 33551 35139
rect 33551 35105 33560 35139
rect 33508 35096 33560 35105
rect 2688 34892 2740 34944
rect 33876 35028 33928 35080
rect 37096 35028 37148 35080
rect 33692 34960 33744 35012
rect 33876 34892 33928 34944
rect 34428 34935 34480 34944
rect 34428 34901 34437 34935
rect 34437 34901 34471 34935
rect 34471 34901 34480 34935
rect 34428 34892 34480 34901
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 33968 34688 34020 34740
rect 2596 34484 2648 34536
rect 37464 34527 37516 34536
rect 37464 34493 37473 34527
rect 37473 34493 37507 34527
rect 37507 34493 37516 34527
rect 37464 34484 37516 34493
rect 37924 34527 37976 34536
rect 37924 34493 37933 34527
rect 37933 34493 37967 34527
rect 37967 34493 37976 34527
rect 37924 34484 37976 34493
rect 1860 34459 1912 34468
rect 1860 34425 1869 34459
rect 1869 34425 1903 34459
rect 1903 34425 1912 34459
rect 1860 34416 1912 34425
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 1860 34051 1912 34060
rect 1860 34017 1869 34051
rect 1869 34017 1903 34051
rect 1903 34017 1912 34051
rect 1860 34008 1912 34017
rect 2688 33872 2740 33924
rect 35808 33804 35860 33856
rect 36544 33804 36596 33856
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 36176 33600 36228 33652
rect 36176 33464 36228 33516
rect 36360 33464 36412 33516
rect 28724 33439 28776 33448
rect 28724 33405 28733 33439
rect 28733 33405 28767 33439
rect 28767 33405 28776 33439
rect 28724 33396 28776 33405
rect 33784 33396 33836 33448
rect 37464 33439 37516 33448
rect 37464 33405 37473 33439
rect 37473 33405 37507 33439
rect 37507 33405 37516 33439
rect 37464 33396 37516 33405
rect 37924 33439 37976 33448
rect 37924 33405 37933 33439
rect 37933 33405 37967 33439
rect 37967 33405 37976 33439
rect 37924 33396 37976 33405
rect 33140 33328 33192 33380
rect 32864 33260 32916 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 1860 33031 1912 33040
rect 1860 32997 1869 33031
rect 1869 32997 1903 33031
rect 1903 32997 1912 33031
rect 1860 32988 1912 32997
rect 32404 32988 32456 33040
rect 36820 32988 36872 33040
rect 34704 32920 34756 32972
rect 35808 32920 35860 32972
rect 37188 32963 37240 32972
rect 37188 32929 37197 32963
rect 37197 32929 37231 32963
rect 37231 32929 37240 32963
rect 37188 32920 37240 32929
rect 1952 32759 2004 32768
rect 1952 32725 1961 32759
rect 1961 32725 1995 32759
rect 1995 32725 2004 32759
rect 1952 32716 2004 32725
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 2412 32512 2464 32564
rect 34428 32376 34480 32428
rect 33324 32351 33376 32360
rect 1860 32283 1912 32292
rect 1860 32249 1869 32283
rect 1869 32249 1903 32283
rect 1903 32249 1912 32283
rect 1860 32240 1912 32249
rect 2412 32240 2464 32292
rect 33324 32317 33333 32351
rect 33333 32317 33367 32351
rect 33367 32317 33376 32351
rect 33324 32308 33376 32317
rect 33416 32351 33468 32360
rect 33416 32317 33425 32351
rect 33425 32317 33459 32351
rect 33459 32317 33468 32351
rect 33416 32308 33468 32317
rect 37188 32308 37240 32360
rect 37924 32351 37976 32360
rect 37924 32317 37933 32351
rect 37933 32317 37967 32351
rect 37967 32317 37976 32351
rect 37924 32308 37976 32317
rect 38752 32240 38804 32292
rect 35348 32172 35400 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 33968 31968 34020 32020
rect 37096 31968 37148 32020
rect 33324 31943 33376 31952
rect 33324 31909 33333 31943
rect 33333 31909 33367 31943
rect 33367 31909 33376 31943
rect 33324 31900 33376 31909
rect 33416 31943 33468 31952
rect 33416 31909 33425 31943
rect 33425 31909 33459 31943
rect 33459 31909 33468 31943
rect 33416 31900 33468 31909
rect 33048 31875 33100 31884
rect 33048 31841 33057 31875
rect 33057 31841 33091 31875
rect 33091 31841 33100 31875
rect 33048 31832 33100 31841
rect 2596 31764 2648 31816
rect 36820 31832 36872 31884
rect 37372 31875 37424 31884
rect 37372 31841 37381 31875
rect 37381 31841 37415 31875
rect 37415 31841 37424 31875
rect 37372 31832 37424 31841
rect 36636 31764 36688 31816
rect 37096 31764 37148 31816
rect 35532 31696 35584 31748
rect 36360 31628 36412 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 33324 31424 33376 31476
rect 33508 31424 33560 31476
rect 33692 31424 33744 31476
rect 35532 31424 35584 31476
rect 37740 31424 37792 31476
rect 1860 31263 1912 31272
rect 1860 31229 1869 31263
rect 1869 31229 1903 31263
rect 1903 31229 1912 31263
rect 1860 31220 1912 31229
rect 2688 31220 2740 31272
rect 36728 31356 36780 31408
rect 36912 31356 36964 31408
rect 33324 31263 33376 31272
rect 2596 31152 2648 31204
rect 33324 31229 33333 31263
rect 33333 31229 33367 31263
rect 33367 31229 33376 31263
rect 33324 31220 33376 31229
rect 36912 31220 36964 31272
rect 37280 31263 37332 31272
rect 37280 31229 37289 31263
rect 37289 31229 37323 31263
rect 37323 31229 37332 31263
rect 37280 31220 37332 31229
rect 37924 31263 37976 31272
rect 37924 31229 37933 31263
rect 37933 31229 37967 31263
rect 37967 31229 37976 31263
rect 37924 31220 37976 31229
rect 33324 31084 33376 31136
rect 33508 31084 33560 31136
rect 33784 31084 33836 31136
rect 34060 31084 34112 31136
rect 34612 31084 34664 31136
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 37188 30923 37240 30932
rect 37188 30889 37197 30923
rect 37197 30889 37231 30923
rect 37231 30889 37240 30923
rect 37188 30880 37240 30889
rect 33416 30855 33468 30864
rect 33416 30821 33425 30855
rect 33425 30821 33459 30855
rect 33459 30821 33468 30855
rect 33416 30812 33468 30821
rect 1860 30787 1912 30796
rect 1860 30753 1869 30787
rect 1869 30753 1903 30787
rect 1903 30753 1912 30787
rect 1860 30744 1912 30753
rect 32956 30744 33008 30796
rect 33324 30787 33376 30796
rect 1952 30676 2004 30728
rect 33324 30753 33333 30787
rect 33333 30753 33367 30787
rect 33367 30753 33376 30787
rect 33324 30744 33376 30753
rect 36636 30744 36688 30796
rect 37372 30787 37424 30796
rect 37372 30753 37381 30787
rect 37381 30753 37415 30787
rect 37415 30753 37424 30787
rect 37372 30744 37424 30753
rect 1952 30583 2004 30592
rect 1952 30549 1961 30583
rect 1961 30549 1995 30583
rect 1995 30549 2004 30583
rect 1952 30540 2004 30549
rect 34428 30540 34480 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 1952 30336 2004 30388
rect 27528 30336 27580 30388
rect 32496 30132 32548 30184
rect 33324 30268 33376 30320
rect 33416 30268 33468 30320
rect 37280 30175 37332 30184
rect 2412 29996 2464 30048
rect 33876 29996 33928 30048
rect 37280 30141 37289 30175
rect 37289 30141 37323 30175
rect 37323 30141 37332 30175
rect 37280 30132 37332 30141
rect 37924 30175 37976 30184
rect 37924 30141 37933 30175
rect 37933 30141 37967 30175
rect 37967 30141 37976 30175
rect 37924 30132 37976 30141
rect 37280 29996 37332 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 1860 29767 1912 29776
rect 1860 29733 1869 29767
rect 1869 29733 1903 29767
rect 1903 29733 1912 29767
rect 1860 29724 1912 29733
rect 2688 29520 2740 29572
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 36820 29248 36872 29300
rect 34428 29180 34480 29232
rect 34888 29180 34940 29232
rect 1860 29087 1912 29096
rect 1860 29053 1869 29087
rect 1869 29053 1903 29087
rect 1903 29053 1912 29087
rect 1860 29044 1912 29053
rect 37464 29087 37516 29096
rect 37464 29053 37473 29087
rect 37473 29053 37507 29087
rect 37507 29053 37516 29087
rect 37464 29044 37516 29053
rect 37924 29087 37976 29096
rect 37924 29053 37933 29087
rect 37933 29053 37967 29087
rect 37967 29053 37976 29087
rect 37924 29044 37976 29053
rect 4068 28976 4120 29028
rect 36360 28976 36412 29028
rect 36820 28976 36872 29028
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 32496 28704 32548 28756
rect 37832 28704 37884 28756
rect 34888 28432 34940 28484
rect 38476 28432 38528 28484
rect 33048 28364 33100 28416
rect 38384 28364 38436 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 36912 28160 36964 28212
rect 2596 28024 2648 28076
rect 1860 27999 1912 28008
rect 1860 27965 1869 27999
rect 1869 27965 1903 27999
rect 1903 27965 1912 27999
rect 1860 27956 1912 27965
rect 2412 27888 2464 27940
rect 26976 27956 27028 28008
rect 27160 27956 27212 28008
rect 27804 27956 27856 28008
rect 28540 27956 28592 28008
rect 33140 27999 33192 28008
rect 26884 27820 26936 27872
rect 33140 27965 33149 27999
rect 33149 27965 33183 27999
rect 33183 27965 33192 27999
rect 33140 27956 33192 27965
rect 36912 27956 36964 28008
rect 37464 27999 37516 28008
rect 37464 27965 37473 27999
rect 37473 27965 37507 27999
rect 37507 27965 37516 27999
rect 37464 27956 37516 27965
rect 38016 27956 38068 28008
rect 32956 27888 33008 27940
rect 38936 27888 38988 27940
rect 33508 27820 33560 27872
rect 33600 27820 33652 27872
rect 34152 27820 34204 27872
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 33140 27616 33192 27668
rect 1860 27523 1912 27532
rect 1860 27489 1869 27523
rect 1869 27489 1903 27523
rect 1903 27489 1912 27523
rect 1860 27480 1912 27489
rect 27988 27591 28040 27600
rect 27988 27557 28018 27591
rect 28018 27557 28040 27591
rect 27988 27548 28040 27557
rect 32956 27548 33008 27600
rect 33600 27616 33652 27668
rect 35624 27548 35676 27600
rect 36360 27548 36412 27600
rect 28540 27480 28592 27532
rect 33048 27523 33100 27532
rect 33048 27489 33057 27523
rect 33057 27489 33091 27523
rect 33091 27489 33100 27523
rect 33048 27480 33100 27489
rect 37464 27548 37516 27600
rect 37188 27523 37240 27532
rect 27528 27412 27580 27464
rect 37188 27489 37197 27523
rect 37197 27489 37231 27523
rect 37231 27489 37240 27523
rect 37188 27480 37240 27489
rect 34244 27412 34296 27464
rect 34428 27412 34480 27464
rect 27804 27276 27856 27328
rect 28080 27276 28132 27328
rect 34244 27276 34296 27328
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 27988 27072 28040 27124
rect 31852 27115 31904 27124
rect 31852 27081 31861 27115
rect 31861 27081 31895 27115
rect 31895 27081 31904 27115
rect 31852 27072 31904 27081
rect 2688 26936 2740 26988
rect 26884 26979 26936 26988
rect 26884 26945 26893 26979
rect 26893 26945 26927 26979
rect 26927 26945 26936 26979
rect 26884 26936 26936 26945
rect 29920 26936 29972 26988
rect 36912 27004 36964 27056
rect 37188 27004 37240 27056
rect 9588 26868 9640 26920
rect 25412 26868 25464 26920
rect 1860 26843 1912 26852
rect 1860 26809 1869 26843
rect 1869 26809 1903 26843
rect 1903 26809 1912 26843
rect 1860 26800 1912 26809
rect 2596 26800 2648 26852
rect 26976 26868 27028 26920
rect 27528 26868 27580 26920
rect 31392 26868 31444 26920
rect 32772 26911 32824 26920
rect 32772 26877 32781 26911
rect 32781 26877 32815 26911
rect 32815 26877 32824 26911
rect 32772 26868 32824 26877
rect 33140 26911 33192 26920
rect 33140 26877 33149 26911
rect 33149 26877 33183 26911
rect 33183 26877 33192 26911
rect 33140 26868 33192 26877
rect 37556 26868 37608 26920
rect 37924 26911 37976 26920
rect 37924 26877 37933 26911
rect 37933 26877 37967 26911
rect 37967 26877 37976 26911
rect 37924 26868 37976 26877
rect 27160 26800 27212 26852
rect 32956 26800 33008 26852
rect 32772 26732 32824 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 4068 26528 4120 26580
rect 33140 26528 33192 26580
rect 28080 26392 28132 26444
rect 32680 26392 32732 26444
rect 36176 26460 36228 26512
rect 36636 26528 36688 26580
rect 37832 26460 37884 26512
rect 25228 26324 25280 26376
rect 25412 26324 25464 26376
rect 26056 26324 26108 26376
rect 32956 26324 33008 26376
rect 34244 26435 34296 26444
rect 34244 26401 34254 26435
rect 34254 26401 34288 26435
rect 34288 26401 34296 26435
rect 34244 26392 34296 26401
rect 37372 26435 37424 26444
rect 33416 26256 33468 26308
rect 33324 26188 33376 26240
rect 34336 26324 34388 26376
rect 34152 26256 34204 26308
rect 34796 26324 34848 26376
rect 37372 26401 37381 26435
rect 37381 26401 37415 26435
rect 37415 26401 37424 26435
rect 37372 26392 37424 26401
rect 38660 26324 38712 26376
rect 34612 26256 34664 26308
rect 34796 26231 34848 26240
rect 34796 26197 34805 26231
rect 34805 26197 34839 26231
rect 34839 26197 34848 26231
rect 34796 26188 34848 26197
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 32312 25916 32364 25968
rect 32680 25916 32732 25968
rect 33048 25916 33100 25968
rect 32220 25848 32272 25900
rect 34428 25848 34480 25900
rect 1860 25823 1912 25832
rect 1860 25789 1869 25823
rect 1869 25789 1903 25823
rect 1903 25789 1912 25823
rect 1860 25780 1912 25789
rect 32496 25780 32548 25832
rect 33140 25823 33192 25832
rect 2688 25712 2740 25764
rect 33140 25789 33149 25823
rect 33149 25789 33183 25823
rect 33183 25789 33192 25823
rect 33140 25780 33192 25789
rect 34980 25780 35032 25832
rect 36176 25823 36228 25832
rect 2412 25644 2464 25696
rect 32956 25712 33008 25764
rect 35164 25712 35216 25764
rect 36176 25789 36185 25823
rect 36185 25789 36219 25823
rect 36219 25789 36228 25823
rect 36176 25780 36228 25789
rect 36360 25780 36412 25832
rect 37280 25823 37332 25832
rect 37280 25789 37289 25823
rect 37289 25789 37323 25823
rect 37323 25789 37332 25823
rect 37280 25780 37332 25789
rect 37924 25823 37976 25832
rect 37924 25789 37933 25823
rect 37933 25789 37967 25823
rect 37967 25789 37976 25823
rect 37924 25780 37976 25789
rect 35624 25644 35676 25696
rect 36636 25712 36688 25764
rect 36912 25712 36964 25764
rect 37096 25712 37148 25764
rect 38384 25644 38436 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 37372 25483 37424 25492
rect 32956 25372 33008 25424
rect 33324 25415 33376 25424
rect 33324 25381 33333 25415
rect 33333 25381 33367 25415
rect 33367 25381 33376 25415
rect 33324 25372 33376 25381
rect 34244 25372 34296 25424
rect 1860 25347 1912 25356
rect 1860 25313 1869 25347
rect 1869 25313 1903 25347
rect 1903 25313 1912 25347
rect 1860 25304 1912 25313
rect 32588 25304 32640 25356
rect 10324 25236 10376 25288
rect 34152 25304 34204 25356
rect 35164 25372 35216 25424
rect 34428 25347 34480 25356
rect 34428 25313 34437 25347
rect 34437 25313 34471 25347
rect 34471 25313 34480 25347
rect 34428 25304 34480 25313
rect 34704 25347 34756 25356
rect 34704 25313 34713 25347
rect 34713 25313 34747 25347
rect 34747 25313 34756 25347
rect 34704 25304 34756 25313
rect 35716 25347 35768 25356
rect 35716 25313 35725 25347
rect 35725 25313 35759 25347
rect 35759 25313 35768 25347
rect 36360 25347 36412 25356
rect 35716 25304 35768 25313
rect 36360 25313 36369 25347
rect 36369 25313 36403 25347
rect 36403 25313 36412 25347
rect 36360 25304 36412 25313
rect 36544 25372 36596 25424
rect 37372 25449 37381 25483
rect 37381 25449 37415 25483
rect 37415 25449 37424 25483
rect 37372 25440 37424 25449
rect 38752 25372 38804 25424
rect 37188 25347 37240 25356
rect 2596 25100 2648 25152
rect 33140 25168 33192 25220
rect 33324 25168 33376 25220
rect 34428 25168 34480 25220
rect 35900 25236 35952 25288
rect 36544 25236 36596 25288
rect 35716 25168 35768 25220
rect 37188 25313 37197 25347
rect 37197 25313 37231 25347
rect 37231 25313 37240 25347
rect 37188 25304 37240 25313
rect 34244 25100 34296 25152
rect 34520 25100 34572 25152
rect 35900 25100 35952 25152
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 32864 24828 32916 24880
rect 33692 24828 33744 24880
rect 35716 24828 35768 24880
rect 27160 24803 27212 24812
rect 27160 24769 27169 24803
rect 27169 24769 27203 24803
rect 27203 24769 27212 24803
rect 27160 24760 27212 24769
rect 27620 24692 27672 24744
rect 27896 24692 27948 24744
rect 32404 24692 32456 24744
rect 32956 24735 33008 24744
rect 32956 24701 32966 24735
rect 32966 24701 33000 24735
rect 33000 24701 33008 24735
rect 34152 24760 34204 24812
rect 32956 24692 33008 24701
rect 33692 24692 33744 24744
rect 2688 24624 2740 24676
rect 34520 24624 34572 24676
rect 35256 24624 35308 24676
rect 27528 24556 27580 24608
rect 32588 24556 32640 24608
rect 34152 24556 34204 24608
rect 36176 24828 36228 24880
rect 36268 24735 36320 24744
rect 36268 24701 36277 24735
rect 36277 24701 36311 24735
rect 36311 24701 36320 24735
rect 37280 24735 37332 24744
rect 36268 24692 36320 24701
rect 37280 24701 37289 24735
rect 37289 24701 37323 24735
rect 37323 24701 37332 24735
rect 37280 24692 37332 24701
rect 37924 24735 37976 24744
rect 37924 24701 37933 24735
rect 37933 24701 37967 24735
rect 37967 24701 37976 24735
rect 37924 24692 37976 24701
rect 37096 24624 37148 24676
rect 36176 24556 36228 24608
rect 36268 24556 36320 24608
rect 36820 24556 36872 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 29920 24352 29972 24404
rect 34244 24352 34296 24404
rect 35256 24352 35308 24404
rect 37188 24395 37240 24404
rect 37188 24361 37197 24395
rect 37197 24361 37231 24395
rect 37231 24361 37240 24395
rect 37188 24352 37240 24361
rect 27620 24284 27672 24336
rect 1860 24259 1912 24268
rect 1860 24225 1869 24259
rect 1869 24225 1903 24259
rect 1903 24225 1912 24259
rect 1860 24216 1912 24225
rect 27160 24216 27212 24268
rect 31852 24284 31904 24336
rect 32404 24284 32456 24336
rect 27896 24148 27948 24200
rect 28632 24216 28684 24268
rect 32956 24216 33008 24268
rect 38292 24284 38344 24336
rect 29092 24191 29144 24200
rect 29092 24157 29101 24191
rect 29101 24157 29135 24191
rect 29135 24157 29144 24191
rect 29092 24148 29144 24157
rect 33140 24148 33192 24200
rect 35716 24216 35768 24268
rect 36084 24216 36136 24268
rect 37372 24259 37424 24268
rect 37372 24225 37381 24259
rect 37381 24225 37415 24259
rect 37415 24225 37424 24259
rect 37372 24216 37424 24225
rect 27528 24080 27580 24132
rect 32128 24080 32180 24132
rect 34336 24080 34388 24132
rect 35164 24080 35216 24132
rect 36084 24080 36136 24132
rect 20996 24012 21048 24064
rect 27252 24012 27304 24064
rect 31944 24012 31996 24064
rect 33692 24012 33744 24064
rect 38016 24012 38068 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 9036 23808 9088 23860
rect 31852 23808 31904 23860
rect 34428 23808 34480 23860
rect 35716 23808 35768 23860
rect 37188 23808 37240 23860
rect 28540 23740 28592 23792
rect 32956 23740 33008 23792
rect 28724 23672 28776 23724
rect 27252 23647 27304 23656
rect 27252 23613 27261 23647
rect 27261 23613 27295 23647
rect 27295 23613 27304 23647
rect 27252 23604 27304 23613
rect 27896 23647 27948 23656
rect 1860 23579 1912 23588
rect 1860 23545 1869 23579
rect 1869 23545 1903 23579
rect 1903 23545 1912 23579
rect 1860 23536 1912 23545
rect 26148 23536 26200 23588
rect 27896 23613 27905 23647
rect 27905 23613 27939 23647
rect 27939 23613 27948 23647
rect 27896 23604 27948 23613
rect 29092 23604 29144 23656
rect 35900 23740 35952 23792
rect 34244 23672 34296 23724
rect 34980 23672 35032 23724
rect 35256 23604 35308 23656
rect 36084 23672 36136 23724
rect 35624 23536 35676 23588
rect 26700 23468 26752 23520
rect 27988 23511 28040 23520
rect 27988 23477 27997 23511
rect 27997 23477 28031 23511
rect 28031 23477 28040 23511
rect 27988 23468 28040 23477
rect 33140 23511 33192 23520
rect 33140 23477 33149 23511
rect 33149 23477 33183 23511
rect 33183 23477 33192 23511
rect 33140 23468 33192 23477
rect 35716 23511 35768 23520
rect 35716 23477 35725 23511
rect 35725 23477 35759 23511
rect 35759 23477 35768 23511
rect 35716 23468 35768 23477
rect 36176 23647 36228 23656
rect 36176 23613 36185 23647
rect 36185 23613 36219 23647
rect 36219 23613 36228 23647
rect 36176 23604 36228 23613
rect 36452 23604 36504 23656
rect 37280 23647 37332 23656
rect 37280 23613 37289 23647
rect 37289 23613 37323 23647
rect 37323 23613 37332 23647
rect 37280 23604 37332 23613
rect 37924 23647 37976 23656
rect 37924 23613 37933 23647
rect 37933 23613 37967 23647
rect 37967 23613 37976 23647
rect 37924 23604 37976 23613
rect 36820 23536 36872 23588
rect 35900 23468 35952 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 27896 23264 27948 23316
rect 30288 23264 30340 23316
rect 27988 23196 28040 23248
rect 32496 23196 32548 23248
rect 34152 23196 34204 23248
rect 28356 23128 28408 23180
rect 33324 23171 33376 23180
rect 33324 23137 33333 23171
rect 33333 23137 33367 23171
rect 33367 23137 33376 23171
rect 33324 23128 33376 23137
rect 27436 23060 27488 23112
rect 32956 23060 33008 23112
rect 33692 23128 33744 23180
rect 34980 23196 35032 23248
rect 34612 23171 34664 23180
rect 34612 23137 34621 23171
rect 34621 23137 34655 23171
rect 34655 23137 34664 23171
rect 34612 23128 34664 23137
rect 27804 22924 27856 22976
rect 31484 22992 31536 23044
rect 33324 22992 33376 23044
rect 35348 22992 35400 23044
rect 32956 22924 33008 22976
rect 33692 22924 33744 22976
rect 33876 22924 33928 22976
rect 34612 22924 34664 22976
rect 36176 23060 36228 23112
rect 36084 22992 36136 23044
rect 37372 22924 37424 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 27436 22720 27488 22772
rect 32220 22720 32272 22772
rect 31852 22652 31904 22704
rect 32496 22652 32548 22704
rect 1860 22559 1912 22568
rect 1860 22525 1869 22559
rect 1869 22525 1903 22559
rect 1903 22525 1912 22559
rect 1860 22516 1912 22525
rect 26700 22559 26752 22568
rect 26700 22525 26734 22559
rect 26734 22525 26752 22559
rect 26700 22516 26752 22525
rect 31852 22516 31904 22568
rect 32036 22559 32088 22568
rect 32036 22525 32045 22559
rect 32045 22525 32079 22559
rect 32079 22525 32088 22559
rect 32036 22516 32088 22525
rect 32680 22584 32732 22636
rect 36544 22720 36596 22772
rect 37464 22763 37516 22772
rect 32496 22516 32548 22568
rect 33324 22516 33376 22568
rect 34060 22652 34112 22704
rect 34152 22652 34204 22704
rect 35072 22652 35124 22704
rect 35716 22652 35768 22704
rect 34428 22559 34480 22568
rect 34428 22525 34437 22559
rect 34437 22525 34471 22559
rect 34471 22525 34480 22559
rect 34428 22516 34480 22525
rect 35256 22516 35308 22568
rect 35716 22516 35768 22568
rect 36084 22584 36136 22636
rect 36544 22584 36596 22636
rect 36176 22559 36228 22568
rect 36176 22525 36185 22559
rect 36185 22525 36219 22559
rect 36219 22525 36228 22559
rect 36176 22516 36228 22525
rect 36728 22516 36780 22568
rect 14556 22380 14608 22432
rect 27620 22380 27672 22432
rect 32404 22380 32456 22432
rect 32864 22423 32916 22432
rect 32864 22389 32873 22423
rect 32873 22389 32907 22423
rect 32907 22389 32916 22423
rect 32864 22380 32916 22389
rect 36452 22448 36504 22500
rect 34336 22380 34388 22432
rect 34704 22380 34756 22432
rect 34888 22380 34940 22432
rect 36728 22380 36780 22432
rect 37464 22729 37473 22763
rect 37473 22729 37507 22763
rect 37507 22729 37516 22763
rect 37464 22720 37516 22729
rect 37280 22559 37332 22568
rect 37280 22525 37289 22559
rect 37289 22525 37323 22559
rect 37323 22525 37332 22559
rect 37280 22516 37332 22525
rect 37924 22559 37976 22568
rect 37924 22525 37933 22559
rect 37933 22525 37967 22559
rect 37967 22525 37976 22559
rect 37924 22516 37976 22525
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 1860 22151 1912 22160
rect 1860 22117 1869 22151
rect 1869 22117 1903 22151
rect 1903 22117 1912 22151
rect 1860 22108 1912 22117
rect 32496 22108 32548 22160
rect 33232 22083 33284 22092
rect 33232 22049 33241 22083
rect 33241 22049 33275 22083
rect 33275 22049 33284 22083
rect 33232 22040 33284 22049
rect 34428 22108 34480 22160
rect 30380 21972 30432 22024
rect 30564 21972 30616 22024
rect 34612 22040 34664 22092
rect 35072 22083 35124 22092
rect 35072 22049 35081 22083
rect 35081 22049 35115 22083
rect 35115 22049 35124 22083
rect 35072 22040 35124 22049
rect 36084 22176 36136 22228
rect 32128 21904 32180 21956
rect 34060 21904 34112 21956
rect 34612 21904 34664 21956
rect 35624 22040 35676 22092
rect 36728 22040 36780 22092
rect 38568 21972 38620 22024
rect 16672 21836 16724 21888
rect 33048 21879 33100 21888
rect 33048 21845 33057 21879
rect 33057 21845 33091 21879
rect 33091 21845 33100 21879
rect 33048 21836 33100 21845
rect 33692 21836 33744 21888
rect 35900 21879 35952 21888
rect 35900 21845 35909 21879
rect 35909 21845 35943 21879
rect 35943 21845 35952 21879
rect 35900 21836 35952 21845
rect 36176 21904 36228 21956
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 31392 21632 31444 21684
rect 32772 21632 32824 21684
rect 37556 21632 37608 21684
rect 32312 21564 32364 21616
rect 34612 21564 34664 21616
rect 32036 21496 32088 21548
rect 37188 21564 37240 21616
rect 35256 21496 35308 21548
rect 38476 21496 38528 21548
rect 31760 21428 31812 21480
rect 32220 21471 32272 21480
rect 32220 21437 32229 21471
rect 32229 21437 32263 21471
rect 32263 21437 32272 21471
rect 32220 21428 32272 21437
rect 32496 21428 32548 21480
rect 37280 21471 37332 21480
rect 37280 21437 37289 21471
rect 37289 21437 37323 21471
rect 37323 21437 37332 21471
rect 37280 21428 37332 21437
rect 37924 21471 37976 21480
rect 37924 21437 37933 21471
rect 37933 21437 37967 21471
rect 37967 21437 37976 21471
rect 37924 21428 37976 21437
rect 34060 21360 34112 21412
rect 36728 21360 36780 21412
rect 31484 21292 31536 21344
rect 31760 21292 31812 21344
rect 33324 21292 33376 21344
rect 34336 21292 34388 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 1860 20995 1912 21004
rect 1860 20961 1869 20995
rect 1869 20961 1903 20995
rect 1903 20961 1912 20995
rect 1860 20952 1912 20961
rect 35900 21088 35952 21140
rect 31392 20952 31444 21004
rect 31668 21020 31720 21072
rect 32312 21020 32364 21072
rect 33140 21020 33192 21072
rect 32220 20952 32272 21004
rect 31024 20884 31076 20936
rect 32496 20952 32548 21004
rect 32772 20952 32824 21004
rect 35348 20995 35400 21004
rect 30472 20816 30524 20868
rect 31392 20816 31444 20868
rect 32220 20816 32272 20868
rect 32312 20816 32364 20868
rect 17132 20748 17184 20800
rect 30288 20791 30340 20800
rect 30288 20757 30297 20791
rect 30297 20757 30331 20791
rect 30331 20757 30340 20791
rect 30288 20748 30340 20757
rect 31024 20748 31076 20800
rect 31760 20791 31812 20800
rect 31760 20757 31769 20791
rect 31769 20757 31803 20791
rect 31803 20757 31812 20791
rect 31760 20748 31812 20757
rect 32496 20748 32548 20800
rect 32956 20748 33008 20800
rect 34244 20748 34296 20800
rect 34520 20748 34572 20800
rect 35348 20961 35357 20995
rect 35357 20961 35391 20995
rect 35391 20961 35400 20995
rect 35348 20952 35400 20961
rect 35440 20995 35492 21004
rect 35440 20961 35449 20995
rect 35449 20961 35483 20995
rect 35483 20961 35492 20995
rect 35440 20952 35492 20961
rect 36176 20995 36228 21004
rect 36176 20961 36185 20995
rect 36185 20961 36219 20995
rect 36219 20961 36228 20995
rect 36176 20952 36228 20961
rect 36912 20952 36964 21004
rect 37188 20995 37240 21004
rect 37188 20961 37197 20995
rect 37197 20961 37231 20995
rect 37231 20961 37240 20995
rect 37188 20952 37240 20961
rect 35900 20859 35952 20868
rect 35900 20825 35909 20859
rect 35909 20825 35943 20859
rect 35943 20825 35952 20859
rect 35900 20816 35952 20825
rect 38476 20884 38528 20936
rect 36176 20816 36228 20868
rect 37464 20748 37516 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 27160 20544 27212 20596
rect 27436 20544 27488 20596
rect 29552 20476 29604 20528
rect 27436 20383 27488 20392
rect 27436 20349 27445 20383
rect 27445 20349 27479 20383
rect 27479 20349 27488 20383
rect 27436 20340 27488 20349
rect 27896 20383 27948 20392
rect 27896 20349 27905 20383
rect 27905 20349 27939 20383
rect 27939 20349 27948 20383
rect 27896 20340 27948 20349
rect 1860 20315 1912 20324
rect 1860 20281 1869 20315
rect 1869 20281 1903 20315
rect 1903 20281 1912 20315
rect 1860 20272 1912 20281
rect 28540 20340 28592 20392
rect 30932 20476 30984 20528
rect 34520 20544 34572 20596
rect 31208 20476 31260 20528
rect 33232 20476 33284 20528
rect 36084 20476 36136 20528
rect 31668 20451 31720 20460
rect 31668 20417 31677 20451
rect 31677 20417 31711 20451
rect 31711 20417 31720 20451
rect 31668 20408 31720 20417
rect 31392 20340 31444 20392
rect 28816 20315 28868 20324
rect 17224 20204 17276 20256
rect 23572 20204 23624 20256
rect 25504 20204 25556 20256
rect 28816 20281 28825 20315
rect 28825 20281 28859 20315
rect 28859 20281 28868 20315
rect 28816 20272 28868 20281
rect 34244 20408 34296 20460
rect 31944 20383 31996 20392
rect 31944 20349 31978 20383
rect 31978 20349 31996 20383
rect 31944 20340 31996 20349
rect 33232 20340 33284 20392
rect 36176 20408 36228 20460
rect 34796 20383 34848 20392
rect 32220 20272 32272 20324
rect 29460 20204 29512 20256
rect 30380 20204 30432 20256
rect 31392 20204 31444 20256
rect 31668 20204 31720 20256
rect 31944 20204 31996 20256
rect 32312 20204 32364 20256
rect 32772 20204 32824 20256
rect 33324 20204 33376 20256
rect 34244 20247 34296 20256
rect 34244 20213 34253 20247
rect 34253 20213 34287 20247
rect 34287 20213 34296 20247
rect 34244 20204 34296 20213
rect 34796 20349 34805 20383
rect 34805 20349 34839 20383
rect 34839 20349 34848 20383
rect 34796 20340 34848 20349
rect 36084 20340 36136 20392
rect 36728 20340 36780 20392
rect 37924 20383 37976 20392
rect 37924 20349 37933 20383
rect 37933 20349 37967 20383
rect 37967 20349 37976 20383
rect 37924 20340 37976 20349
rect 35348 20272 35400 20324
rect 34796 20204 34848 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 26056 19932 26108 19984
rect 25780 19864 25832 19916
rect 27620 19864 27672 19916
rect 27896 19907 27948 19916
rect 27896 19873 27905 19907
rect 27905 19873 27939 19907
rect 27939 19873 27948 19907
rect 27896 19864 27948 19873
rect 28264 19864 28316 19916
rect 37832 20000 37884 20052
rect 29644 19932 29696 19984
rect 26976 19796 27028 19848
rect 29736 19907 29788 19916
rect 29736 19873 29745 19907
rect 29745 19873 29779 19907
rect 29779 19873 29788 19907
rect 29736 19864 29788 19873
rect 34244 19932 34296 19984
rect 34520 19932 34572 19984
rect 30748 19907 30800 19916
rect 27528 19728 27580 19780
rect 29000 19796 29052 19848
rect 29644 19796 29696 19848
rect 30748 19873 30757 19907
rect 30757 19873 30791 19907
rect 30791 19873 30800 19907
rect 30748 19864 30800 19873
rect 30932 19864 30984 19916
rect 31392 19864 31444 19916
rect 28908 19728 28960 19780
rect 32220 19864 32272 19916
rect 33876 19864 33928 19916
rect 28540 19703 28592 19712
rect 28540 19669 28549 19703
rect 28549 19669 28583 19703
rect 28583 19669 28592 19703
rect 28540 19660 28592 19669
rect 28632 19660 28684 19712
rect 29460 19660 29512 19712
rect 29736 19660 29788 19712
rect 31668 19728 31720 19780
rect 35348 19907 35400 19916
rect 34520 19796 34572 19848
rect 35348 19873 35357 19907
rect 35357 19873 35391 19907
rect 35391 19873 35400 19907
rect 35348 19864 35400 19873
rect 35808 19864 35860 19916
rect 35900 19864 35952 19916
rect 36544 19932 36596 19984
rect 37188 19907 37240 19916
rect 37188 19873 37197 19907
rect 37197 19873 37231 19907
rect 37231 19873 37240 19907
rect 37188 19864 37240 19873
rect 37832 19796 37884 19848
rect 30564 19703 30616 19712
rect 30564 19669 30573 19703
rect 30573 19669 30607 19703
rect 30607 19669 30616 19703
rect 30564 19660 30616 19669
rect 31024 19703 31076 19712
rect 31024 19669 31033 19703
rect 31033 19669 31067 19703
rect 31067 19669 31076 19703
rect 31024 19660 31076 19669
rect 32864 19660 32916 19712
rect 33232 19660 33284 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 26792 19456 26844 19508
rect 27068 19499 27120 19508
rect 27068 19465 27077 19499
rect 27077 19465 27111 19499
rect 27111 19465 27120 19499
rect 27068 19456 27120 19465
rect 27436 19456 27488 19508
rect 31944 19456 31996 19508
rect 31668 19388 31720 19440
rect 32128 19388 32180 19440
rect 35072 19388 35124 19440
rect 1860 19295 1912 19304
rect 1860 19261 1869 19295
rect 1869 19261 1903 19295
rect 1903 19261 1912 19295
rect 1860 19252 1912 19261
rect 24124 19295 24176 19304
rect 9128 19184 9180 19236
rect 24124 19261 24133 19295
rect 24133 19261 24167 19295
rect 24167 19261 24176 19295
rect 24124 19252 24176 19261
rect 27344 19320 27396 19372
rect 32220 19320 32272 19372
rect 26148 19295 26200 19304
rect 26148 19261 26157 19295
rect 26157 19261 26191 19295
rect 26191 19261 26200 19295
rect 26148 19252 26200 19261
rect 26240 19252 26292 19304
rect 26976 19295 27028 19304
rect 26976 19261 26985 19295
rect 26985 19261 27019 19295
rect 27019 19261 27028 19295
rect 26976 19252 27028 19261
rect 30104 19252 30156 19304
rect 31852 19252 31904 19304
rect 25964 19227 26016 19236
rect 25964 19193 25973 19227
rect 25973 19193 26007 19227
rect 26007 19193 26016 19227
rect 25964 19184 26016 19193
rect 26056 19184 26108 19236
rect 27896 19184 27948 19236
rect 28448 19116 28500 19168
rect 29460 19184 29512 19236
rect 34520 19252 34572 19304
rect 33048 19184 33100 19236
rect 34704 19295 34756 19304
rect 34704 19261 34713 19295
rect 34713 19261 34747 19295
rect 34747 19261 34756 19295
rect 34704 19252 34756 19261
rect 35164 19252 35216 19304
rect 36084 19388 36136 19440
rect 37280 19295 37332 19304
rect 37280 19261 37289 19295
rect 37289 19261 37323 19295
rect 37323 19261 37332 19295
rect 37280 19252 37332 19261
rect 37924 19295 37976 19304
rect 37924 19261 37933 19295
rect 37933 19261 37967 19295
rect 37967 19261 37976 19295
rect 37924 19252 37976 19261
rect 31392 19116 31444 19168
rect 33692 19159 33744 19168
rect 33692 19125 33701 19159
rect 33701 19125 33735 19159
rect 33735 19125 33744 19159
rect 33692 19116 33744 19125
rect 35348 19116 35400 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 24124 18912 24176 18964
rect 28356 18912 28408 18964
rect 31760 18912 31812 18964
rect 31944 18955 31996 18964
rect 31944 18921 31953 18955
rect 31953 18921 31987 18955
rect 31987 18921 31996 18955
rect 31944 18912 31996 18921
rect 25504 18844 25556 18896
rect 1860 18819 1912 18828
rect 1860 18785 1869 18819
rect 1869 18785 1903 18819
rect 1903 18785 1912 18819
rect 1860 18776 1912 18785
rect 1308 18708 1360 18760
rect 26056 18776 26108 18828
rect 26332 18819 26384 18828
rect 26332 18785 26341 18819
rect 26341 18785 26375 18819
rect 26375 18785 26384 18819
rect 26332 18776 26384 18785
rect 26608 18776 26660 18828
rect 26884 18776 26936 18828
rect 28080 18819 28132 18828
rect 28080 18785 28089 18819
rect 28089 18785 28123 18819
rect 28123 18785 28132 18819
rect 28080 18776 28132 18785
rect 28448 18819 28500 18828
rect 24676 18751 24728 18760
rect 24676 18717 24685 18751
rect 24685 18717 24719 18751
rect 24719 18717 24728 18751
rect 24676 18708 24728 18717
rect 28448 18785 28457 18819
rect 28457 18785 28491 18819
rect 28491 18785 28500 18819
rect 28448 18776 28500 18785
rect 30472 18844 30524 18896
rect 33140 18912 33192 18964
rect 34152 18912 34204 18964
rect 34888 18912 34940 18964
rect 36084 18912 36136 18964
rect 37740 18912 37792 18964
rect 32956 18844 33008 18896
rect 34520 18844 34572 18896
rect 34704 18844 34756 18896
rect 29920 18776 29972 18828
rect 30196 18776 30248 18828
rect 28724 18708 28776 18760
rect 27160 18640 27212 18692
rect 30472 18708 30524 18760
rect 31392 18776 31444 18828
rect 32220 18776 32272 18828
rect 32680 18708 32732 18760
rect 34060 18776 34112 18828
rect 35900 18844 35952 18896
rect 36176 18887 36228 18896
rect 36176 18853 36185 18887
rect 36185 18853 36219 18887
rect 36219 18853 36228 18887
rect 36176 18844 36228 18853
rect 35348 18819 35400 18828
rect 35348 18785 35357 18819
rect 35357 18785 35391 18819
rect 35391 18785 35400 18819
rect 35348 18776 35400 18785
rect 35532 18776 35584 18828
rect 37188 18819 37240 18828
rect 37188 18785 37197 18819
rect 37197 18785 37231 18819
rect 37231 18785 37240 18819
rect 37188 18776 37240 18785
rect 36912 18708 36964 18760
rect 18328 18572 18380 18624
rect 24768 18572 24820 18624
rect 24952 18572 25004 18624
rect 26424 18572 26476 18624
rect 26608 18615 26660 18624
rect 26608 18581 26617 18615
rect 26617 18581 26651 18615
rect 26651 18581 26660 18615
rect 26608 18572 26660 18581
rect 27252 18572 27304 18624
rect 30104 18572 30156 18624
rect 30932 18572 30984 18624
rect 31392 18572 31444 18624
rect 34060 18640 34112 18692
rect 35164 18640 35216 18692
rect 31944 18572 31996 18624
rect 35440 18572 35492 18624
rect 35808 18572 35860 18624
rect 37556 18572 37608 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 26424 18368 26476 18420
rect 28356 18368 28408 18420
rect 28264 18300 28316 18352
rect 31944 18368 31996 18420
rect 29552 18300 29604 18352
rect 25228 18275 25280 18284
rect 25228 18241 25237 18275
rect 25237 18241 25271 18275
rect 25271 18241 25280 18275
rect 25228 18232 25280 18241
rect 23388 18096 23440 18148
rect 26608 18164 26660 18216
rect 27160 18164 27212 18216
rect 27620 18164 27672 18216
rect 28724 18164 28776 18216
rect 29368 18232 29420 18284
rect 25504 18139 25556 18148
rect 25504 18105 25538 18139
rect 25538 18105 25556 18139
rect 25504 18096 25556 18105
rect 26792 18096 26844 18148
rect 27436 18096 27488 18148
rect 29644 18164 29696 18216
rect 32220 18300 32272 18352
rect 33324 18300 33376 18352
rect 33876 18300 33928 18352
rect 32404 18164 32456 18216
rect 33876 18164 33928 18216
rect 34704 18300 34756 18352
rect 29460 18096 29512 18148
rect 23848 18028 23900 18080
rect 28080 18028 28132 18080
rect 29092 18028 29144 18080
rect 30932 18096 30984 18148
rect 34520 18164 34572 18216
rect 35348 18232 35400 18284
rect 34704 18207 34756 18216
rect 34704 18173 34713 18207
rect 34713 18173 34747 18207
rect 34747 18173 34756 18207
rect 34704 18164 34756 18173
rect 34888 18164 34940 18216
rect 37280 18207 37332 18216
rect 37280 18173 37289 18207
rect 37289 18173 37323 18207
rect 37323 18173 37332 18207
rect 37280 18164 37332 18173
rect 37924 18207 37976 18216
rect 37924 18173 37933 18207
rect 37933 18173 37967 18207
rect 37967 18173 37976 18207
rect 37924 18164 37976 18173
rect 31484 18028 31536 18080
rect 32036 18028 32088 18080
rect 32588 18028 32640 18080
rect 33048 18028 33100 18080
rect 34704 18028 34756 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 24768 17824 24820 17876
rect 28264 17824 28316 17876
rect 28908 17824 28960 17876
rect 29368 17824 29420 17876
rect 1860 17799 1912 17808
rect 1860 17765 1869 17799
rect 1869 17765 1903 17799
rect 1903 17765 1912 17799
rect 1860 17756 1912 17765
rect 23848 17799 23900 17808
rect 23848 17765 23882 17799
rect 23882 17765 23900 17799
rect 23848 17756 23900 17765
rect 23940 17756 23992 17808
rect 25228 17756 25280 17808
rect 26884 17756 26936 17808
rect 29000 17756 29052 17808
rect 30380 17756 30432 17808
rect 31852 17756 31904 17808
rect 25228 17620 25280 17672
rect 16304 17484 16356 17536
rect 24308 17484 24360 17536
rect 30748 17688 30800 17740
rect 34060 17824 34112 17876
rect 34428 17867 34480 17876
rect 34428 17833 34437 17867
rect 34437 17833 34471 17867
rect 34471 17833 34480 17867
rect 34428 17824 34480 17833
rect 32496 17756 32548 17808
rect 34612 17756 34664 17808
rect 27160 17620 27212 17672
rect 27804 17663 27856 17672
rect 27804 17629 27813 17663
rect 27813 17629 27847 17663
rect 27847 17629 27856 17663
rect 27804 17620 27856 17629
rect 27804 17484 27856 17536
rect 32220 17688 32272 17740
rect 33140 17688 33192 17740
rect 34888 17688 34940 17740
rect 35072 17731 35124 17740
rect 35072 17697 35081 17731
rect 35081 17697 35115 17731
rect 35115 17697 35124 17731
rect 35072 17688 35124 17697
rect 29644 17484 29696 17536
rect 34520 17620 34572 17672
rect 35716 17688 35768 17740
rect 31392 17552 31444 17604
rect 30748 17484 30800 17536
rect 31208 17484 31260 17536
rect 31760 17484 31812 17536
rect 35072 17552 35124 17604
rect 35348 17552 35400 17604
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 24676 17280 24728 17332
rect 27436 17280 27488 17332
rect 25228 17187 25280 17196
rect 25228 17153 25237 17187
rect 25237 17153 25271 17187
rect 25271 17153 25280 17187
rect 25228 17144 25280 17153
rect 25136 17076 25188 17128
rect 25964 17076 26016 17128
rect 27160 17076 27212 17128
rect 29000 17076 29052 17128
rect 29276 17212 29328 17264
rect 31484 17280 31536 17332
rect 38660 17280 38712 17332
rect 29460 17187 29512 17196
rect 29460 17153 29469 17187
rect 29469 17153 29503 17187
rect 29503 17153 29512 17187
rect 29460 17144 29512 17153
rect 1860 17051 1912 17060
rect 1860 17017 1869 17051
rect 1869 17017 1903 17051
rect 1903 17017 1912 17051
rect 1860 17008 1912 17017
rect 24124 17051 24176 17060
rect 24124 17017 24133 17051
rect 24133 17017 24167 17051
rect 24167 17017 24176 17051
rect 24124 17008 24176 17017
rect 24768 17008 24820 17060
rect 26424 17008 26476 17060
rect 17500 16940 17552 16992
rect 24860 16940 24912 16992
rect 29000 16983 29052 16992
rect 29000 16949 29009 16983
rect 29009 16949 29043 16983
rect 29043 16949 29052 16983
rect 29000 16940 29052 16949
rect 29644 17076 29696 17128
rect 30380 17076 30432 17128
rect 31208 17076 31260 17128
rect 30288 17008 30340 17060
rect 30932 16940 30984 16992
rect 36544 17212 36596 17264
rect 37096 17212 37148 17264
rect 32128 17144 32180 17196
rect 32312 17119 32364 17128
rect 32312 17085 32321 17119
rect 32321 17085 32355 17119
rect 32355 17085 32364 17119
rect 32312 17076 32364 17085
rect 31852 17008 31904 17060
rect 33048 17008 33100 17060
rect 34152 17076 34204 17128
rect 34520 17144 34572 17196
rect 36636 17144 36688 17196
rect 36820 17144 36872 17196
rect 34336 17119 34388 17128
rect 34336 17085 34345 17119
rect 34345 17085 34379 17119
rect 34379 17085 34388 17119
rect 37280 17119 37332 17128
rect 34336 17076 34388 17085
rect 37280 17085 37289 17119
rect 37289 17085 37323 17119
rect 37323 17085 37332 17119
rect 37280 17076 37332 17085
rect 37924 17119 37976 17128
rect 37924 17085 37933 17119
rect 37933 17085 37967 17119
rect 37967 17085 37976 17119
rect 37924 17076 37976 17085
rect 34704 17008 34756 17060
rect 37556 16940 37608 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 24676 16668 24728 16720
rect 24032 16643 24084 16652
rect 24032 16609 24041 16643
rect 24041 16609 24075 16643
rect 24075 16609 24084 16643
rect 24032 16600 24084 16609
rect 24216 16643 24268 16652
rect 24216 16609 24225 16643
rect 24225 16609 24259 16643
rect 24259 16609 24268 16643
rect 24216 16600 24268 16609
rect 24308 16643 24360 16652
rect 24308 16609 24317 16643
rect 24317 16609 24351 16643
rect 24351 16609 24360 16643
rect 24308 16600 24360 16609
rect 24860 16600 24912 16652
rect 25504 16736 25556 16788
rect 26240 16668 26292 16720
rect 29276 16736 29328 16788
rect 31024 16779 31076 16788
rect 27896 16668 27948 16720
rect 28356 16668 28408 16720
rect 30564 16668 30616 16720
rect 31024 16745 31033 16779
rect 31033 16745 31067 16779
rect 31067 16745 31076 16779
rect 31024 16736 31076 16745
rect 31208 16736 31260 16788
rect 32220 16736 32272 16788
rect 27804 16643 27856 16652
rect 27804 16609 27813 16643
rect 27813 16609 27847 16643
rect 27847 16609 27856 16643
rect 27804 16600 27856 16609
rect 30380 16600 30432 16652
rect 31576 16600 31628 16652
rect 25044 16575 25096 16584
rect 25044 16541 25053 16575
rect 25053 16541 25087 16575
rect 25087 16541 25096 16575
rect 25044 16532 25096 16541
rect 31208 16532 31260 16584
rect 23480 16464 23532 16516
rect 24124 16464 24176 16516
rect 32312 16600 32364 16652
rect 22928 16396 22980 16448
rect 24676 16396 24728 16448
rect 28724 16396 28776 16448
rect 29644 16396 29696 16448
rect 31944 16439 31996 16448
rect 31944 16405 31953 16439
rect 31953 16405 31987 16439
rect 31987 16405 31996 16439
rect 31944 16396 31996 16405
rect 33324 16668 33376 16720
rect 34612 16736 34664 16788
rect 35716 16736 35768 16788
rect 36084 16736 36136 16788
rect 34152 16668 34204 16720
rect 34336 16600 34388 16652
rect 34612 16600 34664 16652
rect 34152 16532 34204 16584
rect 32588 16464 32640 16516
rect 34612 16396 34664 16448
rect 35256 16600 35308 16652
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 23848 16192 23900 16244
rect 25044 16056 25096 16108
rect 25412 16056 25464 16108
rect 25964 16192 26016 16244
rect 26792 16192 26844 16244
rect 29644 16192 29696 16244
rect 29920 16192 29972 16244
rect 33048 16192 33100 16244
rect 33784 16192 33836 16244
rect 38108 16192 38160 16244
rect 27528 16099 27580 16108
rect 27528 16065 27537 16099
rect 27537 16065 27571 16099
rect 27571 16065 27580 16099
rect 27528 16056 27580 16065
rect 30196 16124 30248 16176
rect 1860 16031 1912 16040
rect 1860 15997 1869 16031
rect 1869 15997 1903 16031
rect 1903 15997 1912 16031
rect 1860 15988 1912 15997
rect 22652 15988 22704 16040
rect 23940 15988 23992 16040
rect 24308 15988 24360 16040
rect 27436 15988 27488 16040
rect 23020 15920 23072 15972
rect 23848 15920 23900 15972
rect 28540 15988 28592 16040
rect 28724 15988 28776 16040
rect 30656 16031 30708 16040
rect 30656 15997 30665 16031
rect 30665 15997 30699 16031
rect 30699 15997 30708 16031
rect 30656 15988 30708 15997
rect 31208 16124 31260 16176
rect 32312 16056 32364 16108
rect 29920 15920 29972 15972
rect 16396 15852 16448 15904
rect 26240 15852 26292 15904
rect 27344 15852 27396 15904
rect 27436 15852 27488 15904
rect 28540 15852 28592 15904
rect 28632 15852 28684 15904
rect 30472 15895 30524 15904
rect 30472 15861 30481 15895
rect 30481 15861 30515 15895
rect 30515 15861 30524 15895
rect 30472 15852 30524 15861
rect 31208 15988 31260 16040
rect 31668 15988 31720 16040
rect 32404 16031 32456 16040
rect 32404 15997 32413 16031
rect 32413 15997 32447 16031
rect 32447 15997 32456 16031
rect 32404 15988 32456 15997
rect 33324 16056 33376 16108
rect 32772 16031 32824 16040
rect 31576 15963 31628 15972
rect 31576 15929 31585 15963
rect 31585 15929 31619 15963
rect 31619 15929 31628 15963
rect 31576 15920 31628 15929
rect 32772 15997 32781 16031
rect 32781 15997 32815 16031
rect 32815 15997 32824 16031
rect 32772 15988 32824 15997
rect 33048 15988 33100 16040
rect 34704 16124 34756 16176
rect 37280 16031 37332 16040
rect 33140 15920 33192 15972
rect 37280 15997 37289 16031
rect 37289 15997 37323 16031
rect 37323 15997 37332 16031
rect 37280 15988 37332 15997
rect 37924 16031 37976 16040
rect 37924 15997 37933 16031
rect 37933 15997 37967 16031
rect 37967 15997 37976 16031
rect 37924 15988 37976 15997
rect 33968 15920 34020 15972
rect 32588 15852 32640 15904
rect 33784 15852 33836 15904
rect 34612 15852 34664 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 22652 15648 22704 15700
rect 23664 15648 23716 15700
rect 1860 15555 1912 15564
rect 1860 15521 1869 15555
rect 1869 15521 1903 15555
rect 1903 15521 1912 15555
rect 1860 15512 1912 15521
rect 22928 15555 22980 15564
rect 22928 15521 22937 15555
rect 22937 15521 22971 15555
rect 22971 15521 22980 15555
rect 22928 15512 22980 15521
rect 23572 15555 23624 15564
rect 23572 15521 23581 15555
rect 23581 15521 23615 15555
rect 23615 15521 23624 15555
rect 23572 15512 23624 15521
rect 23848 15512 23900 15564
rect 32772 15648 32824 15700
rect 33324 15648 33376 15700
rect 24768 15580 24820 15632
rect 27896 15580 27948 15632
rect 29000 15580 29052 15632
rect 25412 15555 25464 15564
rect 24216 15444 24268 15496
rect 16120 15308 16172 15360
rect 23204 15308 23256 15360
rect 23848 15351 23900 15360
rect 23848 15317 23857 15351
rect 23857 15317 23891 15351
rect 23891 15317 23900 15351
rect 23848 15308 23900 15317
rect 24400 15351 24452 15360
rect 24400 15317 24409 15351
rect 24409 15317 24443 15351
rect 24443 15317 24452 15351
rect 24400 15308 24452 15317
rect 24860 15351 24912 15360
rect 24860 15317 24869 15351
rect 24869 15317 24903 15351
rect 24903 15317 24912 15351
rect 24860 15308 24912 15317
rect 25412 15521 25421 15555
rect 25421 15521 25455 15555
rect 25455 15521 25464 15555
rect 25412 15512 25464 15521
rect 28356 15512 28408 15564
rect 29828 15555 29880 15564
rect 29828 15521 29837 15555
rect 29837 15521 29871 15555
rect 29871 15521 29880 15555
rect 29828 15512 29880 15521
rect 31392 15580 31444 15632
rect 30196 15555 30248 15564
rect 30196 15521 30205 15555
rect 30205 15521 30239 15555
rect 30239 15521 30248 15555
rect 30196 15512 30248 15521
rect 30840 15555 30892 15564
rect 30840 15521 30849 15555
rect 30849 15521 30883 15555
rect 30883 15521 30892 15555
rect 30840 15512 30892 15521
rect 27528 15444 27580 15496
rect 27160 15376 27212 15428
rect 26608 15308 26660 15360
rect 28448 15308 28500 15360
rect 31852 15512 31904 15564
rect 32956 15512 33008 15564
rect 34060 15580 34112 15632
rect 34244 15580 34296 15632
rect 34336 15555 34388 15564
rect 32588 15444 32640 15496
rect 28908 15376 28960 15428
rect 31392 15376 31444 15428
rect 29000 15308 29052 15360
rect 29460 15308 29512 15360
rect 29736 15308 29788 15360
rect 33140 15351 33192 15360
rect 33140 15317 33149 15351
rect 33149 15317 33183 15351
rect 33183 15317 33192 15351
rect 33140 15308 33192 15317
rect 34336 15521 34345 15555
rect 34345 15521 34379 15555
rect 34379 15521 34388 15555
rect 34336 15512 34388 15521
rect 34612 15555 34664 15564
rect 34244 15376 34296 15428
rect 34612 15521 34621 15555
rect 34621 15521 34655 15555
rect 34655 15521 34664 15555
rect 34612 15512 34664 15521
rect 35624 15512 35676 15564
rect 37188 15555 37240 15564
rect 37188 15521 37197 15555
rect 37197 15521 37231 15555
rect 37231 15521 37240 15555
rect 37188 15512 37240 15521
rect 35440 15444 35492 15496
rect 35900 15376 35952 15428
rect 33784 15308 33836 15360
rect 33968 15308 34020 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 22836 14900 22888 14952
rect 23296 15036 23348 15088
rect 23940 15036 23992 15088
rect 24308 15036 24360 15088
rect 27896 15104 27948 15156
rect 28908 15104 28960 15156
rect 31668 15104 31720 15156
rect 32588 15104 32640 15156
rect 35900 15147 35952 15156
rect 35900 15113 35909 15147
rect 35909 15113 35943 15147
rect 35943 15113 35952 15147
rect 35900 15104 35952 15113
rect 23572 14900 23624 14952
rect 23756 14900 23808 14952
rect 24492 14968 24544 15020
rect 26608 14968 26660 15020
rect 32128 15036 32180 15088
rect 24216 14900 24268 14952
rect 26976 14900 27028 14952
rect 27344 14900 27396 14952
rect 27436 14900 27488 14952
rect 28908 14900 28960 14952
rect 29184 14943 29236 14952
rect 29184 14909 29193 14943
rect 29193 14909 29227 14943
rect 29227 14909 29236 14943
rect 29184 14900 29236 14909
rect 32772 14968 32824 15020
rect 36084 15036 36136 15088
rect 30196 14900 30248 14952
rect 14096 14832 14148 14884
rect 25320 14832 25372 14884
rect 30472 14832 30524 14884
rect 22744 14807 22796 14816
rect 22744 14773 22753 14807
rect 22753 14773 22787 14807
rect 22787 14773 22796 14807
rect 22744 14764 22796 14773
rect 23756 14807 23808 14816
rect 23756 14773 23765 14807
rect 23765 14773 23799 14807
rect 23799 14773 23808 14807
rect 23756 14764 23808 14773
rect 25688 14764 25740 14816
rect 26792 14764 26844 14816
rect 28356 14764 28408 14816
rect 31944 14807 31996 14816
rect 31944 14773 31953 14807
rect 31953 14773 31987 14807
rect 31987 14773 31996 14807
rect 31944 14764 31996 14773
rect 32312 14900 32364 14952
rect 32864 14900 32916 14952
rect 33324 14900 33376 14952
rect 33508 14943 33560 14952
rect 33508 14909 33517 14943
rect 33517 14909 33551 14943
rect 33551 14909 33560 14943
rect 35900 14968 35952 15020
rect 33508 14900 33560 14909
rect 34244 14943 34296 14952
rect 34244 14909 34253 14943
rect 34253 14909 34287 14943
rect 34287 14909 34296 14943
rect 34244 14900 34296 14909
rect 33784 14832 33836 14884
rect 35532 14900 35584 14952
rect 37924 14943 37976 14952
rect 37924 14909 37933 14943
rect 37933 14909 37967 14943
rect 37967 14909 37976 14943
rect 37924 14900 37976 14909
rect 34612 14832 34664 14884
rect 33508 14764 33560 14816
rect 34336 14764 34388 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 23480 14603 23532 14612
rect 23480 14569 23489 14603
rect 23489 14569 23523 14603
rect 23523 14569 23532 14603
rect 23480 14560 23532 14569
rect 23572 14560 23624 14612
rect 1860 14535 1912 14544
rect 1860 14501 1869 14535
rect 1869 14501 1903 14535
rect 1903 14501 1912 14535
rect 1860 14492 1912 14501
rect 14924 14492 14976 14544
rect 3056 14424 3108 14476
rect 23020 14424 23072 14476
rect 23480 14424 23532 14476
rect 18696 14356 18748 14408
rect 23664 14356 23716 14408
rect 15476 14220 15528 14272
rect 24308 14560 24360 14612
rect 24676 14424 24728 14476
rect 26240 14424 26292 14476
rect 26516 14467 26568 14476
rect 26516 14433 26525 14467
rect 26525 14433 26559 14467
rect 26559 14433 26568 14467
rect 26516 14424 26568 14433
rect 33140 14560 33192 14612
rect 27160 14492 27212 14544
rect 29368 14492 29420 14544
rect 29736 14535 29788 14544
rect 29736 14501 29745 14535
rect 29745 14501 29779 14535
rect 29779 14501 29788 14535
rect 29736 14492 29788 14501
rect 31576 14492 31628 14544
rect 29276 14424 29328 14476
rect 29920 14424 29972 14476
rect 27528 14356 27580 14408
rect 29184 14356 29236 14408
rect 30288 14356 30340 14408
rect 33324 14467 33376 14476
rect 33324 14433 33333 14467
rect 33333 14433 33367 14467
rect 33367 14433 33376 14467
rect 33784 14560 33836 14612
rect 34612 14560 34664 14612
rect 38016 14560 38068 14612
rect 33324 14424 33376 14433
rect 25320 14288 25372 14340
rect 24676 14220 24728 14272
rect 26332 14263 26384 14272
rect 26332 14229 26341 14263
rect 26341 14229 26375 14263
rect 26375 14229 26384 14263
rect 26332 14220 26384 14229
rect 26792 14263 26844 14272
rect 26792 14229 26801 14263
rect 26801 14229 26835 14263
rect 26835 14229 26844 14263
rect 26792 14220 26844 14229
rect 31852 14288 31904 14340
rect 32680 14288 32732 14340
rect 33232 14288 33284 14340
rect 33324 14288 33376 14340
rect 29184 14263 29236 14272
rect 29184 14229 29193 14263
rect 29193 14229 29227 14263
rect 29227 14229 29236 14263
rect 29184 14220 29236 14229
rect 33600 14467 33652 14476
rect 33600 14433 33609 14467
rect 33609 14433 33643 14467
rect 33643 14433 33652 14467
rect 33600 14424 33652 14433
rect 33784 14424 33836 14476
rect 34336 14467 34388 14476
rect 34336 14433 34345 14467
rect 34345 14433 34379 14467
rect 34379 14433 34388 14467
rect 34336 14424 34388 14433
rect 35716 14424 35768 14476
rect 37188 14467 37240 14476
rect 37188 14433 37197 14467
rect 37197 14433 37231 14467
rect 37231 14433 37240 14467
rect 37188 14424 37240 14433
rect 34060 14263 34112 14272
rect 34060 14229 34069 14263
rect 34069 14229 34103 14263
rect 34103 14229 34112 14263
rect 34060 14220 34112 14229
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 2228 14016 2280 14068
rect 22560 13880 22612 13932
rect 23572 14016 23624 14068
rect 23848 14016 23900 14068
rect 24308 14059 24360 14068
rect 24308 14025 24317 14059
rect 24317 14025 24351 14059
rect 24351 14025 24360 14059
rect 24308 14016 24360 14025
rect 24492 14016 24544 14068
rect 28448 14059 28500 14068
rect 26240 13948 26292 14000
rect 28448 14025 28457 14059
rect 28457 14025 28491 14059
rect 28491 14025 28500 14059
rect 28448 14016 28500 14025
rect 28540 14016 28592 14068
rect 33968 14016 34020 14068
rect 34336 14016 34388 14068
rect 38752 14016 38804 14068
rect 24032 13880 24084 13932
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 23204 13855 23256 13864
rect 23204 13821 23238 13855
rect 23238 13821 23256 13855
rect 23204 13812 23256 13821
rect 25228 13855 25280 13864
rect 25228 13821 25237 13855
rect 25237 13821 25271 13855
rect 25271 13821 25280 13855
rect 25228 13812 25280 13821
rect 28816 13880 28868 13932
rect 26240 13812 26292 13864
rect 27896 13812 27948 13864
rect 20904 13744 20956 13796
rect 21088 13676 21140 13728
rect 22284 13676 22336 13728
rect 22376 13676 22428 13728
rect 26516 13676 26568 13728
rect 26884 13744 26936 13796
rect 28264 13676 28316 13728
rect 28448 13676 28500 13728
rect 28724 13676 28776 13728
rect 29736 13812 29788 13864
rect 30288 13812 30340 13864
rect 32312 13812 32364 13864
rect 34612 13948 34664 14000
rect 38384 13948 38436 14000
rect 33048 13855 33100 13864
rect 33048 13821 33057 13855
rect 33057 13821 33091 13855
rect 33091 13821 33100 13855
rect 33048 13812 33100 13821
rect 34336 13880 34388 13932
rect 33416 13855 33468 13864
rect 33416 13821 33425 13855
rect 33425 13821 33459 13855
rect 33459 13821 33468 13855
rect 33968 13855 34020 13864
rect 33416 13812 33468 13821
rect 33968 13821 33977 13855
rect 33977 13821 34011 13855
rect 34011 13821 34020 13855
rect 33968 13812 34020 13821
rect 34244 13812 34296 13864
rect 37280 13855 37332 13864
rect 37280 13821 37289 13855
rect 37289 13821 37323 13855
rect 37323 13821 37332 13855
rect 37280 13812 37332 13821
rect 37924 13855 37976 13864
rect 37924 13821 37933 13855
rect 37933 13821 37967 13855
rect 37967 13821 37976 13855
rect 37924 13812 37976 13821
rect 32312 13676 32364 13728
rect 32496 13676 32548 13728
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 11888 13472 11940 13524
rect 24860 13472 24912 13524
rect 22284 13404 22336 13456
rect 24216 13404 24268 13456
rect 24400 13404 24452 13456
rect 1860 13379 1912 13388
rect 1860 13345 1869 13379
rect 1869 13345 1903 13379
rect 1903 13345 1912 13379
rect 1860 13336 1912 13345
rect 21548 13336 21600 13388
rect 22376 13336 22428 13388
rect 22560 13379 22612 13388
rect 22560 13345 22569 13379
rect 22569 13345 22603 13379
rect 22603 13345 22612 13379
rect 22560 13336 22612 13345
rect 25228 13336 25280 13388
rect 26240 13336 26292 13388
rect 23572 13268 23624 13320
rect 24492 13311 24544 13320
rect 24492 13277 24501 13311
rect 24501 13277 24535 13311
rect 24535 13277 24544 13311
rect 24492 13268 24544 13277
rect 17040 13132 17092 13184
rect 23848 13132 23900 13184
rect 24768 13132 24820 13184
rect 24860 13132 24912 13184
rect 26148 13268 26200 13320
rect 26700 13472 26752 13524
rect 27804 13472 27856 13524
rect 28724 13472 28776 13524
rect 29184 13515 29236 13524
rect 29184 13481 29193 13515
rect 29193 13481 29227 13515
rect 29227 13481 29236 13515
rect 29184 13472 29236 13481
rect 29552 13472 29604 13524
rect 36728 13472 36780 13524
rect 31944 13404 31996 13456
rect 27160 13336 27212 13388
rect 29092 13336 29144 13388
rect 37188 13379 37240 13388
rect 37188 13345 37197 13379
rect 37197 13345 37231 13379
rect 37231 13345 37240 13379
rect 37188 13336 37240 13345
rect 27620 13268 27672 13320
rect 26056 13200 26108 13252
rect 26884 13200 26936 13252
rect 27528 13200 27580 13252
rect 25964 13132 26016 13184
rect 27620 13132 27672 13184
rect 28908 13132 28960 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 19892 12792 19944 12844
rect 21548 12835 21600 12844
rect 21088 12767 21140 12776
rect 21088 12733 21097 12767
rect 21097 12733 21131 12767
rect 21131 12733 21140 12767
rect 21088 12724 21140 12733
rect 21548 12801 21557 12835
rect 21557 12801 21591 12835
rect 21591 12801 21600 12835
rect 21548 12792 21600 12801
rect 24216 12928 24268 12980
rect 26608 12971 26660 12980
rect 23388 12903 23440 12912
rect 23388 12869 23397 12903
rect 23397 12869 23431 12903
rect 23431 12869 23440 12903
rect 23388 12860 23440 12869
rect 26608 12937 26617 12971
rect 26617 12937 26651 12971
rect 26651 12937 26660 12971
rect 26608 12928 26660 12937
rect 26792 12928 26844 12980
rect 28540 12928 28592 12980
rect 30288 12928 30340 12980
rect 36360 12928 36412 12980
rect 38292 12928 38344 12980
rect 24860 12792 24912 12844
rect 25228 12835 25280 12844
rect 25228 12801 25237 12835
rect 25237 12801 25271 12835
rect 25271 12801 25280 12835
rect 25228 12792 25280 12801
rect 26516 12792 26568 12844
rect 27068 12792 27120 12844
rect 24952 12724 25004 12776
rect 26332 12724 26384 12776
rect 26424 12724 26476 12776
rect 34060 12860 34112 12912
rect 22560 12656 22612 12708
rect 23664 12656 23716 12708
rect 37832 12792 37884 12844
rect 38292 12792 38344 12844
rect 27620 12767 27672 12776
rect 27620 12733 27629 12767
rect 27629 12733 27663 12767
rect 27663 12733 27672 12767
rect 28724 12767 28776 12776
rect 27620 12724 27672 12733
rect 28724 12733 28733 12767
rect 28733 12733 28767 12767
rect 28767 12733 28776 12767
rect 28724 12724 28776 12733
rect 37280 12767 37332 12776
rect 37280 12733 37289 12767
rect 37289 12733 37323 12767
rect 37323 12733 37332 12767
rect 37280 12724 37332 12733
rect 37924 12767 37976 12776
rect 37924 12733 37933 12767
rect 37933 12733 37967 12767
rect 37967 12733 37976 12767
rect 37924 12724 37976 12733
rect 24216 12588 24268 12640
rect 24400 12588 24452 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 10324 12384 10376 12436
rect 1860 12291 1912 12300
rect 1860 12257 1869 12291
rect 1869 12257 1903 12291
rect 1903 12257 1912 12291
rect 1860 12248 1912 12257
rect 16948 12112 17000 12164
rect 22192 12384 22244 12436
rect 23296 12384 23348 12436
rect 26240 12384 26292 12436
rect 22744 12316 22796 12368
rect 22928 12316 22980 12368
rect 22560 12291 22612 12300
rect 22560 12257 22569 12291
rect 22569 12257 22603 12291
rect 22603 12257 22612 12291
rect 22560 12248 22612 12257
rect 24492 12291 24544 12300
rect 24492 12257 24501 12291
rect 24501 12257 24535 12291
rect 24535 12257 24544 12291
rect 24492 12248 24544 12257
rect 25964 12316 26016 12368
rect 34704 12316 34756 12368
rect 35348 12316 35400 12368
rect 32956 12248 33008 12300
rect 35624 12248 35676 12300
rect 26056 12044 26108 12096
rect 33324 12044 33376 12096
rect 36820 12044 36872 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 4988 11840 5040 11892
rect 22192 11840 22244 11892
rect 22560 11840 22612 11892
rect 36544 11840 36596 11892
rect 36636 11772 36688 11824
rect 33324 11704 33376 11756
rect 33876 11704 33928 11756
rect 24400 11636 24452 11688
rect 34520 11636 34572 11688
rect 34796 11636 34848 11688
rect 37280 11679 37332 11688
rect 37280 11645 37289 11679
rect 37289 11645 37323 11679
rect 37323 11645 37332 11679
rect 37280 11636 37332 11645
rect 1860 11611 1912 11620
rect 1860 11577 1869 11611
rect 1869 11577 1903 11611
rect 1903 11577 1912 11611
rect 1860 11568 1912 11577
rect 17868 11500 17920 11552
rect 23664 11543 23716 11552
rect 23664 11509 23673 11543
rect 23673 11509 23707 11543
rect 23707 11509 23716 11543
rect 23664 11500 23716 11509
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 31300 11296 31352 11348
rect 37096 11296 37148 11348
rect 23756 11228 23808 11280
rect 22560 11203 22612 11212
rect 22560 11169 22569 11203
rect 22569 11169 22603 11203
rect 22603 11169 22612 11203
rect 22560 11160 22612 11169
rect 30380 11160 30432 11212
rect 30932 11160 30984 11212
rect 37188 11203 37240 11212
rect 37188 11169 37197 11203
rect 37197 11169 37231 11203
rect 37231 11169 37240 11203
rect 37188 11160 37240 11169
rect 30012 11092 30064 11144
rect 30288 11092 30340 11144
rect 31116 11135 31168 11144
rect 31116 11101 31125 11135
rect 31125 11101 31159 11135
rect 31159 11101 31168 11135
rect 31116 11092 31168 11101
rect 23940 11067 23992 11076
rect 23940 11033 23949 11067
rect 23949 11033 23983 11067
rect 23983 11033 23992 11067
rect 23940 11024 23992 11033
rect 32956 11024 33008 11076
rect 38936 11067 38988 11076
rect 38936 11033 38945 11067
rect 38945 11033 38979 11067
rect 38979 11033 38988 11067
rect 38936 11024 38988 11033
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 8944 10752 8996 10804
rect 36452 10752 36504 10804
rect 35808 10684 35860 10736
rect 1860 10591 1912 10600
rect 1860 10557 1869 10591
rect 1869 10557 1903 10591
rect 1903 10557 1912 10591
rect 1860 10548 1912 10557
rect 37280 10591 37332 10600
rect 37280 10557 37289 10591
rect 37289 10557 37323 10591
rect 37323 10557 37332 10591
rect 37280 10548 37332 10557
rect 37924 10591 37976 10600
rect 37924 10557 37933 10591
rect 37933 10557 37967 10591
rect 37967 10557 37976 10591
rect 37924 10548 37976 10557
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 1860 10115 1912 10124
rect 1860 10081 1869 10115
rect 1869 10081 1903 10115
rect 1903 10081 1912 10115
rect 1860 10072 1912 10081
rect 25780 10072 25832 10124
rect 15936 9868 15988 9920
rect 32496 9868 32548 9920
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 38476 9596 38528 9648
rect 37280 9503 37332 9512
rect 37280 9469 37289 9503
rect 37289 9469 37323 9503
rect 37323 9469 37332 9503
rect 37280 9460 37332 9469
rect 37924 9503 37976 9512
rect 37924 9469 37933 9503
rect 37933 9469 37967 9503
rect 37967 9469 37976 9503
rect 37924 9460 37976 9469
rect 38568 9324 38620 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 37372 9163 37424 9172
rect 37372 9129 37381 9163
rect 37381 9129 37415 9163
rect 37415 9129 37424 9163
rect 37372 9120 37424 9129
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 37188 9027 37240 9036
rect 37188 8993 37197 9027
rect 37197 8993 37231 9027
rect 37231 8993 37240 9027
rect 37188 8984 37240 8993
rect 30196 8916 30248 8968
rect 33692 8916 33744 8968
rect 15292 8780 15344 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 34612 8576 34664 8628
rect 35716 8508 35768 8560
rect 37188 8372 37240 8424
rect 37924 8415 37976 8424
rect 37924 8381 37933 8415
rect 37933 8381 37967 8415
rect 37967 8381 37976 8415
rect 37924 8372 37976 8381
rect 1860 8347 1912 8356
rect 1860 8313 1869 8347
rect 1869 8313 1903 8347
rect 1903 8313 1912 8347
rect 1860 8304 1912 8313
rect 17408 8304 17460 8356
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 28540 8032 28592 8084
rect 26516 7964 26568 8016
rect 22744 7896 22796 7948
rect 28448 7896 28500 7948
rect 29552 7896 29604 7948
rect 27620 7828 27672 7880
rect 31300 7896 31352 7948
rect 10876 7760 10928 7812
rect 24308 7760 24360 7812
rect 5172 7692 5224 7744
rect 5356 7692 5408 7744
rect 12808 7692 12860 7744
rect 26608 7692 26660 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 3424 7488 3476 7540
rect 38292 7488 38344 7540
rect 36912 7420 36964 7472
rect 1860 7327 1912 7336
rect 1860 7293 1869 7327
rect 1869 7293 1903 7327
rect 1903 7293 1912 7327
rect 1860 7284 1912 7293
rect 37280 7327 37332 7336
rect 37280 7293 37289 7327
rect 37289 7293 37323 7327
rect 37323 7293 37332 7327
rect 37280 7284 37332 7293
rect 37924 7327 37976 7336
rect 37924 7293 37933 7327
rect 37933 7293 37967 7327
rect 37967 7293 37976 7327
rect 37924 7284 37976 7293
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 1860 6851 1912 6860
rect 1860 6817 1869 6851
rect 1869 6817 1903 6851
rect 1903 6817 1912 6851
rect 1860 6808 1912 6817
rect 19340 6808 19392 6860
rect 31116 6808 31168 6860
rect 37188 6851 37240 6860
rect 37188 6817 37197 6851
rect 37197 6817 37231 6851
rect 37231 6817 37240 6851
rect 37188 6808 37240 6817
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 33324 6672 33376 6724
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 20628 6400 20680 6452
rect 29000 6400 29052 6452
rect 36820 6443 36872 6452
rect 36820 6409 36829 6443
rect 36829 6409 36863 6443
rect 36863 6409 36872 6443
rect 36820 6400 36872 6409
rect 37464 6443 37516 6452
rect 37464 6409 37473 6443
rect 37473 6409 37507 6443
rect 37507 6409 37516 6443
rect 37464 6400 37516 6409
rect 17684 6332 17736 6384
rect 26700 6332 26752 6384
rect 36176 6332 36228 6384
rect 15752 6264 15804 6316
rect 25688 6264 25740 6316
rect 8944 6196 8996 6248
rect 23940 6196 23992 6248
rect 36912 6196 36964 6248
rect 37280 6239 37332 6248
rect 37280 6205 37289 6239
rect 37289 6205 37323 6239
rect 37323 6205 37332 6239
rect 37280 6196 37332 6205
rect 8024 6128 8076 6180
rect 23664 6128 23716 6180
rect 21272 6060 21324 6112
rect 28632 6060 28684 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 35440 5899 35492 5908
rect 35440 5865 35449 5899
rect 35449 5865 35483 5899
rect 35483 5865 35492 5899
rect 35440 5856 35492 5865
rect 35900 5856 35952 5908
rect 36084 5899 36136 5908
rect 36084 5865 36093 5899
rect 36093 5865 36127 5899
rect 36127 5865 36136 5899
rect 36084 5856 36136 5865
rect 1860 5831 1912 5840
rect 1860 5797 1869 5831
rect 1869 5797 1903 5831
rect 1903 5797 1912 5831
rect 1860 5788 1912 5797
rect 2136 5788 2188 5840
rect 6276 5788 6328 5840
rect 2412 5720 2464 5772
rect 34520 5720 34572 5772
rect 35532 5720 35584 5772
rect 35900 5763 35952 5772
rect 35900 5729 35909 5763
rect 35909 5729 35943 5763
rect 35943 5729 35952 5763
rect 35900 5720 35952 5729
rect 37188 5763 37240 5772
rect 2228 5652 2280 5704
rect 6368 5652 6420 5704
rect 35808 5652 35860 5704
rect 37188 5729 37197 5763
rect 37197 5729 37231 5763
rect 37231 5729 37240 5763
rect 37188 5720 37240 5729
rect 3240 5559 3292 5568
rect 3240 5525 3249 5559
rect 3249 5525 3283 5559
rect 3283 5525 3292 5559
rect 3240 5516 3292 5525
rect 12624 5584 12676 5636
rect 34704 5584 34756 5636
rect 14464 5516 14516 5568
rect 31760 5516 31812 5568
rect 38936 5559 38988 5568
rect 38936 5525 38945 5559
rect 38945 5525 38979 5559
rect 38979 5525 38988 5559
rect 38936 5516 38988 5525
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 2136 5355 2188 5364
rect 2136 5321 2145 5355
rect 2145 5321 2179 5355
rect 2179 5321 2188 5355
rect 2136 5312 2188 5321
rect 24676 5312 24728 5364
rect 30748 5312 30800 5364
rect 34796 5355 34848 5364
rect 34796 5321 34805 5355
rect 34805 5321 34839 5355
rect 34839 5321 34848 5355
rect 34796 5312 34848 5321
rect 35348 5312 35400 5364
rect 23572 5244 23624 5296
rect 31024 5244 31076 5296
rect 33784 5244 33836 5296
rect 2780 5176 2832 5228
rect 18236 5176 18288 5228
rect 30288 5176 30340 5228
rect 16764 5108 16816 5160
rect 28356 5108 28408 5160
rect 34612 5151 34664 5160
rect 34612 5117 34621 5151
rect 34621 5117 34655 5151
rect 34655 5117 34664 5151
rect 34612 5108 34664 5117
rect 36084 5108 36136 5160
rect 36728 5108 36780 5160
rect 37096 5108 37148 5160
rect 1860 5083 1912 5092
rect 1860 5049 1869 5083
rect 1869 5049 1903 5083
rect 1903 5049 1912 5083
rect 1860 5040 1912 5049
rect 4344 5040 4396 5092
rect 16396 5040 16448 5092
rect 30932 5040 30984 5092
rect 34704 5040 34756 5092
rect 39396 5040 39448 5092
rect 6920 4972 6972 5024
rect 23848 4972 23900 5024
rect 32404 4972 32456 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 4620 4768 4672 4820
rect 23388 4768 23440 4820
rect 33048 4768 33100 4820
rect 35716 4768 35768 4820
rect 2228 4743 2280 4752
rect 2228 4709 2237 4743
rect 2237 4709 2271 4743
rect 2271 4709 2280 4743
rect 2228 4700 2280 4709
rect 3148 4700 3200 4752
rect 3240 4700 3292 4752
rect 34428 4700 34480 4752
rect 36360 4700 36412 4752
rect 1860 4675 1912 4684
rect 1860 4641 1869 4675
rect 1869 4641 1903 4675
rect 1903 4641 1912 4675
rect 1860 4632 1912 4641
rect 4344 4675 4396 4684
rect 4344 4641 4353 4675
rect 4353 4641 4387 4675
rect 4387 4641 4396 4675
rect 4344 4632 4396 4641
rect 5172 4632 5224 4684
rect 31944 4632 31996 4684
rect 33600 4632 33652 4684
rect 35624 4632 35676 4684
rect 36452 4675 36504 4684
rect 36452 4641 36461 4675
rect 36461 4641 36495 4675
rect 36495 4641 36504 4675
rect 36452 4632 36504 4641
rect 3148 4496 3200 4548
rect 34796 4496 34848 4548
rect 39764 4496 39816 4548
rect 3608 4471 3660 4480
rect 3608 4437 3617 4471
rect 3617 4437 3651 4471
rect 3651 4437 3660 4471
rect 3608 4428 3660 4437
rect 12440 4428 12492 4480
rect 29276 4428 29328 4480
rect 31852 4428 31904 4480
rect 32036 4428 32088 4480
rect 35256 4428 35308 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 2872 4267 2924 4276
rect 2872 4233 2881 4267
rect 2881 4233 2915 4267
rect 2915 4233 2924 4267
rect 2872 4224 2924 4233
rect 27988 4224 28040 4276
rect 2044 4088 2096 4140
rect 27896 4156 27948 4208
rect 20720 4088 20772 4140
rect 1492 4020 1544 4072
rect 3608 4020 3660 4072
rect 4620 4020 4672 4072
rect 4712 4020 4764 4072
rect 5264 4020 5316 4072
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 11888 4063 11940 4072
rect 11888 4029 11897 4063
rect 11897 4029 11931 4063
rect 11931 4029 11940 4063
rect 11888 4020 11940 4029
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 14372 4020 14424 4072
rect 18696 4063 18748 4072
rect 1860 3995 1912 4004
rect 1860 3961 1869 3995
rect 1869 3961 1903 3995
rect 1903 3961 1912 3995
rect 1860 3952 1912 3961
rect 2688 3952 2740 4004
rect 3608 3884 3660 3936
rect 11796 3884 11848 3936
rect 12716 3884 12768 3936
rect 16764 3995 16816 4004
rect 16764 3961 16773 3995
rect 16773 3961 16807 3995
rect 16807 3961 16816 3995
rect 16764 3952 16816 3961
rect 17684 3995 17736 4004
rect 17684 3961 17693 3995
rect 17693 3961 17727 3995
rect 17727 3961 17736 3995
rect 17684 3952 17736 3961
rect 18696 4029 18705 4063
rect 18705 4029 18739 4063
rect 18739 4029 18748 4063
rect 18696 4020 18748 4029
rect 19984 4020 20036 4072
rect 21824 4020 21876 4072
rect 22836 4020 22888 4072
rect 23204 4020 23256 4072
rect 24124 4020 24176 4072
rect 24768 4020 24820 4072
rect 20076 3952 20128 4004
rect 20996 3952 21048 4004
rect 31668 4088 31720 4140
rect 31760 4088 31812 4140
rect 32956 4156 33008 4208
rect 32128 4088 32180 4140
rect 33140 4088 33192 4140
rect 34336 4088 34388 4140
rect 25964 4063 26016 4072
rect 25964 4029 25973 4063
rect 25973 4029 26007 4063
rect 26007 4029 26016 4063
rect 25964 4020 26016 4029
rect 25780 3952 25832 4004
rect 26884 4020 26936 4072
rect 28908 4063 28960 4072
rect 28908 4029 28917 4063
rect 28917 4029 28951 4063
rect 28951 4029 28960 4063
rect 28908 4020 28960 4029
rect 29552 4063 29604 4072
rect 29552 4029 29561 4063
rect 29561 4029 29595 4063
rect 29595 4029 29604 4063
rect 29552 4020 29604 4029
rect 29644 4020 29696 4072
rect 30748 4020 30800 4072
rect 27528 3952 27580 4004
rect 29276 3952 29328 4004
rect 31852 4020 31904 4072
rect 32588 4020 32640 4072
rect 33416 4063 33468 4072
rect 33416 4029 33425 4063
rect 33425 4029 33459 4063
rect 33459 4029 33468 4063
rect 33416 4020 33468 4029
rect 34796 4020 34848 4072
rect 16672 3884 16724 3936
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 18696 3884 18748 3936
rect 20260 3884 20312 3936
rect 20444 3884 20496 3936
rect 21916 3884 21968 3936
rect 25136 3884 25188 3936
rect 25596 3884 25648 3936
rect 26240 3884 26292 3936
rect 26700 3884 26752 3936
rect 28080 3884 28132 3936
rect 34612 3952 34664 4004
rect 29460 3884 29512 3936
rect 30564 3884 30616 3936
rect 31760 3927 31812 3936
rect 31760 3893 31769 3927
rect 31769 3893 31803 3927
rect 31803 3893 31812 3927
rect 31760 3884 31812 3893
rect 31852 3884 31904 3936
rect 33508 3884 33560 3936
rect 34704 3884 34756 3936
rect 36360 3884 36412 3936
rect 36636 3952 36688 4004
rect 39120 4020 39172 4072
rect 38476 3952 38528 4004
rect 38752 3884 38804 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 1032 3680 1084 3732
rect 2780 3680 2832 3732
rect 3516 3723 3568 3732
rect 3516 3689 3525 3723
rect 3525 3689 3559 3723
rect 3559 3689 3568 3723
rect 3516 3680 3568 3689
rect 2504 3612 2556 3664
rect 6644 3612 6696 3664
rect 6920 3655 6972 3664
rect 6920 3621 6929 3655
rect 6929 3621 6963 3655
rect 6963 3621 6972 3655
rect 6920 3612 6972 3621
rect 8944 3655 8996 3664
rect 8944 3621 8953 3655
rect 8953 3621 8987 3655
rect 8987 3621 8996 3655
rect 8944 3612 8996 3621
rect 10876 3655 10928 3664
rect 10876 3621 10885 3655
rect 10885 3621 10919 3655
rect 10919 3621 10928 3655
rect 10876 3612 10928 3621
rect 12624 3612 12676 3664
rect 13268 3612 13320 3664
rect 14096 3655 14148 3664
rect 14096 3621 14105 3655
rect 14105 3621 14139 3655
rect 14139 3621 14148 3655
rect 14096 3612 14148 3621
rect 19248 3680 19300 3732
rect 19432 3723 19484 3732
rect 19432 3689 19441 3723
rect 19441 3689 19475 3723
rect 19475 3689 19484 3723
rect 19432 3680 19484 3689
rect 20076 3680 20128 3732
rect 25964 3680 26016 3732
rect 27896 3680 27948 3732
rect 1400 3544 1452 3596
rect 3332 3544 3384 3596
rect 4988 3544 5040 3596
rect 112 3476 164 3528
rect 1308 3476 1360 3528
rect 3976 3476 4028 3528
rect 7840 3544 7892 3596
rect 8484 3544 8536 3596
rect 9496 3544 9548 3596
rect 12808 3544 12860 3596
rect 14924 3544 14976 3596
rect 15752 3587 15804 3596
rect 15752 3553 15761 3587
rect 15761 3553 15795 3587
rect 15795 3553 15804 3587
rect 15752 3544 15804 3553
rect 17960 3587 18012 3596
rect 17960 3553 17969 3587
rect 17969 3553 18003 3587
rect 18003 3553 18012 3587
rect 17960 3544 18012 3553
rect 19248 3587 19300 3596
rect 19248 3553 19257 3587
rect 19257 3553 19291 3587
rect 19291 3553 19300 3587
rect 19248 3544 19300 3553
rect 20628 3544 20680 3596
rect 20720 3587 20772 3596
rect 20720 3553 20729 3587
rect 20729 3553 20763 3587
rect 20763 3553 20772 3587
rect 20720 3544 20772 3553
rect 20904 3544 20956 3596
rect 25320 3612 25372 3664
rect 26700 3612 26752 3664
rect 27988 3612 28040 3664
rect 29368 3612 29420 3664
rect 30196 3612 30248 3664
rect 16580 3476 16632 3528
rect 1676 3340 1728 3392
rect 23848 3544 23900 3596
rect 24676 3544 24728 3596
rect 26332 3544 26384 3596
rect 24216 3476 24268 3528
rect 27528 3476 27580 3528
rect 27804 3476 27856 3528
rect 28816 3476 28868 3528
rect 29460 3476 29512 3528
rect 31576 3612 31628 3664
rect 36268 3655 36320 3664
rect 36268 3621 36277 3655
rect 36277 3621 36311 3655
rect 36311 3621 36320 3655
rect 36268 3612 36320 3621
rect 31024 3587 31076 3596
rect 31024 3553 31033 3587
rect 31033 3553 31067 3587
rect 31067 3553 31076 3587
rect 31024 3544 31076 3553
rect 31116 3544 31168 3596
rect 31760 3544 31812 3596
rect 34336 3587 34388 3596
rect 34336 3553 34345 3587
rect 34345 3553 34379 3587
rect 34379 3553 34388 3587
rect 34336 3544 34388 3553
rect 4988 3340 5040 3392
rect 6276 3340 6328 3392
rect 8852 3340 8904 3392
rect 10784 3340 10836 3392
rect 12440 3383 12492 3392
rect 12440 3349 12449 3383
rect 12449 3349 12483 3383
rect 12483 3349 12492 3383
rect 12440 3340 12492 3349
rect 13360 3340 13412 3392
rect 13636 3340 13688 3392
rect 14740 3340 14792 3392
rect 15660 3340 15712 3392
rect 19892 3340 19944 3392
rect 20996 3340 21048 3392
rect 21364 3383 21416 3392
rect 21364 3349 21373 3383
rect 21373 3349 21407 3383
rect 21407 3349 21416 3383
rect 21364 3340 21416 3349
rect 25044 3408 25096 3460
rect 25136 3408 25188 3460
rect 30012 3408 30064 3460
rect 30380 3408 30432 3460
rect 23756 3340 23808 3392
rect 24400 3340 24452 3392
rect 24492 3340 24544 3392
rect 25412 3340 25464 3392
rect 26608 3383 26660 3392
rect 26608 3349 26617 3383
rect 26617 3349 26651 3383
rect 26651 3349 26660 3383
rect 26608 3340 26660 3349
rect 27436 3340 27488 3392
rect 28540 3383 28592 3392
rect 28540 3349 28549 3383
rect 28549 3349 28583 3383
rect 28583 3349 28592 3383
rect 28540 3340 28592 3349
rect 29368 3340 29420 3392
rect 30840 3476 30892 3528
rect 31484 3476 31536 3528
rect 36636 3544 36688 3596
rect 34612 3408 34664 3460
rect 36820 3408 36872 3460
rect 37832 3408 37884 3460
rect 32312 3340 32364 3392
rect 33692 3383 33744 3392
rect 33692 3349 33701 3383
rect 33701 3349 33735 3383
rect 33735 3349 33744 3383
rect 33692 3340 33744 3349
rect 34244 3340 34296 3392
rect 36176 3340 36228 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 2320 3136 2372 3188
rect 3056 3179 3108 3188
rect 3056 3145 3065 3179
rect 3065 3145 3099 3179
rect 3099 3145 3108 3179
rect 3056 3136 3108 3145
rect 7380 3179 7432 3188
rect 7380 3145 7389 3179
rect 7389 3145 7423 3179
rect 7423 3145 7432 3179
rect 7380 3136 7432 3145
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 16488 3179 16540 3188
rect 2044 3068 2096 3120
rect 5172 3068 5224 3120
rect 7564 3068 7616 3120
rect 10508 3068 10560 3120
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 6184 3043 6236 3052
rect 6184 3009 6193 3043
rect 6193 3009 6227 3043
rect 6227 3009 6236 3043
rect 6184 3000 6236 3009
rect 11428 3043 11480 3052
rect 11428 3009 11437 3043
rect 11437 3009 11471 3043
rect 11471 3009 11480 3043
rect 11428 3000 11480 3009
rect 12348 3043 12400 3052
rect 12348 3009 12357 3043
rect 12357 3009 12391 3043
rect 12391 3009 12400 3043
rect 12348 3000 12400 3009
rect 12532 3000 12584 3052
rect 12808 3000 12860 3052
rect 13360 3000 13412 3052
rect 16488 3145 16497 3179
rect 16497 3145 16531 3179
rect 16531 3145 16540 3179
rect 16488 3136 16540 3145
rect 20260 3179 20312 3188
rect 20260 3145 20269 3179
rect 20269 3145 20303 3179
rect 20303 3145 20312 3179
rect 20260 3136 20312 3145
rect 20352 3136 20404 3188
rect 24216 3136 24268 3188
rect 24400 3136 24452 3188
rect 27528 3136 27580 3188
rect 28540 3136 28592 3188
rect 28632 3136 28684 3188
rect 30656 3136 30708 3188
rect 30840 3179 30892 3188
rect 30840 3145 30849 3179
rect 30849 3145 30883 3179
rect 30883 3145 30892 3179
rect 30840 3136 30892 3145
rect 33692 3136 33744 3188
rect 38200 3136 38252 3188
rect 388 2932 440 2984
rect 4620 2975 4672 2984
rect 4620 2941 4629 2975
rect 4629 2941 4663 2975
rect 4663 2941 4672 2975
rect 4620 2932 4672 2941
rect 5908 2975 5960 2984
rect 5908 2941 5917 2975
rect 5917 2941 5951 2975
rect 5951 2941 5960 2975
rect 5908 2932 5960 2941
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 7196 2932 7248 2941
rect 8024 2975 8076 2984
rect 8024 2941 8033 2975
rect 8033 2941 8067 2975
rect 8067 2941 8076 2975
rect 8024 2932 8076 2941
rect 9220 2932 9272 2984
rect 10324 2975 10376 2984
rect 10324 2941 10333 2975
rect 10333 2941 10367 2975
rect 10367 2941 10376 2975
rect 10324 2932 10376 2941
rect 11152 2975 11204 2984
rect 11152 2941 11161 2975
rect 11161 2941 11195 2975
rect 11195 2941 11204 2975
rect 11152 2932 11204 2941
rect 13084 2975 13136 2984
rect 13084 2941 13093 2975
rect 13093 2941 13127 2975
rect 13127 2941 13136 2975
rect 13084 2932 13136 2941
rect 15016 2932 15068 2984
rect 15384 2975 15436 2984
rect 15384 2941 15393 2975
rect 15393 2941 15427 2975
rect 15427 2941 15436 2975
rect 15384 2932 15436 2941
rect 19800 3068 19852 3120
rect 21916 3068 21968 3120
rect 25320 3068 25372 3120
rect 29000 3068 29052 3120
rect 17592 3043 17644 3052
rect 17592 3009 17601 3043
rect 17601 3009 17635 3043
rect 17635 3009 17644 3043
rect 17592 3000 17644 3009
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 21364 3000 21416 3052
rect 25596 3043 25648 3052
rect 25596 3009 25602 3043
rect 25602 3009 25636 3043
rect 25636 3009 25648 3043
rect 25596 3000 25648 3009
rect 28080 3000 28132 3052
rect 29736 3000 29788 3052
rect 31760 3068 31812 3120
rect 32128 3068 32180 3120
rect 37188 3068 37240 3120
rect 32036 3000 32088 3052
rect 16304 2975 16356 2984
rect 16304 2941 16313 2975
rect 16313 2941 16347 2975
rect 16347 2941 16356 2975
rect 16304 2932 16356 2941
rect 17316 2975 17368 2984
rect 17316 2941 17325 2975
rect 17325 2941 17359 2975
rect 17359 2941 17368 2975
rect 17316 2932 17368 2941
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 20444 2932 20496 2984
rect 20536 2932 20588 2984
rect 22744 2975 22796 2984
rect 22744 2941 22753 2975
rect 22753 2941 22787 2975
rect 22787 2941 22796 2975
rect 22744 2932 22796 2941
rect 23572 2975 23624 2984
rect 23572 2941 23581 2975
rect 23581 2941 23615 2975
rect 23615 2941 23624 2975
rect 23572 2932 23624 2941
rect 23756 2932 23808 2984
rect 1860 2907 1912 2916
rect 1860 2873 1869 2907
rect 1869 2873 1903 2907
rect 1903 2873 1912 2907
rect 1860 2864 1912 2873
rect 11428 2864 11480 2916
rect 16580 2864 16632 2916
rect 21272 2907 21324 2916
rect 756 2796 808 2848
rect 3148 2796 3200 2848
rect 7564 2796 7616 2848
rect 9864 2796 9916 2848
rect 20352 2796 20404 2848
rect 21272 2873 21281 2907
rect 21281 2873 21315 2907
rect 21315 2873 21324 2907
rect 21272 2864 21324 2873
rect 26240 2932 26292 2984
rect 26792 2932 26844 2984
rect 28540 2932 28592 2984
rect 31208 2932 31260 2984
rect 31300 2932 31352 2984
rect 32220 2932 32272 2984
rect 33232 2932 33284 2984
rect 34152 2932 34204 2984
rect 21548 2796 21600 2848
rect 22560 2796 22612 2848
rect 23480 2796 23532 2848
rect 34796 2932 34848 2984
rect 37924 2975 37976 2984
rect 37924 2941 37933 2975
rect 37933 2941 37967 2975
rect 37967 2941 37976 2975
rect 37924 2932 37976 2941
rect 38108 2907 38160 2916
rect 38108 2873 38117 2907
rect 38117 2873 38151 2907
rect 38151 2873 38160 2907
rect 38108 2864 38160 2873
rect 26332 2796 26384 2848
rect 26424 2796 26476 2848
rect 28356 2796 28408 2848
rect 31300 2796 31352 2848
rect 32312 2796 32364 2848
rect 33232 2796 33284 2848
rect 36544 2796 36596 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 2964 2592 3016 2644
rect 4896 2592 4948 2644
rect 11244 2635 11296 2644
rect 2872 2524 2924 2576
rect 5356 2524 5408 2576
rect 8392 2524 8444 2576
rect 9956 2524 10008 2576
rect 11244 2601 11253 2635
rect 11253 2601 11287 2635
rect 11287 2601 11296 2635
rect 11244 2592 11296 2601
rect 12900 2592 12952 2644
rect 23112 2635 23164 2644
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 2964 2456 3016 2508
rect 5632 2456 5684 2508
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 8208 2499 8260 2508
rect 6920 2456 6972 2465
rect 8208 2465 8217 2499
rect 8217 2465 8251 2499
rect 8251 2465 8260 2499
rect 8208 2456 8260 2465
rect 10140 2499 10192 2508
rect 10140 2465 10149 2499
rect 10149 2465 10183 2499
rect 10183 2465 10192 2499
rect 10140 2456 10192 2465
rect 13728 2567 13780 2576
rect 12072 2456 12124 2508
rect 1584 2388 1636 2440
rect 5448 2388 5500 2440
rect 10508 2388 10560 2440
rect 13728 2533 13737 2567
rect 13737 2533 13771 2567
rect 13771 2533 13780 2567
rect 13728 2524 13780 2533
rect 16396 2567 16448 2576
rect 16396 2533 16405 2567
rect 16405 2533 16439 2567
rect 16439 2533 16448 2567
rect 16396 2524 16448 2533
rect 23112 2601 23121 2635
rect 23121 2601 23155 2635
rect 23155 2601 23164 2635
rect 23112 2592 23164 2601
rect 24584 2635 24636 2644
rect 24584 2601 24593 2635
rect 24593 2601 24627 2635
rect 24627 2601 24636 2635
rect 24584 2592 24636 2601
rect 27712 2592 27764 2644
rect 33416 2592 33468 2644
rect 34612 2592 34664 2644
rect 32496 2567 32548 2576
rect 32496 2533 32505 2567
rect 32505 2533 32539 2567
rect 32539 2533 32548 2567
rect 32496 2524 32548 2533
rect 35992 2524 36044 2576
rect 37648 2524 37700 2576
rect 13452 2456 13504 2508
rect 14096 2456 14148 2508
rect 16028 2499 16080 2508
rect 5080 2320 5132 2372
rect 6460 2252 6512 2304
rect 7012 2252 7064 2304
rect 16028 2465 16037 2499
rect 16037 2465 16071 2499
rect 16071 2465 16080 2499
rect 16028 2456 16080 2465
rect 16948 2456 17000 2508
rect 18236 2499 18288 2508
rect 18236 2465 18245 2499
rect 18245 2465 18279 2499
rect 18279 2465 18288 2499
rect 18236 2456 18288 2465
rect 18972 2499 19024 2508
rect 18972 2465 18981 2499
rect 18981 2465 19015 2499
rect 19015 2465 19024 2499
rect 18972 2456 19024 2465
rect 20260 2499 20312 2508
rect 20260 2465 20269 2499
rect 20269 2465 20303 2499
rect 20303 2465 20312 2499
rect 20260 2456 20312 2465
rect 21180 2499 21232 2508
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 21456 2499 21508 2508
rect 21456 2465 21465 2499
rect 21465 2465 21499 2499
rect 21499 2465 21508 2499
rect 21456 2456 21508 2465
rect 22192 2456 22244 2508
rect 25136 2456 25188 2508
rect 26056 2499 26108 2508
rect 26056 2465 26065 2499
rect 26065 2465 26099 2499
rect 26099 2465 26108 2499
rect 26056 2456 26108 2465
rect 27068 2499 27120 2508
rect 27068 2465 27077 2499
rect 27077 2465 27111 2499
rect 27111 2465 27120 2499
rect 27068 2456 27120 2465
rect 28080 2456 28132 2508
rect 30012 2456 30064 2508
rect 30932 2456 30984 2508
rect 32956 2456 33008 2508
rect 33876 2456 33928 2508
rect 35900 2456 35952 2508
rect 37464 2499 37516 2508
rect 37464 2465 37473 2499
rect 37473 2465 37507 2499
rect 37507 2465 37516 2499
rect 37464 2456 37516 2465
rect 29736 2431 29788 2440
rect 29736 2397 29745 2431
rect 29745 2397 29779 2431
rect 29779 2397 29788 2431
rect 29736 2388 29788 2397
rect 33968 2388 34020 2440
rect 28172 2320 28224 2372
rect 35532 2320 35584 2372
rect 27344 2252 27396 2304
rect 31116 2295 31168 2304
rect 31116 2261 31125 2295
rect 31125 2261 31159 2295
rect 31159 2261 31168 2295
rect 31116 2252 31168 2261
rect 37004 2252 37056 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 4252 1980 4304 2032
rect 4712 1980 4764 2032
rect 15476 1980 15528 2032
rect 31116 1980 31168 2032
rect 14832 1912 14884 1964
rect 29736 1912 29788 1964
rect 29000 1504 29052 1556
rect 29552 1504 29604 1556
<< metal2 >>
rect 110 119200 166 120800
rect 294 119200 350 120800
rect 570 119200 626 120800
rect 754 119200 810 120800
rect 1030 119200 1086 120800
rect 1214 119200 1270 120800
rect 1490 119200 1546 120800
rect 1674 119200 1730 120800
rect 1950 119200 2006 120800
rect 2134 119200 2190 120800
rect 2410 119200 2466 120800
rect 2594 119200 2650 120800
rect 2870 119200 2926 120800
rect 3054 119200 3110 120800
rect 3330 119200 3386 120800
rect 3422 119504 3478 119513
rect 3422 119439 3478 119448
rect 124 117298 152 119200
rect 308 117434 336 119200
rect 296 117428 348 117434
rect 296 117370 348 117376
rect 112 117292 164 117298
rect 112 117234 164 117240
rect 584 115802 612 119200
rect 768 117230 796 119200
rect 756 117224 808 117230
rect 756 117166 808 117172
rect 1044 117094 1072 119200
rect 1228 117366 1256 119200
rect 1398 117872 1454 117881
rect 1398 117807 1454 117816
rect 1216 117360 1268 117366
rect 1216 117302 1268 117308
rect 1032 117088 1084 117094
rect 1032 117030 1084 117036
rect 572 115796 624 115802
rect 572 115738 624 115744
rect 1412 115258 1440 117807
rect 1504 115530 1532 119200
rect 1688 116890 1716 119200
rect 1860 117156 1912 117162
rect 1860 117098 1912 117104
rect 1676 116884 1728 116890
rect 1676 116826 1728 116832
rect 1872 116278 1900 117098
rect 1964 116362 1992 119200
rect 2148 116822 2176 119200
rect 2136 116816 2188 116822
rect 2136 116758 2188 116764
rect 1964 116334 2176 116362
rect 2424 116346 2452 119200
rect 1860 116272 1912 116278
rect 1860 116214 1912 116220
rect 2042 116240 2098 116249
rect 2042 116175 2044 116184
rect 2096 116175 2098 116184
rect 2044 116146 2096 116152
rect 1768 116068 1820 116074
rect 1768 116010 1820 116016
rect 1492 115524 1544 115530
rect 1492 115466 1544 115472
rect 1400 115252 1452 115258
rect 1400 115194 1452 115200
rect 1398 105904 1454 105913
rect 1398 105839 1400 105848
rect 1452 105839 1454 105848
rect 1400 105810 1452 105816
rect 1584 105800 1636 105806
rect 1584 105742 1636 105748
rect 1490 104272 1546 104281
rect 1490 104207 1546 104216
rect 1504 104174 1532 104207
rect 1492 104168 1544 104174
rect 1492 104110 1544 104116
rect 1492 102604 1544 102610
rect 1492 102546 1544 102552
rect 1400 101992 1452 101998
rect 1400 101934 1452 101940
rect 1412 101833 1440 101934
rect 1398 101824 1454 101833
rect 1398 101759 1454 101768
rect 1398 101008 1454 101017
rect 1398 100943 1454 100952
rect 1412 100910 1440 100943
rect 1400 100904 1452 100910
rect 1400 100846 1452 100852
rect 1400 100428 1452 100434
rect 1400 100370 1452 100376
rect 1412 100337 1440 100370
rect 1398 100328 1454 100337
rect 1398 100263 1454 100272
rect 1398 99512 1454 99521
rect 1398 99447 1454 99456
rect 1412 99346 1440 99447
rect 1400 99340 1452 99346
rect 1400 99282 1452 99288
rect 1400 98728 1452 98734
rect 1398 98696 1400 98705
rect 1452 98696 1454 98705
rect 1398 98631 1454 98640
rect 1398 97880 1454 97889
rect 1398 97815 1454 97824
rect 1412 97646 1440 97815
rect 1400 97640 1452 97646
rect 1400 97582 1452 97588
rect 1400 97164 1452 97170
rect 1400 97106 1452 97112
rect 1412 97073 1440 97106
rect 1398 97064 1454 97073
rect 1398 96999 1454 97008
rect 1398 96248 1454 96257
rect 1398 96183 1454 96192
rect 1412 96082 1440 96183
rect 1400 96076 1452 96082
rect 1400 96018 1452 96024
rect 1400 95464 1452 95470
rect 1398 95432 1400 95441
rect 1452 95432 1454 95441
rect 1398 95367 1454 95376
rect 1398 94616 1454 94625
rect 1398 94551 1454 94560
rect 1412 94382 1440 94551
rect 1400 94376 1452 94382
rect 1400 94318 1452 94324
rect 1400 93900 1452 93906
rect 1400 93842 1452 93848
rect 1412 93809 1440 93842
rect 1398 93800 1454 93809
rect 1398 93735 1454 93744
rect 1400 93288 1452 93294
rect 1400 93230 1452 93236
rect 1412 93129 1440 93230
rect 1398 93120 1454 93129
rect 1398 93055 1454 93064
rect 1398 92304 1454 92313
rect 1398 92239 1454 92248
rect 1412 92206 1440 92239
rect 1400 92200 1452 92206
rect 1400 92142 1452 92148
rect 1400 91724 1452 91730
rect 1400 91666 1452 91672
rect 1412 91497 1440 91666
rect 1398 91488 1454 91497
rect 1398 91423 1454 91432
rect 1400 91112 1452 91118
rect 1400 91054 1452 91060
rect 1412 90114 1440 91054
rect 1504 90778 1532 102546
rect 1492 90772 1544 90778
rect 1492 90714 1544 90720
rect 1412 90086 1532 90114
rect 1400 90024 1452 90030
rect 1400 89966 1452 89972
rect 1412 89865 1440 89966
rect 1398 89856 1454 89865
rect 1398 89791 1454 89800
rect 1398 89040 1454 89049
rect 1398 88975 1454 88984
rect 1412 88942 1440 88975
rect 1400 88936 1452 88942
rect 1400 88878 1452 88884
rect 1400 88460 1452 88466
rect 1400 88402 1452 88408
rect 1412 88233 1440 88402
rect 1398 88224 1454 88233
rect 1398 88159 1454 88168
rect 1398 87408 1454 87417
rect 1398 87343 1400 87352
rect 1452 87343 1454 87352
rect 1400 87314 1452 87320
rect 1400 86760 1452 86766
rect 1398 86728 1400 86737
rect 1452 86728 1454 86737
rect 1398 86663 1454 86672
rect 1398 85912 1454 85921
rect 1398 85847 1454 85856
rect 1412 85678 1440 85847
rect 1400 85672 1452 85678
rect 1400 85614 1452 85620
rect 1400 85196 1452 85202
rect 1400 85138 1452 85144
rect 1412 85105 1440 85138
rect 1398 85096 1454 85105
rect 1398 85031 1454 85040
rect 1398 84280 1454 84289
rect 1398 84215 1454 84224
rect 1412 84114 1440 84215
rect 1400 84108 1452 84114
rect 1400 84050 1452 84056
rect 1400 83496 1452 83502
rect 1398 83464 1400 83473
rect 1452 83464 1454 83473
rect 1398 83399 1454 83408
rect 1398 82648 1454 82657
rect 1398 82583 1454 82592
rect 1412 82414 1440 82583
rect 1400 82408 1452 82414
rect 1400 82350 1452 82356
rect 1400 81932 1452 81938
rect 1400 81874 1452 81880
rect 1412 81841 1440 81874
rect 1398 81832 1454 81841
rect 1398 81767 1454 81776
rect 1398 81016 1454 81025
rect 1398 80951 1454 80960
rect 1412 80850 1440 80951
rect 1400 80844 1452 80850
rect 1400 80786 1452 80792
rect 1398 80336 1454 80345
rect 1398 80271 1454 80280
rect 1412 80238 1440 80271
rect 1400 80232 1452 80238
rect 1400 80174 1452 80180
rect 1400 79756 1452 79762
rect 1400 79698 1452 79704
rect 1412 79529 1440 79698
rect 1398 79520 1454 79529
rect 1398 79455 1454 79464
rect 1398 78704 1454 78713
rect 1398 78639 1400 78648
rect 1452 78639 1454 78648
rect 1400 78610 1452 78616
rect 1400 78056 1452 78062
rect 1400 77998 1452 78004
rect 1412 77897 1440 77998
rect 1398 77888 1454 77897
rect 1398 77823 1454 77832
rect 1398 77072 1454 77081
rect 1398 77007 1454 77016
rect 1412 76974 1440 77007
rect 1400 76968 1452 76974
rect 1400 76910 1452 76916
rect 1400 76492 1452 76498
rect 1400 76434 1452 76440
rect 1412 76265 1440 76434
rect 1398 76256 1454 76265
rect 1398 76191 1454 76200
rect 1398 75440 1454 75449
rect 1398 75375 1400 75384
rect 1452 75375 1454 75384
rect 1400 75346 1452 75352
rect 1400 74792 1452 74798
rect 1400 74734 1452 74740
rect 1412 74633 1440 74734
rect 1398 74624 1454 74633
rect 1398 74559 1454 74568
rect 1398 73808 1454 73817
rect 1398 73743 1454 73752
rect 1412 73710 1440 73743
rect 1400 73704 1452 73710
rect 1400 73646 1452 73652
rect 1400 73228 1452 73234
rect 1400 73170 1452 73176
rect 1412 73137 1440 73170
rect 1398 73128 1454 73137
rect 1398 73063 1454 73072
rect 1398 72312 1454 72321
rect 1398 72247 1454 72256
rect 1412 72146 1440 72247
rect 1400 72140 1452 72146
rect 1400 72082 1452 72088
rect 1400 71528 1452 71534
rect 1398 71496 1400 71505
rect 1452 71496 1454 71505
rect 1398 71431 1454 71440
rect 1398 70680 1454 70689
rect 1398 70615 1454 70624
rect 1412 70446 1440 70615
rect 1400 70440 1452 70446
rect 1400 70382 1452 70388
rect 1400 69964 1452 69970
rect 1400 69906 1452 69912
rect 1412 69873 1440 69906
rect 1398 69864 1454 69873
rect 1398 69799 1454 69808
rect 1398 69048 1454 69057
rect 1398 68983 1454 68992
rect 1412 68882 1440 68983
rect 1400 68876 1452 68882
rect 1400 68818 1452 68824
rect 1400 68264 1452 68270
rect 1398 68232 1400 68241
rect 1452 68232 1454 68241
rect 1398 68167 1454 68176
rect 1398 67416 1454 67425
rect 1398 67351 1454 67360
rect 1412 67182 1440 67351
rect 1400 67176 1452 67182
rect 1400 67118 1452 67124
rect 1398 66736 1454 66745
rect 1398 66671 1400 66680
rect 1452 66671 1454 66680
rect 1400 66642 1452 66648
rect 1400 66088 1452 66094
rect 1400 66030 1452 66036
rect 1412 65929 1440 66030
rect 1398 65920 1454 65929
rect 1398 65855 1454 65864
rect 1398 65104 1454 65113
rect 1398 65039 1454 65048
rect 1412 65006 1440 65039
rect 1400 65000 1452 65006
rect 1400 64942 1452 64948
rect 1400 64524 1452 64530
rect 1400 64466 1452 64472
rect 1412 64297 1440 64466
rect 1398 64288 1454 64297
rect 1398 64223 1454 64232
rect 1398 63472 1454 63481
rect 1398 63407 1400 63416
rect 1452 63407 1454 63416
rect 1400 63378 1452 63384
rect 1400 62824 1452 62830
rect 1400 62766 1452 62772
rect 1412 62665 1440 62766
rect 1398 62656 1454 62665
rect 1398 62591 1454 62600
rect 1398 61840 1454 61849
rect 1398 61775 1454 61784
rect 1412 61742 1440 61775
rect 1400 61736 1452 61742
rect 1400 61678 1452 61684
rect 1400 61260 1452 61266
rect 1400 61202 1452 61208
rect 1412 61033 1440 61202
rect 1398 61024 1454 61033
rect 1398 60959 1454 60968
rect 1398 60344 1454 60353
rect 1398 60279 1454 60288
rect 1412 60178 1440 60279
rect 1400 60172 1452 60178
rect 1400 60114 1452 60120
rect 1400 59560 1452 59566
rect 1398 59528 1400 59537
rect 1452 59528 1454 59537
rect 1398 59463 1454 59472
rect 1398 58712 1454 58721
rect 1398 58647 1454 58656
rect 1412 58478 1440 58647
rect 1400 58472 1452 58478
rect 1400 58414 1452 58420
rect 1400 57996 1452 58002
rect 1400 57938 1452 57944
rect 1412 57905 1440 57938
rect 1398 57896 1454 57905
rect 1398 57831 1454 57840
rect 1398 57080 1454 57089
rect 1398 57015 1454 57024
rect 1412 56914 1440 57015
rect 1400 56908 1452 56914
rect 1400 56850 1452 56856
rect 1400 56296 1452 56302
rect 1398 56264 1400 56273
rect 1452 56264 1454 56273
rect 1398 56199 1454 56208
rect 1398 55448 1454 55457
rect 1398 55383 1454 55392
rect 1412 55214 1440 55383
rect 1400 55208 1452 55214
rect 1400 55150 1452 55156
rect 1400 54732 1452 54738
rect 1400 54674 1452 54680
rect 1412 54641 1440 54674
rect 1398 54632 1454 54641
rect 1398 54567 1454 54576
rect 1398 53816 1454 53825
rect 1398 53751 1454 53760
rect 1412 53650 1440 53751
rect 1400 53644 1452 53650
rect 1400 53586 1452 53592
rect 1398 53136 1454 53145
rect 1398 53071 1454 53080
rect 1412 53038 1440 53071
rect 1400 53032 1452 53038
rect 1400 52974 1452 52980
rect 1400 52556 1452 52562
rect 1400 52498 1452 52504
rect 1412 52329 1440 52498
rect 1398 52320 1454 52329
rect 1398 52255 1454 52264
rect 1398 51504 1454 51513
rect 1398 51439 1400 51448
rect 1452 51439 1454 51448
rect 1400 51410 1452 51416
rect 1504 45554 1532 90086
rect 1596 68202 1624 105742
rect 1676 103692 1728 103698
rect 1676 103634 1728 103640
rect 1688 91322 1716 103634
rect 1780 103514 1808 116010
rect 1952 115456 2004 115462
rect 1950 115424 1952 115433
rect 2004 115424 2006 115433
rect 1950 115359 2006 115368
rect 2042 114608 2098 114617
rect 2042 114543 2098 114552
rect 2056 114510 2084 114543
rect 2044 114504 2096 114510
rect 2044 114446 2096 114452
rect 1860 113892 1912 113898
rect 1860 113834 1912 113840
rect 1872 113801 1900 113834
rect 1858 113792 1914 113801
rect 1858 113727 1914 113736
rect 2148 113490 2176 116334
rect 2412 116340 2464 116346
rect 2412 116282 2464 116288
rect 2608 114900 2636 119200
rect 2884 118810 2912 119200
rect 2884 118782 3004 118810
rect 2870 118688 2926 118697
rect 2870 118623 2926 118632
rect 2778 117056 2834 117065
rect 2778 116991 2834 117000
rect 2792 115190 2820 116991
rect 2780 115184 2832 115190
rect 2780 115126 2832 115132
rect 2608 114872 2820 114900
rect 2596 114572 2648 114578
rect 2596 114514 2648 114520
rect 2136 113484 2188 113490
rect 2136 113426 2188 113432
rect 1950 113112 2006 113121
rect 1950 113047 1952 113056
rect 2004 113047 2006 113056
rect 1952 113018 2004 113024
rect 2228 112804 2280 112810
rect 2228 112746 2280 112752
rect 2044 112328 2096 112334
rect 2042 112296 2044 112305
rect 2096 112296 2098 112305
rect 2042 112231 2098 112240
rect 1950 111480 2006 111489
rect 1950 111415 1952 111424
rect 2004 111415 2006 111424
rect 1952 111386 2004 111392
rect 2136 110696 2188 110702
rect 2042 110664 2098 110673
rect 2136 110638 2188 110644
rect 2042 110599 2044 110608
rect 2096 110599 2098 110608
rect 2044 110570 2096 110576
rect 1950 109848 2006 109857
rect 1950 109783 1952 109792
rect 2004 109783 2006 109792
rect 1952 109754 2004 109760
rect 1952 109540 2004 109546
rect 1952 109482 2004 109488
rect 1860 109132 1912 109138
rect 1860 109074 1912 109080
rect 1872 109041 1900 109074
rect 1858 109032 1914 109041
rect 1858 108967 1914 108976
rect 1964 108338 1992 109482
rect 1872 108310 1992 108338
rect 1872 104938 1900 108310
rect 1950 108216 2006 108225
rect 1950 108151 1952 108160
rect 2004 108151 2006 108160
rect 1952 108122 2004 108128
rect 2042 107400 2098 107409
rect 2042 107335 2044 107344
rect 2096 107335 2098 107344
rect 2044 107306 2096 107312
rect 1952 106752 2004 106758
rect 1950 106720 1952 106729
rect 2004 106720 2006 106729
rect 1950 106655 2006 106664
rect 1952 105120 2004 105126
rect 1950 105088 1952 105097
rect 2004 105088 2006 105097
rect 1950 105023 2006 105032
rect 1872 104910 1992 104938
rect 1780 103486 1900 103514
rect 1872 101862 1900 103486
rect 1860 101856 1912 101862
rect 1860 101798 1912 101804
rect 1964 97850 1992 104910
rect 2044 103556 2096 103562
rect 2044 103498 2096 103504
rect 2056 103465 2084 103498
rect 2042 103456 2098 103465
rect 2042 103391 2098 103400
rect 2042 102640 2098 102649
rect 2042 102575 2044 102584
rect 2096 102575 2098 102584
rect 2044 102546 2096 102552
rect 2148 98394 2176 110638
rect 2240 101114 2268 112746
rect 2504 111308 2556 111314
rect 2504 111250 2556 111256
rect 2412 107432 2464 107438
rect 2412 107374 2464 107380
rect 2320 105188 2372 105194
rect 2320 105130 2372 105136
rect 2228 101108 2280 101114
rect 2228 101050 2280 101056
rect 2136 98388 2188 98394
rect 2136 98330 2188 98336
rect 1952 97844 2004 97850
rect 1952 97786 2004 97792
rect 2332 92954 2360 105130
rect 2424 95674 2452 107374
rect 2516 99210 2544 111250
rect 2504 99204 2556 99210
rect 2504 99146 2556 99152
rect 2412 95668 2464 95674
rect 2412 95610 2464 95616
rect 2320 92948 2372 92954
rect 2320 92890 2372 92896
rect 1676 91316 1728 91322
rect 1676 91258 1728 91264
rect 2042 90672 2098 90681
rect 2042 90607 2044 90616
rect 2096 90607 2098 90616
rect 2044 90578 2096 90584
rect 2608 79558 2636 114514
rect 2688 113892 2740 113898
rect 2688 113834 2740 113840
rect 2700 109614 2728 113834
rect 2792 113490 2820 114872
rect 2884 114510 2912 118623
rect 2976 117434 3004 118782
rect 2964 117428 3016 117434
rect 2964 117370 3016 117376
rect 2964 116544 3016 116550
rect 2964 116486 3016 116492
rect 2976 115802 3004 116486
rect 3068 115802 3096 119200
rect 3240 116748 3292 116754
rect 3240 116690 3292 116696
rect 3148 116068 3200 116074
rect 3148 116010 3200 116016
rect 2964 115796 3016 115802
rect 2964 115738 3016 115744
rect 3056 115796 3108 115802
rect 3056 115738 3108 115744
rect 2872 114504 2924 114510
rect 2872 114446 2924 114452
rect 3160 114170 3188 116010
rect 3252 115598 3280 116690
rect 3240 115592 3292 115598
rect 3240 115534 3292 115540
rect 3148 114164 3200 114170
rect 3148 114106 3200 114112
rect 3344 113490 3372 119200
rect 3436 114714 3464 119439
rect 3514 119200 3570 120800
rect 3790 119200 3846 120800
rect 3974 119200 4030 120800
rect 4250 119200 4306 120800
rect 4434 119200 4490 120800
rect 4710 119200 4766 120800
rect 4894 119200 4950 120800
rect 5170 119200 5226 120800
rect 5354 119200 5410 120800
rect 5630 119200 5686 120800
rect 5814 119200 5870 120800
rect 6090 119200 6146 120800
rect 6274 119200 6330 120800
rect 6550 119200 6606 120800
rect 6734 119200 6790 120800
rect 7010 119200 7066 120800
rect 7194 119200 7250 120800
rect 7470 119200 7526 120800
rect 7654 119200 7710 120800
rect 7930 119200 7986 120800
rect 8206 119200 8262 120800
rect 8390 119200 8446 120800
rect 8666 119200 8722 120800
rect 8850 119200 8906 120800
rect 9126 119200 9182 120800
rect 9310 119200 9366 120800
rect 9586 119200 9642 120800
rect 9770 119200 9826 120800
rect 10046 119200 10102 120800
rect 10230 119200 10286 120800
rect 10506 119200 10562 120800
rect 10690 119200 10746 120800
rect 10966 119200 11022 120800
rect 11150 119200 11206 120800
rect 11426 119200 11482 120800
rect 11610 119200 11666 120800
rect 11886 119200 11942 120800
rect 12070 119200 12126 120800
rect 12346 119200 12402 120800
rect 12530 119200 12586 120800
rect 12806 119200 12862 120800
rect 12990 119200 13046 120800
rect 13266 119200 13322 120800
rect 13450 119200 13506 120800
rect 13726 119200 13782 120800
rect 13910 119200 13966 120800
rect 14186 119200 14242 120800
rect 14370 119200 14426 120800
rect 14646 119200 14702 120800
rect 14830 119200 14886 120800
rect 15106 119200 15162 120800
rect 15290 119200 15346 120800
rect 15566 119200 15622 120800
rect 15750 119200 15806 120800
rect 16026 119200 16082 120800
rect 16302 119200 16358 120800
rect 16486 119200 16542 120800
rect 16762 119200 16818 120800
rect 16946 119200 17002 120800
rect 17222 119200 17278 120800
rect 17406 119200 17462 120800
rect 17682 119200 17738 120800
rect 17866 119200 17922 120800
rect 18142 119200 18198 120800
rect 18326 119200 18382 120800
rect 18602 119200 18658 120800
rect 18786 119200 18842 120800
rect 19062 119200 19118 120800
rect 19246 119200 19302 120800
rect 19522 119200 19578 120800
rect 19706 119200 19762 120800
rect 19982 119200 20038 120800
rect 20166 119200 20222 120800
rect 20442 119200 20498 120800
rect 20626 119200 20682 120800
rect 20902 119200 20958 120800
rect 21086 119200 21142 120800
rect 21362 119200 21418 120800
rect 21546 119200 21602 120800
rect 21822 119200 21878 120800
rect 22006 119200 22062 120800
rect 22282 119200 22338 120800
rect 22466 119200 22522 120800
rect 22742 119200 22798 120800
rect 22926 119200 22982 120800
rect 23202 119200 23258 120800
rect 23386 119200 23442 120800
rect 23662 119200 23718 120800
rect 23846 119200 23902 120800
rect 24122 119200 24178 120800
rect 24398 119200 24454 120800
rect 24582 119200 24638 120800
rect 24858 119200 24914 120800
rect 25042 119200 25098 120800
rect 25318 119200 25374 120800
rect 25502 119200 25558 120800
rect 25778 119200 25834 120800
rect 25962 119200 26018 120800
rect 26238 119200 26294 120800
rect 26422 119200 26478 120800
rect 26698 119200 26754 120800
rect 26882 119200 26938 120800
rect 27158 119200 27214 120800
rect 27342 119200 27398 120800
rect 27618 119200 27674 120800
rect 27802 119200 27858 120800
rect 28078 119200 28134 120800
rect 28262 119200 28318 120800
rect 28538 119200 28594 120800
rect 28722 119200 28778 120800
rect 28998 119200 29054 120800
rect 29182 119200 29238 120800
rect 29458 119200 29514 120800
rect 29642 119200 29698 120800
rect 29918 119200 29974 120800
rect 30102 119200 30158 120800
rect 30378 119200 30434 120800
rect 30562 119200 30618 120800
rect 30838 119200 30894 120800
rect 31022 119200 31078 120800
rect 31298 119200 31354 120800
rect 31482 119200 31538 120800
rect 31758 119200 31814 120800
rect 31942 119200 31998 120800
rect 32218 119200 32274 120800
rect 32494 119200 32550 120800
rect 32678 119200 32734 120800
rect 32954 119200 33010 120800
rect 33138 119200 33194 120800
rect 33414 119200 33470 120800
rect 33598 119200 33654 120800
rect 33874 119200 33930 120800
rect 34058 119200 34114 120800
rect 34334 119200 34390 120800
rect 34518 119200 34574 120800
rect 34794 119200 34850 120800
rect 34978 119200 35034 120800
rect 35254 119200 35310 120800
rect 35438 119200 35494 120800
rect 35714 119200 35770 120800
rect 35898 119200 35954 120800
rect 36082 119640 36138 119649
rect 36082 119575 36138 119584
rect 3528 115802 3556 119200
rect 3804 116346 3832 119200
rect 3884 116748 3936 116754
rect 3884 116690 3936 116696
rect 3792 116340 3844 116346
rect 3792 116282 3844 116288
rect 3516 115796 3568 115802
rect 3516 115738 3568 115744
rect 3424 114708 3476 114714
rect 3424 114650 3476 114656
rect 3700 114572 3752 114578
rect 3700 114514 3752 114520
rect 2780 113484 2832 113490
rect 2780 113426 2832 113432
rect 3332 113484 3384 113490
rect 3332 113426 3384 113432
rect 2688 109608 2740 109614
rect 2688 109550 2740 109556
rect 3516 108044 3568 108050
rect 3516 107986 3568 107992
rect 2872 106956 2924 106962
rect 2872 106898 2924 106904
rect 2884 94586 2912 106898
rect 3528 96218 3556 107986
rect 3608 104100 3660 104106
rect 3608 104042 3660 104048
rect 3516 96212 3568 96218
rect 3516 96154 3568 96160
rect 2872 94580 2924 94586
rect 2872 94522 2924 94528
rect 2872 90568 2924 90574
rect 2872 90510 2924 90516
rect 2596 79552 2648 79558
rect 2596 79494 2648 79500
rect 2228 72140 2280 72146
rect 2228 72082 2280 72088
rect 2136 70644 2188 70650
rect 2136 70586 2188 70592
rect 2044 69352 2096 69358
rect 2044 69294 2096 69300
rect 1584 68196 1636 68202
rect 1584 68138 1636 68144
rect 1860 50788 1912 50794
rect 1860 50730 1912 50736
rect 1872 50697 1900 50730
rect 1858 50688 1914 50697
rect 1858 50623 1914 50632
rect 1858 49872 1914 49881
rect 1858 49807 1914 49816
rect 1872 49774 1900 49807
rect 1860 49768 1912 49774
rect 1860 49710 1912 49716
rect 1860 49292 1912 49298
rect 1860 49234 1912 49240
rect 1872 49065 1900 49234
rect 1858 49056 1914 49065
rect 1858 48991 1914 49000
rect 1858 48240 1914 48249
rect 1858 48175 1860 48184
rect 1912 48175 1914 48184
rect 1860 48146 1912 48152
rect 1860 47524 1912 47530
rect 1860 47466 1912 47472
rect 1872 47433 1900 47466
rect 1952 47456 2004 47462
rect 1858 47424 1914 47433
rect 1952 47398 2004 47404
rect 1858 47359 1914 47368
rect 1964 47258 1992 47398
rect 1952 47252 2004 47258
rect 1952 47194 2004 47200
rect 1858 46744 1914 46753
rect 1858 46679 1914 46688
rect 1872 46510 1900 46679
rect 1860 46504 1912 46510
rect 1860 46446 1912 46452
rect 1860 46028 1912 46034
rect 1860 45970 1912 45976
rect 1872 45937 1900 45970
rect 1858 45928 1914 45937
rect 1858 45863 1914 45872
rect 1412 45526 1532 45554
rect 1308 18760 1360 18766
rect 1308 18702 1360 18708
rect 1032 3732 1084 3738
rect 1032 3674 1084 3680
rect 112 3528 164 3534
rect 112 3470 164 3476
rect 124 800 152 3470
rect 388 2984 440 2990
rect 388 2926 440 2932
rect 400 800 428 2926
rect 756 2848 808 2854
rect 756 2790 808 2796
rect 768 800 796 2790
rect 1044 800 1072 3674
rect 1320 3534 1348 18702
rect 1412 16574 1440 45526
rect 1858 45112 1914 45121
rect 1858 45047 1914 45056
rect 1872 45014 1900 45047
rect 1860 45008 1912 45014
rect 1860 44950 1912 44956
rect 1858 44296 1914 44305
rect 1858 44231 1860 44240
rect 1912 44231 1914 44240
rect 1860 44202 1912 44208
rect 1858 43480 1914 43489
rect 1858 43415 1914 43424
rect 1872 43246 1900 43415
rect 1860 43240 1912 43246
rect 1860 43182 1912 43188
rect 1952 43104 2004 43110
rect 1952 43046 2004 43052
rect 1964 42906 1992 43046
rect 1952 42900 2004 42906
rect 1952 42842 2004 42848
rect 1860 42764 1912 42770
rect 1860 42706 1912 42712
rect 1872 42673 1900 42706
rect 1858 42664 1914 42673
rect 1858 42599 1914 42608
rect 1858 41848 1914 41857
rect 1858 41783 1914 41792
rect 1872 41750 1900 41783
rect 1860 41744 1912 41750
rect 1860 41686 1912 41692
rect 1858 41032 1914 41041
rect 1858 40967 1860 40976
rect 1912 40967 1914 40976
rect 1860 40938 1912 40944
rect 1860 40588 1912 40594
rect 1860 40530 1912 40536
rect 1872 40361 1900 40530
rect 1858 40352 1914 40361
rect 1858 40287 1914 40296
rect 1858 39536 1914 39545
rect 1858 39471 1860 39480
rect 1912 39471 1914 39480
rect 1860 39442 1912 39448
rect 1860 38820 1912 38826
rect 1860 38762 1912 38768
rect 1872 38729 1900 38762
rect 1858 38720 1914 38729
rect 1858 38655 1914 38664
rect 1858 37904 1914 37913
rect 1858 37839 1914 37848
rect 1872 37806 1900 37839
rect 1860 37800 1912 37806
rect 1860 37742 1912 37748
rect 1860 37324 1912 37330
rect 1860 37266 1912 37272
rect 1872 37097 1900 37266
rect 1858 37088 1914 37097
rect 1858 37023 1914 37032
rect 1858 36272 1914 36281
rect 1858 36207 1860 36216
rect 1912 36207 1914 36216
rect 1860 36178 1912 36184
rect 1860 35556 1912 35562
rect 1860 35498 1912 35504
rect 1872 35465 1900 35498
rect 1858 35456 1914 35465
rect 1858 35391 1914 35400
rect 1858 34640 1914 34649
rect 1858 34575 1914 34584
rect 1872 34474 1900 34575
rect 1860 34468 1912 34474
rect 1860 34410 1912 34416
rect 1860 34060 1912 34066
rect 1860 34002 1912 34008
rect 1872 33833 1900 34002
rect 1858 33824 1914 33833
rect 1858 33759 1914 33768
rect 1858 33144 1914 33153
rect 1858 33079 1914 33088
rect 1872 33046 1900 33079
rect 1860 33040 1912 33046
rect 1860 32982 1912 32988
rect 1952 32768 2004 32774
rect 1952 32710 2004 32716
rect 1858 32328 1914 32337
rect 1858 32263 1860 32272
rect 1912 32263 1914 32272
rect 1860 32234 1912 32240
rect 1858 31512 1914 31521
rect 1858 31447 1914 31456
rect 1872 31278 1900 31447
rect 1860 31272 1912 31278
rect 1860 31214 1912 31220
rect 1860 30796 1912 30802
rect 1860 30738 1912 30744
rect 1872 30705 1900 30738
rect 1964 30734 1992 32710
rect 1952 30728 2004 30734
rect 1858 30696 1914 30705
rect 1952 30670 2004 30676
rect 1858 30631 1914 30640
rect 1952 30592 2004 30598
rect 1952 30534 2004 30540
rect 1964 30394 1992 30534
rect 1952 30388 2004 30394
rect 1952 30330 2004 30336
rect 1858 29880 1914 29889
rect 1858 29815 1914 29824
rect 1872 29782 1900 29815
rect 1860 29776 1912 29782
rect 1860 29718 1912 29724
rect 1860 29096 1912 29102
rect 1858 29064 1860 29073
rect 1912 29064 1914 29073
rect 1858 28999 1914 29008
rect 1858 28248 1914 28257
rect 1858 28183 1914 28192
rect 1872 28014 1900 28183
rect 1860 28008 1912 28014
rect 1860 27950 1912 27956
rect 1860 27532 1912 27538
rect 1860 27474 1912 27480
rect 1872 27441 1900 27474
rect 1858 27432 1914 27441
rect 1858 27367 1914 27376
rect 1860 26852 1912 26858
rect 1860 26794 1912 26800
rect 1872 26761 1900 26794
rect 1858 26752 1914 26761
rect 1858 26687 1914 26696
rect 1858 25936 1914 25945
rect 1858 25871 1914 25880
rect 1872 25838 1900 25871
rect 1860 25832 1912 25838
rect 1860 25774 1912 25780
rect 1860 25356 1912 25362
rect 1860 25298 1912 25304
rect 1872 25129 1900 25298
rect 1858 25120 1914 25129
rect 1858 25055 1914 25064
rect 1858 24304 1914 24313
rect 1858 24239 1860 24248
rect 1912 24239 1914 24248
rect 1860 24210 1912 24216
rect 1860 23588 1912 23594
rect 1860 23530 1912 23536
rect 1872 23497 1900 23530
rect 1858 23488 1914 23497
rect 1858 23423 1914 23432
rect 1858 22672 1914 22681
rect 1858 22607 1914 22616
rect 1872 22574 1900 22607
rect 1860 22568 1912 22574
rect 1860 22510 1912 22516
rect 1860 22160 1912 22166
rect 1860 22102 1912 22108
rect 1872 21865 1900 22102
rect 1858 21856 1914 21865
rect 1858 21791 1914 21800
rect 1858 21040 1914 21049
rect 1858 20975 1860 20984
rect 1912 20975 1914 20984
rect 1860 20946 1912 20952
rect 1858 20360 1914 20369
rect 1858 20295 1860 20304
rect 1912 20295 1914 20304
rect 1860 20266 1912 20272
rect 1858 19544 1914 19553
rect 1858 19479 1914 19488
rect 1872 19310 1900 19479
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 1860 18828 1912 18834
rect 1860 18770 1912 18776
rect 1872 18737 1900 18770
rect 1858 18728 1914 18737
rect 1858 18663 1914 18672
rect 1858 17912 1914 17921
rect 1858 17847 1914 17856
rect 1872 17814 1900 17847
rect 1860 17808 1912 17814
rect 1860 17750 1912 17756
rect 1858 17096 1914 17105
rect 1858 17031 1860 17040
rect 1912 17031 1914 17040
rect 1860 17002 1912 17008
rect 1412 16546 1624 16574
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1412 2689 1440 3538
rect 1398 2680 1454 2689
rect 1398 2615 1454 2624
rect 1504 2258 1532 4014
rect 1596 2446 1624 16546
rect 1858 16280 1914 16289
rect 1858 16215 1914 16224
rect 1872 16046 1900 16215
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 1872 15473 1900 15506
rect 1858 15464 1914 15473
rect 1858 15399 1914 15408
rect 1858 14648 1914 14657
rect 1858 14583 1914 14592
rect 1872 14550 1900 14583
rect 1860 14544 1912 14550
rect 1860 14486 1912 14492
rect 1860 13864 1912 13870
rect 1858 13832 1860 13841
rect 1912 13832 1914 13841
rect 1858 13767 1914 13776
rect 1860 13388 1912 13394
rect 1860 13330 1912 13336
rect 1872 13161 1900 13330
rect 1858 13152 1914 13161
rect 1858 13087 1914 13096
rect 1858 12336 1914 12345
rect 1858 12271 1860 12280
rect 1912 12271 1914 12280
rect 1860 12242 1912 12248
rect 1860 11620 1912 11626
rect 1860 11562 1912 11568
rect 1872 11529 1900 11562
rect 1858 11520 1914 11529
rect 1858 11455 1914 11464
rect 1858 10704 1914 10713
rect 1858 10639 1914 10648
rect 1872 10606 1900 10639
rect 1860 10600 1912 10606
rect 1860 10542 1912 10548
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1872 9897 1900 10066
rect 1858 9888 1914 9897
rect 1858 9823 1914 9832
rect 1858 9072 1914 9081
rect 1858 9007 1860 9016
rect 1912 9007 1914 9016
rect 1860 8978 1912 8984
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 1872 8265 1900 8298
rect 1858 8256 1914 8265
rect 1858 8191 1914 8200
rect 1858 7440 1914 7449
rect 1858 7375 1914 7384
rect 1872 7342 1900 7375
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1872 6769 1900 6802
rect 1858 6760 1914 6769
rect 1858 6695 1914 6704
rect 1858 5944 1914 5953
rect 1858 5879 1914 5888
rect 1872 5846 1900 5879
rect 1860 5840 1912 5846
rect 1860 5782 1912 5788
rect 1858 5128 1914 5137
rect 1858 5063 1860 5072
rect 1912 5063 1914 5072
rect 1860 5034 1912 5040
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 1872 4321 1900 4626
rect 1858 4312 1914 4321
rect 1858 4247 1914 4256
rect 2056 4146 2084 69294
rect 2148 6798 2176 70586
rect 2240 14074 2268 72082
rect 2504 71052 2556 71058
rect 2504 70994 2556 71000
rect 2412 55956 2464 55962
rect 2412 55898 2464 55904
rect 2320 51264 2372 51270
rect 2320 51206 2372 51212
rect 2332 49910 2360 51206
rect 2320 49904 2372 49910
rect 2320 49846 2372 49852
rect 2320 49224 2372 49230
rect 2320 49166 2372 49172
rect 2332 48278 2360 49166
rect 2320 48272 2372 48278
rect 2320 48214 2372 48220
rect 2424 45554 2452 55898
rect 2332 45526 2452 45554
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2136 5840 2188 5846
rect 2136 5782 2188 5788
rect 2148 5370 2176 5782
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2240 4758 2268 5646
rect 2228 4752 2280 4758
rect 2228 4694 2280 4700
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1872 3505 1900 3946
rect 1858 3496 1914 3505
rect 1858 3431 1914 3440
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 1412 2230 1532 2258
rect 1412 800 1440 2230
rect 1688 800 1716 3334
rect 2332 3194 2360 45526
rect 2412 35556 2464 35562
rect 2412 35498 2464 35504
rect 2424 32570 2452 35498
rect 2412 32564 2464 32570
rect 2412 32506 2464 32512
rect 2412 32292 2464 32298
rect 2412 32234 2464 32240
rect 2424 30054 2452 32234
rect 2412 30048 2464 30054
rect 2412 29990 2464 29996
rect 2412 27940 2464 27946
rect 2412 27882 2464 27888
rect 2424 25702 2452 27882
rect 2412 25696 2464 25702
rect 2412 25638 2464 25644
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2044 3120 2096 3126
rect 2044 3062 2096 3068
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 1872 1057 1900 2858
rect 1858 1048 1914 1057
rect 1858 983 1914 992
rect 2056 800 2084 3062
rect 2424 2938 2452 5714
rect 2516 3670 2544 70994
rect 2688 41540 2740 41546
rect 2688 41482 2740 41488
rect 2700 41070 2728 41482
rect 2688 41064 2740 41070
rect 2688 41006 2740 41012
rect 2596 40996 2648 41002
rect 2596 40938 2648 40944
rect 2608 40050 2636 40938
rect 2688 40452 2740 40458
rect 2688 40394 2740 40400
rect 2596 40044 2648 40050
rect 2596 39986 2648 39992
rect 2700 39506 2728 40394
rect 2688 39500 2740 39506
rect 2688 39442 2740 39448
rect 2688 39364 2740 39370
rect 2688 39306 2740 39312
rect 2596 38820 2648 38826
rect 2596 38762 2648 38768
rect 2608 36582 2636 38762
rect 2700 37670 2728 39306
rect 2688 37664 2740 37670
rect 2688 37606 2740 37612
rect 2688 37324 2740 37330
rect 2688 37266 2740 37272
rect 2596 36576 2648 36582
rect 2596 36518 2648 36524
rect 2700 36394 2728 37266
rect 2608 36366 2728 36394
rect 2608 35630 2636 36366
rect 2688 36100 2740 36106
rect 2688 36042 2740 36048
rect 2596 35624 2648 35630
rect 2596 35566 2648 35572
rect 2700 34950 2728 36042
rect 2688 34944 2740 34950
rect 2688 34886 2740 34892
rect 2596 34536 2648 34542
rect 2596 34478 2648 34484
rect 2608 31822 2636 34478
rect 2688 33924 2740 33930
rect 2688 33866 2740 33872
rect 2596 31816 2648 31822
rect 2596 31758 2648 31764
rect 2700 31278 2728 33866
rect 2688 31272 2740 31278
rect 2688 31214 2740 31220
rect 2596 31204 2648 31210
rect 2596 31146 2648 31152
rect 2608 28082 2636 31146
rect 2688 29572 2740 29578
rect 2688 29514 2740 29520
rect 2596 28076 2648 28082
rect 2596 28018 2648 28024
rect 2700 26994 2728 29514
rect 2688 26988 2740 26994
rect 2688 26930 2740 26936
rect 2596 26852 2648 26858
rect 2596 26794 2648 26800
rect 2608 25158 2636 26794
rect 2688 25764 2740 25770
rect 2688 25706 2740 25712
rect 2596 25152 2648 25158
rect 2596 25094 2648 25100
rect 2700 24682 2728 25706
rect 2688 24676 2740 24682
rect 2688 24618 2740 24624
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2504 3664 2556 3670
rect 2504 3606 2556 3612
rect 2332 2910 2452 2938
rect 2332 800 2360 2910
rect 2700 800 2728 3946
rect 2792 3738 2820 5170
rect 2884 4282 2912 90510
rect 3424 71120 3476 71126
rect 3424 71062 3476 71068
rect 3148 64388 3200 64394
rect 3148 64330 3200 64336
rect 2964 56228 3016 56234
rect 2964 56170 3016 56176
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2976 2650 3004 56170
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3068 3194 3096 14418
rect 3160 4758 3188 64330
rect 3436 7546 3464 71062
rect 3516 53644 3568 53650
rect 3516 53586 3568 53592
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3252 4758 3280 5510
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 3160 2854 3188 4490
rect 3528 3738 3556 53586
rect 3620 50386 3648 104042
rect 3712 62150 3740 114514
rect 3896 114102 3924 116690
rect 3884 114096 3936 114102
rect 3884 114038 3936 114044
rect 3988 113490 4016 119200
rect 4264 117858 4292 119200
rect 4448 118130 4476 119200
rect 4724 118250 4752 119200
rect 4712 118244 4764 118250
rect 4712 118186 4764 118192
rect 4448 118102 4844 118130
rect 4712 117972 4764 117978
rect 4712 117914 4764 117920
rect 4264 117830 4660 117858
rect 4220 117532 4516 117552
rect 4276 117530 4300 117532
rect 4356 117530 4380 117532
rect 4436 117530 4460 117532
rect 4298 117478 4300 117530
rect 4362 117478 4374 117530
rect 4436 117478 4438 117530
rect 4276 117476 4300 117478
rect 4356 117476 4380 117478
rect 4436 117476 4460 117478
rect 4220 117456 4516 117476
rect 4068 117156 4120 117162
rect 4068 117098 4120 117104
rect 4528 117156 4580 117162
rect 4528 117098 4580 117104
rect 4080 116890 4108 117098
rect 4068 116884 4120 116890
rect 4068 116826 4120 116832
rect 4540 116634 4568 117098
rect 4632 116822 4660 117830
rect 4620 116816 4672 116822
rect 4620 116758 4672 116764
rect 4540 116606 4660 116634
rect 4220 116444 4516 116464
rect 4276 116442 4300 116444
rect 4356 116442 4380 116444
rect 4436 116442 4460 116444
rect 4298 116390 4300 116442
rect 4362 116390 4374 116442
rect 4436 116390 4438 116442
rect 4276 116388 4300 116390
rect 4356 116388 4380 116390
rect 4436 116388 4460 116390
rect 4220 116368 4516 116388
rect 4632 115818 4660 116606
rect 4448 115790 4660 115818
rect 4068 115660 4120 115666
rect 4068 115602 4120 115608
rect 4080 114510 4108 115602
rect 4448 115598 4476 115790
rect 4620 115660 4672 115666
rect 4620 115602 4672 115608
rect 4436 115592 4488 115598
rect 4436 115534 4488 115540
rect 4220 115356 4516 115376
rect 4276 115354 4300 115356
rect 4356 115354 4380 115356
rect 4436 115354 4460 115356
rect 4298 115302 4300 115354
rect 4362 115302 4374 115354
rect 4436 115302 4438 115354
rect 4276 115300 4300 115302
rect 4356 115300 4380 115302
rect 4436 115300 4460 115302
rect 4220 115280 4516 115300
rect 4068 114504 4120 114510
rect 4068 114446 4120 114452
rect 4220 114268 4516 114288
rect 4276 114266 4300 114268
rect 4356 114266 4380 114268
rect 4436 114266 4460 114268
rect 4298 114214 4300 114266
rect 4362 114214 4374 114266
rect 4436 114214 4438 114266
rect 4276 114212 4300 114214
rect 4356 114212 4380 114214
rect 4436 114212 4460 114214
rect 4220 114192 4516 114212
rect 4632 114170 4660 115602
rect 4620 114164 4672 114170
rect 4620 114106 4672 114112
rect 4724 113490 4752 117914
rect 4816 115734 4844 118102
rect 4908 116890 4936 119200
rect 4896 116884 4948 116890
rect 4896 116826 4948 116832
rect 5080 116748 5132 116754
rect 5080 116690 5132 116696
rect 4988 116680 5040 116686
rect 4988 116622 5040 116628
rect 4896 116068 4948 116074
rect 4896 116010 4948 116016
rect 4804 115728 4856 115734
rect 4804 115670 4856 115676
rect 4804 115592 4856 115598
rect 4804 115534 4856 115540
rect 4816 113898 4844 115534
rect 4908 114510 4936 116010
rect 5000 115122 5028 116622
rect 5092 115258 5120 116690
rect 5184 115802 5212 119200
rect 5172 115796 5224 115802
rect 5172 115738 5224 115744
rect 5264 115660 5316 115666
rect 5264 115602 5316 115608
rect 5172 115592 5224 115598
rect 5172 115534 5224 115540
rect 5080 115252 5132 115258
rect 5080 115194 5132 115200
rect 4988 115116 5040 115122
rect 4988 115058 5040 115064
rect 5184 114918 5212 115534
rect 5172 114912 5224 114918
rect 5172 114854 5224 114860
rect 5276 114578 5304 115602
rect 5264 114572 5316 114578
rect 5264 114514 5316 114520
rect 4896 114504 4948 114510
rect 4896 114446 4948 114452
rect 4804 113892 4856 113898
rect 4804 113834 4856 113840
rect 5368 113490 5396 119200
rect 5448 117224 5500 117230
rect 5448 117166 5500 117172
rect 5460 116346 5488 117166
rect 5540 116680 5592 116686
rect 5540 116622 5592 116628
rect 5448 116340 5500 116346
rect 5448 116282 5500 116288
rect 5448 116204 5500 116210
rect 5448 116146 5500 116152
rect 5460 114170 5488 116146
rect 5552 115190 5580 116622
rect 5644 116346 5672 119200
rect 5724 116544 5776 116550
rect 5724 116486 5776 116492
rect 5632 116340 5684 116346
rect 5632 116282 5684 116288
rect 5736 116142 5764 116486
rect 5828 116328 5856 119200
rect 6000 116816 6052 116822
rect 6000 116758 6052 116764
rect 5908 116340 5960 116346
rect 5828 116300 5908 116328
rect 5908 116282 5960 116288
rect 5724 116136 5776 116142
rect 5724 116078 5776 116084
rect 5540 115184 5592 115190
rect 5540 115126 5592 115132
rect 5540 114912 5592 114918
rect 5540 114854 5592 114860
rect 5448 114164 5500 114170
rect 5448 114106 5500 114112
rect 5552 113966 5580 114854
rect 5540 113960 5592 113966
rect 5540 113902 5592 113908
rect 6012 113830 6040 116758
rect 6000 113824 6052 113830
rect 6000 113766 6052 113772
rect 6104 113490 6132 119200
rect 6184 117292 6236 117298
rect 6184 117234 6236 117240
rect 6196 115530 6224 117234
rect 6288 116890 6316 119200
rect 6276 116884 6328 116890
rect 6276 116826 6328 116832
rect 6276 116612 6328 116618
rect 6276 116554 6328 116560
rect 6184 115524 6236 115530
rect 6184 115466 6236 115472
rect 6288 114578 6316 116554
rect 6564 116362 6592 119200
rect 6564 116346 6684 116362
rect 6564 116340 6696 116346
rect 6564 116334 6644 116340
rect 6644 116282 6696 116288
rect 6460 116068 6512 116074
rect 6460 116010 6512 116016
rect 6276 114572 6328 114578
rect 6276 114514 6328 114520
rect 6472 114170 6500 116010
rect 6460 114164 6512 114170
rect 6460 114106 6512 114112
rect 6748 113558 6776 119200
rect 6828 117156 6880 117162
rect 6828 117098 6880 117104
rect 6840 114714 6868 117098
rect 7024 116872 7052 119200
rect 7104 116884 7156 116890
rect 7024 116844 7104 116872
rect 7104 116826 7156 116832
rect 6920 116748 6972 116754
rect 6920 116690 6972 116696
rect 7104 116748 7156 116754
rect 7104 116690 7156 116696
rect 6932 115258 6960 116690
rect 7012 116068 7064 116074
rect 7012 116010 7064 116016
rect 6920 115252 6972 115258
rect 6920 115194 6972 115200
rect 6920 115116 6972 115122
rect 6920 115058 6972 115064
rect 6828 114708 6880 114714
rect 6828 114650 6880 114656
rect 6932 113966 6960 115058
rect 7024 114510 7052 116010
rect 7116 115258 7144 116690
rect 7208 116278 7236 119200
rect 7380 117088 7432 117094
rect 7380 117030 7432 117036
rect 7196 116272 7248 116278
rect 7196 116214 7248 116220
rect 7104 115252 7156 115258
rect 7104 115194 7156 115200
rect 7196 114640 7248 114646
rect 7196 114582 7248 114588
rect 7012 114504 7064 114510
rect 7012 114446 7064 114452
rect 6920 113960 6972 113966
rect 6920 113902 6972 113908
rect 6736 113552 6788 113558
rect 6736 113494 6788 113500
rect 3976 113484 4028 113490
rect 3976 113426 4028 113432
rect 4712 113484 4764 113490
rect 4712 113426 4764 113432
rect 5356 113484 5408 113490
rect 5356 113426 5408 113432
rect 6092 113484 6144 113490
rect 6092 113426 6144 113432
rect 4220 113180 4516 113200
rect 4276 113178 4300 113180
rect 4356 113178 4380 113180
rect 4436 113178 4460 113180
rect 4298 113126 4300 113178
rect 4362 113126 4374 113178
rect 4436 113126 4438 113178
rect 4276 113124 4300 113126
rect 4356 113124 4380 113126
rect 4436 113124 4460 113126
rect 4220 113104 4516 113124
rect 6276 112396 6328 112402
rect 6276 112338 6328 112344
rect 4220 112092 4516 112112
rect 4276 112090 4300 112092
rect 4356 112090 4380 112092
rect 4436 112090 4460 112092
rect 4298 112038 4300 112090
rect 4362 112038 4374 112090
rect 4436 112038 4438 112090
rect 4276 112036 4300 112038
rect 4356 112036 4380 112038
rect 4436 112036 4460 112038
rect 4220 112016 4516 112036
rect 4220 111004 4516 111024
rect 4276 111002 4300 111004
rect 4356 111002 4380 111004
rect 4436 111002 4460 111004
rect 4298 110950 4300 111002
rect 4362 110950 4374 111002
rect 4436 110950 4438 111002
rect 4276 110948 4300 110950
rect 4356 110948 4380 110950
rect 4436 110948 4460 110950
rect 4220 110928 4516 110948
rect 4220 109916 4516 109936
rect 4276 109914 4300 109916
rect 4356 109914 4380 109916
rect 4436 109914 4460 109916
rect 4298 109862 4300 109914
rect 4362 109862 4374 109914
rect 4436 109862 4438 109914
rect 4276 109860 4300 109862
rect 4356 109860 4380 109862
rect 4436 109860 4460 109862
rect 4220 109840 4516 109860
rect 4220 108828 4516 108848
rect 4276 108826 4300 108828
rect 4356 108826 4380 108828
rect 4436 108826 4460 108828
rect 4298 108774 4300 108826
rect 4362 108774 4374 108826
rect 4436 108774 4438 108826
rect 4276 108772 4300 108774
rect 4356 108772 4380 108774
rect 4436 108772 4460 108774
rect 4220 108752 4516 108772
rect 4220 107740 4516 107760
rect 4276 107738 4300 107740
rect 4356 107738 4380 107740
rect 4436 107738 4460 107740
rect 4298 107686 4300 107738
rect 4362 107686 4374 107738
rect 4436 107686 4438 107738
rect 4276 107684 4300 107686
rect 4356 107684 4380 107686
rect 4436 107684 4460 107686
rect 4220 107664 4516 107684
rect 4220 106652 4516 106672
rect 4276 106650 4300 106652
rect 4356 106650 4380 106652
rect 4436 106650 4460 106652
rect 4298 106598 4300 106650
rect 4362 106598 4374 106650
rect 4436 106598 4438 106650
rect 4276 106596 4300 106598
rect 4356 106596 4380 106598
rect 4436 106596 4460 106598
rect 4220 106576 4516 106596
rect 4220 105564 4516 105584
rect 4276 105562 4300 105564
rect 4356 105562 4380 105564
rect 4436 105562 4460 105564
rect 4298 105510 4300 105562
rect 4362 105510 4374 105562
rect 4436 105510 4438 105562
rect 4276 105508 4300 105510
rect 4356 105508 4380 105510
rect 4436 105508 4460 105510
rect 4220 105488 4516 105508
rect 4220 104476 4516 104496
rect 4276 104474 4300 104476
rect 4356 104474 4380 104476
rect 4436 104474 4460 104476
rect 4298 104422 4300 104474
rect 4362 104422 4374 104474
rect 4436 104422 4438 104474
rect 4276 104420 4300 104422
rect 4356 104420 4380 104422
rect 4436 104420 4460 104422
rect 4220 104400 4516 104420
rect 4220 103388 4516 103408
rect 4276 103386 4300 103388
rect 4356 103386 4380 103388
rect 4436 103386 4460 103388
rect 4298 103334 4300 103386
rect 4362 103334 4374 103386
rect 4436 103334 4438 103386
rect 4276 103332 4300 103334
rect 4356 103332 4380 103334
rect 4436 103332 4460 103334
rect 4220 103312 4516 103332
rect 4220 102300 4516 102320
rect 4276 102298 4300 102300
rect 4356 102298 4380 102300
rect 4436 102298 4460 102300
rect 4298 102246 4300 102298
rect 4362 102246 4374 102298
rect 4436 102246 4438 102298
rect 4276 102244 4300 102246
rect 4356 102244 4380 102246
rect 4436 102244 4460 102246
rect 4220 102224 4516 102244
rect 4220 101212 4516 101232
rect 4276 101210 4300 101212
rect 4356 101210 4380 101212
rect 4436 101210 4460 101212
rect 4298 101158 4300 101210
rect 4362 101158 4374 101210
rect 4436 101158 4438 101210
rect 4276 101156 4300 101158
rect 4356 101156 4380 101158
rect 4436 101156 4460 101158
rect 4220 101136 4516 101156
rect 4220 100124 4516 100144
rect 4276 100122 4300 100124
rect 4356 100122 4380 100124
rect 4436 100122 4460 100124
rect 4298 100070 4300 100122
rect 4362 100070 4374 100122
rect 4436 100070 4438 100122
rect 4276 100068 4300 100070
rect 4356 100068 4380 100070
rect 4436 100068 4460 100070
rect 4220 100048 4516 100068
rect 6288 100026 6316 112338
rect 7208 103514 7236 114582
rect 7392 114578 7420 117030
rect 7380 114572 7432 114578
rect 7380 114514 7432 114520
rect 7484 113506 7512 119200
rect 7564 117156 7616 117162
rect 7564 117098 7616 117104
rect 7576 114170 7604 117098
rect 7668 116550 7696 119200
rect 7748 117156 7800 117162
rect 7748 117098 7800 117104
rect 7760 116686 7788 117098
rect 7840 117088 7892 117094
rect 7840 117030 7892 117036
rect 7748 116680 7800 116686
rect 7748 116622 7800 116628
rect 7656 116544 7708 116550
rect 7656 116486 7708 116492
rect 7852 115802 7880 117030
rect 7944 116226 7972 119200
rect 7944 116198 8064 116226
rect 7932 116068 7984 116074
rect 7932 116010 7984 116016
rect 7840 115796 7892 115802
rect 7840 115738 7892 115744
rect 7748 115456 7800 115462
rect 7748 115398 7800 115404
rect 7656 114980 7708 114986
rect 7656 114922 7708 114928
rect 7668 114578 7696 114922
rect 7656 114572 7708 114578
rect 7656 114514 7708 114520
rect 7564 114164 7616 114170
rect 7564 114106 7616 114112
rect 7484 113490 7604 113506
rect 7484 113484 7616 113490
rect 7484 113478 7564 113484
rect 7564 113426 7616 113432
rect 7116 103486 7236 103514
rect 7116 103290 7144 103486
rect 7104 103284 7156 103290
rect 7104 103226 7156 103232
rect 7012 103080 7064 103086
rect 7012 103022 7064 103028
rect 6276 100020 6328 100026
rect 6276 99962 6328 99968
rect 5080 99340 5132 99346
rect 5080 99282 5132 99288
rect 4220 99036 4516 99056
rect 4276 99034 4300 99036
rect 4356 99034 4380 99036
rect 4436 99034 4460 99036
rect 4298 98982 4300 99034
rect 4362 98982 4374 99034
rect 4436 98982 4438 99034
rect 4276 98980 4300 98982
rect 4356 98980 4380 98982
rect 4436 98980 4460 98982
rect 4220 98960 4516 98980
rect 4896 98252 4948 98258
rect 4896 98194 4948 98200
rect 4220 97948 4516 97968
rect 4276 97946 4300 97948
rect 4356 97946 4380 97948
rect 4436 97946 4460 97948
rect 4298 97894 4300 97946
rect 4362 97894 4374 97946
rect 4436 97894 4438 97946
rect 4276 97892 4300 97894
rect 4356 97892 4380 97894
rect 4436 97892 4460 97894
rect 4220 97872 4516 97892
rect 4220 96860 4516 96880
rect 4276 96858 4300 96860
rect 4356 96858 4380 96860
rect 4436 96858 4460 96860
rect 4298 96806 4300 96858
rect 4362 96806 4374 96858
rect 4436 96806 4438 96858
rect 4276 96804 4300 96806
rect 4356 96804 4380 96806
rect 4436 96804 4460 96806
rect 4220 96784 4516 96804
rect 4220 95772 4516 95792
rect 4276 95770 4300 95772
rect 4356 95770 4380 95772
rect 4436 95770 4460 95772
rect 4298 95718 4300 95770
rect 4362 95718 4374 95770
rect 4436 95718 4438 95770
rect 4276 95716 4300 95718
rect 4356 95716 4380 95718
rect 4436 95716 4460 95718
rect 4220 95696 4516 95716
rect 4220 94684 4516 94704
rect 4276 94682 4300 94684
rect 4356 94682 4380 94684
rect 4436 94682 4460 94684
rect 4298 94630 4300 94682
rect 4362 94630 4374 94682
rect 4436 94630 4438 94682
rect 4276 94628 4300 94630
rect 4356 94628 4380 94630
rect 4436 94628 4460 94630
rect 4220 94608 4516 94628
rect 4220 93596 4516 93616
rect 4276 93594 4300 93596
rect 4356 93594 4380 93596
rect 4436 93594 4460 93596
rect 4298 93542 4300 93594
rect 4362 93542 4374 93594
rect 4436 93542 4438 93594
rect 4276 93540 4300 93542
rect 4356 93540 4380 93542
rect 4436 93540 4460 93542
rect 4220 93520 4516 93540
rect 4804 92812 4856 92818
rect 4804 92754 4856 92760
rect 4220 92508 4516 92528
rect 4276 92506 4300 92508
rect 4356 92506 4380 92508
rect 4436 92506 4460 92508
rect 4298 92454 4300 92506
rect 4362 92454 4374 92506
rect 4436 92454 4438 92506
rect 4276 92452 4300 92454
rect 4356 92452 4380 92454
rect 4436 92452 4460 92454
rect 4220 92432 4516 92452
rect 4220 91420 4516 91440
rect 4276 91418 4300 91420
rect 4356 91418 4380 91420
rect 4436 91418 4460 91420
rect 4298 91366 4300 91418
rect 4362 91366 4374 91418
rect 4436 91366 4438 91418
rect 4276 91364 4300 91366
rect 4356 91364 4380 91366
rect 4436 91364 4460 91366
rect 4220 91344 4516 91364
rect 4220 90332 4516 90352
rect 4276 90330 4300 90332
rect 4356 90330 4380 90332
rect 4436 90330 4460 90332
rect 4298 90278 4300 90330
rect 4362 90278 4374 90330
rect 4436 90278 4438 90330
rect 4276 90276 4300 90278
rect 4356 90276 4380 90278
rect 4436 90276 4460 90278
rect 4220 90256 4516 90276
rect 4220 89244 4516 89264
rect 4276 89242 4300 89244
rect 4356 89242 4380 89244
rect 4436 89242 4460 89244
rect 4298 89190 4300 89242
rect 4362 89190 4374 89242
rect 4436 89190 4438 89242
rect 4276 89188 4300 89190
rect 4356 89188 4380 89190
rect 4436 89188 4460 89190
rect 4220 89168 4516 89188
rect 4220 88156 4516 88176
rect 4276 88154 4300 88156
rect 4356 88154 4380 88156
rect 4436 88154 4460 88156
rect 4298 88102 4300 88154
rect 4362 88102 4374 88154
rect 4436 88102 4438 88154
rect 4276 88100 4300 88102
rect 4356 88100 4380 88102
rect 4436 88100 4460 88102
rect 4220 88080 4516 88100
rect 4220 87068 4516 87088
rect 4276 87066 4300 87068
rect 4356 87066 4380 87068
rect 4436 87066 4460 87068
rect 4298 87014 4300 87066
rect 4362 87014 4374 87066
rect 4436 87014 4438 87066
rect 4276 87012 4300 87014
rect 4356 87012 4380 87014
rect 4436 87012 4460 87014
rect 4220 86992 4516 87012
rect 4220 85980 4516 86000
rect 4276 85978 4300 85980
rect 4356 85978 4380 85980
rect 4436 85978 4460 85980
rect 4298 85926 4300 85978
rect 4362 85926 4374 85978
rect 4436 85926 4438 85978
rect 4276 85924 4300 85926
rect 4356 85924 4380 85926
rect 4436 85924 4460 85926
rect 4220 85904 4516 85924
rect 4220 84892 4516 84912
rect 4276 84890 4300 84892
rect 4356 84890 4380 84892
rect 4436 84890 4460 84892
rect 4298 84838 4300 84890
rect 4362 84838 4374 84890
rect 4436 84838 4438 84890
rect 4276 84836 4300 84838
rect 4356 84836 4380 84838
rect 4436 84836 4460 84838
rect 4220 84816 4516 84836
rect 4220 83804 4516 83824
rect 4276 83802 4300 83804
rect 4356 83802 4380 83804
rect 4436 83802 4460 83804
rect 4298 83750 4300 83802
rect 4362 83750 4374 83802
rect 4436 83750 4438 83802
rect 4276 83748 4300 83750
rect 4356 83748 4380 83750
rect 4436 83748 4460 83750
rect 4220 83728 4516 83748
rect 4220 82716 4516 82736
rect 4276 82714 4300 82716
rect 4356 82714 4380 82716
rect 4436 82714 4460 82716
rect 4298 82662 4300 82714
rect 4362 82662 4374 82714
rect 4436 82662 4438 82714
rect 4276 82660 4300 82662
rect 4356 82660 4380 82662
rect 4436 82660 4460 82662
rect 4220 82640 4516 82660
rect 4220 81628 4516 81648
rect 4276 81626 4300 81628
rect 4356 81626 4380 81628
rect 4436 81626 4460 81628
rect 4298 81574 4300 81626
rect 4362 81574 4374 81626
rect 4436 81574 4438 81626
rect 4276 81572 4300 81574
rect 4356 81572 4380 81574
rect 4436 81572 4460 81574
rect 4220 81552 4516 81572
rect 4220 80540 4516 80560
rect 4276 80538 4300 80540
rect 4356 80538 4380 80540
rect 4436 80538 4460 80540
rect 4298 80486 4300 80538
rect 4362 80486 4374 80538
rect 4436 80486 4438 80538
rect 4276 80484 4300 80486
rect 4356 80484 4380 80486
rect 4436 80484 4460 80486
rect 4220 80464 4516 80484
rect 4220 79452 4516 79472
rect 4276 79450 4300 79452
rect 4356 79450 4380 79452
rect 4436 79450 4460 79452
rect 4298 79398 4300 79450
rect 4362 79398 4374 79450
rect 4436 79398 4438 79450
rect 4276 79396 4300 79398
rect 4356 79396 4380 79398
rect 4436 79396 4460 79398
rect 4220 79376 4516 79396
rect 4220 78364 4516 78384
rect 4276 78362 4300 78364
rect 4356 78362 4380 78364
rect 4436 78362 4460 78364
rect 4298 78310 4300 78362
rect 4362 78310 4374 78362
rect 4436 78310 4438 78362
rect 4276 78308 4300 78310
rect 4356 78308 4380 78310
rect 4436 78308 4460 78310
rect 4220 78288 4516 78308
rect 4220 77276 4516 77296
rect 4276 77274 4300 77276
rect 4356 77274 4380 77276
rect 4436 77274 4460 77276
rect 4298 77222 4300 77274
rect 4362 77222 4374 77274
rect 4436 77222 4438 77274
rect 4276 77220 4300 77222
rect 4356 77220 4380 77222
rect 4436 77220 4460 77222
rect 4220 77200 4516 77220
rect 4220 76188 4516 76208
rect 4276 76186 4300 76188
rect 4356 76186 4380 76188
rect 4436 76186 4460 76188
rect 4298 76134 4300 76186
rect 4362 76134 4374 76186
rect 4436 76134 4438 76186
rect 4276 76132 4300 76134
rect 4356 76132 4380 76134
rect 4436 76132 4460 76134
rect 4220 76112 4516 76132
rect 4220 75100 4516 75120
rect 4276 75098 4300 75100
rect 4356 75098 4380 75100
rect 4436 75098 4460 75100
rect 4298 75046 4300 75098
rect 4362 75046 4374 75098
rect 4436 75046 4438 75098
rect 4276 75044 4300 75046
rect 4356 75044 4380 75046
rect 4436 75044 4460 75046
rect 4220 75024 4516 75044
rect 4220 74012 4516 74032
rect 4276 74010 4300 74012
rect 4356 74010 4380 74012
rect 4436 74010 4460 74012
rect 4298 73958 4300 74010
rect 4362 73958 4374 74010
rect 4436 73958 4438 74010
rect 4276 73956 4300 73958
rect 4356 73956 4380 73958
rect 4436 73956 4460 73958
rect 4220 73936 4516 73956
rect 4220 72924 4516 72944
rect 4276 72922 4300 72924
rect 4356 72922 4380 72924
rect 4436 72922 4460 72924
rect 4298 72870 4300 72922
rect 4362 72870 4374 72922
rect 4436 72870 4438 72922
rect 4276 72868 4300 72870
rect 4356 72868 4380 72870
rect 4436 72868 4460 72870
rect 4220 72848 4516 72868
rect 4220 71836 4516 71856
rect 4276 71834 4300 71836
rect 4356 71834 4380 71836
rect 4436 71834 4460 71836
rect 4298 71782 4300 71834
rect 4362 71782 4374 71834
rect 4436 71782 4438 71834
rect 4276 71780 4300 71782
rect 4356 71780 4380 71782
rect 4436 71780 4460 71782
rect 4220 71760 4516 71780
rect 4220 70748 4516 70768
rect 4276 70746 4300 70748
rect 4356 70746 4380 70748
rect 4436 70746 4460 70748
rect 4298 70694 4300 70746
rect 4362 70694 4374 70746
rect 4436 70694 4438 70746
rect 4276 70692 4300 70694
rect 4356 70692 4380 70694
rect 4436 70692 4460 70694
rect 4220 70672 4516 70692
rect 4220 69660 4516 69680
rect 4276 69658 4300 69660
rect 4356 69658 4380 69660
rect 4436 69658 4460 69660
rect 4298 69606 4300 69658
rect 4362 69606 4374 69658
rect 4436 69606 4438 69658
rect 4276 69604 4300 69606
rect 4356 69604 4380 69606
rect 4436 69604 4460 69606
rect 4220 69584 4516 69604
rect 4220 68572 4516 68592
rect 4276 68570 4300 68572
rect 4356 68570 4380 68572
rect 4436 68570 4460 68572
rect 4298 68518 4300 68570
rect 4362 68518 4374 68570
rect 4436 68518 4438 68570
rect 4276 68516 4300 68518
rect 4356 68516 4380 68518
rect 4436 68516 4460 68518
rect 4220 68496 4516 68516
rect 4220 67484 4516 67504
rect 4276 67482 4300 67484
rect 4356 67482 4380 67484
rect 4436 67482 4460 67484
rect 4298 67430 4300 67482
rect 4362 67430 4374 67482
rect 4436 67430 4438 67482
rect 4276 67428 4300 67430
rect 4356 67428 4380 67430
rect 4436 67428 4460 67430
rect 4220 67408 4516 67428
rect 4220 66396 4516 66416
rect 4276 66394 4300 66396
rect 4356 66394 4380 66396
rect 4436 66394 4460 66396
rect 4298 66342 4300 66394
rect 4362 66342 4374 66394
rect 4436 66342 4438 66394
rect 4276 66340 4300 66342
rect 4356 66340 4380 66342
rect 4436 66340 4460 66342
rect 4220 66320 4516 66340
rect 4220 65308 4516 65328
rect 4276 65306 4300 65308
rect 4356 65306 4380 65308
rect 4436 65306 4460 65308
rect 4298 65254 4300 65306
rect 4362 65254 4374 65306
rect 4436 65254 4438 65306
rect 4276 65252 4300 65254
rect 4356 65252 4380 65254
rect 4436 65252 4460 65254
rect 4220 65232 4516 65252
rect 4220 64220 4516 64240
rect 4276 64218 4300 64220
rect 4356 64218 4380 64220
rect 4436 64218 4460 64220
rect 4298 64166 4300 64218
rect 4362 64166 4374 64218
rect 4436 64166 4438 64218
rect 4276 64164 4300 64166
rect 4356 64164 4380 64166
rect 4436 64164 4460 64166
rect 4220 64144 4516 64164
rect 4220 63132 4516 63152
rect 4276 63130 4300 63132
rect 4356 63130 4380 63132
rect 4436 63130 4460 63132
rect 4298 63078 4300 63130
rect 4362 63078 4374 63130
rect 4436 63078 4438 63130
rect 4276 63076 4300 63078
rect 4356 63076 4380 63078
rect 4436 63076 4460 63078
rect 4220 63056 4516 63076
rect 3700 62144 3752 62150
rect 3700 62086 3752 62092
rect 4220 62044 4516 62064
rect 4276 62042 4300 62044
rect 4356 62042 4380 62044
rect 4436 62042 4460 62044
rect 4298 61990 4300 62042
rect 4362 61990 4374 62042
rect 4436 61990 4438 62042
rect 4276 61988 4300 61990
rect 4356 61988 4380 61990
rect 4436 61988 4460 61990
rect 4220 61968 4516 61988
rect 4220 60956 4516 60976
rect 4276 60954 4300 60956
rect 4356 60954 4380 60956
rect 4436 60954 4460 60956
rect 4298 60902 4300 60954
rect 4362 60902 4374 60954
rect 4436 60902 4438 60954
rect 4276 60900 4300 60902
rect 4356 60900 4380 60902
rect 4436 60900 4460 60902
rect 4220 60880 4516 60900
rect 4220 59868 4516 59888
rect 4276 59866 4300 59868
rect 4356 59866 4380 59868
rect 4436 59866 4460 59868
rect 4298 59814 4300 59866
rect 4362 59814 4374 59866
rect 4436 59814 4438 59866
rect 4276 59812 4300 59814
rect 4356 59812 4380 59814
rect 4436 59812 4460 59814
rect 4220 59792 4516 59812
rect 4220 58780 4516 58800
rect 4276 58778 4300 58780
rect 4356 58778 4380 58780
rect 4436 58778 4460 58780
rect 4298 58726 4300 58778
rect 4362 58726 4374 58778
rect 4436 58726 4438 58778
rect 4276 58724 4300 58726
rect 4356 58724 4380 58726
rect 4436 58724 4460 58726
rect 4220 58704 4516 58724
rect 4220 57692 4516 57712
rect 4276 57690 4300 57692
rect 4356 57690 4380 57692
rect 4436 57690 4460 57692
rect 4298 57638 4300 57690
rect 4362 57638 4374 57690
rect 4436 57638 4438 57690
rect 4276 57636 4300 57638
rect 4356 57636 4380 57638
rect 4436 57636 4460 57638
rect 4220 57616 4516 57636
rect 4220 56604 4516 56624
rect 4276 56602 4300 56604
rect 4356 56602 4380 56604
rect 4436 56602 4460 56604
rect 4298 56550 4300 56602
rect 4362 56550 4374 56602
rect 4436 56550 4438 56602
rect 4276 56548 4300 56550
rect 4356 56548 4380 56550
rect 4436 56548 4460 56550
rect 4220 56528 4516 56548
rect 4220 55516 4516 55536
rect 4276 55514 4300 55516
rect 4356 55514 4380 55516
rect 4436 55514 4460 55516
rect 4298 55462 4300 55514
rect 4362 55462 4374 55514
rect 4436 55462 4438 55514
rect 4276 55460 4300 55462
rect 4356 55460 4380 55462
rect 4436 55460 4460 55462
rect 4220 55440 4516 55460
rect 4220 54428 4516 54448
rect 4276 54426 4300 54428
rect 4356 54426 4380 54428
rect 4436 54426 4460 54428
rect 4298 54374 4300 54426
rect 4362 54374 4374 54426
rect 4436 54374 4438 54426
rect 4276 54372 4300 54374
rect 4356 54372 4380 54374
rect 4436 54372 4460 54374
rect 4220 54352 4516 54372
rect 4220 53340 4516 53360
rect 4276 53338 4300 53340
rect 4356 53338 4380 53340
rect 4436 53338 4460 53340
rect 4298 53286 4300 53338
rect 4362 53286 4374 53338
rect 4436 53286 4438 53338
rect 4276 53284 4300 53286
rect 4356 53284 4380 53286
rect 4436 53284 4460 53286
rect 4220 53264 4516 53284
rect 4220 52252 4516 52272
rect 4276 52250 4300 52252
rect 4356 52250 4380 52252
rect 4436 52250 4460 52252
rect 4298 52198 4300 52250
rect 4362 52198 4374 52250
rect 4436 52198 4438 52250
rect 4276 52196 4300 52198
rect 4356 52196 4380 52198
rect 4436 52196 4460 52198
rect 4220 52176 4516 52196
rect 4220 51164 4516 51184
rect 4276 51162 4300 51164
rect 4356 51162 4380 51164
rect 4436 51162 4460 51164
rect 4298 51110 4300 51162
rect 4362 51110 4374 51162
rect 4436 51110 4438 51162
rect 4276 51108 4300 51110
rect 4356 51108 4380 51110
rect 4436 51108 4460 51110
rect 4220 51088 4516 51108
rect 3608 50380 3660 50386
rect 3608 50322 3660 50328
rect 4220 50076 4516 50096
rect 4276 50074 4300 50076
rect 4356 50074 4380 50076
rect 4436 50074 4460 50076
rect 4298 50022 4300 50074
rect 4362 50022 4374 50074
rect 4436 50022 4438 50074
rect 4276 50020 4300 50022
rect 4356 50020 4380 50022
rect 4436 50020 4460 50022
rect 4220 50000 4516 50020
rect 4220 48988 4516 49008
rect 4276 48986 4300 48988
rect 4356 48986 4380 48988
rect 4436 48986 4460 48988
rect 4298 48934 4300 48986
rect 4362 48934 4374 48986
rect 4436 48934 4438 48986
rect 4276 48932 4300 48934
rect 4356 48932 4380 48934
rect 4436 48932 4460 48934
rect 4220 48912 4516 48932
rect 4220 47900 4516 47920
rect 4276 47898 4300 47900
rect 4356 47898 4380 47900
rect 4436 47898 4460 47900
rect 4298 47846 4300 47898
rect 4362 47846 4374 47898
rect 4436 47846 4438 47898
rect 4276 47844 4300 47846
rect 4356 47844 4380 47846
rect 4436 47844 4460 47846
rect 4220 47824 4516 47844
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4220 45648 4516 45668
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 4068 37732 4120 37738
rect 4068 37674 4120 37680
rect 4080 36310 4108 37674
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4068 36304 4120 36310
rect 4068 36246 4120 36252
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4068 29028 4120 29034
rect 4068 28970 4120 28976
rect 4080 26586 4108 28970
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4068 26580 4120 26586
rect 4068 26522 4120 26528
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4356 4690 4384 5034
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3620 4078 3648 4422
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4632 4078 4660 4762
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 2872 2576 2924 2582
rect 2872 2518 2924 2524
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2792 1873 2820 2450
rect 2778 1864 2834 1873
rect 2778 1799 2834 1808
rect 110 -800 166 800
rect 386 -800 442 800
rect 754 -800 810 800
rect 1030 -800 1086 800
rect 1398 -800 1454 800
rect 1674 -800 1730 800
rect 2042 -800 2098 800
rect 2318 -800 2374 800
rect 2686 -800 2742 800
rect 2884 377 2912 2518
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 2976 800 3004 2450
rect 3344 800 3372 3538
rect 3620 800 3648 3878
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3988 800 4016 3470
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4252 2032 4304 2038
rect 4252 1974 4304 1980
rect 4264 800 4292 1974
rect 4632 800 4660 2926
rect 4724 2038 4752 4014
rect 4816 3058 4844 92754
rect 4908 16574 4936 98194
rect 4908 16546 5028 16574
rect 5000 12434 5028 16546
rect 4908 12406 5028 12434
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4908 2650 4936 12406
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5000 3602 5028 11834
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 4712 2032 4764 2038
rect 4712 1974 4764 1980
rect 5000 800 5028 3334
rect 5092 2378 5120 99282
rect 5264 96076 5316 96082
rect 5264 96018 5316 96024
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5184 7426 5212 7686
rect 5276 7562 5304 96018
rect 6184 95464 6236 95470
rect 6184 95406 6236 95412
rect 5356 94376 5408 94382
rect 5356 94318 5408 94324
rect 5368 7750 5396 94318
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5276 7534 5488 7562
rect 5184 7398 5396 7426
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5184 3126 5212 4626
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 5080 2372 5132 2378
rect 5080 2314 5132 2320
rect 5276 800 5304 4014
rect 5368 2582 5396 7398
rect 5356 2576 5408 2582
rect 5356 2518 5408 2524
rect 5460 2446 5488 7534
rect 6196 3058 6224 95406
rect 6276 70508 6328 70514
rect 6276 70450 6328 70456
rect 6288 5846 6316 70450
rect 6368 69964 6420 69970
rect 6368 69906 6420 69912
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6380 5710 6408 69906
rect 6460 56160 6512 56166
rect 6460 56102 6512 56108
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5644 800 5672 2450
rect 5920 800 5948 2926
rect 6288 800 6316 3334
rect 6472 2310 6500 56102
rect 6644 48612 6696 48618
rect 6644 48554 6696 48560
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6564 800 6592 4014
rect 6656 3670 6684 48554
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 3670 6960 4966
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 6932 800 6960 2450
rect 7024 2310 7052 103022
rect 7760 102746 7788 115398
rect 7944 115258 7972 116010
rect 8036 115802 8064 116198
rect 8024 115796 8076 115802
rect 8024 115738 8076 115744
rect 7932 115252 7984 115258
rect 7932 115194 7984 115200
rect 8220 113558 8248 119200
rect 8404 116890 8432 119200
rect 8392 116884 8444 116890
rect 8392 116826 8444 116832
rect 8392 116748 8444 116754
rect 8392 116690 8444 116696
rect 8404 115734 8432 116690
rect 8680 116346 8708 119200
rect 8668 116340 8720 116346
rect 8668 116282 8720 116288
rect 8392 115728 8444 115734
rect 8392 115670 8444 115676
rect 8300 115660 8352 115666
rect 8300 115602 8352 115608
rect 8312 115258 8340 115602
rect 8484 115592 8536 115598
rect 8484 115534 8536 115540
rect 8300 115252 8352 115258
rect 8300 115194 8352 115200
rect 8300 114708 8352 114714
rect 8300 114650 8352 114656
rect 8312 113898 8340 114650
rect 8300 113892 8352 113898
rect 8300 113834 8352 113840
rect 8208 113552 8260 113558
rect 8208 113494 8260 113500
rect 8496 108730 8524 115534
rect 8760 115116 8812 115122
rect 8760 115058 8812 115064
rect 8668 115048 8720 115054
rect 8668 114990 8720 114996
rect 8484 108724 8536 108730
rect 8484 108666 8536 108672
rect 8680 106010 8708 114990
rect 8772 114578 8800 115058
rect 8864 114578 8892 119200
rect 9140 117298 9168 119200
rect 9128 117292 9180 117298
rect 9128 117234 9180 117240
rect 9324 116890 9352 119200
rect 9312 116884 9364 116890
rect 9312 116826 9364 116832
rect 9128 116748 9180 116754
rect 9128 116690 9180 116696
rect 9140 115802 9168 116690
rect 9600 116498 9628 119200
rect 9784 117230 9812 119200
rect 9772 117224 9824 117230
rect 9772 117166 9824 117172
rect 9680 117156 9732 117162
rect 9680 117098 9732 117104
rect 9508 116470 9628 116498
rect 9128 115796 9180 115802
rect 9128 115738 9180 115744
rect 9508 114578 9536 116470
rect 9588 116068 9640 116074
rect 9588 116010 9640 116016
rect 8760 114572 8812 114578
rect 8760 114514 8812 114520
rect 8852 114572 8904 114578
rect 8852 114514 8904 114520
rect 9496 114572 9548 114578
rect 9496 114514 9548 114520
rect 8668 106004 8720 106010
rect 8668 105946 8720 105952
rect 7748 102740 7800 102746
rect 7748 102682 7800 102688
rect 7564 102604 7616 102610
rect 7564 102546 7616 102552
rect 7380 54052 7432 54058
rect 7380 53994 7432 54000
rect 7392 3194 7420 53994
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7576 3126 7604 102546
rect 8392 97640 8444 97646
rect 8392 97582 8444 97588
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 7840 3596 7892 3602
rect 7840 3538 7892 3544
rect 7564 3120 7616 3126
rect 7564 3062 7616 3068
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7208 800 7236 2926
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7576 800 7604 2790
rect 7852 800 7880 3538
rect 8036 2990 8064 6122
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 8404 2582 8432 97582
rect 9036 75812 9088 75818
rect 9036 75754 9088 75760
rect 8944 72140 8996 72146
rect 8944 72082 8996 72088
rect 8956 10810 8984 72082
rect 9048 23866 9076 75754
rect 9128 40044 9180 40050
rect 9128 39986 9180 39992
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 9140 19242 9168 39986
rect 9600 26926 9628 116010
rect 9692 115666 9720 117098
rect 10060 116890 10088 119200
rect 10048 116884 10100 116890
rect 10048 116826 10100 116832
rect 9864 116748 9916 116754
rect 9864 116690 9916 116696
rect 9680 115660 9732 115666
rect 9680 115602 9732 115608
rect 9876 115258 9904 116690
rect 9864 115252 9916 115258
rect 9864 115194 9916 115200
rect 10244 114578 10272 119200
rect 10520 117298 10548 119200
rect 10508 117292 10560 117298
rect 10508 117234 10560 117240
rect 10416 117156 10468 117162
rect 10416 117098 10468 117104
rect 10428 115666 10456 117098
rect 10600 116748 10652 116754
rect 10600 116690 10652 116696
rect 10416 115660 10468 115666
rect 10416 115602 10468 115608
rect 10612 115258 10640 116690
rect 10704 116346 10732 119200
rect 10692 116340 10744 116346
rect 10692 116282 10744 116288
rect 10784 116068 10836 116074
rect 10784 116010 10836 116016
rect 10796 115258 10824 116010
rect 10600 115252 10652 115258
rect 10600 115194 10652 115200
rect 10784 115252 10836 115258
rect 10784 115194 10836 115200
rect 10980 115054 11008 119200
rect 11164 117434 11192 119200
rect 11152 117428 11204 117434
rect 11152 117370 11204 117376
rect 11152 117156 11204 117162
rect 11152 117098 11204 117104
rect 11164 115666 11192 117098
rect 11440 116890 11468 119200
rect 11624 117314 11652 119200
rect 11624 117286 11744 117314
rect 11900 117298 11928 119200
rect 11612 117156 11664 117162
rect 11612 117098 11664 117104
rect 11428 116884 11480 116890
rect 11428 116826 11480 116832
rect 11624 116346 11652 117098
rect 11612 116340 11664 116346
rect 11612 116282 11664 116288
rect 11152 115660 11204 115666
rect 11152 115602 11204 115608
rect 10968 115048 11020 115054
rect 10968 114990 11020 114996
rect 10692 114912 10744 114918
rect 10692 114854 10744 114860
rect 10232 114572 10284 114578
rect 10232 114514 10284 114520
rect 10704 114442 10732 114854
rect 11716 114578 11744 117286
rect 11888 117292 11940 117298
rect 11888 117234 11940 117240
rect 12084 116822 12112 119200
rect 12072 116816 12124 116822
rect 12072 116758 12124 116764
rect 12164 116748 12216 116754
rect 12164 116690 12216 116696
rect 12176 115666 12204 116690
rect 12164 115660 12216 115666
rect 12164 115602 12216 115608
rect 12360 114578 12388 119200
rect 12544 117094 12572 119200
rect 12532 117088 12584 117094
rect 12532 117030 12584 117036
rect 12820 116890 12848 119200
rect 13004 117314 13032 119200
rect 13280 117314 13308 119200
rect 13004 117286 13216 117314
rect 13280 117298 13400 117314
rect 13280 117292 13412 117298
rect 13280 117286 13360 117292
rect 13084 117156 13136 117162
rect 13084 117098 13136 117104
rect 12808 116884 12860 116890
rect 12808 116826 12860 116832
rect 12900 116748 12952 116754
rect 12900 116690 12952 116696
rect 12992 116748 13044 116754
rect 12992 116690 13044 116696
rect 12912 115666 12940 116690
rect 12900 115660 12952 115666
rect 12900 115602 12952 115608
rect 13004 115258 13032 116690
rect 13096 116346 13124 117098
rect 13084 116340 13136 116346
rect 13084 116282 13136 116288
rect 12992 115252 13044 115258
rect 12992 115194 13044 115200
rect 13188 114578 13216 117286
rect 13360 117234 13412 117240
rect 13464 116822 13492 119200
rect 13452 116816 13504 116822
rect 13452 116758 13504 116764
rect 13360 114980 13412 114986
rect 13360 114922 13412 114928
rect 13372 114714 13400 114922
rect 13360 114708 13412 114714
rect 13360 114650 13412 114656
rect 13740 114578 13768 119200
rect 13924 117230 13952 119200
rect 13912 117224 13964 117230
rect 13912 117166 13964 117172
rect 13820 117156 13872 117162
rect 13820 117098 13872 117104
rect 14004 117156 14056 117162
rect 14004 117098 14056 117104
rect 13832 116278 13860 117098
rect 14016 116346 14044 117098
rect 14200 116890 14228 119200
rect 14188 116884 14240 116890
rect 14384 116872 14412 119200
rect 14660 117094 14688 119200
rect 14648 117088 14700 117094
rect 14648 117030 14700 117036
rect 14384 116844 14504 116872
rect 14188 116826 14240 116832
rect 14372 116748 14424 116754
rect 14372 116690 14424 116696
rect 14004 116340 14056 116346
rect 14004 116282 14056 116288
rect 13820 116272 13872 116278
rect 13820 116214 13872 116220
rect 14384 115258 14412 116690
rect 14372 115252 14424 115258
rect 14372 115194 14424 115200
rect 14476 114578 14504 116844
rect 14844 116346 14872 119200
rect 15120 116872 15148 119200
rect 15200 117156 15252 117162
rect 15200 117098 15252 117104
rect 15028 116844 15148 116872
rect 14832 116340 14884 116346
rect 14832 116282 14884 116288
rect 14924 116068 14976 116074
rect 14924 116010 14976 116016
rect 14936 115258 14964 116010
rect 14924 115252 14976 115258
rect 14924 115194 14976 115200
rect 15028 114578 15056 116844
rect 15108 116748 15160 116754
rect 15108 116690 15160 116696
rect 15120 115666 15148 116690
rect 15108 115660 15160 115666
rect 15108 115602 15160 115608
rect 15212 115598 15240 117098
rect 15304 116142 15332 119200
rect 15580 116890 15608 119200
rect 15568 116884 15620 116890
rect 15568 116826 15620 116832
rect 15292 116136 15344 116142
rect 15292 116078 15344 116084
rect 15200 115592 15252 115598
rect 15200 115534 15252 115540
rect 15292 115116 15344 115122
rect 15292 115058 15344 115064
rect 15304 114714 15332 115058
rect 15292 114708 15344 114714
rect 15292 114650 15344 114656
rect 15764 114578 15792 119200
rect 15844 116748 15896 116754
rect 15844 116690 15896 116696
rect 15856 115258 15884 116690
rect 16040 115682 16068 119200
rect 16316 117366 16344 119200
rect 16500 117450 16528 119200
rect 16408 117422 16528 117450
rect 16304 117360 16356 117366
rect 16304 117302 16356 117308
rect 16212 117156 16264 117162
rect 16212 117098 16264 117104
rect 16040 115654 16160 115682
rect 16132 115598 16160 115654
rect 16120 115592 16172 115598
rect 16120 115534 16172 115540
rect 16224 115530 16252 117098
rect 16408 116226 16436 117422
rect 16776 117366 16804 119200
rect 16488 117360 16540 117366
rect 16764 117360 16816 117366
rect 16540 117308 16620 117314
rect 16488 117302 16620 117308
rect 16764 117302 16816 117308
rect 16500 117286 16620 117302
rect 16592 116278 16620 117286
rect 16960 116890 16988 119200
rect 17040 117088 17092 117094
rect 17040 117030 17092 117036
rect 16948 116884 17000 116890
rect 16948 116826 17000 116832
rect 16580 116272 16632 116278
rect 16408 116198 16528 116226
rect 16580 116214 16632 116220
rect 16396 116068 16448 116074
rect 16396 116010 16448 116016
rect 16212 115524 16264 115530
rect 16212 115466 16264 115472
rect 16408 115258 16436 116010
rect 15844 115252 15896 115258
rect 15844 115194 15896 115200
rect 16396 115252 16448 115258
rect 16396 115194 16448 115200
rect 16500 115054 16528 116198
rect 17052 116142 17080 117030
rect 17040 116136 17092 116142
rect 17040 116078 17092 116084
rect 17236 115054 17264 119200
rect 17420 117434 17448 119200
rect 17408 117428 17460 117434
rect 17408 117370 17460 117376
rect 17696 117314 17724 119200
rect 17592 117292 17644 117298
rect 17696 117286 17816 117314
rect 17592 117234 17644 117240
rect 17316 117224 17368 117230
rect 17316 117166 17368 117172
rect 17328 115666 17356 117166
rect 17408 116748 17460 116754
rect 17408 116690 17460 116696
rect 17420 115666 17448 116690
rect 17316 115660 17368 115666
rect 17316 115602 17368 115608
rect 17408 115660 17460 115666
rect 17408 115602 17460 115608
rect 17604 115598 17632 117234
rect 17684 117156 17736 117162
rect 17684 117098 17736 117104
rect 17696 116346 17724 117098
rect 17788 116890 17816 117286
rect 17776 116884 17828 116890
rect 17776 116826 17828 116832
rect 17684 116340 17736 116346
rect 17684 116282 17736 116288
rect 17592 115592 17644 115598
rect 17592 115534 17644 115540
rect 17776 115524 17828 115530
rect 17776 115466 17828 115472
rect 16488 115048 16540 115054
rect 16488 114990 16540 114996
rect 17224 115048 17276 115054
rect 17224 114990 17276 114996
rect 17788 114714 17816 115466
rect 17776 114708 17828 114714
rect 17776 114650 17828 114656
rect 17880 114578 17908 119200
rect 18156 117434 18184 119200
rect 17960 117428 18012 117434
rect 17960 117370 18012 117376
rect 18144 117428 18196 117434
rect 18144 117370 18196 117376
rect 17972 117094 18000 117370
rect 17960 117088 18012 117094
rect 17960 117030 18012 117036
rect 18340 116890 18368 119200
rect 18328 116884 18380 116890
rect 18328 116826 18380 116832
rect 18144 116748 18196 116754
rect 18144 116690 18196 116696
rect 18156 115666 18184 116690
rect 18144 115660 18196 115666
rect 18144 115602 18196 115608
rect 18616 115054 18644 119200
rect 18800 116686 18828 119200
rect 19076 116890 19104 119200
rect 19156 117156 19208 117162
rect 19156 117098 19208 117104
rect 19064 116884 19116 116890
rect 19064 116826 19116 116832
rect 18880 116748 18932 116754
rect 18880 116690 18932 116696
rect 18788 116680 18840 116686
rect 18788 116622 18840 116628
rect 18892 115258 18920 116690
rect 19168 116278 19196 117098
rect 19156 116272 19208 116278
rect 19156 116214 19208 116220
rect 18880 115252 18932 115258
rect 18880 115194 18932 115200
rect 18604 115048 18656 115054
rect 18604 114990 18656 114996
rect 19260 114578 19288 119200
rect 19536 117366 19564 119200
rect 19524 117360 19576 117366
rect 19524 117302 19576 117308
rect 19720 117178 19748 119200
rect 19340 117156 19392 117162
rect 19720 117150 19932 117178
rect 19340 117098 19392 117104
rect 19352 116346 19380 117098
rect 19580 116988 19876 117008
rect 19636 116986 19660 116988
rect 19716 116986 19740 116988
rect 19796 116986 19820 116988
rect 19658 116934 19660 116986
rect 19722 116934 19734 116986
rect 19796 116934 19798 116986
rect 19636 116932 19660 116934
rect 19716 116932 19740 116934
rect 19796 116932 19820 116934
rect 19580 116912 19876 116932
rect 19904 116822 19932 117150
rect 19892 116816 19944 116822
rect 19892 116758 19944 116764
rect 19432 116748 19484 116754
rect 19432 116690 19484 116696
rect 19340 116340 19392 116346
rect 19340 116282 19392 116288
rect 19444 115666 19472 116690
rect 19580 115900 19876 115920
rect 19636 115898 19660 115900
rect 19716 115898 19740 115900
rect 19796 115898 19820 115900
rect 19658 115846 19660 115898
rect 19722 115846 19734 115898
rect 19796 115846 19798 115898
rect 19636 115844 19660 115846
rect 19716 115844 19740 115846
rect 19796 115844 19820 115846
rect 19580 115824 19876 115844
rect 19432 115660 19484 115666
rect 19432 115602 19484 115608
rect 19580 114812 19876 114832
rect 19636 114810 19660 114812
rect 19716 114810 19740 114812
rect 19796 114810 19820 114812
rect 19658 114758 19660 114810
rect 19722 114758 19734 114810
rect 19796 114758 19798 114810
rect 19636 114756 19660 114758
rect 19716 114756 19740 114758
rect 19796 114756 19820 114758
rect 19580 114736 19876 114756
rect 19996 114578 20024 119200
rect 20180 117314 20208 119200
rect 20180 117286 20300 117314
rect 20272 116618 20300 117286
rect 20456 116890 20484 119200
rect 20536 117156 20588 117162
rect 20536 117098 20588 117104
rect 20444 116884 20496 116890
rect 20444 116826 20496 116832
rect 20352 116748 20404 116754
rect 20352 116690 20404 116696
rect 20444 116748 20496 116754
rect 20444 116690 20496 116696
rect 20260 116612 20312 116618
rect 20260 116554 20312 116560
rect 20364 115258 20392 116690
rect 20456 115598 20484 116690
rect 20548 116210 20576 117098
rect 20536 116204 20588 116210
rect 20536 116146 20588 116152
rect 20444 115592 20496 115598
rect 20444 115534 20496 115540
rect 20352 115252 20404 115258
rect 20352 115194 20404 115200
rect 20640 115054 20668 119200
rect 20916 117434 20944 119200
rect 20904 117428 20956 117434
rect 20904 117370 20956 117376
rect 21100 116872 21128 119200
rect 21272 117156 21324 117162
rect 21272 117098 21324 117104
rect 21100 116844 21220 116872
rect 21088 116748 21140 116754
rect 21088 116690 21140 116696
rect 20720 116544 20772 116550
rect 20720 116486 20772 116492
rect 20732 115666 20760 116486
rect 20720 115660 20772 115666
rect 20720 115602 20772 115608
rect 20996 115456 21048 115462
rect 20996 115398 21048 115404
rect 20628 115048 20680 115054
rect 20628 114990 20680 114996
rect 21008 114578 21036 115398
rect 21100 115258 21128 116690
rect 21192 116346 21220 116844
rect 21284 116822 21312 117098
rect 21272 116816 21324 116822
rect 21272 116758 21324 116764
rect 21180 116340 21232 116346
rect 21180 116282 21232 116288
rect 21180 116068 21232 116074
rect 21180 116010 21232 116016
rect 21192 115666 21220 116010
rect 21376 115734 21404 119200
rect 21560 116278 21588 119200
rect 21836 116890 21864 119200
rect 21916 117088 21968 117094
rect 21916 117030 21968 117036
rect 21824 116884 21876 116890
rect 21824 116826 21876 116832
rect 21928 116686 21956 117030
rect 21916 116680 21968 116686
rect 21916 116622 21968 116628
rect 21548 116272 21600 116278
rect 21548 116214 21600 116220
rect 21364 115728 21416 115734
rect 21364 115670 21416 115676
rect 21916 115728 21968 115734
rect 21916 115670 21968 115676
rect 21180 115660 21232 115666
rect 21180 115602 21232 115608
rect 21088 115252 21140 115258
rect 21088 115194 21140 115200
rect 21456 115184 21508 115190
rect 21454 115152 21456 115161
rect 21508 115152 21510 115161
rect 21454 115087 21510 115096
rect 21824 115116 21876 115122
rect 21824 115058 21876 115064
rect 21088 114912 21140 114918
rect 21088 114854 21140 114860
rect 21100 114578 21128 114854
rect 21836 114714 21864 115058
rect 21928 115054 21956 115670
rect 21916 115048 21968 115054
rect 21916 114990 21968 114996
rect 21824 114708 21876 114714
rect 21824 114650 21876 114656
rect 11704 114572 11756 114578
rect 11704 114514 11756 114520
rect 12348 114572 12400 114578
rect 12348 114514 12400 114520
rect 13176 114572 13228 114578
rect 13176 114514 13228 114520
rect 13728 114572 13780 114578
rect 13728 114514 13780 114520
rect 14464 114572 14516 114578
rect 14464 114514 14516 114520
rect 15016 114572 15068 114578
rect 15016 114514 15068 114520
rect 15752 114572 15804 114578
rect 15752 114514 15804 114520
rect 17868 114572 17920 114578
rect 17868 114514 17920 114520
rect 19248 114572 19300 114578
rect 19248 114514 19300 114520
rect 19984 114572 20036 114578
rect 19984 114514 20036 114520
rect 20996 114572 21048 114578
rect 20996 114514 21048 114520
rect 21088 114572 21140 114578
rect 21088 114514 21140 114520
rect 10692 114436 10744 114442
rect 10692 114378 10744 114384
rect 12716 114368 12768 114374
rect 12716 114310 12768 114316
rect 14648 114368 14700 114374
rect 14648 114310 14700 114316
rect 12728 114034 12756 114310
rect 12716 114028 12768 114034
rect 12716 113970 12768 113976
rect 14660 113966 14688 114310
rect 22020 113966 22048 119200
rect 22296 117366 22324 119200
rect 22284 117360 22336 117366
rect 22284 117302 22336 117308
rect 22480 116822 22508 119200
rect 22468 116816 22520 116822
rect 22468 116758 22520 116764
rect 22652 116748 22704 116754
rect 22652 116690 22704 116696
rect 22376 116680 22428 116686
rect 22376 116622 22428 116628
rect 22388 115598 22416 116622
rect 22664 116385 22692 116690
rect 22650 116376 22706 116385
rect 22650 116311 22706 116320
rect 22466 116240 22522 116249
rect 22466 116175 22468 116184
rect 22520 116175 22522 116184
rect 22468 116146 22520 116152
rect 22376 115592 22428 115598
rect 22376 115534 22428 115540
rect 22756 115172 22784 119200
rect 22940 117434 22968 119200
rect 22928 117428 22980 117434
rect 22928 117370 22980 117376
rect 22928 117224 22980 117230
rect 23216 117178 23244 119200
rect 22928 117166 22980 117172
rect 22940 116278 22968 117166
rect 23020 117156 23072 117162
rect 23020 117098 23072 117104
rect 23124 117150 23244 117178
rect 23296 117156 23348 117162
rect 23032 116346 23060 117098
rect 23124 116890 23152 117150
rect 23296 117098 23348 117104
rect 23204 117088 23256 117094
rect 23204 117030 23256 117036
rect 23112 116884 23164 116890
rect 23112 116826 23164 116832
rect 23110 116784 23166 116793
rect 23110 116719 23166 116728
rect 23020 116340 23072 116346
rect 23020 116282 23072 116288
rect 22928 116272 22980 116278
rect 22928 116214 22980 116220
rect 22756 115144 22968 115172
rect 22468 115048 22520 115054
rect 22468 114990 22520 114996
rect 22480 114578 22508 114990
rect 22836 114980 22888 114986
rect 22836 114922 22888 114928
rect 22848 114578 22876 114922
rect 22940 114578 22968 115144
rect 23018 115152 23074 115161
rect 23018 115087 23074 115096
rect 23032 115054 23060 115087
rect 23020 115048 23072 115054
rect 23020 114990 23072 114996
rect 22468 114572 22520 114578
rect 22468 114514 22520 114520
rect 22836 114572 22888 114578
rect 22836 114514 22888 114520
rect 22928 114572 22980 114578
rect 22928 114514 22980 114520
rect 14648 113960 14700 113966
rect 14648 113902 14700 113908
rect 22008 113960 22060 113966
rect 22008 113902 22060 113908
rect 19580 113724 19876 113744
rect 19636 113722 19660 113724
rect 19716 113722 19740 113724
rect 19796 113722 19820 113724
rect 19658 113670 19660 113722
rect 19722 113670 19734 113722
rect 19796 113670 19798 113722
rect 19636 113668 19660 113670
rect 19716 113668 19740 113670
rect 19796 113668 19820 113670
rect 19580 113648 19876 113668
rect 19580 112636 19876 112656
rect 19636 112634 19660 112636
rect 19716 112634 19740 112636
rect 19796 112634 19820 112636
rect 19658 112582 19660 112634
rect 19722 112582 19734 112634
rect 19796 112582 19798 112634
rect 19636 112580 19660 112582
rect 19716 112580 19740 112582
rect 19796 112580 19820 112582
rect 19580 112560 19876 112580
rect 19580 111548 19876 111568
rect 19636 111546 19660 111548
rect 19716 111546 19740 111548
rect 19796 111546 19820 111548
rect 19658 111494 19660 111546
rect 19722 111494 19734 111546
rect 19796 111494 19798 111546
rect 19636 111492 19660 111494
rect 19716 111492 19740 111494
rect 19796 111492 19820 111494
rect 19580 111472 19876 111492
rect 13728 110696 13780 110702
rect 13728 110638 13780 110644
rect 12900 108520 12952 108526
rect 12900 108462 12952 108468
rect 9956 105868 10008 105874
rect 9956 105810 10008 105816
rect 9680 53508 9732 53514
rect 9680 53450 9732 53456
rect 9588 26920 9640 26926
rect 9588 26862 9640 26868
rect 9128 19236 9180 19242
rect 9128 19178 9180 19184
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8956 3670 8984 6190
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 8392 2576 8444 2582
rect 8392 2518 8444 2524
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8220 800 8248 2450
rect 8496 800 8524 3538
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8864 800 8892 3334
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9232 800 9260 2926
rect 9508 800 9536 3538
rect 9692 3194 9720 53450
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9876 800 9904 2790
rect 9968 2582 9996 105810
rect 11428 103012 11480 103018
rect 11428 102954 11480 102960
rect 10508 100904 10560 100910
rect 10508 100846 10560 100852
rect 10324 75404 10376 75410
rect 10324 75346 10376 75352
rect 10336 25294 10364 75346
rect 10324 25288 10376 25294
rect 10324 25230 10376 25236
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10336 2990 10364 12378
rect 10520 3126 10548 100846
rect 11244 53576 11296 53582
rect 11244 53518 11296 53524
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10888 3670 10916 7754
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10324 2984 10376 2990
rect 10324 2926 10376 2932
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10152 800 10180 2450
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10520 800 10548 2382
rect 10796 800 10824 3334
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 11164 800 11192 2926
rect 11256 2650 11284 53518
rect 11440 3058 11468 102954
rect 12348 101924 12400 101930
rect 12348 101866 12400 101872
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11900 4078 11928 13466
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 11428 2916 11480 2922
rect 11428 2858 11480 2864
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11440 800 11468 2858
rect 11808 800 11836 3878
rect 12360 3058 12388 101866
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12452 3398 12480 4422
rect 12636 3670 12664 5578
rect 12820 4078 12848 7686
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 12084 800 12112 2450
rect 12544 1850 12572 2994
rect 12452 1822 12572 1850
rect 12452 800 12480 1822
rect 12728 800 12756 3878
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12820 3058 12848 3538
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 12912 2650 12940 108462
rect 13268 99816 13320 99822
rect 13268 99758 13320 99764
rect 13280 3670 13308 99758
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13372 3058 13400 3334
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13096 800 13124 2926
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 13464 800 13492 2450
rect 13648 1714 13676 3334
rect 13740 2582 13768 110638
rect 19580 110460 19876 110480
rect 19636 110458 19660 110460
rect 19716 110458 19740 110460
rect 19796 110458 19820 110460
rect 19658 110406 19660 110458
rect 19722 110406 19734 110458
rect 19796 110406 19798 110458
rect 19636 110404 19660 110406
rect 19716 110404 19740 110406
rect 19796 110404 19820 110406
rect 19580 110384 19876 110404
rect 19580 109372 19876 109392
rect 19636 109370 19660 109372
rect 19716 109370 19740 109372
rect 19796 109370 19820 109372
rect 19658 109318 19660 109370
rect 19722 109318 19734 109370
rect 19796 109318 19798 109370
rect 19636 109316 19660 109318
rect 19716 109316 19740 109318
rect 19796 109316 19820 109318
rect 19580 109296 19876 109316
rect 23124 109034 23152 116719
rect 23216 116618 23244 117030
rect 23204 116612 23256 116618
rect 23204 116554 23256 116560
rect 23308 116550 23336 117098
rect 23296 116544 23348 116550
rect 23296 116486 23348 116492
rect 23400 113966 23428 119200
rect 23480 116136 23532 116142
rect 23480 116078 23532 116084
rect 23492 115802 23520 116078
rect 23480 115796 23532 115802
rect 23480 115738 23532 115744
rect 23676 115666 23704 119200
rect 23860 116346 23888 119200
rect 23848 116340 23900 116346
rect 23848 116282 23900 116288
rect 23664 115660 23716 115666
rect 23664 115602 23716 115608
rect 23480 115524 23532 115530
rect 23480 115466 23532 115472
rect 23492 114918 23520 115466
rect 24032 115184 24084 115190
rect 24030 115152 24032 115161
rect 24084 115152 24086 115161
rect 24030 115087 24086 115096
rect 23480 114912 23532 114918
rect 23480 114854 23532 114860
rect 23572 114912 23624 114918
rect 23572 114854 23624 114860
rect 23584 114714 23612 114854
rect 24136 114714 24164 119200
rect 24412 117638 24440 119200
rect 24400 117632 24452 117638
rect 24400 117574 24452 117580
rect 24492 117156 24544 117162
rect 24492 117098 24544 117104
rect 24504 116618 24532 117098
rect 24596 116890 24624 119200
rect 24676 117156 24728 117162
rect 24676 117098 24728 117104
rect 24584 116884 24636 116890
rect 24584 116826 24636 116832
rect 24492 116612 24544 116618
rect 24492 116554 24544 116560
rect 24688 116006 24716 117098
rect 24768 116748 24820 116754
rect 24768 116690 24820 116696
rect 24780 116346 24808 116690
rect 24768 116340 24820 116346
rect 24768 116282 24820 116288
rect 24766 116104 24822 116113
rect 24766 116039 24822 116048
rect 24676 116000 24728 116006
rect 24676 115942 24728 115948
rect 24780 115802 24808 116039
rect 24768 115796 24820 115802
rect 24768 115738 24820 115744
rect 24216 115456 24268 115462
rect 24216 115398 24268 115404
rect 24228 115190 24256 115398
rect 24216 115184 24268 115190
rect 24216 115126 24268 115132
rect 24400 115116 24452 115122
rect 24400 115058 24452 115064
rect 24412 115002 24440 115058
rect 24320 114974 24440 115002
rect 24320 114918 24348 114974
rect 24308 114912 24360 114918
rect 24308 114854 24360 114860
rect 24400 114912 24452 114918
rect 24400 114854 24452 114860
rect 23572 114708 23624 114714
rect 23572 114650 23624 114656
rect 24124 114708 24176 114714
rect 24124 114650 24176 114656
rect 24412 114578 24440 114854
rect 24872 114646 24900 119200
rect 25056 117706 25084 119200
rect 25044 117700 25096 117706
rect 25044 117642 25096 117648
rect 24950 117056 25006 117065
rect 24950 116991 25006 117000
rect 24964 115598 24992 116991
rect 25332 116890 25360 119200
rect 25320 116884 25372 116890
rect 25320 116826 25372 116832
rect 25410 116376 25466 116385
rect 25410 116311 25466 116320
rect 25228 115728 25280 115734
rect 25228 115670 25280 115676
rect 24952 115592 25004 115598
rect 24952 115534 25004 115540
rect 25240 115530 25268 115670
rect 25228 115524 25280 115530
rect 25228 115466 25280 115472
rect 25424 115258 25452 116311
rect 25412 115252 25464 115258
rect 25412 115194 25464 115200
rect 25516 114714 25544 119200
rect 25792 117337 25820 119200
rect 25778 117328 25834 117337
rect 25778 117263 25834 117272
rect 25976 116890 26004 119200
rect 25964 116884 26016 116890
rect 25964 116826 26016 116832
rect 25688 116680 25740 116686
rect 25688 116622 25740 116628
rect 25700 115530 25728 116622
rect 25872 116544 25924 116550
rect 25872 116486 25924 116492
rect 25884 116006 25912 116486
rect 25872 116000 25924 116006
rect 25872 115942 25924 115948
rect 25688 115524 25740 115530
rect 25688 115466 25740 115472
rect 25504 114708 25556 114714
rect 25504 114650 25556 114656
rect 24860 114640 24912 114646
rect 24860 114582 24912 114588
rect 24400 114572 24452 114578
rect 24400 114514 24452 114520
rect 26252 113966 26280 119200
rect 26436 117366 26464 119200
rect 26424 117360 26476 117366
rect 26424 117302 26476 117308
rect 26424 117156 26476 117162
rect 26424 117098 26476 117104
rect 26436 116249 26464 117098
rect 26712 116346 26740 119200
rect 26608 116340 26660 116346
rect 26608 116282 26660 116288
rect 26700 116340 26752 116346
rect 26700 116282 26752 116288
rect 26422 116240 26478 116249
rect 26422 116175 26478 116184
rect 26424 115048 26476 115054
rect 26422 115016 26424 115025
rect 26476 115016 26478 115025
rect 26422 114951 26478 114960
rect 26620 114714 26648 116282
rect 26700 116068 26752 116074
rect 26700 116010 26752 116016
rect 26712 114918 26740 116010
rect 26700 114912 26752 114918
rect 26700 114854 26752 114860
rect 26608 114708 26660 114714
rect 26608 114650 26660 114656
rect 26896 113966 26924 119200
rect 26974 117328 27030 117337
rect 27172 117298 27200 119200
rect 27356 117434 27384 119200
rect 27344 117428 27396 117434
rect 27344 117370 27396 117376
rect 26974 117263 27030 117272
rect 27160 117292 27212 117298
rect 26988 116346 27016 117263
rect 27160 117234 27212 117240
rect 27160 117156 27212 117162
rect 27160 117098 27212 117104
rect 26976 116340 27028 116346
rect 26976 116282 27028 116288
rect 27172 116278 27200 117098
rect 27160 116272 27212 116278
rect 27160 116214 27212 116220
rect 26976 116136 27028 116142
rect 26976 116078 27028 116084
rect 26988 115734 27016 116078
rect 26976 115728 27028 115734
rect 26976 115670 27028 115676
rect 27068 115728 27120 115734
rect 27068 115670 27120 115676
rect 27080 115122 27108 115670
rect 27068 115116 27120 115122
rect 27068 115058 27120 115064
rect 27632 113966 27660 119200
rect 27712 117224 27764 117230
rect 27712 117166 27764 117172
rect 27724 116346 27752 117166
rect 27816 116890 27844 119200
rect 28092 116890 28120 119200
rect 28172 117088 28224 117094
rect 28172 117030 28224 117036
rect 27804 116884 27856 116890
rect 27804 116826 27856 116832
rect 28080 116884 28132 116890
rect 28080 116826 28132 116832
rect 27896 116748 27948 116754
rect 27896 116690 27948 116696
rect 27712 116340 27764 116346
rect 27712 116282 27764 116288
rect 27908 115666 27936 116690
rect 27896 115660 27948 115666
rect 27896 115602 27948 115608
rect 28080 115660 28132 115666
rect 28080 115602 28132 115608
rect 27712 115592 27764 115598
rect 28092 115546 28120 115602
rect 27764 115540 28120 115546
rect 27712 115534 28120 115540
rect 27724 115518 28120 115534
rect 28184 115530 28212 117030
rect 28276 116346 28304 119200
rect 28356 117156 28408 117162
rect 28356 117098 28408 117104
rect 28264 116340 28316 116346
rect 28264 116282 28316 116288
rect 28368 116113 28396 117098
rect 28552 116822 28580 119200
rect 28632 117156 28684 117162
rect 28632 117098 28684 117104
rect 28644 117065 28672 117098
rect 28630 117056 28686 117065
rect 28630 116991 28686 117000
rect 28448 116816 28500 116822
rect 28448 116758 28500 116764
rect 28540 116816 28592 116822
rect 28540 116758 28592 116764
rect 28354 116104 28410 116113
rect 28354 116039 28410 116048
rect 28172 115524 28224 115530
rect 28172 115466 28224 115472
rect 28460 114714 28488 116758
rect 28632 116748 28684 116754
rect 28632 116690 28684 116696
rect 28540 116680 28592 116686
rect 28540 116622 28592 116628
rect 28552 114714 28580 116622
rect 28644 115258 28672 116690
rect 28736 116346 28764 119200
rect 28816 117632 28868 117638
rect 28816 117574 28868 117580
rect 28828 117094 28856 117574
rect 28908 117360 28960 117366
rect 28908 117302 28960 117308
rect 28816 117088 28868 117094
rect 28816 117030 28868 117036
rect 28920 116890 28948 117302
rect 28908 116884 28960 116890
rect 28908 116826 28960 116832
rect 28816 116748 28868 116754
rect 28816 116690 28868 116696
rect 28724 116340 28776 116346
rect 28724 116282 28776 116288
rect 28724 116068 28776 116074
rect 28724 116010 28776 116016
rect 28632 115252 28684 115258
rect 28632 115194 28684 115200
rect 28448 114708 28500 114714
rect 28448 114650 28500 114656
rect 28540 114708 28592 114714
rect 28540 114650 28592 114656
rect 23388 113960 23440 113966
rect 23388 113902 23440 113908
rect 26240 113960 26292 113966
rect 26240 113902 26292 113908
rect 26884 113960 26936 113966
rect 26884 113902 26936 113908
rect 27620 113960 27672 113966
rect 27620 113902 27672 113908
rect 25780 113892 25832 113898
rect 25780 113834 25832 113840
rect 25044 113552 25096 113558
rect 25044 113494 25096 113500
rect 23032 109006 23152 109034
rect 17592 108520 17644 108526
rect 17592 108462 17644 108468
rect 16948 85808 17000 85814
rect 16948 85750 17000 85756
rect 16488 84040 16540 84046
rect 16488 83982 16540 83988
rect 16028 82952 16080 82958
rect 16028 82894 16080 82900
rect 15844 81796 15896 81802
rect 15844 81738 15896 81744
rect 15568 81388 15620 81394
rect 15568 81330 15620 81336
rect 14832 79756 14884 79762
rect 14832 79698 14884 79704
rect 14556 74724 14608 74730
rect 14556 74666 14608 74672
rect 14464 70440 14516 70446
rect 14464 70382 14516 70388
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14108 3670 14136 14826
rect 14476 5574 14504 70382
rect 14568 22438 14596 74666
rect 14556 22432 14608 22438
rect 14556 22374 14608 22380
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 13648 1686 13768 1714
rect 13740 800 13768 1686
rect 14108 800 14136 2450
rect 14384 800 14412 4014
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14752 800 14780 3334
rect 14844 1970 14872 79698
rect 15292 71528 15344 71534
rect 15292 71470 15344 71476
rect 14924 14544 14976 14550
rect 14924 14486 14976 14492
rect 14936 3602 14964 14486
rect 15304 8838 15332 71470
rect 15580 71194 15608 81330
rect 15752 71460 15804 71466
rect 15752 71402 15804 71408
rect 15568 71188 15620 71194
rect 15568 71130 15620 71136
rect 15476 70984 15528 70990
rect 15476 70926 15528 70932
rect 15488 70854 15516 70926
rect 15476 70848 15528 70854
rect 15476 70790 15528 70796
rect 15488 70446 15516 70790
rect 15476 70440 15528 70446
rect 15476 70382 15528 70388
rect 15488 69902 15516 70382
rect 15476 69896 15528 69902
rect 15476 69838 15528 69844
rect 15384 62348 15436 62354
rect 15384 62290 15436 62296
rect 15396 12434 15424 62290
rect 15660 58472 15712 58478
rect 15660 58414 15712 58420
rect 15672 43450 15700 58414
rect 15764 56506 15792 71402
rect 15856 70650 15884 81738
rect 15936 72616 15988 72622
rect 15936 72558 15988 72564
rect 15844 70644 15896 70650
rect 15844 70586 15896 70592
rect 15752 56500 15804 56506
rect 15752 56442 15804 56448
rect 15660 43444 15712 43450
rect 15660 43386 15712 43392
rect 15476 43240 15528 43246
rect 15476 43182 15528 43188
rect 15488 14278 15516 43182
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15396 12406 15516 12434
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 14832 1964 14884 1970
rect 14832 1906 14884 1912
rect 15028 800 15056 2926
rect 15396 800 15424 2926
rect 15488 2038 15516 12406
rect 15948 9926 15976 72558
rect 16040 71670 16068 82894
rect 16212 80232 16264 80238
rect 16212 80174 16264 80180
rect 16120 73840 16172 73846
rect 16120 73782 16172 73788
rect 16132 72826 16160 73782
rect 16120 72820 16172 72826
rect 16120 72762 16172 72768
rect 16028 71664 16080 71670
rect 16028 71606 16080 71612
rect 16224 70106 16252 80174
rect 16304 79348 16356 79354
rect 16304 79290 16356 79296
rect 16212 70100 16264 70106
rect 16212 70042 16264 70048
rect 16120 69896 16172 69902
rect 16120 69838 16172 69844
rect 16132 69426 16160 69838
rect 16316 69562 16344 79290
rect 16396 77988 16448 77994
rect 16396 77930 16448 77936
rect 16408 71194 16436 77930
rect 16500 72282 16528 83982
rect 16672 81864 16724 81870
rect 16672 81806 16724 81812
rect 16488 72276 16540 72282
rect 16488 72218 16540 72224
rect 16580 72072 16632 72078
rect 16580 72014 16632 72020
rect 16592 71602 16620 72014
rect 16580 71596 16632 71602
rect 16580 71538 16632 71544
rect 16396 71188 16448 71194
rect 16396 71130 16448 71136
rect 16580 70984 16632 70990
rect 16580 70926 16632 70932
rect 16592 70530 16620 70926
rect 16684 70650 16712 81806
rect 16960 72826 16988 85750
rect 17500 80776 17552 80782
rect 17500 80718 17552 80724
rect 17132 79552 17184 79558
rect 17132 79494 17184 79500
rect 16948 72820 17000 72826
rect 16948 72762 17000 72768
rect 17040 72616 17092 72622
rect 17040 72558 17092 72564
rect 16948 72548 17000 72554
rect 16948 72490 17000 72496
rect 16856 71732 16908 71738
rect 16856 71674 16908 71680
rect 16868 71602 16896 71674
rect 16856 71596 16908 71602
rect 16856 71538 16908 71544
rect 16764 71188 16816 71194
rect 16764 71130 16816 71136
rect 16672 70644 16724 70650
rect 16672 70586 16724 70592
rect 16408 70514 16620 70530
rect 16396 70508 16620 70514
rect 16448 70502 16620 70508
rect 16396 70450 16448 70456
rect 16304 69556 16356 69562
rect 16304 69498 16356 69504
rect 16120 69420 16172 69426
rect 16120 69362 16172 69368
rect 16776 64874 16804 71130
rect 16868 70990 16896 71538
rect 16856 70984 16908 70990
rect 16856 70926 16908 70932
rect 16776 64846 16896 64874
rect 16580 60172 16632 60178
rect 16580 60114 16632 60120
rect 16028 55888 16080 55894
rect 16028 55830 16080 55836
rect 16040 40050 16068 55830
rect 16488 53236 16540 53242
rect 16488 53178 16540 53184
rect 16304 43444 16356 43450
rect 16304 43386 16356 43392
rect 16316 42770 16344 43386
rect 16396 43240 16448 43246
rect 16396 43182 16448 43188
rect 16120 42764 16172 42770
rect 16120 42706 16172 42712
rect 16304 42764 16356 42770
rect 16304 42706 16356 42712
rect 16028 40044 16080 40050
rect 16028 39986 16080 39992
rect 16132 15366 16160 42706
rect 16304 42152 16356 42158
rect 16304 42094 16356 42100
rect 16316 17542 16344 42094
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16408 15910 16436 43182
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15764 3602 15792 6258
rect 16396 5092 16448 5098
rect 16396 5034 16448 5040
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15476 2032 15528 2038
rect 15476 1974 15528 1980
rect 15672 800 15700 3334
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 16040 800 16068 2450
rect 16316 800 16344 2926
rect 16408 2582 16436 5034
rect 16500 3194 16528 53178
rect 16592 42362 16620 60114
rect 16868 56506 16896 64846
rect 16856 56500 16908 56506
rect 16856 56442 16908 56448
rect 16764 56228 16816 56234
rect 16764 56170 16816 56176
rect 16776 48686 16804 56170
rect 16856 56160 16908 56166
rect 16856 56102 16908 56108
rect 16868 55962 16896 56102
rect 16856 55956 16908 55962
rect 16856 55898 16908 55904
rect 16764 48680 16816 48686
rect 16764 48622 16816 48628
rect 16776 47598 16804 48622
rect 16856 48544 16908 48550
rect 16856 48486 16908 48492
rect 16764 47592 16816 47598
rect 16764 47534 16816 47540
rect 16868 43314 16896 48486
rect 16856 43308 16908 43314
rect 16856 43250 16908 43256
rect 16868 42702 16896 43250
rect 16856 42696 16908 42702
rect 16856 42638 16908 42644
rect 16580 42356 16632 42362
rect 16580 42298 16632 42304
rect 16868 42226 16896 42638
rect 16856 42220 16908 42226
rect 16856 42162 16908 42168
rect 16672 39976 16724 39982
rect 16672 39918 16724 39924
rect 16684 21894 16712 39918
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16960 12170 16988 72490
rect 17052 13190 17080 72558
rect 17144 71738 17172 79494
rect 17316 73636 17368 73642
rect 17316 73578 17368 73584
rect 17328 72758 17356 73578
rect 17408 73568 17460 73574
rect 17408 73510 17460 73516
rect 17316 72752 17368 72758
rect 17316 72694 17368 72700
rect 17224 72480 17276 72486
rect 17224 72422 17276 72428
rect 17132 71732 17184 71738
rect 17132 71674 17184 71680
rect 17236 70854 17264 72422
rect 17328 71602 17356 72694
rect 17420 72690 17448 73510
rect 17408 72684 17460 72690
rect 17408 72626 17460 72632
rect 17420 72146 17448 72626
rect 17408 72140 17460 72146
rect 17408 72082 17460 72088
rect 17316 71596 17368 71602
rect 17316 71538 17368 71544
rect 17408 71392 17460 71398
rect 17408 71334 17460 71340
rect 17224 70848 17276 70854
rect 17224 70790 17276 70796
rect 17236 70446 17264 70790
rect 17224 70440 17276 70446
rect 17224 70382 17276 70388
rect 17316 64320 17368 64326
rect 17316 64262 17368 64268
rect 17328 56302 17356 64262
rect 17316 56296 17368 56302
rect 17316 56238 17368 56244
rect 17316 47456 17368 47462
rect 17316 47398 17368 47404
rect 17224 40588 17276 40594
rect 17224 40530 17276 40536
rect 17132 39908 17184 39914
rect 17132 39850 17184 39856
rect 17144 20806 17172 39850
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 17236 20262 17264 40530
rect 17328 40526 17356 47398
rect 17316 40520 17368 40526
rect 17316 40462 17368 40468
rect 17328 40118 17356 40462
rect 17316 40112 17368 40118
rect 17316 40054 17368 40060
rect 17328 39982 17356 40054
rect 17316 39976 17368 39982
rect 17316 39918 17368 39924
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17040 13184 17092 13190
rect 17040 13126 17092 13132
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 17420 8362 17448 71334
rect 17512 70650 17540 80718
rect 17500 70644 17552 70650
rect 17500 70586 17552 70592
rect 17500 42764 17552 42770
rect 17500 42706 17552 42712
rect 17512 16998 17540 42706
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16776 4010 16804 5102
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16592 2922 16620 3470
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 16684 800 16712 3878
rect 17604 3058 17632 108462
rect 19580 108284 19876 108304
rect 19636 108282 19660 108284
rect 19716 108282 19740 108284
rect 19796 108282 19820 108284
rect 19658 108230 19660 108282
rect 19722 108230 19734 108282
rect 19796 108230 19798 108282
rect 19636 108228 19660 108230
rect 19716 108228 19740 108230
rect 19796 108228 19820 108230
rect 19580 108208 19876 108228
rect 19580 107196 19876 107216
rect 19636 107194 19660 107196
rect 19716 107194 19740 107196
rect 19796 107194 19820 107196
rect 19658 107142 19660 107194
rect 19722 107142 19734 107194
rect 19796 107142 19798 107194
rect 19636 107140 19660 107142
rect 19716 107140 19740 107142
rect 19796 107140 19820 107142
rect 19580 107120 19876 107140
rect 19580 106108 19876 106128
rect 19636 106106 19660 106108
rect 19716 106106 19740 106108
rect 19796 106106 19820 106108
rect 19658 106054 19660 106106
rect 19722 106054 19734 106106
rect 19796 106054 19798 106106
rect 19636 106052 19660 106054
rect 19716 106052 19740 106054
rect 19796 106052 19820 106054
rect 19580 106032 19876 106052
rect 19580 105020 19876 105040
rect 19636 105018 19660 105020
rect 19716 105018 19740 105020
rect 19796 105018 19820 105020
rect 19658 104966 19660 105018
rect 19722 104966 19734 105018
rect 19796 104966 19798 105018
rect 19636 104964 19660 104966
rect 19716 104964 19740 104966
rect 19796 104964 19820 104966
rect 19580 104944 19876 104964
rect 19580 103932 19876 103952
rect 19636 103930 19660 103932
rect 19716 103930 19740 103932
rect 19796 103930 19820 103932
rect 19658 103878 19660 103930
rect 19722 103878 19734 103930
rect 19796 103878 19798 103930
rect 19636 103876 19660 103878
rect 19716 103876 19740 103878
rect 19796 103876 19820 103878
rect 19580 103856 19876 103876
rect 23032 103514 23060 109006
rect 22940 103486 23060 103514
rect 19580 102844 19876 102864
rect 19636 102842 19660 102844
rect 19716 102842 19740 102844
rect 19796 102842 19820 102844
rect 19658 102790 19660 102842
rect 19722 102790 19734 102842
rect 19796 102790 19798 102842
rect 19636 102788 19660 102790
rect 19716 102788 19740 102790
rect 19796 102788 19820 102790
rect 19580 102768 19876 102788
rect 18604 101992 18656 101998
rect 18604 101934 18656 101940
rect 17684 84652 17736 84658
rect 17684 84594 17736 84600
rect 17696 72282 17724 84594
rect 17776 83564 17828 83570
rect 17776 83506 17828 83512
rect 17684 72276 17736 72282
rect 17684 72218 17736 72224
rect 17788 71738 17816 83506
rect 17868 83496 17920 83502
rect 17868 83438 17920 83444
rect 17880 72826 17908 83438
rect 17868 72820 17920 72826
rect 17868 72762 17920 72768
rect 17776 71732 17828 71738
rect 17776 71674 17828 71680
rect 17868 71664 17920 71670
rect 17868 71606 17920 71612
rect 17776 70984 17828 70990
rect 17776 70926 17828 70932
rect 17788 56506 17816 70926
rect 17776 56500 17828 56506
rect 17776 56442 17828 56448
rect 17684 55820 17736 55826
rect 17684 55762 17736 55768
rect 17696 40186 17724 55762
rect 17684 40180 17736 40186
rect 17684 40122 17736 40128
rect 17880 11558 17908 71606
rect 18512 55140 18564 55146
rect 18512 55082 18564 55088
rect 18524 40050 18552 55082
rect 18512 40044 18564 40050
rect 18512 39986 18564 39992
rect 18328 39976 18380 39982
rect 18328 39918 18380 39924
rect 18340 18630 18368 39918
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17696 4010 17724 6326
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 16960 800 16988 2450
rect 17328 800 17356 2926
rect 17788 2774 17816 3878
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 17696 2746 17816 2774
rect 17696 1986 17724 2746
rect 17604 1958 17724 1986
rect 17604 800 17632 1958
rect 17972 800 18000 3538
rect 18248 2514 18276 5170
rect 18616 3058 18644 101934
rect 19580 101756 19876 101776
rect 19636 101754 19660 101756
rect 19716 101754 19740 101756
rect 19796 101754 19820 101756
rect 19658 101702 19660 101754
rect 19722 101702 19734 101754
rect 19796 101702 19798 101754
rect 19636 101700 19660 101702
rect 19716 101700 19740 101702
rect 19796 101700 19820 101702
rect 19580 101680 19876 101700
rect 19580 100668 19876 100688
rect 19636 100666 19660 100668
rect 19716 100666 19740 100668
rect 19796 100666 19820 100668
rect 19658 100614 19660 100666
rect 19722 100614 19734 100666
rect 19796 100614 19798 100666
rect 19636 100612 19660 100614
rect 19716 100612 19740 100614
rect 19796 100612 19820 100614
rect 19580 100592 19876 100612
rect 19580 99580 19876 99600
rect 19636 99578 19660 99580
rect 19716 99578 19740 99580
rect 19796 99578 19820 99580
rect 19658 99526 19660 99578
rect 19722 99526 19734 99578
rect 19796 99526 19798 99578
rect 19636 99524 19660 99526
rect 19716 99524 19740 99526
rect 19796 99524 19820 99526
rect 19580 99504 19876 99524
rect 19580 98492 19876 98512
rect 19636 98490 19660 98492
rect 19716 98490 19740 98492
rect 19796 98490 19820 98492
rect 19658 98438 19660 98490
rect 19722 98438 19734 98490
rect 19796 98438 19798 98490
rect 19636 98436 19660 98438
rect 19716 98436 19740 98438
rect 19796 98436 19820 98438
rect 19580 98416 19876 98436
rect 19580 97404 19876 97424
rect 19636 97402 19660 97404
rect 19716 97402 19740 97404
rect 19796 97402 19820 97404
rect 19658 97350 19660 97402
rect 19722 97350 19734 97402
rect 19796 97350 19798 97402
rect 19636 97348 19660 97350
rect 19716 97348 19740 97350
rect 19796 97348 19820 97350
rect 19580 97328 19876 97348
rect 19580 96316 19876 96336
rect 19636 96314 19660 96316
rect 19716 96314 19740 96316
rect 19796 96314 19820 96316
rect 19658 96262 19660 96314
rect 19722 96262 19734 96314
rect 19796 96262 19798 96314
rect 19636 96260 19660 96262
rect 19716 96260 19740 96262
rect 19796 96260 19820 96262
rect 19580 96240 19876 96260
rect 19580 95228 19876 95248
rect 19636 95226 19660 95228
rect 19716 95226 19740 95228
rect 19796 95226 19820 95228
rect 19658 95174 19660 95226
rect 19722 95174 19734 95226
rect 19796 95174 19798 95226
rect 19636 95172 19660 95174
rect 19716 95172 19740 95174
rect 19796 95172 19820 95174
rect 19580 95152 19876 95172
rect 19580 94140 19876 94160
rect 19636 94138 19660 94140
rect 19716 94138 19740 94140
rect 19796 94138 19820 94140
rect 19658 94086 19660 94138
rect 19722 94086 19734 94138
rect 19796 94086 19798 94138
rect 19636 94084 19660 94086
rect 19716 94084 19740 94086
rect 19796 94084 19820 94086
rect 19580 94064 19876 94084
rect 19580 93052 19876 93072
rect 19636 93050 19660 93052
rect 19716 93050 19740 93052
rect 19796 93050 19820 93052
rect 19658 92998 19660 93050
rect 19722 92998 19734 93050
rect 19796 92998 19798 93050
rect 19636 92996 19660 92998
rect 19716 92996 19740 92998
rect 19796 92996 19820 92998
rect 19580 92976 19876 92996
rect 21364 92812 21416 92818
rect 21364 92754 21416 92760
rect 19580 91964 19876 91984
rect 19636 91962 19660 91964
rect 19716 91962 19740 91964
rect 19796 91962 19820 91964
rect 19658 91910 19660 91962
rect 19722 91910 19734 91962
rect 19796 91910 19798 91962
rect 19636 91908 19660 91910
rect 19716 91908 19740 91910
rect 19796 91908 19820 91910
rect 19580 91888 19876 91908
rect 19340 91792 19392 91798
rect 19340 91734 19392 91740
rect 18788 58132 18840 58138
rect 18788 58074 18840 58080
rect 18696 54800 18748 54806
rect 18696 54742 18748 54748
rect 18708 39914 18736 54742
rect 18800 43382 18828 58074
rect 19352 53786 19380 91734
rect 19580 90876 19876 90896
rect 19636 90874 19660 90876
rect 19716 90874 19740 90876
rect 19796 90874 19820 90876
rect 19658 90822 19660 90874
rect 19722 90822 19734 90874
rect 19796 90822 19798 90874
rect 19636 90820 19660 90822
rect 19716 90820 19740 90822
rect 19796 90820 19820 90822
rect 19580 90800 19876 90820
rect 19580 89788 19876 89808
rect 19636 89786 19660 89788
rect 19716 89786 19740 89788
rect 19796 89786 19820 89788
rect 19658 89734 19660 89786
rect 19722 89734 19734 89786
rect 19796 89734 19798 89786
rect 19636 89732 19660 89734
rect 19716 89732 19740 89734
rect 19796 89732 19820 89734
rect 19580 89712 19876 89732
rect 19580 88700 19876 88720
rect 19636 88698 19660 88700
rect 19716 88698 19740 88700
rect 19796 88698 19820 88700
rect 19658 88646 19660 88698
rect 19722 88646 19734 88698
rect 19796 88646 19798 88698
rect 19636 88644 19660 88646
rect 19716 88644 19740 88646
rect 19796 88644 19820 88646
rect 19580 88624 19876 88644
rect 19580 87612 19876 87632
rect 19636 87610 19660 87612
rect 19716 87610 19740 87612
rect 19796 87610 19820 87612
rect 19658 87558 19660 87610
rect 19722 87558 19734 87610
rect 19796 87558 19798 87610
rect 19636 87556 19660 87558
rect 19716 87556 19740 87558
rect 19796 87556 19820 87558
rect 19580 87536 19876 87556
rect 21180 87372 21232 87378
rect 21180 87314 21232 87320
rect 20352 87236 20404 87242
rect 20352 87178 20404 87184
rect 19580 86524 19876 86544
rect 19636 86522 19660 86524
rect 19716 86522 19740 86524
rect 19796 86522 19820 86524
rect 19658 86470 19660 86522
rect 19722 86470 19734 86522
rect 19796 86470 19798 86522
rect 19636 86468 19660 86470
rect 19716 86468 19740 86470
rect 19796 86468 19820 86470
rect 19580 86448 19876 86468
rect 19580 85436 19876 85456
rect 19636 85434 19660 85436
rect 19716 85434 19740 85436
rect 19796 85434 19820 85436
rect 19658 85382 19660 85434
rect 19722 85382 19734 85434
rect 19796 85382 19798 85434
rect 19636 85380 19660 85382
rect 19716 85380 19740 85382
rect 19796 85380 19820 85382
rect 19580 85360 19876 85380
rect 19580 84348 19876 84368
rect 19636 84346 19660 84348
rect 19716 84346 19740 84348
rect 19796 84346 19820 84348
rect 19658 84294 19660 84346
rect 19722 84294 19734 84346
rect 19796 84294 19798 84346
rect 19636 84292 19660 84294
rect 19716 84292 19740 84294
rect 19796 84292 19820 84294
rect 19580 84272 19876 84292
rect 19580 83260 19876 83280
rect 19636 83258 19660 83260
rect 19716 83258 19740 83260
rect 19796 83258 19820 83260
rect 19658 83206 19660 83258
rect 19722 83206 19734 83258
rect 19796 83206 19798 83258
rect 19636 83204 19660 83206
rect 19716 83204 19740 83206
rect 19796 83204 19820 83206
rect 19580 83184 19876 83204
rect 19580 82172 19876 82192
rect 19636 82170 19660 82172
rect 19716 82170 19740 82172
rect 19796 82170 19820 82172
rect 19658 82118 19660 82170
rect 19722 82118 19734 82170
rect 19796 82118 19798 82170
rect 19636 82116 19660 82118
rect 19716 82116 19740 82118
rect 19796 82116 19820 82118
rect 19580 82096 19876 82116
rect 19580 81084 19876 81104
rect 19636 81082 19660 81084
rect 19716 81082 19740 81084
rect 19796 81082 19820 81084
rect 19658 81030 19660 81082
rect 19722 81030 19734 81082
rect 19796 81030 19798 81082
rect 19636 81028 19660 81030
rect 19716 81028 19740 81030
rect 19796 81028 19820 81030
rect 19580 81008 19876 81028
rect 19580 79996 19876 80016
rect 19636 79994 19660 79996
rect 19716 79994 19740 79996
rect 19796 79994 19820 79996
rect 19658 79942 19660 79994
rect 19722 79942 19734 79994
rect 19796 79942 19798 79994
rect 19636 79940 19660 79942
rect 19716 79940 19740 79942
rect 19796 79940 19820 79942
rect 19580 79920 19876 79940
rect 19580 78908 19876 78928
rect 19636 78906 19660 78908
rect 19716 78906 19740 78908
rect 19796 78906 19820 78908
rect 19658 78854 19660 78906
rect 19722 78854 19734 78906
rect 19796 78854 19798 78906
rect 19636 78852 19660 78854
rect 19716 78852 19740 78854
rect 19796 78852 19820 78854
rect 19580 78832 19876 78852
rect 19580 77820 19876 77840
rect 19636 77818 19660 77820
rect 19716 77818 19740 77820
rect 19796 77818 19820 77820
rect 19658 77766 19660 77818
rect 19722 77766 19734 77818
rect 19796 77766 19798 77818
rect 19636 77764 19660 77766
rect 19716 77764 19740 77766
rect 19796 77764 19820 77766
rect 19580 77744 19876 77764
rect 19580 76732 19876 76752
rect 19636 76730 19660 76732
rect 19716 76730 19740 76732
rect 19796 76730 19820 76732
rect 19658 76678 19660 76730
rect 19722 76678 19734 76730
rect 19796 76678 19798 76730
rect 19636 76676 19660 76678
rect 19716 76676 19740 76678
rect 19796 76676 19820 76678
rect 19580 76656 19876 76676
rect 20076 75880 20128 75886
rect 20076 75822 20128 75828
rect 19580 75644 19876 75664
rect 19636 75642 19660 75644
rect 19716 75642 19740 75644
rect 19796 75642 19820 75644
rect 19658 75590 19660 75642
rect 19722 75590 19734 75642
rect 19796 75590 19798 75642
rect 19636 75588 19660 75590
rect 19716 75588 19740 75590
rect 19796 75588 19820 75590
rect 19580 75568 19876 75588
rect 20088 75342 20116 75822
rect 20076 75336 20128 75342
rect 20076 75278 20128 75284
rect 20088 74866 20116 75278
rect 20364 75002 20392 87178
rect 20536 86284 20588 86290
rect 20536 86226 20588 86232
rect 20444 86148 20496 86154
rect 20444 86090 20496 86096
rect 20456 75546 20484 86090
rect 20548 75886 20576 86226
rect 20536 75880 20588 75886
rect 20536 75822 20588 75828
rect 21192 75546 21220 87314
rect 20444 75540 20496 75546
rect 20444 75482 20496 75488
rect 21180 75540 21232 75546
rect 21180 75482 21232 75488
rect 20996 75404 21048 75410
rect 20996 75346 21048 75352
rect 20352 74996 20404 75002
rect 20352 74938 20404 74944
rect 20076 74860 20128 74866
rect 20076 74802 20128 74808
rect 19580 74556 19876 74576
rect 19636 74554 19660 74556
rect 19716 74554 19740 74556
rect 19796 74554 19820 74556
rect 19658 74502 19660 74554
rect 19722 74502 19734 74554
rect 19796 74502 19798 74554
rect 19636 74500 19660 74502
rect 19716 74500 19740 74502
rect 19796 74500 19820 74502
rect 19580 74480 19876 74500
rect 20168 73704 20220 73710
rect 20168 73646 20220 73652
rect 19580 73468 19876 73488
rect 19636 73466 19660 73468
rect 19716 73466 19740 73468
rect 19796 73466 19820 73468
rect 19658 73414 19660 73466
rect 19722 73414 19734 73466
rect 19796 73414 19798 73466
rect 19636 73412 19660 73414
rect 19716 73412 19740 73414
rect 19796 73412 19820 73414
rect 19580 73392 19876 73412
rect 20180 72622 20208 73646
rect 20168 72616 20220 72622
rect 20168 72558 20220 72564
rect 19580 72380 19876 72400
rect 19636 72378 19660 72380
rect 19716 72378 19740 72380
rect 19796 72378 19820 72380
rect 19658 72326 19660 72378
rect 19722 72326 19734 72378
rect 19796 72326 19798 72378
rect 19636 72324 19660 72326
rect 19716 72324 19740 72326
rect 19796 72324 19820 72326
rect 19580 72304 19876 72324
rect 19580 71292 19876 71312
rect 19636 71290 19660 71292
rect 19716 71290 19740 71292
rect 19796 71290 19820 71292
rect 19658 71238 19660 71290
rect 19722 71238 19734 71290
rect 19796 71238 19798 71290
rect 19636 71236 19660 71238
rect 19716 71236 19740 71238
rect 19796 71236 19820 71238
rect 19580 71216 19876 71236
rect 19580 70204 19876 70224
rect 19636 70202 19660 70204
rect 19716 70202 19740 70204
rect 19796 70202 19820 70204
rect 19658 70150 19660 70202
rect 19722 70150 19734 70202
rect 19796 70150 19798 70202
rect 19636 70148 19660 70150
rect 19716 70148 19740 70150
rect 19796 70148 19820 70150
rect 19580 70128 19876 70148
rect 19580 69116 19876 69136
rect 19636 69114 19660 69116
rect 19716 69114 19740 69116
rect 19796 69114 19820 69116
rect 19658 69062 19660 69114
rect 19722 69062 19734 69114
rect 19796 69062 19798 69114
rect 19636 69060 19660 69062
rect 19716 69060 19740 69062
rect 19796 69060 19820 69062
rect 19580 69040 19876 69060
rect 19580 68028 19876 68048
rect 19636 68026 19660 68028
rect 19716 68026 19740 68028
rect 19796 68026 19820 68028
rect 19658 67974 19660 68026
rect 19722 67974 19734 68026
rect 19796 67974 19798 68026
rect 19636 67972 19660 67974
rect 19716 67972 19740 67974
rect 19796 67972 19820 67974
rect 19580 67952 19876 67972
rect 19580 66940 19876 66960
rect 19636 66938 19660 66940
rect 19716 66938 19740 66940
rect 19796 66938 19820 66940
rect 19658 66886 19660 66938
rect 19722 66886 19734 66938
rect 19796 66886 19798 66938
rect 19636 66884 19660 66886
rect 19716 66884 19740 66886
rect 19796 66884 19820 66886
rect 19580 66864 19876 66884
rect 19580 65852 19876 65872
rect 19636 65850 19660 65852
rect 19716 65850 19740 65852
rect 19796 65850 19820 65852
rect 19658 65798 19660 65850
rect 19722 65798 19734 65850
rect 19796 65798 19798 65850
rect 19636 65796 19660 65798
rect 19716 65796 19740 65798
rect 19796 65796 19820 65798
rect 19580 65776 19876 65796
rect 19580 64764 19876 64784
rect 19636 64762 19660 64764
rect 19716 64762 19740 64764
rect 19796 64762 19820 64764
rect 19658 64710 19660 64762
rect 19722 64710 19734 64762
rect 19796 64710 19798 64762
rect 19636 64708 19660 64710
rect 19716 64708 19740 64710
rect 19796 64708 19820 64710
rect 19580 64688 19876 64708
rect 20180 64598 20208 72558
rect 20168 64592 20220 64598
rect 20168 64534 20220 64540
rect 19580 63676 19876 63696
rect 19636 63674 19660 63676
rect 19716 63674 19740 63676
rect 19796 63674 19820 63676
rect 19658 63622 19660 63674
rect 19722 63622 19734 63674
rect 19796 63622 19798 63674
rect 19636 63620 19660 63622
rect 19716 63620 19740 63622
rect 19796 63620 19820 63622
rect 19580 63600 19876 63620
rect 19580 62588 19876 62608
rect 19636 62586 19660 62588
rect 19716 62586 19740 62588
rect 19796 62586 19820 62588
rect 19658 62534 19660 62586
rect 19722 62534 19734 62586
rect 19796 62534 19798 62586
rect 19636 62532 19660 62534
rect 19716 62532 19740 62534
rect 19796 62532 19820 62534
rect 19580 62512 19876 62532
rect 19580 61500 19876 61520
rect 19636 61498 19660 61500
rect 19716 61498 19740 61500
rect 19796 61498 19820 61500
rect 19658 61446 19660 61498
rect 19722 61446 19734 61498
rect 19796 61446 19798 61498
rect 19636 61444 19660 61446
rect 19716 61444 19740 61446
rect 19796 61444 19820 61446
rect 19580 61424 19876 61444
rect 19580 60412 19876 60432
rect 19636 60410 19660 60412
rect 19716 60410 19740 60412
rect 19796 60410 19820 60412
rect 19658 60358 19660 60410
rect 19722 60358 19734 60410
rect 19796 60358 19798 60410
rect 19636 60356 19660 60358
rect 19716 60356 19740 60358
rect 19796 60356 19820 60358
rect 19580 60336 19876 60356
rect 19580 59324 19876 59344
rect 19636 59322 19660 59324
rect 19716 59322 19740 59324
rect 19796 59322 19820 59324
rect 19658 59270 19660 59322
rect 19722 59270 19734 59322
rect 19796 59270 19798 59322
rect 19636 59268 19660 59270
rect 19716 59268 19740 59270
rect 19796 59268 19820 59270
rect 19580 59248 19876 59268
rect 19580 58236 19876 58256
rect 19636 58234 19660 58236
rect 19716 58234 19740 58236
rect 19796 58234 19820 58236
rect 19658 58182 19660 58234
rect 19722 58182 19734 58234
rect 19796 58182 19798 58234
rect 19636 58180 19660 58182
rect 19716 58180 19740 58182
rect 19796 58180 19820 58182
rect 19580 58160 19876 58180
rect 19580 57148 19876 57168
rect 19636 57146 19660 57148
rect 19716 57146 19740 57148
rect 19796 57146 19820 57148
rect 19658 57094 19660 57146
rect 19722 57094 19734 57146
rect 19796 57094 19798 57146
rect 19636 57092 19660 57094
rect 19716 57092 19740 57094
rect 19796 57092 19820 57094
rect 19580 57072 19876 57092
rect 19580 56060 19876 56080
rect 19636 56058 19660 56060
rect 19716 56058 19740 56060
rect 19796 56058 19820 56060
rect 19658 56006 19660 56058
rect 19722 56006 19734 56058
rect 19796 56006 19798 56058
rect 19636 56004 19660 56006
rect 19716 56004 19740 56006
rect 19796 56004 19820 56006
rect 19580 55984 19876 56004
rect 19580 54972 19876 54992
rect 19636 54970 19660 54972
rect 19716 54970 19740 54972
rect 19796 54970 19820 54972
rect 19658 54918 19660 54970
rect 19722 54918 19734 54970
rect 19796 54918 19798 54970
rect 19636 54916 19660 54918
rect 19716 54916 19740 54918
rect 19796 54916 19820 54918
rect 19580 54896 19876 54916
rect 19580 53884 19876 53904
rect 19636 53882 19660 53884
rect 19716 53882 19740 53884
rect 19796 53882 19820 53884
rect 19658 53830 19660 53882
rect 19722 53830 19734 53882
rect 19796 53830 19798 53882
rect 19636 53828 19660 53830
rect 19716 53828 19740 53830
rect 19796 53828 19820 53830
rect 19580 53808 19876 53828
rect 19340 53780 19392 53786
rect 19340 53722 19392 53728
rect 19432 53440 19484 53446
rect 19432 53382 19484 53388
rect 18788 43376 18840 43382
rect 18788 43318 18840 43324
rect 18696 39908 18748 39914
rect 18696 39850 18748 39856
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18708 4078 18736 14350
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 18340 800 18368 2926
rect 18708 1986 18736 3878
rect 19352 3754 19380 6802
rect 19260 3738 19380 3754
rect 19444 3738 19472 53382
rect 19580 52796 19876 52816
rect 19636 52794 19660 52796
rect 19716 52794 19740 52796
rect 19796 52794 19820 52796
rect 19658 52742 19660 52794
rect 19722 52742 19734 52794
rect 19796 52742 19798 52794
rect 19636 52740 19660 52742
rect 19716 52740 19740 52742
rect 19796 52740 19820 52742
rect 19580 52720 19876 52740
rect 19580 51708 19876 51728
rect 19636 51706 19660 51708
rect 19716 51706 19740 51708
rect 19796 51706 19820 51708
rect 19658 51654 19660 51706
rect 19722 51654 19734 51706
rect 19796 51654 19798 51706
rect 19636 51652 19660 51654
rect 19716 51652 19740 51654
rect 19796 51652 19820 51654
rect 19580 51632 19876 51652
rect 19580 50620 19876 50640
rect 19636 50618 19660 50620
rect 19716 50618 19740 50620
rect 19796 50618 19820 50620
rect 19658 50566 19660 50618
rect 19722 50566 19734 50618
rect 19796 50566 19798 50618
rect 19636 50564 19660 50566
rect 19716 50564 19740 50566
rect 19796 50564 19820 50566
rect 19580 50544 19876 50564
rect 19580 49532 19876 49552
rect 19636 49530 19660 49532
rect 19716 49530 19740 49532
rect 19796 49530 19820 49532
rect 19658 49478 19660 49530
rect 19722 49478 19734 49530
rect 19796 49478 19798 49530
rect 19636 49476 19660 49478
rect 19716 49476 19740 49478
rect 19796 49476 19820 49478
rect 19580 49456 19876 49476
rect 19580 48444 19876 48464
rect 19636 48442 19660 48444
rect 19716 48442 19740 48444
rect 19796 48442 19820 48444
rect 19658 48390 19660 48442
rect 19722 48390 19734 48442
rect 19796 48390 19798 48442
rect 19636 48388 19660 48390
rect 19716 48388 19740 48390
rect 19796 48388 19820 48390
rect 19580 48368 19876 48388
rect 19580 47356 19876 47376
rect 19636 47354 19660 47356
rect 19716 47354 19740 47356
rect 19796 47354 19820 47356
rect 19658 47302 19660 47354
rect 19722 47302 19734 47354
rect 19796 47302 19798 47354
rect 19636 47300 19660 47302
rect 19716 47300 19740 47302
rect 19796 47300 19820 47302
rect 19580 47280 19876 47300
rect 19580 46268 19876 46288
rect 19636 46266 19660 46268
rect 19716 46266 19740 46268
rect 19796 46266 19820 46268
rect 19658 46214 19660 46266
rect 19722 46214 19734 46266
rect 19796 46214 19798 46266
rect 19636 46212 19660 46214
rect 19716 46212 19740 46214
rect 19796 46212 19820 46214
rect 19580 46192 19876 46212
rect 19580 45180 19876 45200
rect 19636 45178 19660 45180
rect 19716 45178 19740 45180
rect 19796 45178 19820 45180
rect 19658 45126 19660 45178
rect 19722 45126 19734 45178
rect 19796 45126 19798 45178
rect 19636 45124 19660 45126
rect 19716 45124 19740 45126
rect 19796 45124 19820 45126
rect 19580 45104 19876 45124
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19580 42928 19876 42948
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 19580 40828 19876 40848
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 21008 24070 21036 75346
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 21376 16574 21404 92754
rect 21548 91860 21600 91866
rect 21548 91802 21600 91808
rect 21560 54330 21588 91802
rect 22836 70848 22888 70854
rect 22836 70790 22888 70796
rect 21548 54324 21600 54330
rect 21548 54266 21600 54272
rect 21376 16546 21496 16574
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 20916 12986 20944 13738
rect 21088 13728 21140 13734
rect 21088 13670 21140 13676
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19248 3732 19380 3738
rect 19300 3726 19380 3732
rect 19432 3732 19484 3738
rect 19248 3674 19300 3680
rect 19432 3674 19484 3680
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 18972 2508 19024 2514
rect 18972 2450 19024 2456
rect 18616 1958 18736 1986
rect 18616 800 18644 1958
rect 18984 800 19012 2450
rect 19260 800 19288 3538
rect 19904 3482 19932 12786
rect 21100 12782 21128 13670
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 19984 4072 20036 4078
rect 19984 4014 20036 4020
rect 19812 3454 19932 3482
rect 19812 3126 19840 3454
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19800 3120 19852 3126
rect 19800 3062 19852 3068
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19904 1714 19932 3334
rect 19628 1686 19932 1714
rect 19628 800 19656 1686
rect 19996 1578 20024 4014
rect 20076 4004 20128 4010
rect 20076 3946 20128 3952
rect 20088 3738 20116 3946
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 20272 3194 20300 3878
rect 20260 3188 20312 3194
rect 20260 3130 20312 3136
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20364 2854 20392 3130
rect 20456 2990 20484 3878
rect 20640 3602 20668 6394
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20732 3602 20760 4082
rect 20996 4004 21048 4010
rect 20996 3946 21048 3952
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 20260 2508 20312 2514
rect 20260 2450 20312 2456
rect 19904 1550 20024 1578
rect 19904 800 19932 1550
rect 20272 800 20300 2450
rect 20548 800 20576 2926
rect 20916 800 20944 3538
rect 21008 3398 21036 3946
rect 20996 3392 21048 3398
rect 20996 3334 21048 3340
rect 21284 2922 21312 6054
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 21376 3058 21404 3334
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 21272 2916 21324 2922
rect 21272 2858 21324 2864
rect 21468 2514 21496 16546
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22664 15706 22692 15982
rect 22652 15700 22704 15706
rect 22652 15642 22704 15648
rect 22848 14958 22876 70790
rect 22940 53786 22968 103486
rect 23480 95940 23532 95946
rect 23480 95882 23532 95888
rect 23492 76566 23520 95882
rect 24216 82884 24268 82890
rect 24216 82826 24268 82832
rect 23572 81524 23624 81530
rect 23572 81466 23624 81472
rect 23584 80054 23612 81466
rect 23756 80708 23808 80714
rect 23756 80650 23808 80656
rect 23584 80026 23704 80054
rect 23480 76560 23532 76566
rect 23480 76502 23532 76508
rect 23112 76492 23164 76498
rect 23112 76434 23164 76440
rect 22928 53780 22980 53786
rect 22928 53722 22980 53728
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 22940 15570 22968 16390
rect 23020 15972 23072 15978
rect 23020 15914 23072 15920
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22744 14816 22796 14822
rect 22744 14758 22796 14764
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22296 13462 22324 13670
rect 22284 13456 22336 13462
rect 22284 13398 22336 13404
rect 22388 13394 22416 13670
rect 22572 13394 22600 13874
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22560 13388 22612 13394
rect 22560 13330 22612 13336
rect 21560 12850 21588 13330
rect 21548 12844 21600 12850
rect 21548 12786 21600 12792
rect 22572 12714 22600 13330
rect 22560 12708 22612 12714
rect 22560 12650 22612 12656
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 22204 11898 22232 12378
rect 22572 12306 22600 12650
rect 22756 12374 22784 14758
rect 22940 12374 22968 15506
rect 23032 14482 23060 15914
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 22744 12368 22796 12374
rect 22744 12310 22796 12316
rect 22928 12368 22980 12374
rect 22928 12310 22980 12316
rect 22560 12300 22612 12306
rect 22560 12242 22612 12248
rect 22572 11898 22600 12242
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22560 11892 22612 11898
rect 22560 11834 22612 11840
rect 22572 11218 22600 11834
rect 22560 11212 22612 11218
rect 22560 11154 22612 11160
rect 22744 7948 22796 7954
rect 22744 7890 22796 7896
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21456 2508 21508 2514
rect 21456 2450 21508 2456
rect 21192 800 21220 2450
rect 21560 800 21588 2790
rect 21836 800 21864 4014
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 21928 3126 21956 3878
rect 21916 3120 21968 3126
rect 21916 3062 21968 3068
rect 22756 2990 22784 7890
rect 22836 4072 22888 4078
rect 22836 4014 22888 4020
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22204 800 22232 2450
rect 22572 800 22600 2790
rect 22848 800 22876 4014
rect 23124 2650 23152 76434
rect 23492 73710 23520 76502
rect 23480 73704 23532 73710
rect 23480 73646 23532 73652
rect 23572 20256 23624 20262
rect 23572 20198 23624 20204
rect 23388 18148 23440 18154
rect 23388 18090 23440 18096
rect 23204 15360 23256 15366
rect 23204 15302 23256 15308
rect 23216 13870 23244 15302
rect 23296 15088 23348 15094
rect 23296 15030 23348 15036
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 23308 12442 23336 15030
rect 23400 12918 23428 18090
rect 23480 16516 23532 16522
rect 23480 16458 23532 16464
rect 23492 14618 23520 16458
rect 23584 15570 23612 20198
rect 23676 15706 23704 80026
rect 23664 15700 23716 15706
rect 23664 15642 23716 15648
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 23768 14958 23796 80650
rect 23848 76356 23900 76362
rect 23848 76298 23900 76304
rect 23860 75478 23888 76298
rect 23848 75472 23900 75478
rect 23848 75414 23900 75420
rect 24124 19304 24176 19310
rect 24124 19246 24176 19252
rect 24136 18970 24164 19246
rect 24124 18964 24176 18970
rect 24124 18906 24176 18912
rect 23848 18080 23900 18086
rect 23848 18022 23900 18028
rect 23860 17814 23888 18022
rect 23848 17808 23900 17814
rect 23848 17750 23900 17756
rect 23940 17808 23992 17814
rect 23940 17750 23992 17756
rect 23860 16250 23888 17750
rect 23848 16244 23900 16250
rect 23848 16186 23900 16192
rect 23952 16046 23980 17750
rect 24124 17060 24176 17066
rect 24124 17002 24176 17008
rect 24032 16652 24084 16658
rect 24032 16594 24084 16600
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 23848 15972 23900 15978
rect 23848 15914 23900 15920
rect 23860 15570 23888 15914
rect 23848 15564 23900 15570
rect 23848 15506 23900 15512
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 23572 14952 23624 14958
rect 23572 14894 23624 14900
rect 23756 14952 23808 14958
rect 23756 14894 23808 14900
rect 23584 14793 23612 14894
rect 23756 14816 23808 14822
rect 23570 14784 23626 14793
rect 23756 14758 23808 14764
rect 23570 14719 23626 14728
rect 23480 14612 23532 14618
rect 23480 14554 23532 14560
rect 23572 14612 23624 14618
rect 23572 14554 23624 14560
rect 23478 14512 23534 14521
rect 23478 14447 23480 14456
rect 23532 14447 23534 14456
rect 23480 14418 23532 14424
rect 23584 14074 23612 14554
rect 23664 14408 23716 14414
rect 23662 14376 23664 14385
rect 23716 14376 23718 14385
rect 23662 14311 23718 14320
rect 23572 14068 23624 14074
rect 23572 14010 23624 14016
rect 23584 13326 23612 14010
rect 23572 13320 23624 13326
rect 23572 13262 23624 13268
rect 23388 12912 23440 12918
rect 23388 12854 23440 12860
rect 23296 12436 23348 12442
rect 23296 12378 23348 12384
rect 23400 4826 23428 12854
rect 23664 12708 23716 12714
rect 23664 12650 23716 12656
rect 23676 11558 23704 12650
rect 23664 11552 23716 11558
rect 23664 11494 23716 11500
rect 23676 6186 23704 11494
rect 23768 11286 23796 14758
rect 23860 14074 23888 15302
rect 23940 15088 23992 15094
rect 23940 15030 23992 15036
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 23756 11280 23808 11286
rect 23756 11222 23808 11228
rect 23664 6180 23716 6186
rect 23664 6122 23716 6128
rect 23572 5296 23624 5302
rect 23572 5238 23624 5244
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 23216 800 23244 4014
rect 23584 2990 23612 5238
rect 23860 5030 23888 13126
rect 23952 11082 23980 15030
rect 24044 13938 24072 16594
rect 24136 16522 24164 17002
rect 24228 16658 24256 82826
rect 24400 54052 24452 54058
rect 24400 53994 24452 54000
rect 24412 22094 24440 53994
rect 25056 53786 25084 113494
rect 25792 102134 25820 113834
rect 27160 109064 27212 109070
rect 27160 109006 27212 109012
rect 27068 105800 27120 105806
rect 27068 105742 27120 105748
rect 25780 102128 25832 102134
rect 25780 102070 25832 102076
rect 26976 84584 27028 84590
rect 26976 84526 27028 84532
rect 26516 81728 26568 81734
rect 26516 81670 26568 81676
rect 25596 81456 25648 81462
rect 25596 81398 25648 81404
rect 25504 80640 25556 80646
rect 25504 80582 25556 80588
rect 25044 53780 25096 53786
rect 25044 53722 25096 53728
rect 25044 53644 25096 53650
rect 25044 53586 25096 53592
rect 25056 53242 25084 53586
rect 25044 53236 25096 53242
rect 25044 53178 25096 53184
rect 24860 50312 24912 50318
rect 24860 50254 24912 50260
rect 24872 49230 24900 50254
rect 24860 49224 24912 49230
rect 24860 49166 24912 49172
rect 24860 42900 24912 42906
rect 24860 42842 24912 42848
rect 24872 42158 24900 42842
rect 24860 42152 24912 42158
rect 24860 42094 24912 42100
rect 25412 26920 25464 26926
rect 25412 26862 25464 26868
rect 25424 26382 25452 26862
rect 25228 26376 25280 26382
rect 25228 26318 25280 26324
rect 25412 26376 25464 26382
rect 25412 26318 25464 26324
rect 24412 22066 24624 22094
rect 24308 17536 24360 17542
rect 24308 17478 24360 17484
rect 24320 16658 24348 17478
rect 24216 16652 24268 16658
rect 24216 16594 24268 16600
rect 24308 16652 24360 16658
rect 24308 16594 24360 16600
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 24308 16040 24360 16046
rect 24308 15982 24360 15988
rect 24216 15496 24268 15502
rect 24216 15438 24268 15444
rect 24228 14958 24256 15438
rect 24320 15094 24348 15982
rect 24400 15360 24452 15366
rect 24400 15302 24452 15308
rect 24308 15088 24360 15094
rect 24308 15030 24360 15036
rect 24216 14952 24268 14958
rect 24216 14894 24268 14900
rect 24320 14618 24348 15030
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 24214 13560 24270 13569
rect 24214 13495 24270 13504
rect 24228 13462 24256 13495
rect 24216 13456 24268 13462
rect 24216 13398 24268 13404
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 24228 12646 24256 12922
rect 24216 12640 24268 12646
rect 24216 12582 24268 12588
rect 23940 11076 23992 11082
rect 23940 11018 23992 11024
rect 23952 6254 23980 11018
rect 24320 7818 24348 14010
rect 24412 13462 24440 15302
rect 24492 15020 24544 15026
rect 24492 14962 24544 14968
rect 24504 14074 24532 14962
rect 24492 14068 24544 14074
rect 24492 14010 24544 14016
rect 24400 13456 24452 13462
rect 24400 13398 24452 13404
rect 24492 13320 24544 13326
rect 24492 13262 24544 13268
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 24412 11694 24440 12582
rect 24504 12306 24532 13262
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24400 11688 24452 11694
rect 24400 11630 24452 11636
rect 24308 7812 24360 7818
rect 24308 7754 24360 7760
rect 23940 6248 23992 6254
rect 23940 6190 23992 6196
rect 23848 5024 23900 5030
rect 23848 4966 23900 4972
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 23848 3596 23900 3602
rect 23848 3538 23900 3544
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23768 2990 23796 3334
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23756 2984 23808 2990
rect 23756 2926 23808 2932
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 23492 800 23520 2790
rect 23860 800 23888 3538
rect 24136 800 24164 4014
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24228 3194 24256 3470
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24412 3194 24440 3334
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24400 3188 24452 3194
rect 24400 3130 24452 3136
rect 24504 800 24532 3334
rect 24596 2650 24624 22066
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 25134 18728 25190 18737
rect 24688 17338 24716 18702
rect 25134 18663 25190 18672
rect 24768 18624 24820 18630
rect 24768 18566 24820 18572
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24780 17882 24808 18566
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24688 16726 24716 17274
rect 24780 17066 24808 17818
rect 24768 17060 24820 17066
rect 24768 17002 24820 17008
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 24676 16720 24728 16726
rect 24676 16662 24728 16668
rect 24872 16658 24900 16934
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24688 14482 24716 16390
rect 24768 15632 24820 15638
rect 24768 15574 24820 15580
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24688 14278 24716 14418
rect 24676 14272 24728 14278
rect 24676 14214 24728 14220
rect 24780 13190 24808 15574
rect 24860 15360 24912 15366
rect 24860 15302 24912 15308
rect 24872 13530 24900 15302
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 24768 13184 24820 13190
rect 24768 13126 24820 13132
rect 24860 13184 24912 13190
rect 24860 13126 24912 13132
rect 24872 12850 24900 13126
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24964 12782 24992 18566
rect 25148 17134 25176 18663
rect 25240 18290 25268 26318
rect 25516 20262 25544 80582
rect 25608 73846 25636 81398
rect 26424 80980 26476 80986
rect 26424 80922 26476 80928
rect 25596 73840 25648 73846
rect 25596 73782 25648 73788
rect 26332 70372 26384 70378
rect 26332 70314 26384 70320
rect 26148 65068 26200 65074
rect 26148 65010 26200 65016
rect 25688 59628 25740 59634
rect 25688 59570 25740 59576
rect 25596 59016 25648 59022
rect 25596 58958 25648 58964
rect 25608 42770 25636 58958
rect 25700 43450 25728 59570
rect 25688 43444 25740 43450
rect 25688 43386 25740 43392
rect 25596 42764 25648 42770
rect 25596 42706 25648 42712
rect 26160 41138 26188 65010
rect 26148 41132 26200 41138
rect 26148 41074 26200 41080
rect 26056 26376 26108 26382
rect 26056 26318 26108 26324
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 26068 19990 26096 26318
rect 26148 23588 26200 23594
rect 26148 23530 26200 23536
rect 26056 19984 26108 19990
rect 26056 19926 26108 19932
rect 25780 19916 25832 19922
rect 25780 19858 25832 19864
rect 25504 18896 25556 18902
rect 25504 18838 25556 18844
rect 25228 18284 25280 18290
rect 25228 18226 25280 18232
rect 25240 17814 25268 18226
rect 25516 18154 25544 18838
rect 25504 18148 25556 18154
rect 25504 18090 25556 18096
rect 25228 17808 25280 17814
rect 25228 17750 25280 17756
rect 25240 17678 25268 17750
rect 25228 17672 25280 17678
rect 25228 17614 25280 17620
rect 25240 17202 25268 17614
rect 25228 17196 25280 17202
rect 25228 17138 25280 17144
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 25056 16114 25084 16526
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 25148 14793 25176 17070
rect 25516 16794 25544 18090
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 25412 16108 25464 16114
rect 25412 16050 25464 16056
rect 25424 15570 25452 16050
rect 25412 15564 25464 15570
rect 25240 15524 25412 15552
rect 25134 14784 25190 14793
rect 25134 14719 25190 14728
rect 25240 13870 25268 15524
rect 25412 15506 25464 15512
rect 25320 14884 25372 14890
rect 25320 14826 25372 14832
rect 25332 14346 25360 14826
rect 25688 14816 25740 14822
rect 25688 14758 25740 14764
rect 25320 14340 25372 14346
rect 25320 14282 25372 14288
rect 25228 13864 25280 13870
rect 25228 13806 25280 13812
rect 25240 13394 25268 13806
rect 25228 13388 25280 13394
rect 25228 13330 25280 13336
rect 25240 12850 25268 13330
rect 25228 12844 25280 12850
rect 25228 12786 25280 12792
rect 24952 12776 25004 12782
rect 24952 12718 25004 12724
rect 25700 6322 25728 14758
rect 25792 10130 25820 19858
rect 26160 19310 26188 23530
rect 26148 19304 26200 19310
rect 26148 19246 26200 19252
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 25964 19236 26016 19242
rect 25964 19178 26016 19184
rect 26056 19236 26108 19242
rect 26056 19178 26108 19184
rect 25976 17218 26004 19178
rect 26068 18834 26096 19178
rect 26056 18828 26108 18834
rect 26056 18770 26108 18776
rect 25976 17190 26096 17218
rect 25964 17128 26016 17134
rect 25964 17070 26016 17076
rect 25976 16250 26004 17070
rect 25964 16244 26016 16250
rect 25964 16186 26016 16192
rect 26068 14521 26096 17190
rect 26252 16726 26280 19246
rect 26344 18834 26372 70314
rect 26332 18828 26384 18834
rect 26332 18770 26384 18776
rect 26436 18714 26464 80922
rect 26344 18686 26464 18714
rect 26344 16946 26372 18686
rect 26424 18624 26476 18630
rect 26424 18566 26476 18572
rect 26436 18426 26464 18566
rect 26424 18420 26476 18426
rect 26424 18362 26476 18368
rect 26436 17066 26464 18362
rect 26424 17060 26476 17066
rect 26424 17002 26476 17008
rect 26344 16918 26464 16946
rect 26240 16720 26292 16726
rect 26240 16662 26292 16668
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26252 14634 26280 15846
rect 26160 14606 26280 14634
rect 26054 14512 26110 14521
rect 26054 14447 26110 14456
rect 26160 13326 26188 14606
rect 26240 14476 26292 14482
rect 26240 14418 26292 14424
rect 26252 14006 26280 14418
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 26240 14000 26292 14006
rect 26240 13942 26292 13948
rect 26240 13864 26292 13870
rect 26240 13806 26292 13812
rect 26252 13394 26280 13806
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 26148 13320 26200 13326
rect 26148 13262 26200 13268
rect 26056 13252 26108 13258
rect 26056 13194 26108 13200
rect 25964 13184 26016 13190
rect 25964 13126 26016 13132
rect 25976 12374 26004 13126
rect 25964 12368 26016 12374
rect 25964 12310 26016 12316
rect 26068 12102 26096 13194
rect 26252 12442 26280 13330
rect 26344 12782 26372 14214
rect 26436 12782 26464 16918
rect 26528 14482 26556 81670
rect 26792 80164 26844 80170
rect 26792 80106 26844 80112
rect 26608 71596 26660 71602
rect 26608 71538 26660 71544
rect 26620 70446 26648 71538
rect 26608 70440 26660 70446
rect 26608 70382 26660 70388
rect 26700 23520 26752 23526
rect 26700 23462 26752 23468
rect 26712 22574 26740 23462
rect 26700 22568 26752 22574
rect 26700 22510 26752 22516
rect 26804 22094 26832 80106
rect 26988 78674 27016 84526
rect 26976 78668 27028 78674
rect 26976 78610 27028 78616
rect 26976 28008 27028 28014
rect 26976 27950 27028 27956
rect 26884 27872 26936 27878
rect 26884 27814 26936 27820
rect 26896 26994 26924 27814
rect 26884 26988 26936 26994
rect 26884 26930 26936 26936
rect 26988 26926 27016 27950
rect 26976 26920 27028 26926
rect 26976 26862 27028 26868
rect 26712 22066 26832 22094
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26620 18737 26648 18770
rect 26606 18728 26662 18737
rect 26606 18663 26662 18672
rect 26608 18624 26660 18630
rect 26608 18566 26660 18572
rect 26620 18222 26648 18566
rect 26608 18216 26660 18222
rect 26608 18158 26660 18164
rect 26608 15360 26660 15366
rect 26608 15302 26660 15308
rect 26620 15026 26648 15302
rect 26608 15020 26660 15026
rect 26608 14962 26660 14968
rect 26516 14476 26568 14482
rect 26516 14418 26568 14424
rect 26516 13728 26568 13734
rect 26516 13670 26568 13676
rect 26528 12850 26556 13670
rect 26620 13410 26648 14962
rect 26712 13530 26740 22066
rect 26976 19848 27028 19854
rect 26976 19790 27028 19796
rect 26792 19508 26844 19514
rect 26792 19450 26844 19456
rect 26804 18154 26832 19450
rect 26988 19394 27016 19790
rect 27080 19514 27108 105742
rect 27172 86766 27200 109006
rect 27620 105664 27672 105670
rect 27620 105606 27672 105612
rect 27160 86760 27212 86766
rect 27160 86702 27212 86708
rect 27172 85678 27200 86702
rect 27160 85672 27212 85678
rect 27160 85614 27212 85620
rect 27172 84590 27200 85614
rect 27160 84584 27212 84590
rect 27160 84526 27212 84532
rect 27528 67924 27580 67930
rect 27528 67866 27580 67872
rect 27540 50862 27568 67866
rect 27528 50856 27580 50862
rect 27528 50798 27580 50804
rect 27632 48686 27660 105606
rect 28736 103514 28764 116010
rect 28828 115666 28856 116690
rect 28908 116612 28960 116618
rect 28908 116554 28960 116560
rect 28816 115660 28868 115666
rect 28816 115602 28868 115608
rect 28920 115258 28948 116554
rect 29012 115957 29040 119200
rect 28998 115948 29054 115957
rect 28998 115883 29054 115892
rect 29196 115841 29224 119200
rect 29276 117700 29328 117706
rect 29276 117642 29328 117648
rect 29288 117094 29316 117642
rect 29276 117088 29328 117094
rect 29276 117030 29328 117036
rect 29368 116748 29420 116754
rect 29368 116690 29420 116696
rect 29276 116340 29328 116346
rect 29276 116282 29328 116288
rect 29182 115832 29238 115841
rect 29182 115767 29238 115776
rect 29184 115524 29236 115530
rect 29184 115466 29236 115472
rect 29196 115297 29224 115466
rect 29182 115288 29238 115297
rect 28908 115252 28960 115258
rect 29182 115223 29238 115232
rect 28908 115194 28960 115200
rect 28816 115048 28868 115054
rect 28814 115016 28816 115025
rect 29184 115048 29236 115054
rect 28868 115016 28870 115025
rect 29184 114990 29236 114996
rect 28814 114951 28870 114960
rect 29196 113354 29224 114990
rect 29184 113348 29236 113354
rect 29184 113290 29236 113296
rect 29288 113014 29316 116282
rect 29380 115161 29408 116690
rect 29472 115734 29500 119200
rect 29550 115832 29606 115841
rect 29550 115767 29552 115776
rect 29604 115767 29606 115776
rect 29552 115738 29604 115744
rect 29460 115728 29512 115734
rect 29460 115670 29512 115676
rect 29550 115696 29606 115705
rect 29550 115631 29606 115640
rect 29564 115598 29592 115631
rect 29552 115592 29604 115598
rect 29552 115534 29604 115540
rect 29656 115258 29684 119200
rect 29828 117156 29880 117162
rect 29828 117098 29880 117104
rect 29840 116210 29868 117098
rect 29828 116204 29880 116210
rect 29828 116146 29880 116152
rect 29644 115252 29696 115258
rect 29644 115194 29696 115200
rect 29366 115152 29422 115161
rect 29366 115087 29422 115096
rect 29368 115048 29420 115054
rect 29368 114990 29420 114996
rect 29380 114102 29408 114990
rect 29932 114714 29960 119200
rect 30012 117156 30064 117162
rect 30012 117098 30064 117104
rect 30024 116550 30052 117098
rect 30012 116544 30064 116550
rect 30012 116486 30064 116492
rect 30012 115184 30064 115190
rect 30012 115126 30064 115132
rect 29920 114708 29972 114714
rect 29920 114650 29972 114656
rect 30024 114578 30052 115126
rect 30116 114578 30144 119200
rect 30392 116872 30420 119200
rect 30576 117042 30604 119200
rect 30576 117014 30696 117042
rect 30392 116844 30604 116872
rect 30472 116748 30524 116754
rect 30472 116690 30524 116696
rect 30288 116000 30340 116006
rect 30288 115942 30340 115948
rect 30378 115968 30434 115977
rect 30300 115802 30328 115942
rect 30378 115903 30434 115912
rect 30288 115796 30340 115802
rect 30288 115738 30340 115744
rect 30392 115682 30420 115903
rect 30208 115654 30420 115682
rect 30012 114572 30064 114578
rect 30012 114514 30064 114520
rect 30104 114572 30156 114578
rect 30104 114514 30156 114520
rect 29368 114096 29420 114102
rect 29368 114038 29420 114044
rect 30208 114050 30236 115654
rect 30286 115288 30342 115297
rect 30286 115223 30342 115232
rect 30300 114714 30328 115223
rect 30380 114980 30432 114986
rect 30380 114922 30432 114928
rect 30288 114708 30340 114714
rect 30288 114650 30340 114656
rect 30392 114170 30420 114922
rect 30380 114164 30432 114170
rect 30380 114106 30432 114112
rect 30208 114022 30420 114050
rect 29276 113008 29328 113014
rect 29276 112950 29328 112956
rect 30392 112878 30420 114022
rect 30380 112872 30432 112878
rect 30380 112814 30432 112820
rect 29000 112736 29052 112742
rect 29000 112678 29052 112684
rect 28552 103486 28764 103514
rect 27988 91180 28040 91186
rect 27988 91122 28040 91128
rect 27896 87780 27948 87786
rect 27896 87722 27948 87728
rect 27712 53984 27764 53990
rect 27712 53926 27764 53932
rect 27620 48680 27672 48686
rect 27620 48622 27672 48628
rect 27528 30388 27580 30394
rect 27528 30330 27580 30336
rect 27160 28008 27212 28014
rect 27160 27950 27212 27956
rect 27172 26858 27200 27950
rect 27540 27470 27568 30330
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27528 26920 27580 26926
rect 27528 26862 27580 26868
rect 27160 26852 27212 26858
rect 27160 26794 27212 26800
rect 27172 24818 27200 26794
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 27172 24274 27200 24754
rect 27540 24614 27568 26862
rect 27620 24744 27672 24750
rect 27620 24686 27672 24692
rect 27528 24608 27580 24614
rect 27528 24550 27580 24556
rect 27160 24268 27212 24274
rect 27160 24210 27212 24216
rect 27540 24138 27568 24550
rect 27632 24342 27660 24686
rect 27620 24336 27672 24342
rect 27620 24278 27672 24284
rect 27528 24132 27580 24138
rect 27528 24074 27580 24080
rect 27252 24064 27304 24070
rect 27252 24006 27304 24012
rect 27264 23662 27292 24006
rect 27252 23656 27304 23662
rect 27252 23598 27304 23604
rect 27436 23112 27488 23118
rect 27436 23054 27488 23060
rect 27448 22778 27476 23054
rect 27436 22772 27488 22778
rect 27436 22714 27488 22720
rect 27448 20602 27476 22714
rect 27160 20596 27212 20602
rect 27160 20538 27212 20544
rect 27436 20596 27488 20602
rect 27436 20538 27488 20544
rect 27068 19508 27120 19514
rect 27068 19450 27120 19456
rect 26988 19366 27108 19394
rect 26976 19304 27028 19310
rect 26976 19246 27028 19252
rect 26884 18828 26936 18834
rect 26884 18770 26936 18776
rect 26792 18148 26844 18154
rect 26792 18090 26844 18096
rect 26896 17814 26924 18770
rect 26884 17808 26936 17814
rect 26884 17750 26936 17756
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 26804 14822 26832 16186
rect 26988 14958 27016 19246
rect 26976 14952 27028 14958
rect 26976 14894 27028 14900
rect 26792 14816 26844 14822
rect 26792 14758 26844 14764
rect 26792 14272 26844 14278
rect 26792 14214 26844 14220
rect 26700 13524 26752 13530
rect 26700 13466 26752 13472
rect 26620 13382 26740 13410
rect 26608 12980 26660 12986
rect 26608 12922 26660 12928
rect 26516 12844 26568 12850
rect 26516 12786 26568 12792
rect 26332 12776 26384 12782
rect 26332 12718 26384 12724
rect 26424 12776 26476 12782
rect 26424 12718 26476 12724
rect 26240 12436 26292 12442
rect 26240 12378 26292 12384
rect 26056 12096 26108 12102
rect 26056 12038 26108 12044
rect 25780 10124 25832 10130
rect 25780 10066 25832 10072
rect 26528 8022 26556 12786
rect 26516 8016 26568 8022
rect 26516 7958 26568 7964
rect 26620 7750 26648 12922
rect 26608 7744 26660 7750
rect 26608 7686 26660 7692
rect 26712 6390 26740 13382
rect 26804 12986 26832 14214
rect 26884 13796 26936 13802
rect 26884 13738 26936 13744
rect 26896 13258 26924 13738
rect 26884 13252 26936 13258
rect 26884 13194 26936 13200
rect 26792 12980 26844 12986
rect 26792 12922 26844 12928
rect 27080 12850 27108 19366
rect 27172 18698 27200 20538
rect 27436 20392 27488 20398
rect 27436 20334 27488 20340
rect 27448 19514 27476 20334
rect 27540 19786 27568 24074
rect 27632 22438 27660 24278
rect 27620 22432 27672 22438
rect 27620 22374 27672 22380
rect 27632 19922 27660 22374
rect 27620 19916 27672 19922
rect 27620 19858 27672 19864
rect 27528 19780 27580 19786
rect 27528 19722 27580 19728
rect 27436 19508 27488 19514
rect 27436 19450 27488 19456
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27160 18692 27212 18698
rect 27160 18634 27212 18640
rect 27172 18222 27200 18634
rect 27252 18624 27304 18630
rect 27252 18566 27304 18572
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 27172 17678 27200 18158
rect 27160 17672 27212 17678
rect 27160 17614 27212 17620
rect 27160 17128 27212 17134
rect 27160 17070 27212 17076
rect 27172 15434 27200 17070
rect 27160 15428 27212 15434
rect 27160 15370 27212 15376
rect 27172 14550 27200 15370
rect 27160 14544 27212 14550
rect 27160 14486 27212 14492
rect 27172 13394 27200 14486
rect 27160 13388 27212 13394
rect 27160 13330 27212 13336
rect 27068 12844 27120 12850
rect 27068 12786 27120 12792
rect 27264 12730 27292 18566
rect 27356 15910 27384 19314
rect 27620 18216 27672 18222
rect 27620 18158 27672 18164
rect 27436 18148 27488 18154
rect 27436 18090 27488 18096
rect 27448 17338 27476 18090
rect 27436 17332 27488 17338
rect 27436 17274 27488 17280
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 27436 16040 27488 16046
rect 27436 15982 27488 15988
rect 27448 15910 27476 15982
rect 27344 15904 27396 15910
rect 27344 15846 27396 15852
rect 27436 15904 27488 15910
rect 27436 15846 27488 15852
rect 27356 15042 27384 15846
rect 27540 15502 27568 16050
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 27356 15014 27476 15042
rect 27448 14958 27476 15014
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 26896 12702 27292 12730
rect 26896 12434 26924 12702
rect 26804 12406 26924 12434
rect 26700 6384 26752 6390
rect 26700 6326 26752 6332
rect 25688 6316 25740 6322
rect 25688 6258 25740 6264
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 24688 3602 24716 5306
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 25964 4072 26016 4078
rect 25964 4014 26016 4020
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 24780 800 24808 4014
rect 25780 4004 25832 4010
rect 25780 3946 25832 3952
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 25596 3936 25648 3942
rect 25596 3878 25648 3884
rect 25042 3496 25098 3505
rect 25148 3466 25176 3878
rect 25320 3664 25372 3670
rect 25320 3606 25372 3612
rect 25042 3431 25044 3440
rect 25096 3431 25098 3440
rect 25136 3460 25188 3466
rect 25044 3402 25096 3408
rect 25136 3402 25188 3408
rect 25332 3126 25360 3606
rect 25412 3392 25464 3398
rect 25412 3334 25464 3340
rect 25320 3120 25372 3126
rect 25320 3062 25372 3068
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 25148 800 25176 2450
rect 25424 800 25452 3334
rect 25608 3058 25636 3878
rect 25596 3052 25648 3058
rect 25596 2994 25648 3000
rect 25792 800 25820 3946
rect 25976 3738 26004 4014
rect 26240 3936 26292 3942
rect 26240 3878 26292 3884
rect 26700 3936 26752 3942
rect 26700 3878 26752 3884
rect 25964 3732 26016 3738
rect 25964 3674 26016 3680
rect 26252 2990 26280 3878
rect 26330 3768 26386 3777
rect 26330 3703 26386 3712
rect 26344 3602 26372 3703
rect 26712 3670 26740 3878
rect 26700 3664 26752 3670
rect 26700 3606 26752 3612
rect 26332 3596 26384 3602
rect 26332 3538 26384 3544
rect 26608 3392 26660 3398
rect 26608 3334 26660 3340
rect 26620 3233 26648 3334
rect 26606 3224 26662 3233
rect 26606 3159 26662 3168
rect 26804 2990 26832 12406
rect 26884 4072 26936 4078
rect 26884 4014 26936 4020
rect 26240 2984 26292 2990
rect 26792 2984 26844 2990
rect 26240 2926 26292 2932
rect 26330 2952 26386 2961
rect 26792 2926 26844 2932
rect 26330 2887 26386 2896
rect 26344 2854 26372 2887
rect 26332 2848 26384 2854
rect 26332 2790 26384 2796
rect 26424 2848 26476 2854
rect 26424 2790 26476 2796
rect 26056 2508 26108 2514
rect 26056 2450 26108 2456
rect 26068 800 26096 2450
rect 26436 800 26464 2790
rect 26896 2774 26924 4014
rect 26804 2746 26924 2774
rect 26804 800 26832 2746
rect 27068 2508 27120 2514
rect 27068 2450 27120 2456
rect 27080 800 27108 2450
rect 27356 2310 27384 14894
rect 27434 14784 27490 14793
rect 27434 14719 27490 14728
rect 27448 12764 27476 14719
rect 27528 14408 27580 14414
rect 27528 14350 27580 14356
rect 27540 13258 27568 14350
rect 27632 13569 27660 18158
rect 27618 13560 27674 13569
rect 27618 13495 27674 13504
rect 27620 13320 27672 13326
rect 27620 13262 27672 13268
rect 27528 13252 27580 13258
rect 27528 13194 27580 13200
rect 27632 13190 27660 13262
rect 27620 13184 27672 13190
rect 27620 13126 27672 13132
rect 27620 12776 27672 12782
rect 27448 12736 27620 12764
rect 27620 12718 27672 12724
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 27528 4004 27580 4010
rect 27528 3946 27580 3952
rect 27540 3534 27568 3946
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 27436 3392 27488 3398
rect 27436 3334 27488 3340
rect 27344 2304 27396 2310
rect 27344 2246 27396 2252
rect 27448 800 27476 3334
rect 27632 3210 27660 7822
rect 27540 3194 27660 3210
rect 27528 3188 27660 3194
rect 27580 3182 27660 3188
rect 27528 3130 27580 3136
rect 27724 2650 27752 53926
rect 27804 28008 27856 28014
rect 27804 27950 27856 27956
rect 27816 27334 27844 27950
rect 27804 27328 27856 27334
rect 27804 27270 27856 27276
rect 27908 26234 27936 87722
rect 28000 53786 28028 91122
rect 28356 86692 28408 86698
rect 28356 86634 28408 86640
rect 28264 85604 28316 85610
rect 28264 85546 28316 85552
rect 28172 54120 28224 54126
rect 28172 54062 28224 54068
rect 27988 53780 28040 53786
rect 27988 53722 28040 53728
rect 27988 27600 28040 27606
rect 27988 27542 28040 27548
rect 28000 27130 28028 27542
rect 28080 27328 28132 27334
rect 28080 27270 28132 27276
rect 27988 27124 28040 27130
rect 27988 27066 28040 27072
rect 28092 26450 28120 27270
rect 28080 26444 28132 26450
rect 28080 26386 28132 26392
rect 27816 26206 27936 26234
rect 27816 22982 27844 26206
rect 27896 24744 27948 24750
rect 27896 24686 27948 24692
rect 27908 24206 27936 24686
rect 27896 24200 27948 24206
rect 27896 24142 27948 24148
rect 27908 23662 27936 24142
rect 27896 23656 27948 23662
rect 27896 23598 27948 23604
rect 27908 23322 27936 23598
rect 27988 23520 28040 23526
rect 27988 23462 28040 23468
rect 27896 23316 27948 23322
rect 27896 23258 27948 23264
rect 28000 23254 28028 23462
rect 27988 23248 28040 23254
rect 27988 23190 28040 23196
rect 27804 22976 27856 22982
rect 27804 22918 27856 22924
rect 27896 20392 27948 20398
rect 27896 20334 27948 20340
rect 27908 19922 27936 20334
rect 27896 19916 27948 19922
rect 27896 19858 27948 19864
rect 27896 19236 27948 19242
rect 27896 19178 27948 19184
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 27816 17542 27844 17614
rect 27804 17536 27856 17542
rect 27804 17478 27856 17484
rect 27816 16658 27844 17478
rect 27908 16726 27936 19178
rect 28080 18828 28132 18834
rect 28080 18770 28132 18776
rect 28092 18086 28120 18770
rect 28080 18080 28132 18086
rect 28080 18022 28132 18028
rect 27896 16720 27948 16726
rect 27896 16662 27948 16668
rect 27804 16652 27856 16658
rect 27804 16594 27856 16600
rect 27896 15632 27948 15638
rect 27896 15574 27948 15580
rect 27908 15473 27936 15574
rect 27894 15464 27950 15473
rect 27894 15399 27950 15408
rect 27896 15156 27948 15162
rect 27896 15098 27948 15104
rect 27802 14512 27858 14521
rect 27802 14447 27858 14456
rect 27816 13530 27844 14447
rect 27908 13870 27936 15098
rect 27896 13864 27948 13870
rect 27896 13806 27948 13812
rect 27804 13524 27856 13530
rect 27804 13466 27856 13472
rect 27988 4276 28040 4282
rect 27988 4218 28040 4224
rect 27896 4208 27948 4214
rect 27896 4150 27948 4156
rect 27908 3738 27936 4150
rect 27896 3732 27948 3738
rect 27896 3674 27948 3680
rect 28000 3670 28028 4218
rect 28080 3936 28132 3942
rect 28080 3878 28132 3884
rect 27988 3664 28040 3670
rect 27988 3606 28040 3612
rect 27804 3528 27856 3534
rect 27804 3470 27856 3476
rect 27712 2644 27764 2650
rect 27712 2586 27764 2592
rect 27816 1442 27844 3470
rect 28092 3058 28120 3878
rect 28080 3052 28132 3058
rect 28080 2994 28132 3000
rect 28080 2508 28132 2514
rect 28080 2450 28132 2456
rect 27724 1414 27844 1442
rect 27724 800 27752 1414
rect 28092 800 28120 2450
rect 28184 2378 28212 54062
rect 28276 19922 28304 85546
rect 28368 23186 28396 86634
rect 28552 60790 28580 103486
rect 28632 87168 28684 87174
rect 28632 87110 28684 87116
rect 28540 60784 28592 60790
rect 28540 60726 28592 60732
rect 28540 48680 28592 48686
rect 28540 48622 28592 48628
rect 28552 28014 28580 48622
rect 28540 28008 28592 28014
rect 28540 27950 28592 27956
rect 28540 27532 28592 27538
rect 28540 27474 28592 27480
rect 28552 23798 28580 27474
rect 28644 26234 28672 87110
rect 29012 64394 29040 112678
rect 29460 112464 29512 112470
rect 29460 112406 29512 112412
rect 29368 84516 29420 84522
rect 29368 84458 29420 84464
rect 29184 83904 29236 83910
rect 29184 83846 29236 83852
rect 29000 64388 29052 64394
rect 29000 64330 29052 64336
rect 28908 50380 28960 50386
rect 28908 50322 28960 50328
rect 28920 50250 28948 50322
rect 28908 50244 28960 50250
rect 28908 50186 28960 50192
rect 28920 38486 28948 50186
rect 28908 38480 28960 38486
rect 28908 38422 28960 38428
rect 28920 36310 28948 38422
rect 28724 36304 28776 36310
rect 28724 36246 28776 36252
rect 28908 36304 28960 36310
rect 28908 36246 28960 36252
rect 28736 35562 28764 36246
rect 28724 35556 28776 35562
rect 28724 35498 28776 35504
rect 28736 33454 28764 35498
rect 28724 33448 28776 33454
rect 28724 33390 28776 33396
rect 28644 26206 28764 26234
rect 28632 24268 28684 24274
rect 28632 24210 28684 24216
rect 28540 23792 28592 23798
rect 28540 23734 28592 23740
rect 28356 23180 28408 23186
rect 28356 23122 28408 23128
rect 28552 20398 28580 23734
rect 28644 22094 28672 24210
rect 28736 23730 28764 26206
rect 29092 24200 29144 24206
rect 29092 24142 29144 24148
rect 28724 23724 28776 23730
rect 28724 23666 28776 23672
rect 29104 23662 29132 24142
rect 29092 23656 29144 23662
rect 29092 23598 29144 23604
rect 28644 22066 28764 22094
rect 28540 20392 28592 20398
rect 28540 20334 28592 20340
rect 28264 19916 28316 19922
rect 28264 19858 28316 19864
rect 28540 19712 28592 19718
rect 28540 19654 28592 19660
rect 28632 19712 28684 19718
rect 28632 19654 28684 19660
rect 28448 19168 28500 19174
rect 28448 19110 28500 19116
rect 28356 18964 28408 18970
rect 28356 18906 28408 18912
rect 28262 18728 28318 18737
rect 28262 18663 28318 18672
rect 28276 18358 28304 18663
rect 28368 18426 28396 18906
rect 28460 18834 28488 19110
rect 28448 18828 28500 18834
rect 28448 18770 28500 18776
rect 28356 18420 28408 18426
rect 28356 18362 28408 18368
rect 28264 18352 28316 18358
rect 28264 18294 28316 18300
rect 28264 17876 28316 17882
rect 28264 17818 28316 17824
rect 28276 13734 28304 17818
rect 28368 16726 28396 18362
rect 28356 16720 28408 16726
rect 28356 16662 28408 16668
rect 28552 16046 28580 19654
rect 28540 16040 28592 16046
rect 28540 15982 28592 15988
rect 28644 15910 28672 19654
rect 28736 18766 28764 22066
rect 28816 20324 28868 20330
rect 28816 20266 28868 20272
rect 28724 18760 28776 18766
rect 28724 18702 28776 18708
rect 28736 18222 28764 18702
rect 28724 18216 28776 18222
rect 28724 18158 28776 18164
rect 28724 16448 28776 16454
rect 28724 16390 28776 16396
rect 28736 16046 28764 16390
rect 28724 16040 28776 16046
rect 28724 15982 28776 15988
rect 28540 15904 28592 15910
rect 28540 15846 28592 15852
rect 28632 15904 28684 15910
rect 28632 15846 28684 15852
rect 28356 15564 28408 15570
rect 28356 15506 28408 15512
rect 28368 14822 28396 15506
rect 28448 15360 28500 15366
rect 28448 15302 28500 15308
rect 28356 14816 28408 14822
rect 28356 14758 28408 14764
rect 28460 14074 28488 15302
rect 28552 14074 28580 15846
rect 28448 14068 28500 14074
rect 28448 14010 28500 14016
rect 28540 14068 28592 14074
rect 28540 14010 28592 14016
rect 28460 13818 28488 14010
rect 28368 13790 28488 13818
rect 28264 13728 28316 13734
rect 28264 13670 28316 13676
rect 28368 5166 28396 13790
rect 28448 13728 28500 13734
rect 28448 13670 28500 13676
rect 28460 7954 28488 13670
rect 28540 12980 28592 12986
rect 28540 12922 28592 12928
rect 28552 8090 28580 12922
rect 28540 8084 28592 8090
rect 28540 8026 28592 8032
rect 28448 7948 28500 7954
rect 28448 7890 28500 7896
rect 28644 6118 28672 15846
rect 28828 13938 28856 20266
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 28908 19780 28960 19786
rect 28908 19722 28960 19728
rect 28920 17882 28948 19722
rect 28908 17876 28960 17882
rect 28908 17818 28960 17824
rect 29012 17814 29040 19790
rect 29092 18080 29144 18086
rect 29092 18022 29144 18028
rect 29000 17808 29052 17814
rect 29000 17750 29052 17756
rect 28998 17640 29054 17649
rect 28998 17575 29054 17584
rect 29012 17134 29040 17575
rect 29000 17128 29052 17134
rect 29000 17070 29052 17076
rect 29000 16992 29052 16998
rect 29000 16934 29052 16940
rect 29012 15638 29040 16934
rect 29000 15632 29052 15638
rect 29000 15574 29052 15580
rect 28908 15428 28960 15434
rect 28908 15370 28960 15376
rect 28920 15162 28948 15370
rect 29000 15360 29052 15366
rect 29000 15302 29052 15308
rect 28908 15156 28960 15162
rect 28908 15098 28960 15104
rect 28908 14952 28960 14958
rect 28906 14920 28908 14929
rect 28960 14920 28962 14929
rect 28906 14855 28962 14864
rect 28906 14784 28962 14793
rect 28906 14719 28962 14728
rect 28816 13932 28868 13938
rect 28816 13874 28868 13880
rect 28724 13728 28776 13734
rect 28724 13670 28776 13676
rect 28736 13530 28764 13670
rect 28724 13524 28776 13530
rect 28724 13466 28776 13472
rect 28736 12782 28764 13466
rect 28920 13190 28948 14719
rect 28908 13184 28960 13190
rect 28908 13126 28960 13132
rect 28724 12776 28776 12782
rect 28724 12718 28776 12724
rect 29012 6458 29040 15302
rect 29104 13394 29132 18022
rect 29196 14958 29224 83846
rect 29276 83564 29328 83570
rect 29276 83506 29328 83512
rect 29288 83162 29316 83506
rect 29276 83156 29328 83162
rect 29276 83098 29328 83104
rect 29276 83020 29328 83026
rect 29276 82962 29328 82968
rect 29288 17270 29316 82962
rect 29380 18290 29408 84458
rect 29472 53718 29500 112406
rect 30012 103692 30064 103698
rect 30012 103634 30064 103640
rect 29644 86624 29696 86630
rect 29644 86566 29696 86572
rect 29656 86329 29684 86566
rect 29642 86320 29698 86329
rect 29642 86255 29698 86264
rect 29552 83428 29604 83434
rect 29552 83370 29604 83376
rect 29564 83026 29592 83370
rect 29552 83020 29604 83026
rect 29552 82962 29604 82968
rect 29552 75540 29604 75546
rect 29552 75482 29604 75488
rect 29460 53712 29512 53718
rect 29460 53654 29512 53660
rect 29564 48822 29592 75482
rect 29656 75410 29684 86255
rect 29828 82340 29880 82346
rect 29828 82282 29880 82288
rect 29644 75404 29696 75410
rect 29644 75346 29696 75352
rect 29644 59220 29696 59226
rect 29644 59162 29696 59168
rect 29656 58002 29684 59162
rect 29736 58404 29788 58410
rect 29736 58346 29788 58352
rect 29644 57996 29696 58002
rect 29644 57938 29696 57944
rect 29644 54732 29696 54738
rect 29644 54674 29696 54680
rect 29552 48816 29604 48822
rect 29552 48758 29604 48764
rect 29656 40390 29684 54674
rect 29644 40384 29696 40390
rect 29644 40326 29696 40332
rect 29552 20528 29604 20534
rect 29552 20470 29604 20476
rect 29460 20256 29512 20262
rect 29460 20198 29512 20204
rect 29472 19718 29500 20198
rect 29460 19712 29512 19718
rect 29460 19654 29512 19660
rect 29460 19236 29512 19242
rect 29460 19178 29512 19184
rect 29368 18284 29420 18290
rect 29368 18226 29420 18232
rect 29472 18154 29500 19178
rect 29564 18465 29592 20470
rect 29644 19984 29696 19990
rect 29644 19926 29696 19932
rect 29656 19854 29684 19926
rect 29748 19922 29776 58346
rect 29736 19916 29788 19922
rect 29736 19858 29788 19864
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29550 18456 29606 18465
rect 29550 18391 29606 18400
rect 29552 18352 29604 18358
rect 29552 18294 29604 18300
rect 29460 18148 29512 18154
rect 29460 18090 29512 18096
rect 29368 17876 29420 17882
rect 29368 17818 29420 17824
rect 29276 17264 29328 17270
rect 29276 17206 29328 17212
rect 29276 16788 29328 16794
rect 29276 16730 29328 16736
rect 29184 14952 29236 14958
rect 29184 14894 29236 14900
rect 29288 14482 29316 16730
rect 29380 14550 29408 17818
rect 29460 17196 29512 17202
rect 29460 17138 29512 17144
rect 29472 15366 29500 17138
rect 29460 15360 29512 15366
rect 29460 15302 29512 15308
rect 29368 14544 29420 14550
rect 29368 14486 29420 14492
rect 29276 14476 29328 14482
rect 29196 14414 29224 14445
rect 29276 14418 29328 14424
rect 29184 14408 29236 14414
rect 29182 14376 29184 14385
rect 29236 14376 29238 14385
rect 29182 14311 29238 14320
rect 29196 14278 29224 14311
rect 29184 14272 29236 14278
rect 29184 14214 29236 14220
rect 29564 13530 29592 18294
rect 29656 18222 29684 19790
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29644 18216 29696 18222
rect 29644 18158 29696 18164
rect 29656 17542 29684 18158
rect 29644 17536 29696 17542
rect 29644 17478 29696 17484
rect 29656 17134 29684 17478
rect 29644 17128 29696 17134
rect 29644 17070 29696 17076
rect 29644 16448 29696 16454
rect 29748 16436 29776 19654
rect 29696 16408 29776 16436
rect 29644 16390 29696 16396
rect 29656 16250 29684 16390
rect 29644 16244 29696 16250
rect 29644 16186 29696 16192
rect 29840 15570 29868 82282
rect 29920 76900 29972 76906
rect 29920 76842 29972 76848
rect 29932 75410 29960 76842
rect 29920 75404 29972 75410
rect 29920 75346 29972 75352
rect 29920 67856 29972 67862
rect 29920 67798 29972 67804
rect 29932 58342 29960 67798
rect 29920 58336 29972 58342
rect 29920 58278 29972 58284
rect 29920 26988 29972 26994
rect 29920 26930 29972 26936
rect 29932 24410 29960 26930
rect 29920 24404 29972 24410
rect 29920 24346 29972 24352
rect 29920 18828 29972 18834
rect 29920 18770 29972 18776
rect 29932 16250 29960 18770
rect 29920 16244 29972 16250
rect 29920 16186 29972 16192
rect 29920 15972 29972 15978
rect 29920 15914 29972 15920
rect 29828 15564 29880 15570
rect 29828 15506 29880 15512
rect 29736 15360 29788 15366
rect 29736 15302 29788 15308
rect 29748 14793 29776 15302
rect 29734 14784 29790 14793
rect 29734 14719 29790 14728
rect 29736 14544 29788 14550
rect 29736 14486 29788 14492
rect 29748 13870 29776 14486
rect 29932 14482 29960 15914
rect 29920 14476 29972 14482
rect 29920 14418 29972 14424
rect 29736 13864 29788 13870
rect 29736 13806 29788 13812
rect 29184 13524 29236 13530
rect 29184 13466 29236 13472
rect 29552 13524 29604 13530
rect 29552 13466 29604 13472
rect 29092 13388 29144 13394
rect 29092 13330 29144 13336
rect 29000 6452 29052 6458
rect 29000 6394 29052 6400
rect 28632 6112 28684 6118
rect 28632 6054 28684 6060
rect 28356 5160 28408 5166
rect 28356 5102 28408 5108
rect 28908 4072 28960 4078
rect 28908 4014 28960 4020
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 28540 3392 28592 3398
rect 28540 3334 28592 3340
rect 28552 3194 28580 3334
rect 28630 3224 28686 3233
rect 28540 3188 28592 3194
rect 28630 3159 28632 3168
rect 28540 3130 28592 3136
rect 28684 3159 28686 3168
rect 28632 3130 28684 3136
rect 28828 3074 28856 3470
rect 28552 3046 28856 3074
rect 28552 2990 28580 3046
rect 28540 2984 28592 2990
rect 28540 2926 28592 2932
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 28172 2372 28224 2378
rect 28172 2314 28224 2320
rect 28368 800 28396 2790
rect 28920 2774 28948 4014
rect 29000 3120 29052 3126
rect 28998 3088 29000 3097
rect 29052 3088 29054 3097
rect 28998 3023 29054 3032
rect 29196 2961 29224 13466
rect 30024 11150 30052 103634
rect 30380 83972 30432 83978
rect 30380 83914 30432 83920
rect 30104 68400 30156 68406
rect 30104 68342 30156 68348
rect 30116 59226 30144 68342
rect 30196 67584 30248 67590
rect 30196 67526 30248 67532
rect 30104 59220 30156 59226
rect 30104 59162 30156 59168
rect 30104 58948 30156 58954
rect 30104 58890 30156 58896
rect 30116 58138 30144 58890
rect 30208 58138 30236 67526
rect 30288 66020 30340 66026
rect 30288 65962 30340 65968
rect 30104 58132 30156 58138
rect 30104 58074 30156 58080
rect 30196 58132 30248 58138
rect 30196 58074 30248 58080
rect 30300 58070 30328 65962
rect 30288 58064 30340 58070
rect 30288 58006 30340 58012
rect 30288 45892 30340 45898
rect 30288 45834 30340 45840
rect 30300 23322 30328 45834
rect 30288 23316 30340 23322
rect 30288 23258 30340 23264
rect 30392 22030 30420 83914
rect 30484 57934 30512 116690
rect 30576 113966 30604 116844
rect 30668 114918 30696 117014
rect 30656 114912 30708 114918
rect 30656 114854 30708 114860
rect 30656 114504 30708 114510
rect 30656 114446 30708 114452
rect 30564 113960 30616 113966
rect 30564 113902 30616 113908
rect 30668 113082 30696 114446
rect 30748 114436 30800 114442
rect 30748 114378 30800 114384
rect 30656 113076 30708 113082
rect 30656 113018 30708 113024
rect 30760 113014 30788 114378
rect 30852 113490 30880 119200
rect 30932 117088 30984 117094
rect 30932 117030 30984 117036
rect 30944 116278 30972 117030
rect 31036 116872 31064 119200
rect 31208 117088 31260 117094
rect 31208 117030 31260 117036
rect 31220 116890 31248 117030
rect 31208 116884 31260 116890
rect 31036 116844 31156 116872
rect 31024 116748 31076 116754
rect 31024 116690 31076 116696
rect 30932 116272 30984 116278
rect 30932 116214 30984 116220
rect 30930 116104 30986 116113
rect 30930 116039 30932 116048
rect 30984 116039 30986 116048
rect 30932 116010 30984 116016
rect 30932 115660 30984 115666
rect 30932 115602 30984 115608
rect 30944 113626 30972 115602
rect 30932 113620 30984 113626
rect 30932 113562 30984 113568
rect 30840 113484 30892 113490
rect 30840 113426 30892 113432
rect 30748 113008 30800 113014
rect 30748 112950 30800 112956
rect 30564 109064 30616 109070
rect 30564 109006 30616 109012
rect 30472 57928 30524 57934
rect 30472 57870 30524 57876
rect 30576 22114 30604 109006
rect 30656 104168 30708 104174
rect 30656 104110 30708 104116
rect 30668 103086 30696 104110
rect 30656 103080 30708 103086
rect 30656 103022 30708 103028
rect 30668 102202 30696 103022
rect 30656 102196 30708 102202
rect 30656 102138 30708 102144
rect 30748 95668 30800 95674
rect 30748 95610 30800 95616
rect 30760 92886 30788 95610
rect 30840 93356 30892 93362
rect 30840 93298 30892 93304
rect 30748 92880 30800 92886
rect 30748 92822 30800 92828
rect 30748 88324 30800 88330
rect 30748 88266 30800 88272
rect 30760 83026 30788 88266
rect 30852 84114 30880 93298
rect 30932 86896 30984 86902
rect 30932 86838 30984 86844
rect 30840 84108 30892 84114
rect 30840 84050 30892 84056
rect 30656 83020 30708 83026
rect 30656 82962 30708 82968
rect 30748 83020 30800 83026
rect 30748 82962 30800 82968
rect 30484 22086 30604 22114
rect 30380 22024 30432 22030
rect 30380 21966 30432 21972
rect 30484 21026 30512 22086
rect 30564 22024 30616 22030
rect 30564 21966 30616 21972
rect 30392 20998 30512 21026
rect 30392 20890 30420 20998
rect 30208 20862 30420 20890
rect 30472 20868 30524 20874
rect 30104 19304 30156 19310
rect 30104 19246 30156 19252
rect 30116 18630 30144 19246
rect 30208 18834 30236 20862
rect 30472 20810 30524 20816
rect 30288 20800 30340 20806
rect 30288 20742 30340 20748
rect 30196 18828 30248 18834
rect 30196 18770 30248 18776
rect 30104 18624 30156 18630
rect 30104 18566 30156 18572
rect 30194 17640 30250 17649
rect 30194 17575 30250 17584
rect 30208 16182 30236 17575
rect 30300 17066 30328 20742
rect 30380 20256 30432 20262
rect 30380 20198 30432 20204
rect 30392 17814 30420 20198
rect 30484 18902 30512 20810
rect 30576 19825 30604 21966
rect 30562 19816 30618 19825
rect 30562 19751 30618 19760
rect 30564 19712 30616 19718
rect 30564 19654 30616 19660
rect 30472 18896 30524 18902
rect 30472 18838 30524 18844
rect 30472 18760 30524 18766
rect 30472 18702 30524 18708
rect 30380 17808 30432 17814
rect 30380 17750 30432 17756
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30288 17060 30340 17066
rect 30288 17002 30340 17008
rect 30392 16658 30420 17070
rect 30380 16652 30432 16658
rect 30380 16594 30432 16600
rect 30286 16552 30342 16561
rect 30286 16487 30342 16496
rect 30196 16176 30248 16182
rect 30196 16118 30248 16124
rect 30208 15570 30236 16118
rect 30196 15564 30248 15570
rect 30196 15506 30248 15512
rect 30208 14958 30236 15506
rect 30196 14952 30248 14958
rect 30196 14894 30248 14900
rect 30300 14414 30328 16487
rect 30484 15994 30512 18702
rect 30576 16726 30604 19654
rect 30564 16720 30616 16726
rect 30564 16662 30616 16668
rect 30668 16046 30696 82962
rect 30840 81320 30892 81326
rect 30840 81262 30892 81268
rect 30852 80850 30880 81262
rect 30840 80844 30892 80850
rect 30840 80786 30892 80792
rect 30748 79892 30800 79898
rect 30748 79834 30800 79840
rect 30760 71058 30788 79834
rect 30840 78464 30892 78470
rect 30840 78406 30892 78412
rect 30852 71670 30880 78406
rect 30944 76906 30972 86838
rect 30932 76900 30984 76906
rect 30932 76842 30984 76848
rect 31036 76634 31064 116690
rect 31128 113490 31156 116844
rect 31208 116826 31260 116832
rect 31208 116000 31260 116006
rect 31208 115942 31260 115948
rect 31220 114102 31248 115942
rect 31208 114096 31260 114102
rect 31208 114038 31260 114044
rect 31116 113484 31168 113490
rect 31116 113426 31168 113432
rect 31312 112878 31340 119200
rect 31392 117156 31444 117162
rect 31392 117098 31444 117104
rect 31404 116686 31432 117098
rect 31392 116680 31444 116686
rect 31392 116622 31444 116628
rect 31496 116498 31524 119200
rect 31772 116890 31800 119200
rect 31760 116884 31812 116890
rect 31760 116826 31812 116832
rect 31852 116748 31904 116754
rect 31852 116690 31904 116696
rect 31496 116470 31616 116498
rect 31484 116272 31536 116278
rect 31484 116214 31536 116220
rect 31392 116204 31444 116210
rect 31392 116146 31444 116152
rect 31404 115258 31432 116146
rect 31496 115258 31524 116214
rect 31588 116210 31616 116470
rect 31576 116204 31628 116210
rect 31576 116146 31628 116152
rect 31668 116136 31720 116142
rect 31760 116136 31812 116142
rect 31668 116078 31720 116084
rect 31758 116104 31760 116113
rect 31812 116104 31814 116113
rect 31576 115456 31628 115462
rect 31576 115398 31628 115404
rect 31392 115252 31444 115258
rect 31392 115194 31444 115200
rect 31484 115252 31536 115258
rect 31484 115194 31536 115200
rect 31588 115122 31616 115398
rect 31576 115116 31628 115122
rect 31576 115058 31628 115064
rect 31392 114912 31444 114918
rect 31392 114854 31444 114860
rect 31484 114912 31536 114918
rect 31484 114854 31536 114860
rect 31404 113966 31432 114854
rect 31496 114578 31524 114854
rect 31680 114714 31708 116078
rect 31758 116039 31814 116048
rect 31760 115660 31812 115666
rect 31760 115602 31812 115608
rect 31668 114708 31720 114714
rect 31668 114650 31720 114656
rect 31484 114572 31536 114578
rect 31484 114514 31536 114520
rect 31392 113960 31444 113966
rect 31392 113902 31444 113908
rect 31772 113898 31800 115602
rect 31760 113892 31812 113898
rect 31760 113834 31812 113840
rect 31300 112872 31352 112878
rect 31864 112826 31892 116690
rect 31956 115054 31984 119200
rect 32232 116906 32260 119200
rect 32140 116878 32260 116906
rect 32312 116884 32364 116890
rect 32036 116204 32088 116210
rect 32036 116146 32088 116152
rect 31944 115048 31996 115054
rect 31944 114990 31996 114996
rect 32048 114170 32076 116146
rect 32140 115190 32168 116878
rect 32312 116826 32364 116832
rect 32220 116272 32272 116278
rect 32220 116214 32272 116220
rect 32128 115184 32180 115190
rect 32128 115126 32180 115132
rect 32128 114436 32180 114442
rect 32128 114378 32180 114384
rect 32036 114164 32088 114170
rect 32036 114106 32088 114112
rect 32140 113082 32168 114378
rect 32128 113076 32180 113082
rect 32128 113018 32180 113024
rect 32232 112878 32260 116214
rect 32324 112878 32352 116826
rect 32404 116340 32456 116346
rect 32404 116282 32456 116288
rect 32416 115977 32444 116282
rect 32402 115968 32458 115977
rect 32402 115903 32458 115912
rect 32404 115048 32456 115054
rect 32404 114990 32456 114996
rect 31300 112814 31352 112820
rect 31772 112798 31892 112826
rect 32220 112872 32272 112878
rect 32220 112814 32272 112820
rect 32312 112872 32364 112878
rect 32312 112814 32364 112820
rect 31116 107432 31168 107438
rect 31116 107374 31168 107380
rect 31024 76628 31076 76634
rect 31024 76570 31076 76576
rect 30840 71664 30892 71670
rect 30840 71606 30892 71612
rect 31024 71664 31076 71670
rect 31024 71606 31076 71612
rect 30840 71460 30892 71466
rect 30840 71402 30892 71408
rect 30748 71052 30800 71058
rect 30748 70994 30800 71000
rect 30748 59492 30800 59498
rect 30748 59434 30800 59440
rect 30760 19922 30788 59434
rect 30748 19916 30800 19922
rect 30748 19858 30800 19864
rect 30746 19816 30802 19825
rect 30746 19751 30802 19760
rect 30760 17746 30788 19751
rect 30748 17740 30800 17746
rect 30748 17682 30800 17688
rect 30748 17536 30800 17542
rect 30748 17478 30800 17484
rect 30392 15966 30512 15994
rect 30656 16040 30708 16046
rect 30656 15982 30708 15988
rect 30392 14929 30420 15966
rect 30472 15904 30524 15910
rect 30472 15846 30524 15852
rect 30378 14920 30434 14929
rect 30484 14890 30512 15846
rect 30378 14855 30434 14864
rect 30472 14884 30524 14890
rect 30288 14408 30340 14414
rect 30288 14350 30340 14356
rect 30288 13864 30340 13870
rect 30288 13806 30340 13812
rect 30300 12986 30328 13806
rect 30288 12980 30340 12986
rect 30288 12922 30340 12928
rect 30392 11218 30420 14855
rect 30472 14826 30524 14832
rect 30380 11212 30432 11218
rect 30380 11154 30432 11160
rect 30012 11144 30064 11150
rect 30012 11086 30064 11092
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 30196 8968 30248 8974
rect 30196 8910 30248 8916
rect 29552 7948 29604 7954
rect 29604 7908 29776 7936
rect 29552 7890 29604 7896
rect 29276 4480 29328 4486
rect 29276 4422 29328 4428
rect 29288 4010 29316 4422
rect 29552 4072 29604 4078
rect 29552 4014 29604 4020
rect 29644 4072 29696 4078
rect 29644 4014 29696 4020
rect 29276 4004 29328 4010
rect 29276 3946 29328 3952
rect 29460 3936 29512 3942
rect 29366 3904 29422 3913
rect 29460 3878 29512 3884
rect 29366 3839 29422 3848
rect 29380 3670 29408 3839
rect 29368 3664 29420 3670
rect 29368 3606 29420 3612
rect 29472 3534 29500 3878
rect 29460 3528 29512 3534
rect 29460 3470 29512 3476
rect 29368 3392 29420 3398
rect 29368 3334 29420 3340
rect 29182 2952 29238 2961
rect 29182 2887 29238 2896
rect 28736 2746 28948 2774
rect 28736 800 28764 2746
rect 29000 1556 29052 1562
rect 29000 1498 29052 1504
rect 29012 800 29040 1498
rect 29380 800 29408 3334
rect 29564 1562 29592 4014
rect 29552 1556 29604 1562
rect 29552 1498 29604 1504
rect 29656 800 29684 4014
rect 29748 3058 29776 7908
rect 30208 3670 30236 8910
rect 30300 5234 30328 11086
rect 30760 5370 30788 17478
rect 30852 15570 30880 71402
rect 31036 64530 31064 71606
rect 31024 64524 31076 64530
rect 31024 64466 31076 64472
rect 31024 58880 31076 58886
rect 31024 58822 31076 58828
rect 30932 41472 30984 41478
rect 30932 41414 30984 41420
rect 30944 20534 30972 41414
rect 31036 20942 31064 58822
rect 31024 20936 31076 20942
rect 31024 20878 31076 20884
rect 31024 20800 31076 20806
rect 31024 20742 31076 20748
rect 30932 20528 30984 20534
rect 30932 20470 30984 20476
rect 30930 20088 30986 20097
rect 30930 20023 30986 20032
rect 30944 19922 30972 20023
rect 30932 19916 30984 19922
rect 30932 19858 30984 19864
rect 31036 19802 31064 20742
rect 30944 19774 31064 19802
rect 30944 18630 30972 19774
rect 31024 19712 31076 19718
rect 31024 19654 31076 19660
rect 30932 18624 30984 18630
rect 30932 18566 30984 18572
rect 30932 18148 30984 18154
rect 30932 18090 30984 18096
rect 30944 16998 30972 18090
rect 30932 16992 30984 16998
rect 30932 16934 30984 16940
rect 31036 16794 31064 19654
rect 31024 16788 31076 16794
rect 31024 16730 31076 16736
rect 30840 15564 30892 15570
rect 30840 15506 30892 15512
rect 30932 11212 30984 11218
rect 30932 11154 30984 11160
rect 30748 5364 30800 5370
rect 30748 5306 30800 5312
rect 30288 5228 30340 5234
rect 30288 5170 30340 5176
rect 30944 5098 30972 11154
rect 31036 5302 31064 16730
rect 31128 11150 31156 107374
rect 31208 104100 31260 104106
rect 31208 104042 31260 104048
rect 31220 82074 31248 104042
rect 31576 102944 31628 102950
rect 31576 102886 31628 102892
rect 31300 102196 31352 102202
rect 31300 102138 31352 102144
rect 31208 82068 31260 82074
rect 31208 82010 31260 82016
rect 31208 80844 31260 80850
rect 31208 80786 31260 80792
rect 31220 80442 31248 80786
rect 31208 80436 31260 80442
rect 31208 80378 31260 80384
rect 31208 71392 31260 71398
rect 31208 71334 31260 71340
rect 31220 71194 31248 71334
rect 31208 71188 31260 71194
rect 31208 71130 31260 71136
rect 31208 67312 31260 67318
rect 31208 67254 31260 67260
rect 31220 58682 31248 67254
rect 31208 58676 31260 58682
rect 31208 58618 31260 58624
rect 31208 20528 31260 20534
rect 31208 20470 31260 20476
rect 31220 17542 31248 20470
rect 31208 17536 31260 17542
rect 31208 17478 31260 17484
rect 31208 17128 31260 17134
rect 31208 17070 31260 17076
rect 31220 16794 31248 17070
rect 31208 16788 31260 16794
rect 31208 16730 31260 16736
rect 31208 16584 31260 16590
rect 31208 16526 31260 16532
rect 31220 16182 31248 16526
rect 31208 16176 31260 16182
rect 31208 16118 31260 16124
rect 31208 16040 31260 16046
rect 31208 15982 31260 15988
rect 31116 11144 31168 11150
rect 31116 11086 31168 11092
rect 31128 6866 31156 11086
rect 31116 6860 31168 6866
rect 31116 6802 31168 6808
rect 31024 5296 31076 5302
rect 31024 5238 31076 5244
rect 30932 5092 30984 5098
rect 30932 5034 30984 5040
rect 30748 4072 30800 4078
rect 30748 4014 30800 4020
rect 30564 3936 30616 3942
rect 30484 3896 30564 3924
rect 30196 3664 30248 3670
rect 30010 3632 30066 3641
rect 30196 3606 30248 3612
rect 30010 3567 30066 3576
rect 30024 3466 30052 3567
rect 30012 3460 30064 3466
rect 30380 3460 30432 3466
rect 30012 3402 30064 3408
rect 30300 3420 30380 3448
rect 29736 3052 29788 3058
rect 29736 2994 29788 3000
rect 30012 2508 30064 2514
rect 30012 2450 30064 2456
rect 29736 2440 29788 2446
rect 29736 2382 29788 2388
rect 29748 1970 29776 2382
rect 29736 1964 29788 1970
rect 29736 1906 29788 1912
rect 30024 800 30052 2450
rect 30300 800 30328 3420
rect 30380 3402 30432 3408
rect 30484 3097 30512 3896
rect 30564 3878 30616 3884
rect 30656 3188 30708 3194
rect 30656 3130 30708 3136
rect 30668 3097 30696 3130
rect 30470 3088 30526 3097
rect 30470 3023 30526 3032
rect 30654 3088 30710 3097
rect 30654 3023 30710 3032
rect 30760 2774 30788 4014
rect 31022 3904 31078 3913
rect 31022 3839 31078 3848
rect 31036 3602 31064 3839
rect 31114 3632 31170 3641
rect 31024 3596 31076 3602
rect 31114 3567 31116 3576
rect 31024 3538 31076 3544
rect 31168 3567 31170 3576
rect 31116 3538 31168 3544
rect 30840 3528 30892 3534
rect 30840 3470 30892 3476
rect 30852 3194 30880 3470
rect 30840 3188 30892 3194
rect 30840 3130 30892 3136
rect 31220 2990 31248 15982
rect 31312 11354 31340 102138
rect 31392 101312 31444 101318
rect 31392 101254 31444 101260
rect 31404 71602 31432 101254
rect 31484 95464 31536 95470
rect 31484 95406 31536 95412
rect 31392 71596 31444 71602
rect 31392 71538 31444 71544
rect 31392 71052 31444 71058
rect 31392 70994 31444 71000
rect 31404 70582 31432 70994
rect 31392 70576 31444 70582
rect 31392 70518 31444 70524
rect 31404 70446 31432 70518
rect 31392 70440 31444 70446
rect 31392 70382 31444 70388
rect 31392 66564 31444 66570
rect 31392 66506 31444 66512
rect 31404 58614 31432 66506
rect 31496 59090 31524 95406
rect 31588 81326 31616 102886
rect 31772 91186 31800 112798
rect 31852 112736 31904 112742
rect 31852 112678 31904 112684
rect 31760 91180 31812 91186
rect 31760 91122 31812 91128
rect 31668 91112 31720 91118
rect 31668 91054 31720 91060
rect 31576 81320 31628 81326
rect 31576 81262 31628 81268
rect 31576 81184 31628 81190
rect 31576 81126 31628 81132
rect 31484 59084 31536 59090
rect 31484 59026 31536 59032
rect 31392 58608 31444 58614
rect 31392 58550 31444 58556
rect 31392 26920 31444 26926
rect 31392 26862 31444 26868
rect 31404 21690 31432 26862
rect 31482 23080 31538 23089
rect 31482 23015 31484 23024
rect 31536 23015 31538 23024
rect 31484 22986 31536 22992
rect 31392 21684 31444 21690
rect 31392 21626 31444 21632
rect 31484 21344 31536 21350
rect 31484 21286 31536 21292
rect 31392 21004 31444 21010
rect 31392 20946 31444 20952
rect 31404 20874 31432 20946
rect 31392 20868 31444 20874
rect 31392 20810 31444 20816
rect 31404 20398 31432 20810
rect 31392 20392 31444 20398
rect 31392 20334 31444 20340
rect 31404 20262 31432 20334
rect 31392 20256 31444 20262
rect 31392 20198 31444 20204
rect 31404 19922 31432 20198
rect 31392 19916 31444 19922
rect 31392 19858 31444 19864
rect 31392 19168 31444 19174
rect 31392 19110 31444 19116
rect 31404 18834 31432 19110
rect 31392 18828 31444 18834
rect 31392 18770 31444 18776
rect 31392 18624 31444 18630
rect 31392 18566 31444 18572
rect 31404 17762 31432 18566
rect 31496 18086 31524 21286
rect 31484 18080 31536 18086
rect 31484 18022 31536 18028
rect 31404 17734 31524 17762
rect 31392 17604 31444 17610
rect 31392 17546 31444 17552
rect 31404 15638 31432 17546
rect 31496 17338 31524 17734
rect 31484 17332 31536 17338
rect 31484 17274 31536 17280
rect 31392 15632 31444 15638
rect 31392 15574 31444 15580
rect 31390 15464 31446 15473
rect 31390 15399 31392 15408
rect 31444 15399 31446 15408
rect 31392 15370 31444 15376
rect 31496 12434 31524 17274
rect 31588 16658 31616 81126
rect 31680 70446 31708 91054
rect 31760 85876 31812 85882
rect 31760 85818 31812 85824
rect 31772 83026 31800 85818
rect 31760 83020 31812 83026
rect 31760 82962 31812 82968
rect 31772 82278 31800 82962
rect 31760 82272 31812 82278
rect 31760 82214 31812 82220
rect 31772 81938 31800 82214
rect 31760 81932 31812 81938
rect 31760 81874 31812 81880
rect 31760 81728 31812 81734
rect 31760 81670 31812 81676
rect 31772 81326 31800 81670
rect 31760 81320 31812 81326
rect 31760 81262 31812 81268
rect 31760 81184 31812 81190
rect 31760 81126 31812 81132
rect 31772 77994 31800 81126
rect 31760 77988 31812 77994
rect 31760 77930 31812 77936
rect 31760 71596 31812 71602
rect 31760 71538 31812 71544
rect 31772 70582 31800 71538
rect 31760 70576 31812 70582
rect 31760 70518 31812 70524
rect 31668 70440 31720 70446
rect 31668 70382 31720 70388
rect 31760 65612 31812 65618
rect 31760 65554 31812 65560
rect 31668 64524 31720 64530
rect 31668 64466 31720 64472
rect 31680 62830 31708 64466
rect 31668 62824 31720 62830
rect 31668 62766 31720 62772
rect 31668 59968 31720 59974
rect 31668 59910 31720 59916
rect 31680 21078 31708 59910
rect 31772 59566 31800 65554
rect 31760 59560 31812 59566
rect 31760 59502 31812 59508
rect 31760 55072 31812 55078
rect 31760 55014 31812 55020
rect 31772 21486 31800 55014
rect 31864 27130 31892 112678
rect 31944 110016 31996 110022
rect 31944 109958 31996 109964
rect 31956 59090 31984 109958
rect 32220 96484 32272 96490
rect 32220 96426 32272 96432
rect 32036 94852 32088 94858
rect 32036 94794 32088 94800
rect 32048 82550 32076 94794
rect 32128 86760 32180 86766
rect 32128 86702 32180 86708
rect 32140 85202 32168 86702
rect 32128 85196 32180 85202
rect 32128 85138 32180 85144
rect 32140 84590 32168 85138
rect 32128 84584 32180 84590
rect 32128 84526 32180 84532
rect 32140 84250 32168 84526
rect 32128 84244 32180 84250
rect 32128 84186 32180 84192
rect 32128 83360 32180 83366
rect 32128 83302 32180 83308
rect 32140 83094 32168 83302
rect 32128 83088 32180 83094
rect 32128 83030 32180 83036
rect 32036 82544 32088 82550
rect 32036 82486 32088 82492
rect 32140 82482 32168 83030
rect 32128 82476 32180 82482
rect 32128 82418 32180 82424
rect 32140 82006 32168 82418
rect 32128 82000 32180 82006
rect 32128 81942 32180 81948
rect 32036 81320 32088 81326
rect 32140 81308 32168 81942
rect 32088 81280 32168 81308
rect 32036 81262 32088 81268
rect 32036 80776 32088 80782
rect 32036 80718 32088 80724
rect 32048 80238 32076 80718
rect 32036 80232 32088 80238
rect 32036 80174 32088 80180
rect 32036 75540 32088 75546
rect 32036 75482 32088 75488
rect 32048 71058 32076 75482
rect 32128 71664 32180 71670
rect 32128 71606 32180 71612
rect 32140 71534 32168 71606
rect 32128 71528 32180 71534
rect 32128 71470 32180 71476
rect 32140 71126 32168 71470
rect 32128 71120 32180 71126
rect 32128 71062 32180 71068
rect 32036 71052 32088 71058
rect 32036 70994 32088 71000
rect 32128 70984 32180 70990
rect 32128 70926 32180 70932
rect 32036 70916 32088 70922
rect 32036 70858 32088 70864
rect 32048 70446 32076 70858
rect 32036 70440 32088 70446
rect 32036 70382 32088 70388
rect 32036 65544 32088 65550
rect 32036 65486 32088 65492
rect 31944 59084 31996 59090
rect 31944 59026 31996 59032
rect 32048 58018 32076 65486
rect 31956 57990 32076 58018
rect 31956 56710 31984 57990
rect 32036 57928 32088 57934
rect 32036 57870 32088 57876
rect 31944 56704 31996 56710
rect 31944 56646 31996 56652
rect 31944 55684 31996 55690
rect 31944 55626 31996 55632
rect 31956 41414 31984 55626
rect 32048 54262 32076 57870
rect 32140 54330 32168 70926
rect 32232 55214 32260 96426
rect 32416 95674 32444 114990
rect 32508 113966 32536 119200
rect 32588 116204 32640 116210
rect 32588 116146 32640 116152
rect 32496 113960 32548 113966
rect 32496 113902 32548 113908
rect 32600 113626 32628 116146
rect 32692 114578 32720 119200
rect 32772 116544 32824 116550
rect 32772 116486 32824 116492
rect 32784 116346 32812 116486
rect 32772 116340 32824 116346
rect 32772 116282 32824 116288
rect 32864 116272 32916 116278
rect 32864 116214 32916 116220
rect 32772 116000 32824 116006
rect 32772 115942 32824 115948
rect 32680 114572 32732 114578
rect 32680 114514 32732 114520
rect 32588 113620 32640 113626
rect 32588 113562 32640 113568
rect 32784 112742 32812 115942
rect 32876 114170 32904 116214
rect 32864 114164 32916 114170
rect 32864 114106 32916 114112
rect 32968 113966 32996 119200
rect 33048 117088 33100 117094
rect 33048 117030 33100 117036
rect 33060 116006 33088 117030
rect 33048 116000 33100 116006
rect 33048 115942 33100 115948
rect 33048 114572 33100 114578
rect 33048 114514 33100 114520
rect 32956 113960 33008 113966
rect 32956 113902 33008 113908
rect 32772 112736 32824 112742
rect 32772 112678 32824 112684
rect 32588 110560 32640 110566
rect 32588 110502 32640 110508
rect 32496 107908 32548 107914
rect 32496 107850 32548 107856
rect 32404 95668 32456 95674
rect 32404 95610 32456 95616
rect 32404 94512 32456 94518
rect 32404 94454 32456 94460
rect 32312 86624 32364 86630
rect 32312 86566 32364 86572
rect 32324 85882 32352 86566
rect 32312 85876 32364 85882
rect 32312 85818 32364 85824
rect 32324 85746 32352 85818
rect 32312 85740 32364 85746
rect 32312 85682 32364 85688
rect 32416 85678 32444 94454
rect 32404 85672 32456 85678
rect 32404 85614 32456 85620
rect 32404 85536 32456 85542
rect 32324 85484 32404 85490
rect 32324 85478 32456 85484
rect 32324 85462 32444 85478
rect 32324 83502 32352 85462
rect 32508 84590 32536 107850
rect 32496 84584 32548 84590
rect 32496 84526 32548 84532
rect 32496 84244 32548 84250
rect 32496 84186 32548 84192
rect 32404 84176 32456 84182
rect 32404 84118 32456 84124
rect 32416 83502 32444 84118
rect 32312 83496 32364 83502
rect 32312 83438 32364 83444
rect 32404 83496 32456 83502
rect 32404 83438 32456 83444
rect 32312 82408 32364 82414
rect 32312 82350 32364 82356
rect 32324 81462 32352 82350
rect 32404 82272 32456 82278
rect 32404 82214 32456 82220
rect 32312 81456 32364 81462
rect 32312 81398 32364 81404
rect 32416 81326 32444 82214
rect 32404 81320 32456 81326
rect 32404 81262 32456 81268
rect 32508 78062 32536 84186
rect 32496 78056 32548 78062
rect 32496 77998 32548 78004
rect 32496 77920 32548 77926
rect 32496 77862 32548 77868
rect 32312 75268 32364 75274
rect 32312 75210 32364 75216
rect 32220 55208 32272 55214
rect 32220 55150 32272 55156
rect 32128 54324 32180 54330
rect 32128 54266 32180 54272
rect 32036 54256 32088 54262
rect 32036 54198 32088 54204
rect 32128 50244 32180 50250
rect 32128 50186 32180 50192
rect 32140 49842 32168 50186
rect 32128 49836 32180 49842
rect 32128 49778 32180 49784
rect 32220 49768 32272 49774
rect 32220 49710 32272 49716
rect 32036 49632 32088 49638
rect 32036 49574 32088 49580
rect 32048 48754 32076 49574
rect 32036 48748 32088 48754
rect 32036 48690 32088 48696
rect 31956 41386 32076 41414
rect 31852 27124 31904 27130
rect 31852 27066 31904 27072
rect 31864 24342 31892 27066
rect 31852 24336 31904 24342
rect 31852 24278 31904 24284
rect 31944 24064 31996 24070
rect 31944 24006 31996 24012
rect 31852 23860 31904 23866
rect 31852 23802 31904 23808
rect 31864 22710 31892 23802
rect 31852 22704 31904 22710
rect 31852 22646 31904 22652
rect 31852 22568 31904 22574
rect 31852 22510 31904 22516
rect 31760 21480 31812 21486
rect 31760 21422 31812 21428
rect 31760 21344 31812 21350
rect 31760 21286 31812 21292
rect 31668 21072 31720 21078
rect 31668 21014 31720 21020
rect 31772 20924 31800 21286
rect 31680 20896 31800 20924
rect 31680 20466 31708 20896
rect 31760 20800 31812 20806
rect 31760 20742 31812 20748
rect 31668 20460 31720 20466
rect 31668 20402 31720 20408
rect 31668 20256 31720 20262
rect 31668 20198 31720 20204
rect 31680 19786 31708 20198
rect 31668 19780 31720 19786
rect 31668 19722 31720 19728
rect 31668 19440 31720 19446
rect 31668 19382 31720 19388
rect 31576 16652 31628 16658
rect 31576 16594 31628 16600
rect 31680 16046 31708 19382
rect 31772 18970 31800 20742
rect 31864 19310 31892 22510
rect 31956 20398 31984 24006
rect 32048 22574 32076 41386
rect 32232 25906 32260 49710
rect 32324 25974 32352 75210
rect 32404 73160 32456 73166
rect 32404 73102 32456 73108
rect 32416 71534 32444 73102
rect 32508 71602 32536 77862
rect 32496 71596 32548 71602
rect 32496 71538 32548 71544
rect 32404 71528 32456 71534
rect 32404 71470 32456 71476
rect 32404 71120 32456 71126
rect 32404 71062 32456 71068
rect 32416 70446 32444 71062
rect 32404 70440 32456 70446
rect 32404 70382 32456 70388
rect 32404 69488 32456 69494
rect 32404 69430 32456 69436
rect 32416 64938 32444 69430
rect 32404 64932 32456 64938
rect 32404 64874 32456 64880
rect 32508 64598 32536 71538
rect 32496 64592 32548 64598
rect 32496 64534 32548 64540
rect 32508 62898 32536 64534
rect 32496 62892 32548 62898
rect 32496 62834 32548 62840
rect 32496 62756 32548 62762
rect 32496 62698 32548 62704
rect 32404 58880 32456 58886
rect 32404 58822 32456 58828
rect 32416 41478 32444 58822
rect 32508 56234 32536 62698
rect 32496 56228 32548 56234
rect 32496 56170 32548 56176
rect 32508 55758 32536 56170
rect 32496 55752 32548 55758
rect 32496 55694 32548 55700
rect 32496 55616 32548 55622
rect 32496 55558 32548 55564
rect 32404 41472 32456 41478
rect 32404 41414 32456 41420
rect 32404 36372 32456 36378
rect 32404 36314 32456 36320
rect 32416 36145 32444 36314
rect 32402 36136 32458 36145
rect 32402 36071 32458 36080
rect 32404 33040 32456 33046
rect 32404 32982 32456 32988
rect 32312 25968 32364 25974
rect 32312 25910 32364 25916
rect 32220 25900 32272 25906
rect 32220 25842 32272 25848
rect 32128 24132 32180 24138
rect 32128 24074 32180 24080
rect 32036 22568 32088 22574
rect 32036 22510 32088 22516
rect 32140 22094 32168 24074
rect 32232 22964 32260 25842
rect 32416 24750 32444 32982
rect 32508 30190 32536 55558
rect 32600 55214 32628 110502
rect 32680 109608 32732 109614
rect 32680 109550 32732 109556
rect 32692 65550 32720 109550
rect 32864 108656 32916 108662
rect 32864 108598 32916 108604
rect 32772 102196 32824 102202
rect 32772 102138 32824 102144
rect 32784 86766 32812 102138
rect 32772 86760 32824 86766
rect 32772 86702 32824 86708
rect 32772 86624 32824 86630
rect 32772 86566 32824 86572
rect 32784 86154 32812 86566
rect 32772 86148 32824 86154
rect 32772 86090 32824 86096
rect 32772 85876 32824 85882
rect 32772 85818 32824 85824
rect 32784 84590 32812 85818
rect 32772 84584 32824 84590
rect 32772 84526 32824 84532
rect 32784 84182 32812 84526
rect 32772 84176 32824 84182
rect 32772 84118 32824 84124
rect 32772 83700 32824 83706
rect 32772 83642 32824 83648
rect 32784 83026 32812 83642
rect 32772 83020 32824 83026
rect 32772 82962 32824 82968
rect 32772 82816 32824 82822
rect 32772 82758 32824 82764
rect 32784 81734 32812 82758
rect 32772 81728 32824 81734
rect 32772 81670 32824 81676
rect 32770 81560 32826 81569
rect 32770 81495 32826 81504
rect 32784 65618 32812 81495
rect 32876 65618 32904 108598
rect 33060 103514 33088 114514
rect 33152 113490 33180 119200
rect 33324 117156 33376 117162
rect 33324 117098 33376 117104
rect 33232 116068 33284 116074
rect 33232 116010 33284 116016
rect 33140 113484 33192 113490
rect 33140 113426 33192 113432
rect 33244 113082 33272 116010
rect 33336 115462 33364 117098
rect 33324 115456 33376 115462
rect 33324 115398 33376 115404
rect 33324 114572 33376 114578
rect 33324 114514 33376 114520
rect 33232 113076 33284 113082
rect 33232 113018 33284 113024
rect 33232 110084 33284 110090
rect 33232 110026 33284 110032
rect 33244 109614 33272 110026
rect 33232 109608 33284 109614
rect 33232 109550 33284 109556
rect 33140 109472 33192 109478
rect 33140 109414 33192 109420
rect 33152 105942 33180 109414
rect 33232 109132 33284 109138
rect 33232 109074 33284 109080
rect 33244 108050 33272 109074
rect 33232 108044 33284 108050
rect 33232 107986 33284 107992
rect 33140 105936 33192 105942
rect 33140 105878 33192 105884
rect 33244 103834 33272 107986
rect 33232 103828 33284 103834
rect 33232 103770 33284 103776
rect 33336 103514 33364 114514
rect 33428 112878 33456 119200
rect 33612 116362 33640 119200
rect 33888 116550 33916 119200
rect 33968 116748 34020 116754
rect 33968 116690 34020 116696
rect 33876 116544 33928 116550
rect 33876 116486 33928 116492
rect 33612 116334 33916 116362
rect 33692 116272 33744 116278
rect 33692 116214 33744 116220
rect 33508 116204 33560 116210
rect 33508 116146 33560 116152
rect 33520 114170 33548 116146
rect 33600 115660 33652 115666
rect 33600 115602 33652 115608
rect 33508 114164 33560 114170
rect 33508 114106 33560 114112
rect 33416 112872 33468 112878
rect 33416 112814 33468 112820
rect 33508 111240 33560 111246
rect 33508 111182 33560 111188
rect 33416 109200 33468 109206
rect 33416 109142 33468 109148
rect 33428 108526 33456 109142
rect 33416 108520 33468 108526
rect 33416 108462 33468 108468
rect 33428 107438 33456 108462
rect 33520 108458 33548 111182
rect 33508 108452 33560 108458
rect 33508 108394 33560 108400
rect 33416 107432 33468 107438
rect 33416 107374 33468 107380
rect 33520 105806 33548 108394
rect 33508 105800 33560 105806
rect 33508 105742 33560 105748
rect 32968 103486 33088 103514
rect 33244 103486 33364 103514
rect 32968 91866 32996 103486
rect 33048 100224 33100 100230
rect 33048 100166 33100 100172
rect 32956 91860 33008 91866
rect 32956 91802 33008 91808
rect 33060 91118 33088 100166
rect 33140 96960 33192 96966
rect 33140 96902 33192 96908
rect 33048 91112 33100 91118
rect 33048 91054 33100 91060
rect 32956 86080 33008 86086
rect 32956 86022 33008 86028
rect 32968 75274 32996 86022
rect 33048 84788 33100 84794
rect 33048 84730 33100 84736
rect 33060 81977 33088 84730
rect 33046 81968 33102 81977
rect 33046 81903 33102 81912
rect 33152 81818 33180 96902
rect 33060 81790 33180 81818
rect 33060 81410 33088 81790
rect 33140 81728 33192 81734
rect 33140 81670 33192 81676
rect 33152 81530 33180 81670
rect 33140 81524 33192 81530
rect 33140 81466 33192 81472
rect 33060 81382 33180 81410
rect 33048 77376 33100 77382
rect 33048 77318 33100 77324
rect 32956 75268 33008 75274
rect 32956 75210 33008 75216
rect 32956 74996 33008 75002
rect 32956 74938 33008 74944
rect 32968 70990 32996 74938
rect 32956 70984 33008 70990
rect 32956 70926 33008 70932
rect 33060 70922 33088 77318
rect 33048 70916 33100 70922
rect 33048 70858 33100 70864
rect 33048 68196 33100 68202
rect 33048 68138 33100 68144
rect 32956 68128 33008 68134
rect 32956 68070 33008 68076
rect 32772 65612 32824 65618
rect 32772 65554 32824 65560
rect 32864 65612 32916 65618
rect 32864 65554 32916 65560
rect 32680 65544 32732 65550
rect 32968 65498 32996 68070
rect 33060 67182 33088 68138
rect 33048 67176 33100 67182
rect 33048 67118 33100 67124
rect 33060 66094 33088 67118
rect 33048 66088 33100 66094
rect 33048 66030 33100 66036
rect 33060 65618 33088 66030
rect 33048 65612 33100 65618
rect 33048 65554 33100 65560
rect 32680 65486 32732 65492
rect 32784 65470 32996 65498
rect 32680 60716 32732 60722
rect 32680 60658 32732 60664
rect 32692 55622 32720 60658
rect 32680 55616 32732 55622
rect 32680 55558 32732 55564
rect 32588 55208 32640 55214
rect 32588 55150 32640 55156
rect 32680 55208 32732 55214
rect 32680 55150 32732 55156
rect 32692 54806 32720 55150
rect 32680 54800 32732 54806
rect 32680 54742 32732 54748
rect 32680 52420 32732 52426
rect 32680 52362 32732 52368
rect 32588 50992 32640 50998
rect 32588 50934 32640 50940
rect 32496 30184 32548 30190
rect 32496 30126 32548 30132
rect 32496 28756 32548 28762
rect 32496 28698 32548 28704
rect 32508 25838 32536 28698
rect 32496 25832 32548 25838
rect 32496 25774 32548 25780
rect 32600 25362 32628 50934
rect 32692 26450 32720 52362
rect 32784 49774 32812 65470
rect 32864 65408 32916 65414
rect 32864 65350 32916 65356
rect 32876 58478 32904 65350
rect 33060 65006 33088 65554
rect 33152 65482 33180 81382
rect 33140 65476 33192 65482
rect 33140 65418 33192 65424
rect 33048 65000 33100 65006
rect 33048 64942 33100 64948
rect 32956 64932 33008 64938
rect 32956 64874 33008 64880
rect 32864 58472 32916 58478
rect 32864 58414 32916 58420
rect 32864 55752 32916 55758
rect 32864 55694 32916 55700
rect 32876 55282 32904 55694
rect 32864 55276 32916 55282
rect 32864 55218 32916 55224
rect 32876 55146 32904 55218
rect 32864 55140 32916 55146
rect 32864 55082 32916 55088
rect 32876 54670 32904 55082
rect 32864 54664 32916 54670
rect 32864 54606 32916 54612
rect 32968 51950 32996 64874
rect 33140 64320 33192 64326
rect 33140 64262 33192 64268
rect 33048 61056 33100 61062
rect 33048 60998 33100 61004
rect 33060 56386 33088 60998
rect 33152 60314 33180 64262
rect 33140 60308 33192 60314
rect 33140 60250 33192 60256
rect 33152 59634 33180 60250
rect 33140 59628 33192 59634
rect 33140 59570 33192 59576
rect 33152 59158 33180 59570
rect 33140 59152 33192 59158
rect 33140 59094 33192 59100
rect 33152 58478 33180 59094
rect 33140 58472 33192 58478
rect 33140 58414 33192 58420
rect 33060 56358 33180 56386
rect 33048 56296 33100 56302
rect 33048 56238 33100 56244
rect 33060 55894 33088 56238
rect 33048 55888 33100 55894
rect 33048 55830 33100 55836
rect 33152 55706 33180 56358
rect 33060 55678 33180 55706
rect 32956 51944 33008 51950
rect 32956 51886 33008 51892
rect 32864 51808 32916 51814
rect 32864 51750 32916 51756
rect 32876 50726 32904 51750
rect 33060 51074 33088 55678
rect 33140 55616 33192 55622
rect 33140 55558 33192 55564
rect 32968 51046 33088 51074
rect 32864 50720 32916 50726
rect 32864 50662 32916 50668
rect 32772 49768 32824 49774
rect 32772 49710 32824 49716
rect 32772 38752 32824 38758
rect 32772 38694 32824 38700
rect 32784 26926 32812 38694
rect 32864 33312 32916 33318
rect 32864 33254 32916 33260
rect 32876 27962 32904 33254
rect 32968 30802 32996 51046
rect 33152 50386 33180 55558
rect 33244 54330 33272 103486
rect 33416 98048 33468 98054
rect 33416 97990 33468 97996
rect 33324 86828 33376 86834
rect 33324 86770 33376 86776
rect 33336 85814 33364 86770
rect 33324 85808 33376 85814
rect 33324 85750 33376 85756
rect 33336 84590 33364 85750
rect 33324 84584 33376 84590
rect 33324 84526 33376 84532
rect 33336 84250 33364 84526
rect 33324 84244 33376 84250
rect 33324 84186 33376 84192
rect 33336 83910 33364 84186
rect 33324 83904 33376 83910
rect 33324 83846 33376 83852
rect 33336 83570 33364 83846
rect 33324 83564 33376 83570
rect 33324 83506 33376 83512
rect 33324 81184 33376 81190
rect 33324 81126 33376 81132
rect 33336 80714 33364 81126
rect 33324 80708 33376 80714
rect 33324 80650 33376 80656
rect 33324 65544 33376 65550
rect 33324 65486 33376 65492
rect 33336 59702 33364 65486
rect 33324 59696 33376 59702
rect 33324 59638 33376 59644
rect 33324 57996 33376 58002
rect 33324 57938 33376 57944
rect 33232 54324 33284 54330
rect 33232 54266 33284 54272
rect 33336 54210 33364 57938
rect 33428 55214 33456 97990
rect 33508 97504 33560 97510
rect 33508 97446 33560 97452
rect 33520 55962 33548 97446
rect 33612 91798 33640 115602
rect 33704 114646 33732 116214
rect 33784 116204 33836 116210
rect 33784 116146 33836 116152
rect 33692 114640 33744 114646
rect 33692 114582 33744 114588
rect 33796 112538 33824 116146
rect 33888 114034 33916 116334
rect 33876 114028 33928 114034
rect 33876 113970 33928 113976
rect 33980 113830 34008 116690
rect 33968 113824 34020 113830
rect 33968 113766 34020 113772
rect 33784 112532 33836 112538
rect 33784 112474 33836 112480
rect 34072 112402 34100 119200
rect 34152 117156 34204 117162
rect 34152 117098 34204 117104
rect 34164 116822 34192 117098
rect 34152 116816 34204 116822
rect 34152 116758 34204 116764
rect 34244 116612 34296 116618
rect 34244 116554 34296 116560
rect 34152 116544 34204 116550
rect 34152 116486 34204 116492
rect 34164 115122 34192 116486
rect 34256 116278 34284 116554
rect 34244 116272 34296 116278
rect 34244 116214 34296 116220
rect 34348 116124 34376 119200
rect 34532 116260 34560 119200
rect 34610 118824 34666 118833
rect 34610 118759 34666 118768
rect 34624 117162 34652 118759
rect 34808 118250 34836 119200
rect 34796 118244 34848 118250
rect 34796 118186 34848 118192
rect 34796 118040 34848 118046
rect 34796 117982 34848 117988
rect 34704 117700 34756 117706
rect 34704 117642 34756 117648
rect 34716 117314 34744 117642
rect 34808 117434 34836 117982
rect 34992 117706 35020 119200
rect 34980 117700 35032 117706
rect 34980 117642 35032 117648
rect 34940 117532 35236 117552
rect 34996 117530 35020 117532
rect 35076 117530 35100 117532
rect 35156 117530 35180 117532
rect 35018 117478 35020 117530
rect 35082 117478 35094 117530
rect 35156 117478 35158 117530
rect 34996 117476 35020 117478
rect 35076 117476 35100 117478
rect 35156 117476 35180 117478
rect 34940 117456 35236 117476
rect 34796 117428 34848 117434
rect 34796 117370 34848 117376
rect 34716 117286 34836 117314
rect 34612 117156 34664 117162
rect 34612 117098 34664 117104
rect 34704 116748 34756 116754
rect 34704 116690 34756 116696
rect 34532 116232 34652 116260
rect 34520 116136 34572 116142
rect 34348 116096 34520 116124
rect 34520 116078 34572 116084
rect 34336 116000 34388 116006
rect 34336 115942 34388 115948
rect 34152 115116 34204 115122
rect 34152 115058 34204 115064
rect 34244 114980 34296 114986
rect 34244 114922 34296 114928
rect 34152 114436 34204 114442
rect 34152 114378 34204 114384
rect 34164 113626 34192 114378
rect 34152 113620 34204 113626
rect 34152 113562 34204 113568
rect 34152 113416 34204 113422
rect 34152 113358 34204 113364
rect 34164 112878 34192 113358
rect 34152 112872 34204 112878
rect 34152 112814 34204 112820
rect 34060 112396 34112 112402
rect 34060 112338 34112 112344
rect 33784 111648 33836 111654
rect 33784 111590 33836 111596
rect 33796 107846 33824 111590
rect 34060 111308 34112 111314
rect 34060 111250 34112 111256
rect 34072 109478 34100 111250
rect 34164 111246 34192 112814
rect 34152 111240 34204 111246
rect 34152 111182 34204 111188
rect 34152 109540 34204 109546
rect 34152 109482 34204 109488
rect 34060 109472 34112 109478
rect 34060 109414 34112 109420
rect 34072 109034 34100 109414
rect 33888 109006 34100 109034
rect 33784 107840 33836 107846
rect 33784 107782 33836 107788
rect 33888 103766 33916 109006
rect 34164 108526 34192 109482
rect 34152 108520 34204 108526
rect 34152 108462 34204 108468
rect 34060 106412 34112 106418
rect 34060 106354 34112 106360
rect 33968 105120 34020 105126
rect 33968 105062 34020 105068
rect 33876 103760 33928 103766
rect 33876 103702 33928 103708
rect 33692 96416 33744 96422
rect 33692 96358 33744 96364
rect 33600 91792 33652 91798
rect 33600 91734 33652 91740
rect 33600 89956 33652 89962
rect 33600 89898 33652 89904
rect 33612 85542 33640 89898
rect 33600 85536 33652 85542
rect 33600 85478 33652 85484
rect 33600 84992 33652 84998
rect 33600 84934 33652 84940
rect 33612 83434 33640 84934
rect 33600 83428 33652 83434
rect 33600 83370 33652 83376
rect 33612 83026 33640 83370
rect 33600 83020 33652 83026
rect 33600 82962 33652 82968
rect 33600 81932 33652 81938
rect 33600 81874 33652 81880
rect 33612 81734 33640 81874
rect 33600 81728 33652 81734
rect 33600 81670 33652 81676
rect 33600 81388 33652 81394
rect 33600 81330 33652 81336
rect 33612 80986 33640 81330
rect 33600 80980 33652 80986
rect 33600 80922 33652 80928
rect 33600 66020 33652 66026
rect 33600 65962 33652 65968
rect 33612 62937 33640 65962
rect 33598 62928 33654 62937
rect 33598 62863 33654 62872
rect 33600 62756 33652 62762
rect 33600 62698 33652 62704
rect 33612 59770 33640 62698
rect 33600 59764 33652 59770
rect 33600 59706 33652 59712
rect 33600 59424 33652 59430
rect 33600 59366 33652 59372
rect 33612 59090 33640 59366
rect 33600 59084 33652 59090
rect 33600 59026 33652 59032
rect 33600 58336 33652 58342
rect 33600 58278 33652 58284
rect 33508 55956 33560 55962
rect 33508 55898 33560 55904
rect 33612 55622 33640 58278
rect 33704 56370 33732 96358
rect 33876 94784 33928 94790
rect 33876 94726 33928 94732
rect 33888 93362 33916 94726
rect 33980 94602 34008 105062
rect 34072 94790 34100 106354
rect 34164 103290 34192 108462
rect 34256 108118 34284 114922
rect 34348 112878 34376 115942
rect 34520 115728 34572 115734
rect 34518 115696 34520 115705
rect 34572 115696 34574 115705
rect 34518 115631 34574 115640
rect 34520 114980 34572 114986
rect 34520 114922 34572 114928
rect 34428 114368 34480 114374
rect 34428 114310 34480 114316
rect 34440 114102 34468 114310
rect 34428 114096 34480 114102
rect 34428 114038 34480 114044
rect 34428 113416 34480 113422
rect 34428 113358 34480 113364
rect 34336 112872 34388 112878
rect 34336 112814 34388 112820
rect 34336 112736 34388 112742
rect 34336 112678 34388 112684
rect 34348 111654 34376 112678
rect 34336 111648 34388 111654
rect 34336 111590 34388 111596
rect 34440 111314 34468 113358
rect 34428 111308 34480 111314
rect 34428 111250 34480 111256
rect 34428 111104 34480 111110
rect 34428 111046 34480 111052
rect 34336 109472 34388 109478
rect 34336 109414 34388 109420
rect 34348 109206 34376 109414
rect 34336 109200 34388 109206
rect 34336 109142 34388 109148
rect 34440 108474 34468 111046
rect 34532 109274 34560 114922
rect 34624 114034 34652 116232
rect 34612 114028 34664 114034
rect 34612 113970 34664 113976
rect 34612 113892 34664 113898
rect 34612 113834 34664 113840
rect 34520 109268 34572 109274
rect 34520 109210 34572 109216
rect 34348 108446 34468 108474
rect 34244 108112 34296 108118
rect 34244 108054 34296 108060
rect 34348 107386 34376 108446
rect 34520 108384 34572 108390
rect 34520 108326 34572 108332
rect 34428 108112 34480 108118
rect 34428 108054 34480 108060
rect 34256 107358 34376 107386
rect 34152 103284 34204 103290
rect 34152 103226 34204 103232
rect 34152 100496 34204 100502
rect 34152 100438 34204 100444
rect 34060 94784 34112 94790
rect 34060 94726 34112 94732
rect 33980 94574 34100 94602
rect 33968 94036 34020 94042
rect 33968 93978 34020 93984
rect 33876 93356 33928 93362
rect 33876 93298 33928 93304
rect 33980 91746 34008 93978
rect 33888 91718 34008 91746
rect 33784 87848 33836 87854
rect 33784 87790 33836 87796
rect 33796 87378 33824 87790
rect 33784 87372 33836 87378
rect 33784 87314 33836 87320
rect 33796 86902 33824 87314
rect 33784 86896 33836 86902
rect 33784 86838 33836 86844
rect 33796 86766 33824 86838
rect 33784 86760 33836 86766
rect 33784 86702 33836 86708
rect 33796 86290 33824 86702
rect 33784 86284 33836 86290
rect 33784 86226 33836 86232
rect 33888 84590 33916 91718
rect 33968 91588 34020 91594
rect 33968 91530 34020 91536
rect 33980 85678 34008 91530
rect 34072 88330 34100 94574
rect 34060 88324 34112 88330
rect 34060 88266 34112 88272
rect 34164 87922 34192 100438
rect 34152 87916 34204 87922
rect 34152 87858 34204 87864
rect 34060 87848 34112 87854
rect 34060 87790 34112 87796
rect 34072 87242 34100 87790
rect 34152 87440 34204 87446
rect 34152 87382 34204 87388
rect 34060 87236 34112 87242
rect 34060 87178 34112 87184
rect 34164 86086 34192 87382
rect 34152 86080 34204 86086
rect 34152 86022 34204 86028
rect 33968 85672 34020 85678
rect 33968 85614 34020 85620
rect 34152 84720 34204 84726
rect 34152 84662 34204 84668
rect 33876 84584 33928 84590
rect 33876 84526 33928 84532
rect 34060 84516 34112 84522
rect 34060 84458 34112 84464
rect 33784 84448 33836 84454
rect 33784 84390 33836 84396
rect 33796 81734 33824 84390
rect 34072 84182 34100 84458
rect 34060 84176 34112 84182
rect 34060 84118 34112 84124
rect 33968 84108 34020 84114
rect 33888 84068 33968 84096
rect 33784 81728 33836 81734
rect 33784 81670 33836 81676
rect 33796 81326 33824 81670
rect 33784 81320 33836 81326
rect 33784 81262 33836 81268
rect 33796 80850 33824 81262
rect 33784 80844 33836 80850
rect 33784 80786 33836 80792
rect 33796 80442 33824 80786
rect 33784 80436 33836 80442
rect 33784 80378 33836 80384
rect 33888 79558 33916 84068
rect 33968 84050 34020 84056
rect 34164 81938 34192 84662
rect 34152 81932 34204 81938
rect 34152 81874 34204 81880
rect 33968 81388 34020 81394
rect 33968 81330 34020 81336
rect 33980 80986 34008 81330
rect 34164 81326 34192 81874
rect 34060 81320 34112 81326
rect 34060 81262 34112 81268
rect 34152 81320 34204 81326
rect 34152 81262 34204 81268
rect 33968 80980 34020 80986
rect 33968 80922 34020 80928
rect 33876 79552 33928 79558
rect 33876 79494 33928 79500
rect 34072 79354 34100 81262
rect 34164 80850 34192 81262
rect 34152 80844 34204 80850
rect 34152 80786 34204 80792
rect 34164 80714 34192 80786
rect 34152 80708 34204 80714
rect 34152 80650 34204 80656
rect 34060 79348 34112 79354
rect 34060 79290 34112 79296
rect 33784 76016 33836 76022
rect 33784 75958 33836 75964
rect 33796 60042 33824 75958
rect 33876 75268 33928 75274
rect 33876 75210 33928 75216
rect 33784 60036 33836 60042
rect 33784 59978 33836 59984
rect 33888 59922 33916 75210
rect 34060 74452 34112 74458
rect 34060 74394 34112 74400
rect 33968 69216 34020 69222
rect 33968 69158 34020 69164
rect 33796 59894 33916 59922
rect 33796 59022 33824 59894
rect 33876 59764 33928 59770
rect 33876 59706 33928 59712
rect 33784 59016 33836 59022
rect 33784 58958 33836 58964
rect 33784 58676 33836 58682
rect 33784 58618 33836 58624
rect 33692 56364 33744 56370
rect 33692 56306 33744 56312
rect 33600 55616 33652 55622
rect 33600 55558 33652 55564
rect 33508 55276 33560 55282
rect 33508 55218 33560 55224
rect 33416 55208 33468 55214
rect 33416 55150 33468 55156
rect 33520 54738 33548 55218
rect 33692 55072 33744 55078
rect 33692 55014 33744 55020
rect 33508 54732 33560 54738
rect 33508 54674 33560 54680
rect 33416 54528 33468 54534
rect 33416 54470 33468 54476
rect 33244 54182 33364 54210
rect 33244 51474 33272 54182
rect 33232 51468 33284 51474
rect 33232 51410 33284 51416
rect 33428 51074 33456 54470
rect 33508 51808 33560 51814
rect 33508 51750 33560 51756
rect 33600 51808 33652 51814
rect 33600 51750 33652 51756
rect 33520 51474 33548 51750
rect 33612 51610 33640 51750
rect 33600 51604 33652 51610
rect 33600 51546 33652 51552
rect 33508 51468 33560 51474
rect 33508 51410 33560 51416
rect 33244 51046 33456 51074
rect 33140 50380 33192 50386
rect 33140 50322 33192 50328
rect 33048 42764 33100 42770
rect 33048 42706 33100 42712
rect 33060 31890 33088 42706
rect 33140 35828 33192 35834
rect 33140 35770 33192 35776
rect 33152 35154 33180 35770
rect 33140 35148 33192 35154
rect 33140 35090 33192 35096
rect 33140 33380 33192 33386
rect 33140 33322 33192 33328
rect 33048 31884 33100 31890
rect 33048 31826 33100 31832
rect 32956 30796 33008 30802
rect 32956 30738 33008 30744
rect 33048 28416 33100 28422
rect 33048 28358 33100 28364
rect 32876 27946 32996 27962
rect 32876 27940 33008 27946
rect 32876 27934 32956 27940
rect 32956 27882 33008 27888
rect 32968 27606 32996 27882
rect 32956 27600 33008 27606
rect 32956 27542 33008 27548
rect 32772 26920 32824 26926
rect 32772 26862 32824 26868
rect 32968 26858 32996 27542
rect 33060 27538 33088 28358
rect 33152 28014 33180 33322
rect 33140 28008 33192 28014
rect 33140 27950 33192 27956
rect 33152 27674 33180 27950
rect 33140 27668 33192 27674
rect 33140 27610 33192 27616
rect 33048 27532 33100 27538
rect 33048 27474 33100 27480
rect 33152 26926 33180 27610
rect 33140 26920 33192 26926
rect 33140 26862 33192 26868
rect 32956 26852 33008 26858
rect 32956 26794 33008 26800
rect 32772 26784 32824 26790
rect 32772 26726 32824 26732
rect 32680 26444 32732 26450
rect 32680 26386 32732 26392
rect 32680 25968 32732 25974
rect 32680 25910 32732 25916
rect 32588 25356 32640 25362
rect 32588 25298 32640 25304
rect 32404 24744 32456 24750
rect 32404 24686 32456 24692
rect 32588 24608 32640 24614
rect 32588 24550 32640 24556
rect 32404 24336 32456 24342
rect 32404 24278 32456 24284
rect 32232 22936 32352 22964
rect 32220 22772 32272 22778
rect 32220 22714 32272 22720
rect 32048 22066 32168 22094
rect 32048 21729 32076 22066
rect 32128 21956 32180 21962
rect 32128 21898 32180 21904
rect 32034 21720 32090 21729
rect 32034 21655 32090 21664
rect 32036 21548 32088 21554
rect 32036 21490 32088 21496
rect 31944 20392 31996 20398
rect 31944 20334 31996 20340
rect 31944 20256 31996 20262
rect 31944 20198 31996 20204
rect 31956 19514 31984 20198
rect 31944 19508 31996 19514
rect 31944 19450 31996 19456
rect 31852 19304 31904 19310
rect 31852 19246 31904 19252
rect 31956 18970 31984 19450
rect 31760 18964 31812 18970
rect 31760 18906 31812 18912
rect 31944 18964 31996 18970
rect 31944 18906 31996 18912
rect 31944 18624 31996 18630
rect 31944 18566 31996 18572
rect 31956 18426 31984 18566
rect 31944 18420 31996 18426
rect 31944 18362 31996 18368
rect 31852 17808 31904 17814
rect 31852 17750 31904 17756
rect 31760 17536 31812 17542
rect 31760 17478 31812 17484
rect 31772 16561 31800 17478
rect 31864 17066 31892 17750
rect 31852 17060 31904 17066
rect 31852 17002 31904 17008
rect 31956 16946 31984 18362
rect 32048 18086 32076 21490
rect 32140 19446 32168 21898
rect 32232 21593 32260 22714
rect 32324 22273 32352 22936
rect 32416 22556 32444 24278
rect 32496 23248 32548 23254
rect 32496 23190 32548 23196
rect 32508 22710 32536 23190
rect 32496 22704 32548 22710
rect 32496 22646 32548 22652
rect 32496 22568 32548 22574
rect 32416 22528 32496 22556
rect 32496 22510 32548 22516
rect 32404 22432 32456 22438
rect 32404 22374 32456 22380
rect 32310 22264 32366 22273
rect 32310 22199 32366 22208
rect 32312 21616 32364 21622
rect 32218 21584 32274 21593
rect 32312 21558 32364 21564
rect 32218 21519 32274 21528
rect 32220 21480 32272 21486
rect 32220 21422 32272 21428
rect 32232 21010 32260 21422
rect 32324 21078 32352 21558
rect 32312 21072 32364 21078
rect 32312 21014 32364 21020
rect 32220 21004 32272 21010
rect 32220 20946 32272 20952
rect 32232 20874 32260 20946
rect 32220 20868 32272 20874
rect 32220 20810 32272 20816
rect 32312 20868 32364 20874
rect 32312 20810 32364 20816
rect 32220 20324 32272 20330
rect 32220 20266 32272 20272
rect 32232 19922 32260 20266
rect 32324 20262 32352 20810
rect 32312 20256 32364 20262
rect 32312 20198 32364 20204
rect 32220 19916 32272 19922
rect 32220 19858 32272 19864
rect 32128 19440 32180 19446
rect 32128 19382 32180 19388
rect 32232 19378 32260 19858
rect 32310 19408 32366 19417
rect 32220 19372 32272 19378
rect 32310 19343 32366 19352
rect 32220 19314 32272 19320
rect 32232 18834 32260 19314
rect 32220 18828 32272 18834
rect 32220 18770 32272 18776
rect 32232 18358 32260 18770
rect 32220 18352 32272 18358
rect 32220 18294 32272 18300
rect 32036 18080 32088 18086
rect 32036 18022 32088 18028
rect 31864 16918 31984 16946
rect 31758 16552 31814 16561
rect 31758 16487 31814 16496
rect 31668 16040 31720 16046
rect 31668 15982 31720 15988
rect 31576 15972 31628 15978
rect 31576 15914 31628 15920
rect 31588 14550 31616 15914
rect 31864 15570 31892 16918
rect 31944 16448 31996 16454
rect 31944 16390 31996 16396
rect 31852 15564 31904 15570
rect 31852 15506 31904 15512
rect 31666 15328 31722 15337
rect 31666 15263 31722 15272
rect 31680 15162 31708 15263
rect 31668 15156 31720 15162
rect 31668 15098 31720 15104
rect 31956 14906 31984 16390
rect 31864 14878 31984 14906
rect 31576 14544 31628 14550
rect 31576 14486 31628 14492
rect 31864 14346 31892 14878
rect 31944 14816 31996 14822
rect 31944 14758 31996 14764
rect 31852 14340 31904 14346
rect 31852 14282 31904 14288
rect 31956 13462 31984 14758
rect 31944 13456 31996 13462
rect 31944 13398 31996 13404
rect 32048 12434 32076 18022
rect 32232 17746 32260 18294
rect 32324 18034 32352 19343
rect 32416 18222 32444 22374
rect 32508 22166 32536 22510
rect 32496 22160 32548 22166
rect 32496 22102 32548 22108
rect 32508 21593 32536 22102
rect 32494 21584 32550 21593
rect 32494 21519 32550 21528
rect 32496 21480 32548 21486
rect 32496 21422 32548 21428
rect 32508 21010 32536 21422
rect 32496 21004 32548 21010
rect 32496 20946 32548 20952
rect 32496 20800 32548 20806
rect 32496 20742 32548 20748
rect 32404 18216 32456 18222
rect 32404 18158 32456 18164
rect 32324 18006 32444 18034
rect 32220 17740 32272 17746
rect 32220 17682 32272 17688
rect 32128 17196 32180 17202
rect 32128 17138 32180 17144
rect 32140 15094 32168 17138
rect 32232 16794 32260 17682
rect 32312 17128 32364 17134
rect 32312 17070 32364 17076
rect 32220 16788 32272 16794
rect 32220 16730 32272 16736
rect 32324 16658 32352 17070
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 32416 16538 32444 18006
rect 32508 17814 32536 20742
rect 32600 19258 32628 24550
rect 32692 22642 32720 25910
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32784 22522 32812 26726
rect 32968 26382 32996 26794
rect 33152 26586 33180 26862
rect 33140 26580 33192 26586
rect 33140 26522 33192 26528
rect 32956 26376 33008 26382
rect 32956 26318 33008 26324
rect 32968 25770 32996 26318
rect 33048 25968 33100 25974
rect 33048 25910 33100 25916
rect 32956 25764 33008 25770
rect 32956 25706 33008 25712
rect 32956 25424 33008 25430
rect 32956 25366 33008 25372
rect 32864 24880 32916 24886
rect 32864 24822 32916 24828
rect 32876 22545 32904 24822
rect 32968 24750 32996 25366
rect 32956 24744 33008 24750
rect 32956 24686 33008 24692
rect 32954 24576 33010 24585
rect 32954 24511 33010 24520
rect 32968 24274 32996 24511
rect 32956 24268 33008 24274
rect 32956 24210 33008 24216
rect 32956 23792 33008 23798
rect 32956 23734 33008 23740
rect 32968 23118 32996 23734
rect 32956 23112 33008 23118
rect 32956 23054 33008 23060
rect 32956 22976 33008 22982
rect 32956 22918 33008 22924
rect 32692 22494 32812 22522
rect 32862 22536 32918 22545
rect 32692 19394 32720 22494
rect 32862 22471 32918 22480
rect 32864 22432 32916 22438
rect 32864 22374 32916 22380
rect 32772 21684 32824 21690
rect 32772 21626 32824 21632
rect 32784 21010 32812 21626
rect 32772 21004 32824 21010
rect 32772 20946 32824 20952
rect 32770 20904 32826 20913
rect 32770 20839 32826 20848
rect 32784 20262 32812 20839
rect 32876 20448 32904 22374
rect 32968 20806 32996 22918
rect 33060 22137 33088 25910
rect 33152 25838 33180 26522
rect 33140 25832 33192 25838
rect 33140 25774 33192 25780
rect 33140 25220 33192 25226
rect 33140 25162 33192 25168
rect 33152 24206 33180 25162
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 33140 23520 33192 23526
rect 33140 23462 33192 23468
rect 33046 22128 33102 22137
rect 33046 22063 33102 22072
rect 33048 21888 33100 21894
rect 33048 21830 33100 21836
rect 32956 20800 33008 20806
rect 32956 20742 33008 20748
rect 32876 20420 32996 20448
rect 32862 20360 32918 20369
rect 32862 20295 32918 20304
rect 32772 20256 32824 20262
rect 32772 20198 32824 20204
rect 32784 19553 32812 20198
rect 32876 19718 32904 20295
rect 32864 19712 32916 19718
rect 32864 19654 32916 19660
rect 32770 19544 32826 19553
rect 32770 19479 32826 19488
rect 32692 19366 32904 19394
rect 32600 19230 32812 19258
rect 32680 18760 32732 18766
rect 32680 18702 32732 18708
rect 32588 18080 32640 18086
rect 32588 18022 32640 18028
rect 32496 17808 32548 17814
rect 32496 17750 32548 17756
rect 32600 17626 32628 18022
rect 32232 16510 32444 16538
rect 32508 17598 32628 17626
rect 32128 15088 32180 15094
rect 32128 15030 32180 15036
rect 31404 12406 31524 12434
rect 31864 12406 32076 12434
rect 31300 11348 31352 11354
rect 31300 11290 31352 11296
rect 31300 7948 31352 7954
rect 31300 7890 31352 7896
rect 31312 2990 31340 7890
rect 31404 3777 31432 12406
rect 31760 5568 31812 5574
rect 31760 5510 31812 5516
rect 31772 4146 31800 5510
rect 31864 4486 31892 12406
rect 31944 4684 31996 4690
rect 31944 4626 31996 4632
rect 31852 4480 31904 4486
rect 31852 4422 31904 4428
rect 31668 4140 31720 4146
rect 31668 4082 31720 4088
rect 31760 4140 31812 4146
rect 31760 4082 31812 4088
rect 31680 4026 31708 4082
rect 31852 4072 31904 4078
rect 31496 3998 31708 4026
rect 31850 4040 31852 4049
rect 31904 4040 31906 4049
rect 31390 3768 31446 3777
rect 31390 3703 31446 3712
rect 31496 3534 31524 3998
rect 31850 3975 31906 3984
rect 31760 3936 31812 3942
rect 31666 3904 31722 3913
rect 31760 3878 31812 3884
rect 31852 3936 31904 3942
rect 31852 3878 31904 3884
rect 31666 3839 31722 3848
rect 31576 3664 31628 3670
rect 31576 3606 31628 3612
rect 31484 3528 31536 3534
rect 31588 3505 31616 3606
rect 31484 3470 31536 3476
rect 31574 3496 31630 3505
rect 31574 3431 31630 3440
rect 31208 2984 31260 2990
rect 31208 2926 31260 2932
rect 31300 2984 31352 2990
rect 31300 2926 31352 2932
rect 31300 2848 31352 2854
rect 31300 2790 31352 2796
rect 30668 2746 30788 2774
rect 30668 800 30696 2746
rect 30932 2508 30984 2514
rect 30932 2450 30984 2456
rect 30944 800 30972 2450
rect 31116 2304 31168 2310
rect 31116 2246 31168 2252
rect 31128 2038 31156 2246
rect 31116 2032 31168 2038
rect 31116 1974 31168 1980
rect 31312 800 31340 2790
rect 31680 800 31708 3839
rect 31772 3602 31800 3878
rect 31760 3596 31812 3602
rect 31760 3538 31812 3544
rect 31864 3210 31892 3878
rect 31772 3182 31892 3210
rect 31772 3126 31800 3182
rect 31760 3120 31812 3126
rect 31760 3062 31812 3068
rect 31956 800 31984 4626
rect 32036 4480 32088 4486
rect 32036 4422 32088 4428
rect 32048 3058 32076 4422
rect 32128 4140 32180 4146
rect 32128 4082 32180 4088
rect 32140 3126 32168 4082
rect 32128 3120 32180 3126
rect 32128 3062 32180 3068
rect 32036 3052 32088 3058
rect 32036 2994 32088 3000
rect 32232 2990 32260 16510
rect 32312 16108 32364 16114
rect 32312 16050 32364 16056
rect 32324 16017 32352 16050
rect 32404 16040 32456 16046
rect 32310 16008 32366 16017
rect 32404 15982 32456 15988
rect 32310 15943 32366 15952
rect 32312 14952 32364 14958
rect 32312 14894 32364 14900
rect 32324 13870 32352 14894
rect 32312 13864 32364 13870
rect 32312 13806 32364 13812
rect 32312 13728 32364 13734
rect 32312 13670 32364 13676
rect 32324 3398 32352 13670
rect 32416 5030 32444 15982
rect 32508 13734 32536 17598
rect 32588 16516 32640 16522
rect 32588 16458 32640 16464
rect 32600 15910 32628 16458
rect 32588 15904 32640 15910
rect 32588 15846 32640 15852
rect 32588 15496 32640 15502
rect 32588 15438 32640 15444
rect 32600 15162 32628 15438
rect 32588 15156 32640 15162
rect 32588 15098 32640 15104
rect 32692 14346 32720 18702
rect 32784 16046 32812 19230
rect 32772 16040 32824 16046
rect 32772 15982 32824 15988
rect 32772 15700 32824 15706
rect 32772 15642 32824 15648
rect 32784 15026 32812 15642
rect 32772 15020 32824 15026
rect 32772 14962 32824 14968
rect 32876 14958 32904 19366
rect 32968 18902 32996 20420
rect 33060 19242 33088 21830
rect 33152 21078 33180 23462
rect 33244 22098 33272 51046
rect 33520 50862 33548 51410
rect 33508 50856 33560 50862
rect 33508 50798 33560 50804
rect 33324 50720 33376 50726
rect 33324 50662 33376 50668
rect 33336 49094 33364 50662
rect 33520 50182 33548 50798
rect 33612 50726 33640 51546
rect 33704 50930 33732 55014
rect 33692 50924 33744 50930
rect 33692 50866 33744 50872
rect 33600 50720 33652 50726
rect 33600 50662 33652 50668
rect 33612 50250 33640 50662
rect 33692 50516 33744 50522
rect 33692 50458 33744 50464
rect 33600 50244 33652 50250
rect 33600 50186 33652 50192
rect 33704 50182 33732 50458
rect 33508 50176 33560 50182
rect 33508 50118 33560 50124
rect 33692 50176 33744 50182
rect 33692 50118 33744 50124
rect 33520 49910 33548 50118
rect 33508 49904 33560 49910
rect 33508 49846 33560 49852
rect 33324 49088 33376 49094
rect 33324 49030 33376 49036
rect 33796 46510 33824 58618
rect 33888 56234 33916 59706
rect 33876 56228 33928 56234
rect 33876 56170 33928 56176
rect 33888 55894 33916 56170
rect 33876 55888 33928 55894
rect 33876 55830 33928 55836
rect 33888 55282 33916 55830
rect 33876 55276 33928 55282
rect 33876 55218 33928 55224
rect 33980 55214 34008 69158
rect 34072 60178 34100 74394
rect 34152 67108 34204 67114
rect 34152 67050 34204 67056
rect 34164 64530 34192 67050
rect 34152 64524 34204 64530
rect 34152 64466 34204 64472
rect 34152 64388 34204 64394
rect 34152 64330 34204 64336
rect 34060 60172 34112 60178
rect 34060 60114 34112 60120
rect 34164 60110 34192 64330
rect 34152 60104 34204 60110
rect 34152 60046 34204 60052
rect 34164 59498 34192 60046
rect 34152 59492 34204 59498
rect 34152 59434 34204 59440
rect 34164 59226 34192 59434
rect 34152 59220 34204 59226
rect 34152 59162 34204 59168
rect 34164 59090 34192 59162
rect 34152 59084 34204 59090
rect 34152 59026 34204 59032
rect 34060 58608 34112 58614
rect 34060 58550 34112 58556
rect 34072 58426 34100 58550
rect 34164 58546 34192 59026
rect 34152 58540 34204 58546
rect 34152 58482 34204 58488
rect 34072 58398 34192 58426
rect 34060 58132 34112 58138
rect 34060 58074 34112 58080
rect 33968 55208 34020 55214
rect 33968 55150 34020 55156
rect 33876 54868 33928 54874
rect 33876 54810 33928 54816
rect 33784 46504 33836 46510
rect 33784 46446 33836 46452
rect 33784 45076 33836 45082
rect 33784 45018 33836 45024
rect 33416 44464 33468 44470
rect 33416 44406 33468 44412
rect 33428 38486 33456 44406
rect 33692 44396 33744 44402
rect 33692 44338 33744 44344
rect 33704 38554 33732 44338
rect 33796 42158 33824 45018
rect 33888 44334 33916 54810
rect 34072 51074 34100 58074
rect 34164 56250 34192 58398
rect 34256 56370 34284 107358
rect 34336 107296 34388 107302
rect 34336 107238 34388 107244
rect 34348 94518 34376 107238
rect 34336 94512 34388 94518
rect 34336 94454 34388 94460
rect 34336 87848 34388 87854
rect 34336 87790 34388 87796
rect 34348 87378 34376 87790
rect 34336 87372 34388 87378
rect 34336 87314 34388 87320
rect 34348 86766 34376 87314
rect 34336 86760 34388 86766
rect 34336 86702 34388 86708
rect 34348 86329 34376 86702
rect 34334 86320 34390 86329
rect 34334 86255 34336 86264
rect 34388 86255 34390 86264
rect 34336 86226 34388 86232
rect 34336 86080 34388 86086
rect 34336 86022 34388 86028
rect 34348 83706 34376 86022
rect 34336 83700 34388 83706
rect 34336 83642 34388 83648
rect 34336 73092 34388 73098
rect 34336 73034 34388 73040
rect 34348 59090 34376 73034
rect 34440 65754 34468 108054
rect 34532 105874 34560 108326
rect 34520 105868 34572 105874
rect 34520 105810 34572 105816
rect 34520 99952 34572 99958
rect 34520 99894 34572 99900
rect 34532 86290 34560 99894
rect 34520 86284 34572 86290
rect 34520 86226 34572 86232
rect 34520 85604 34572 85610
rect 34520 85546 34572 85552
rect 34532 75546 34560 85546
rect 34520 75540 34572 75546
rect 34520 75482 34572 75488
rect 34520 68672 34572 68678
rect 34520 68614 34572 68620
rect 34532 68406 34560 68614
rect 34520 68400 34572 68406
rect 34520 68342 34572 68348
rect 34520 66496 34572 66502
rect 34520 66438 34572 66444
rect 34428 65748 34480 65754
rect 34428 65690 34480 65696
rect 34532 65686 34560 66438
rect 34520 65680 34572 65686
rect 34520 65622 34572 65628
rect 34428 65476 34480 65482
rect 34428 65418 34480 65424
rect 34336 59084 34388 59090
rect 34336 59026 34388 59032
rect 34336 58064 34388 58070
rect 34336 58006 34388 58012
rect 34244 56364 34296 56370
rect 34244 56306 34296 56312
rect 34164 56222 34284 56250
rect 34152 56160 34204 56166
rect 34152 56102 34204 56108
rect 33980 51046 34100 51074
rect 33980 47122 34008 51046
rect 34060 50924 34112 50930
rect 34060 50866 34112 50872
rect 33968 47116 34020 47122
rect 33968 47058 34020 47064
rect 34072 47002 34100 50866
rect 33980 46974 34100 47002
rect 33876 44328 33928 44334
rect 33876 44270 33928 44276
rect 33980 43994 34008 46974
rect 34060 45416 34112 45422
rect 34060 45358 34112 45364
rect 34072 44742 34100 45358
rect 34060 44736 34112 44742
rect 34060 44678 34112 44684
rect 34060 44464 34112 44470
rect 34060 44406 34112 44412
rect 34072 44266 34100 44406
rect 34060 44260 34112 44266
rect 34060 44202 34112 44208
rect 33968 43988 34020 43994
rect 33968 43930 34020 43936
rect 33876 42628 33928 42634
rect 33876 42570 33928 42576
rect 33784 42152 33836 42158
rect 33784 42094 33836 42100
rect 33888 41682 33916 42570
rect 33968 42152 34020 42158
rect 33968 42094 34020 42100
rect 33876 41676 33928 41682
rect 33876 41618 33928 41624
rect 33980 41562 34008 42094
rect 34060 42084 34112 42090
rect 34060 42026 34112 42032
rect 34072 41750 34100 42026
rect 34060 41744 34112 41750
rect 34060 41686 34112 41692
rect 33980 41546 34100 41562
rect 33876 41540 33928 41546
rect 33980 41540 34112 41546
rect 33980 41534 34060 41540
rect 33876 41482 33928 41488
rect 34060 41482 34112 41488
rect 33888 41070 33916 41482
rect 33876 41064 33928 41070
rect 33876 41006 33928 41012
rect 33888 39982 33916 41006
rect 34072 41002 34100 41482
rect 34060 40996 34112 41002
rect 34060 40938 34112 40944
rect 33876 39976 33928 39982
rect 33876 39918 33928 39924
rect 33888 39574 33916 39918
rect 34072 39914 34100 40938
rect 34060 39908 34112 39914
rect 34060 39850 34112 39856
rect 33876 39568 33928 39574
rect 33876 39510 33928 39516
rect 33692 38548 33744 38554
rect 33692 38490 33744 38496
rect 33416 38480 33468 38486
rect 33416 38422 33468 38428
rect 33508 38480 33560 38486
rect 33508 38422 33560 38428
rect 33520 36174 33548 38422
rect 33784 38412 33836 38418
rect 33784 38354 33836 38360
rect 33692 38276 33744 38282
rect 33692 38218 33744 38224
rect 33600 38208 33652 38214
rect 33600 38150 33652 38156
rect 33612 37806 33640 38150
rect 33704 37806 33732 38218
rect 33600 37800 33652 37806
rect 33600 37742 33652 37748
rect 33692 37800 33744 37806
rect 33692 37742 33744 37748
rect 33612 36786 33640 37742
rect 33600 36780 33652 36786
rect 33600 36722 33652 36728
rect 33612 36378 33640 36722
rect 33704 36582 33732 37742
rect 33692 36576 33744 36582
rect 33692 36518 33744 36524
rect 33704 36378 33732 36518
rect 33600 36372 33652 36378
rect 33600 36314 33652 36320
rect 33692 36372 33744 36378
rect 33692 36314 33744 36320
rect 33508 36168 33560 36174
rect 33508 36110 33560 36116
rect 33612 35698 33640 36314
rect 33600 35692 33652 35698
rect 33600 35634 33652 35640
rect 33416 35488 33468 35494
rect 33416 35430 33468 35436
rect 33508 35488 33560 35494
rect 33508 35430 33560 35436
rect 33428 32366 33456 35430
rect 33520 35154 33548 35430
rect 33612 35290 33640 35634
rect 33704 35494 33732 36314
rect 33796 36145 33824 38354
rect 33888 36922 33916 39510
rect 34072 39506 34100 39850
rect 34060 39500 34112 39506
rect 34060 39442 34112 39448
rect 34072 39386 34100 39442
rect 33980 39358 34100 39386
rect 33876 36916 33928 36922
rect 33876 36858 33928 36864
rect 33876 36576 33928 36582
rect 33876 36518 33928 36524
rect 33888 36310 33916 36518
rect 33980 36378 34008 39358
rect 34060 37664 34112 37670
rect 34060 37606 34112 37612
rect 33968 36372 34020 36378
rect 33968 36314 34020 36320
rect 33876 36304 33928 36310
rect 33876 36246 33928 36252
rect 33968 36236 34020 36242
rect 33968 36178 34020 36184
rect 33782 36136 33838 36145
rect 33782 36071 33838 36080
rect 33692 35488 33744 35494
rect 33692 35430 33744 35436
rect 33796 35306 33824 36071
rect 33876 35488 33928 35494
rect 33876 35430 33928 35436
rect 33600 35284 33652 35290
rect 33600 35226 33652 35232
rect 33704 35278 33824 35306
rect 33704 35170 33732 35278
rect 33508 35148 33560 35154
rect 33508 35090 33560 35096
rect 33612 35142 33732 35170
rect 33784 35216 33836 35222
rect 33784 35158 33836 35164
rect 33324 32360 33376 32366
rect 33324 32302 33376 32308
rect 33416 32360 33468 32366
rect 33416 32302 33468 32308
rect 33336 31958 33364 32302
rect 33428 31958 33456 32302
rect 33324 31952 33376 31958
rect 33324 31894 33376 31900
rect 33416 31952 33468 31958
rect 33416 31894 33468 31900
rect 33336 31482 33364 31894
rect 33324 31476 33376 31482
rect 33324 31418 33376 31424
rect 33428 31362 33456 31894
rect 33508 31476 33560 31482
rect 33508 31418 33560 31424
rect 33336 31334 33456 31362
rect 33336 31278 33364 31334
rect 33324 31272 33376 31278
rect 33324 31214 33376 31220
rect 33324 31136 33376 31142
rect 33324 31078 33376 31084
rect 33336 30802 33364 31078
rect 33428 30870 33456 31334
rect 33520 31142 33548 31418
rect 33508 31136 33560 31142
rect 33508 31078 33560 31084
rect 33416 30864 33468 30870
rect 33416 30806 33468 30812
rect 33324 30796 33376 30802
rect 33324 30738 33376 30744
rect 33336 30326 33364 30738
rect 33428 30326 33456 30806
rect 33324 30320 33376 30326
rect 33324 30262 33376 30268
rect 33416 30320 33468 30326
rect 33416 30262 33468 30268
rect 33612 27878 33640 35142
rect 33692 35012 33744 35018
rect 33692 34954 33744 34960
rect 33704 31482 33732 34954
rect 33796 33454 33824 35158
rect 33888 35086 33916 35430
rect 33876 35080 33928 35086
rect 33876 35022 33928 35028
rect 33876 34944 33928 34950
rect 33876 34886 33928 34892
rect 33784 33448 33836 33454
rect 33784 33390 33836 33396
rect 33692 31476 33744 31482
rect 33692 31418 33744 31424
rect 33888 31226 33916 34886
rect 33980 34746 34008 36178
rect 33968 34740 34020 34746
rect 33968 34682 34020 34688
rect 33968 32020 34020 32026
rect 33968 31962 34020 31968
rect 33704 31198 33916 31226
rect 33508 27872 33560 27878
rect 33508 27814 33560 27820
rect 33600 27872 33652 27878
rect 33600 27814 33652 27820
rect 33416 26308 33468 26314
rect 33416 26250 33468 26256
rect 33324 26240 33376 26246
rect 33324 26182 33376 26188
rect 33336 25430 33364 26182
rect 33324 25424 33376 25430
rect 33324 25366 33376 25372
rect 33324 25220 33376 25226
rect 33324 25162 33376 25168
rect 33336 23186 33364 25162
rect 33324 23180 33376 23186
rect 33324 23122 33376 23128
rect 33324 23044 33376 23050
rect 33324 22986 33376 22992
rect 33336 22574 33364 22986
rect 33324 22568 33376 22574
rect 33324 22510 33376 22516
rect 33322 22400 33378 22409
rect 33322 22335 33378 22344
rect 33232 22092 33284 22098
rect 33232 22034 33284 22040
rect 33230 21992 33286 22001
rect 33230 21927 33286 21936
rect 33140 21072 33192 21078
rect 33140 21014 33192 21020
rect 33138 20768 33194 20777
rect 33138 20703 33194 20712
rect 33048 19236 33100 19242
rect 33048 19178 33100 19184
rect 33152 18970 33180 20703
rect 33244 20534 33272 21927
rect 33336 21350 33364 22335
rect 33324 21344 33376 21350
rect 33324 21286 33376 21292
rect 33322 21176 33378 21185
rect 33322 21111 33378 21120
rect 33232 20528 33284 20534
rect 33232 20470 33284 20476
rect 33232 20392 33284 20398
rect 33336 20369 33364 21111
rect 33232 20334 33284 20340
rect 33322 20360 33378 20369
rect 33244 19802 33272 20334
rect 33322 20295 33378 20304
rect 33324 20256 33376 20262
rect 33324 20198 33376 20204
rect 33336 19961 33364 20198
rect 33322 19952 33378 19961
rect 33322 19887 33378 19896
rect 33244 19774 33364 19802
rect 33232 19712 33284 19718
rect 33232 19654 33284 19660
rect 33140 18964 33192 18970
rect 33140 18906 33192 18912
rect 32956 18896 33008 18902
rect 32956 18838 33008 18844
rect 33244 18816 33272 19654
rect 33060 18788 33272 18816
rect 33060 18086 33088 18788
rect 33336 18442 33364 19774
rect 33244 18414 33364 18442
rect 33048 18080 33100 18086
rect 33048 18022 33100 18028
rect 33140 17740 33192 17746
rect 33140 17682 33192 17688
rect 33048 17060 33100 17066
rect 33048 17002 33100 17008
rect 33060 16250 33088 17002
rect 33048 16244 33100 16250
rect 33048 16186 33100 16192
rect 33048 16040 33100 16046
rect 33048 15982 33100 15988
rect 32956 15564 33008 15570
rect 32956 15506 33008 15512
rect 32864 14952 32916 14958
rect 32864 14894 32916 14900
rect 32968 14385 32996 15506
rect 32954 14376 33010 14385
rect 32680 14340 32732 14346
rect 32954 14311 33010 14320
rect 32680 14282 32732 14288
rect 33060 13954 33088 15982
rect 33152 15978 33180 17682
rect 33140 15972 33192 15978
rect 33140 15914 33192 15920
rect 33140 15360 33192 15366
rect 33140 15302 33192 15308
rect 33152 14618 33180 15302
rect 33140 14612 33192 14618
rect 33140 14554 33192 14560
rect 33244 14498 33272 18414
rect 33324 18352 33376 18358
rect 33324 18294 33376 18300
rect 33336 16969 33364 18294
rect 33322 16960 33378 16969
rect 33322 16895 33378 16904
rect 33324 16720 33376 16726
rect 33324 16662 33376 16668
rect 33336 16114 33364 16662
rect 33324 16108 33376 16114
rect 33324 16050 33376 16056
rect 33336 15706 33364 16050
rect 33324 15700 33376 15706
rect 33324 15642 33376 15648
rect 33324 14952 33376 14958
rect 33324 14894 33376 14900
rect 33336 14521 33364 14894
rect 32968 13926 33088 13954
rect 33152 14470 33272 14498
rect 33322 14512 33378 14521
rect 32496 13728 32548 13734
rect 32496 13670 32548 13676
rect 32968 12306 32996 13926
rect 33048 13864 33100 13870
rect 33048 13806 33100 13812
rect 32956 12300 33008 12306
rect 32956 12242 33008 12248
rect 32956 11076 33008 11082
rect 32956 11018 33008 11024
rect 32496 9920 32548 9926
rect 32496 9862 32548 9868
rect 32404 5024 32456 5030
rect 32404 4966 32456 4972
rect 32312 3392 32364 3398
rect 32312 3334 32364 3340
rect 32220 2984 32272 2990
rect 32220 2926 32272 2932
rect 32312 2848 32364 2854
rect 32312 2790 32364 2796
rect 32324 800 32352 2790
rect 32508 2582 32536 9862
rect 32968 4214 32996 11018
rect 33060 4826 33088 13806
rect 33048 4820 33100 4826
rect 33048 4762 33100 4768
rect 32956 4208 33008 4214
rect 32956 4150 33008 4156
rect 33152 4146 33180 14470
rect 33322 14447 33324 14456
rect 33376 14447 33378 14456
rect 33324 14418 33376 14424
rect 33232 14340 33284 14346
rect 33232 14282 33284 14288
rect 33324 14340 33376 14346
rect 33324 14282 33376 14288
rect 33140 4140 33192 4146
rect 33140 4082 33192 4088
rect 32588 4072 32640 4078
rect 32588 4014 32640 4020
rect 32496 2576 32548 2582
rect 32496 2518 32548 2524
rect 32600 800 32628 4014
rect 33244 2990 33272 14282
rect 33336 12102 33364 14282
rect 33428 13870 33456 26250
rect 33520 14958 33548 27814
rect 33600 27668 33652 27674
rect 33600 27610 33652 27616
rect 33508 14952 33560 14958
rect 33508 14894 33560 14900
rect 33508 14816 33560 14822
rect 33508 14758 33560 14764
rect 33416 13864 33468 13870
rect 33416 13806 33468 13812
rect 33324 12096 33376 12102
rect 33324 12038 33376 12044
rect 33324 11756 33376 11762
rect 33324 11698 33376 11704
rect 33336 6730 33364 11698
rect 33324 6724 33376 6730
rect 33324 6666 33376 6672
rect 33416 4072 33468 4078
rect 33416 4014 33468 4020
rect 33232 2984 33284 2990
rect 33232 2926 33284 2932
rect 33232 2848 33284 2854
rect 33232 2790 33284 2796
rect 32956 2508 33008 2514
rect 32956 2450 33008 2456
rect 32968 800 32996 2450
rect 33244 800 33272 2790
rect 33428 2650 33456 4014
rect 33520 3942 33548 14758
rect 33612 14482 33640 27610
rect 33704 24886 33732 31198
rect 33784 31136 33836 31142
rect 33784 31078 33836 31084
rect 33692 24880 33744 24886
rect 33692 24822 33744 24828
rect 33692 24744 33744 24750
rect 33692 24686 33744 24692
rect 33704 24070 33732 24686
rect 33692 24064 33744 24070
rect 33692 24006 33744 24012
rect 33692 23180 33744 23186
rect 33692 23122 33744 23128
rect 33704 23089 33732 23122
rect 33690 23080 33746 23089
rect 33690 23015 33746 23024
rect 33692 22976 33744 22982
rect 33692 22918 33744 22924
rect 33704 22001 33732 22918
rect 33690 21992 33746 22001
rect 33690 21927 33746 21936
rect 33692 21888 33744 21894
rect 33692 21830 33744 21836
rect 33704 19174 33732 21830
rect 33692 19168 33744 19174
rect 33692 19110 33744 19116
rect 33600 14476 33652 14482
rect 33600 14418 33652 14424
rect 33704 8974 33732 19110
rect 33796 16250 33824 31078
rect 33876 30048 33928 30054
rect 33876 29990 33928 29996
rect 33888 23089 33916 29990
rect 33874 23080 33930 23089
rect 33874 23015 33930 23024
rect 33876 22976 33928 22982
rect 33876 22918 33928 22924
rect 33888 19922 33916 22918
rect 33876 19916 33928 19922
rect 33876 19858 33928 19864
rect 33874 19816 33930 19825
rect 33874 19751 33930 19760
rect 33888 18358 33916 19751
rect 33876 18352 33928 18358
rect 33876 18294 33928 18300
rect 33876 18216 33928 18222
rect 33876 18158 33928 18164
rect 33784 16244 33836 16250
rect 33784 16186 33836 16192
rect 33784 15904 33836 15910
rect 33784 15846 33836 15852
rect 33796 15366 33824 15846
rect 33784 15360 33836 15366
rect 33784 15302 33836 15308
rect 33796 14890 33824 15302
rect 33784 14884 33836 14890
rect 33784 14826 33836 14832
rect 33796 14618 33824 14826
rect 33784 14612 33836 14618
rect 33784 14554 33836 14560
rect 33784 14476 33836 14482
rect 33784 14418 33836 14424
rect 33692 8968 33744 8974
rect 33692 8910 33744 8916
rect 33796 5302 33824 14418
rect 33888 11762 33916 18158
rect 33980 17105 34008 31962
rect 34072 31142 34100 37606
rect 34060 31136 34112 31142
rect 34060 31078 34112 31084
rect 34164 28994 34192 56102
rect 34256 54874 34284 56222
rect 34244 54868 34296 54874
rect 34244 54810 34296 54816
rect 34244 53440 34296 53446
rect 34244 53382 34296 53388
rect 34256 50862 34284 53382
rect 34244 50856 34296 50862
rect 34244 50798 34296 50804
rect 34244 47116 34296 47122
rect 34244 47058 34296 47064
rect 34256 46442 34284 47058
rect 34244 46436 34296 46442
rect 34244 46378 34296 46384
rect 34256 46034 34284 46378
rect 34348 46170 34376 58006
rect 34440 54806 34468 65418
rect 34520 65204 34572 65210
rect 34520 65146 34572 65152
rect 34532 60246 34560 65146
rect 34624 65074 34652 113834
rect 34716 113082 34744 116690
rect 34808 115598 34836 117286
rect 35268 116822 35296 119200
rect 35346 118280 35402 118289
rect 35346 118215 35402 118224
rect 35256 116816 35308 116822
rect 35256 116758 35308 116764
rect 35360 116634 35388 118215
rect 35452 117230 35480 119200
rect 35622 117464 35678 117473
rect 35622 117399 35678 117408
rect 35440 117224 35492 117230
rect 35440 117166 35492 117172
rect 35530 116920 35586 116929
rect 35530 116855 35586 116864
rect 35440 116748 35492 116754
rect 35440 116690 35492 116696
rect 35268 116606 35388 116634
rect 34940 116444 35236 116464
rect 34996 116442 35020 116444
rect 35076 116442 35100 116444
rect 35156 116442 35180 116444
rect 35018 116390 35020 116442
rect 35082 116390 35094 116442
rect 35156 116390 35158 116442
rect 34996 116388 35020 116390
rect 35076 116388 35100 116390
rect 35156 116388 35180 116390
rect 34940 116368 35236 116388
rect 34888 116136 34940 116142
rect 34888 116078 34940 116084
rect 35162 116104 35218 116113
rect 34796 115592 34848 115598
rect 34796 115534 34848 115540
rect 34900 115444 34928 116078
rect 35162 116039 35218 116048
rect 35176 115569 35204 116039
rect 35268 115682 35296 116606
rect 35346 116512 35402 116521
rect 35346 116447 35402 116456
rect 35360 115802 35388 116447
rect 35348 115796 35400 115802
rect 35348 115738 35400 115744
rect 35268 115654 35388 115682
rect 35162 115560 35218 115569
rect 35162 115495 35218 115504
rect 34808 115416 34928 115444
rect 35256 115456 35308 115462
rect 34808 115138 34836 115416
rect 35256 115398 35308 115404
rect 34940 115356 35236 115376
rect 34996 115354 35020 115356
rect 35076 115354 35100 115356
rect 35156 115354 35180 115356
rect 35018 115302 35020 115354
rect 35082 115302 35094 115354
rect 35156 115302 35158 115354
rect 34996 115300 35020 115302
rect 35076 115300 35100 115302
rect 35156 115300 35180 115302
rect 34940 115280 35236 115300
rect 34808 115110 35204 115138
rect 34796 115048 34848 115054
rect 34796 114990 34848 114996
rect 34808 114578 34836 114990
rect 34796 114572 34848 114578
rect 34796 114514 34848 114520
rect 34808 113642 34836 114514
rect 35176 114356 35204 115110
rect 35268 114918 35296 115398
rect 35360 115258 35388 115654
rect 35348 115252 35400 115258
rect 35348 115194 35400 115200
rect 35346 115152 35402 115161
rect 35346 115087 35402 115096
rect 35256 114912 35308 114918
rect 35256 114854 35308 114860
rect 35176 114328 35296 114356
rect 34940 114268 35236 114288
rect 34996 114266 35020 114268
rect 35076 114266 35100 114268
rect 35156 114266 35180 114268
rect 35018 114214 35020 114266
rect 35082 114214 35094 114266
rect 35156 114214 35158 114266
rect 34996 114212 35020 114214
rect 35076 114212 35100 114214
rect 35156 114212 35180 114214
rect 34940 114192 35236 114212
rect 35268 114102 35296 114328
rect 35256 114096 35308 114102
rect 35256 114038 35308 114044
rect 34808 113614 34928 113642
rect 34900 113558 34928 113614
rect 34888 113552 34940 113558
rect 34888 113494 34940 113500
rect 35256 113552 35308 113558
rect 35256 113494 35308 113500
rect 34796 113484 34848 113490
rect 34796 113426 34848 113432
rect 34704 113076 34756 113082
rect 34704 113018 34756 113024
rect 34808 112878 34836 113426
rect 34940 113180 35236 113200
rect 34996 113178 35020 113180
rect 35076 113178 35100 113180
rect 35156 113178 35180 113180
rect 35018 113126 35020 113178
rect 35082 113126 35094 113178
rect 35156 113126 35158 113178
rect 34996 113124 35020 113126
rect 35076 113124 35100 113126
rect 35156 113124 35180 113126
rect 34940 113104 35236 113124
rect 35268 112946 35296 113494
rect 35256 112940 35308 112946
rect 35256 112882 35308 112888
rect 34796 112872 34848 112878
rect 34796 112814 34848 112820
rect 34704 112736 34756 112742
rect 34704 112678 34756 112684
rect 34716 110090 34744 112678
rect 34940 112092 35236 112112
rect 34996 112090 35020 112092
rect 35076 112090 35100 112092
rect 35156 112090 35180 112092
rect 35018 112038 35020 112090
rect 35082 112038 35094 112090
rect 35156 112038 35158 112090
rect 34996 112036 35020 112038
rect 35076 112036 35100 112038
rect 35156 112036 35180 112038
rect 34940 112016 35236 112036
rect 34796 111852 34848 111858
rect 34796 111794 34848 111800
rect 34704 110084 34756 110090
rect 34704 110026 34756 110032
rect 34808 109614 34836 111794
rect 34940 111004 35236 111024
rect 34996 111002 35020 111004
rect 35076 111002 35100 111004
rect 35156 111002 35180 111004
rect 35018 110950 35020 111002
rect 35082 110950 35094 111002
rect 35156 110950 35158 111002
rect 34996 110948 35020 110950
rect 35076 110948 35100 110950
rect 35156 110948 35180 110950
rect 34940 110928 35236 110948
rect 34940 109916 35236 109936
rect 34996 109914 35020 109916
rect 35076 109914 35100 109916
rect 35156 109914 35180 109916
rect 35018 109862 35020 109914
rect 35082 109862 35094 109914
rect 35156 109862 35158 109914
rect 34996 109860 35020 109862
rect 35076 109860 35100 109862
rect 35156 109860 35180 109862
rect 34940 109840 35236 109860
rect 34796 109608 34848 109614
rect 34796 109550 34848 109556
rect 34808 109138 34836 109550
rect 34796 109132 34848 109138
rect 34796 109074 34848 109080
rect 34900 109070 34928 109117
rect 34888 109064 34940 109070
rect 34808 109012 34888 109034
rect 35268 109034 35296 112882
rect 35360 112402 35388 115087
rect 35348 112396 35400 112402
rect 35348 112338 35400 112344
rect 35348 112260 35400 112266
rect 35348 112202 35400 112208
rect 34940 109012 35296 109034
rect 34808 109006 35296 109012
rect 34704 105800 34756 105806
rect 34704 105742 34756 105748
rect 34716 87310 34744 105742
rect 34808 104378 34836 109006
rect 34940 108828 35236 108848
rect 34996 108826 35020 108828
rect 35076 108826 35100 108828
rect 35156 108826 35180 108828
rect 35018 108774 35020 108826
rect 35082 108774 35094 108826
rect 35156 108774 35158 108826
rect 34996 108772 35020 108774
rect 35076 108772 35100 108774
rect 35156 108772 35180 108774
rect 34940 108752 35236 108772
rect 35256 107840 35308 107846
rect 35256 107782 35308 107788
rect 34940 107740 35236 107760
rect 34996 107738 35020 107740
rect 35076 107738 35100 107740
rect 35156 107738 35180 107740
rect 35018 107686 35020 107738
rect 35082 107686 35094 107738
rect 35156 107686 35158 107738
rect 34996 107684 35020 107686
rect 35076 107684 35100 107686
rect 35156 107684 35180 107686
rect 34940 107664 35236 107684
rect 34940 106652 35236 106672
rect 34996 106650 35020 106652
rect 35076 106650 35100 106652
rect 35156 106650 35180 106652
rect 35018 106598 35020 106650
rect 35082 106598 35094 106650
rect 35156 106598 35158 106650
rect 34996 106596 35020 106598
rect 35076 106596 35100 106598
rect 35156 106596 35180 106598
rect 34940 106576 35236 106596
rect 35268 105942 35296 107782
rect 35256 105936 35308 105942
rect 35256 105878 35308 105884
rect 34940 105564 35236 105584
rect 34996 105562 35020 105564
rect 35076 105562 35100 105564
rect 35156 105562 35180 105564
rect 35018 105510 35020 105562
rect 35082 105510 35094 105562
rect 35156 105510 35158 105562
rect 34996 105508 35020 105510
rect 35076 105508 35100 105510
rect 35156 105508 35180 105510
rect 34940 105488 35236 105508
rect 34940 104476 35236 104496
rect 34996 104474 35020 104476
rect 35076 104474 35100 104476
rect 35156 104474 35180 104476
rect 35018 104422 35020 104474
rect 35082 104422 35094 104474
rect 35156 104422 35158 104474
rect 34996 104420 35020 104422
rect 35076 104420 35100 104422
rect 35156 104420 35180 104422
rect 34940 104400 35236 104420
rect 34796 104372 34848 104378
rect 34796 104314 34848 104320
rect 34940 103388 35236 103408
rect 34996 103386 35020 103388
rect 35076 103386 35100 103388
rect 35156 103386 35180 103388
rect 35018 103334 35020 103386
rect 35082 103334 35094 103386
rect 35156 103334 35158 103386
rect 34996 103332 35020 103334
rect 35076 103332 35100 103334
rect 35156 103332 35180 103334
rect 34940 103312 35236 103332
rect 34940 102300 35236 102320
rect 34996 102298 35020 102300
rect 35076 102298 35100 102300
rect 35156 102298 35180 102300
rect 35018 102246 35020 102298
rect 35082 102246 35094 102298
rect 35156 102246 35158 102298
rect 34996 102244 35020 102246
rect 35076 102244 35100 102246
rect 35156 102244 35180 102246
rect 34940 102224 35236 102244
rect 34940 101212 35236 101232
rect 34996 101210 35020 101212
rect 35076 101210 35100 101212
rect 35156 101210 35180 101212
rect 35018 101158 35020 101210
rect 35082 101158 35094 101210
rect 35156 101158 35158 101210
rect 34996 101156 35020 101158
rect 35076 101156 35100 101158
rect 35156 101156 35180 101158
rect 34940 101136 35236 101156
rect 34940 100124 35236 100144
rect 34996 100122 35020 100124
rect 35076 100122 35100 100124
rect 35156 100122 35180 100124
rect 35018 100070 35020 100122
rect 35082 100070 35094 100122
rect 35156 100070 35158 100122
rect 34996 100068 35020 100070
rect 35076 100068 35100 100070
rect 35156 100068 35180 100070
rect 34940 100048 35236 100068
rect 34796 99136 34848 99142
rect 34796 99078 34848 99084
rect 34808 89894 34836 99078
rect 34940 99036 35236 99056
rect 34996 99034 35020 99036
rect 35076 99034 35100 99036
rect 35156 99034 35180 99036
rect 35018 98982 35020 99034
rect 35082 98982 35094 99034
rect 35156 98982 35158 99034
rect 34996 98980 35020 98982
rect 35076 98980 35100 98982
rect 35156 98980 35180 98982
rect 34940 98960 35236 98980
rect 35360 98938 35388 112202
rect 35452 109818 35480 116690
rect 35544 115190 35572 116855
rect 35532 115184 35584 115190
rect 35532 115126 35584 115132
rect 35532 114980 35584 114986
rect 35532 114922 35584 114928
rect 35544 114578 35572 114922
rect 35532 114572 35584 114578
rect 35532 114514 35584 114520
rect 35544 114170 35572 114514
rect 35532 114164 35584 114170
rect 35532 114106 35584 114112
rect 35544 113422 35572 114106
rect 35532 113416 35584 113422
rect 35532 113358 35584 113364
rect 35636 112962 35664 117399
rect 35728 117314 35756 119200
rect 35912 117450 35940 119200
rect 35912 117422 36032 117450
rect 35728 117286 35940 117314
rect 35912 116346 35940 117286
rect 35716 116340 35768 116346
rect 35716 116282 35768 116288
rect 35900 116340 35952 116346
rect 35900 116282 35952 116288
rect 35728 115802 35756 116282
rect 35808 116068 35860 116074
rect 35808 116010 35860 116016
rect 35716 115796 35768 115802
rect 35716 115738 35768 115744
rect 35716 115660 35768 115666
rect 35716 115602 35768 115608
rect 35728 114578 35756 115602
rect 35716 114572 35768 114578
rect 35716 114514 35768 114520
rect 35820 113626 35848 116010
rect 36004 115818 36032 117422
rect 36096 116142 36124 119575
rect 36174 119200 36230 120800
rect 36358 119200 36414 120800
rect 36634 119200 36690 120800
rect 36818 119200 36874 120800
rect 37094 119200 37150 120800
rect 37186 119232 37242 119241
rect 36084 116136 36136 116142
rect 36084 116078 36136 116084
rect 35912 115790 36032 115818
rect 35912 114714 35940 115790
rect 36188 115734 36216 119200
rect 36372 116754 36400 119200
rect 36452 117088 36504 117094
rect 36452 117030 36504 117036
rect 36544 117088 36596 117094
rect 36544 117030 36596 117036
rect 36360 116748 36412 116754
rect 36360 116690 36412 116696
rect 36268 116680 36320 116686
rect 36268 116622 36320 116628
rect 36176 115728 36228 115734
rect 36176 115670 36228 115676
rect 35992 115660 36044 115666
rect 35992 115602 36044 115608
rect 35900 114708 35952 114714
rect 35900 114650 35952 114656
rect 35808 113620 35860 113626
rect 35808 113562 35860 113568
rect 35716 113484 35768 113490
rect 35716 113426 35768 113432
rect 35544 112934 35664 112962
rect 35544 112538 35572 112934
rect 35624 112872 35676 112878
rect 35624 112814 35676 112820
rect 35532 112532 35584 112538
rect 35532 112474 35584 112480
rect 35636 111790 35664 112814
rect 35624 111784 35676 111790
rect 35624 111726 35676 111732
rect 35532 111716 35584 111722
rect 35532 111658 35584 111664
rect 35544 111314 35572 111658
rect 35636 111382 35664 111726
rect 35624 111376 35676 111382
rect 35624 111318 35676 111324
rect 35532 111308 35584 111314
rect 35532 111250 35584 111256
rect 35440 109812 35492 109818
rect 35440 109754 35492 109760
rect 35438 109712 35494 109721
rect 35438 109647 35494 109656
rect 35452 108594 35480 109647
rect 35440 108588 35492 108594
rect 35440 108530 35492 108536
rect 35544 108390 35572 111250
rect 35532 108384 35584 108390
rect 35532 108326 35584 108332
rect 35636 108202 35664 111318
rect 35452 108174 35664 108202
rect 35452 107574 35480 108174
rect 35440 107568 35492 107574
rect 35440 107510 35492 107516
rect 35452 105874 35480 107510
rect 35624 107364 35676 107370
rect 35624 107306 35676 107312
rect 35532 106752 35584 106758
rect 35532 106694 35584 106700
rect 35440 105868 35492 105874
rect 35440 105810 35492 105816
rect 35440 105664 35492 105670
rect 35440 105606 35492 105612
rect 35348 98932 35400 98938
rect 35348 98874 35400 98880
rect 35452 98818 35480 105606
rect 35268 98790 35480 98818
rect 34940 97948 35236 97968
rect 34996 97946 35020 97948
rect 35076 97946 35100 97948
rect 35156 97946 35180 97948
rect 35018 97894 35020 97946
rect 35082 97894 35094 97946
rect 35156 97894 35158 97946
rect 34996 97892 35020 97894
rect 35076 97892 35100 97894
rect 35156 97892 35180 97894
rect 34940 97872 35236 97892
rect 34940 96860 35236 96880
rect 34996 96858 35020 96860
rect 35076 96858 35100 96860
rect 35156 96858 35180 96860
rect 35018 96806 35020 96858
rect 35082 96806 35094 96858
rect 35156 96806 35158 96858
rect 34996 96804 35020 96806
rect 35076 96804 35100 96806
rect 35156 96804 35180 96806
rect 34940 96784 35236 96804
rect 34940 95772 35236 95792
rect 34996 95770 35020 95772
rect 35076 95770 35100 95772
rect 35156 95770 35180 95772
rect 35018 95718 35020 95770
rect 35082 95718 35094 95770
rect 35156 95718 35158 95770
rect 34996 95716 35020 95718
rect 35076 95716 35100 95718
rect 35156 95716 35180 95718
rect 34940 95696 35236 95716
rect 35268 94858 35296 98790
rect 35348 98660 35400 98666
rect 35348 98602 35400 98608
rect 35256 94852 35308 94858
rect 35256 94794 35308 94800
rect 34940 94684 35236 94704
rect 34996 94682 35020 94684
rect 35076 94682 35100 94684
rect 35156 94682 35180 94684
rect 35018 94630 35020 94682
rect 35082 94630 35094 94682
rect 35156 94630 35158 94682
rect 34996 94628 35020 94630
rect 35076 94628 35100 94630
rect 35156 94628 35180 94630
rect 34940 94608 35236 94628
rect 35256 94512 35308 94518
rect 35256 94454 35308 94460
rect 34940 93596 35236 93616
rect 34996 93594 35020 93596
rect 35076 93594 35100 93596
rect 35156 93594 35180 93596
rect 35018 93542 35020 93594
rect 35082 93542 35094 93594
rect 35156 93542 35158 93594
rect 34996 93540 35020 93542
rect 35076 93540 35100 93542
rect 35156 93540 35180 93542
rect 34940 93520 35236 93540
rect 34940 92508 35236 92528
rect 34996 92506 35020 92508
rect 35076 92506 35100 92508
rect 35156 92506 35180 92508
rect 35018 92454 35020 92506
rect 35082 92454 35094 92506
rect 35156 92454 35158 92506
rect 34996 92452 35020 92454
rect 35076 92452 35100 92454
rect 35156 92452 35180 92454
rect 34940 92432 35236 92452
rect 34940 91420 35236 91440
rect 34996 91418 35020 91420
rect 35076 91418 35100 91420
rect 35156 91418 35180 91420
rect 35018 91366 35020 91418
rect 35082 91366 35094 91418
rect 35156 91366 35158 91418
rect 34996 91364 35020 91366
rect 35076 91364 35100 91366
rect 35156 91364 35180 91366
rect 34940 91344 35236 91364
rect 34940 90332 35236 90352
rect 34996 90330 35020 90332
rect 35076 90330 35100 90332
rect 35156 90330 35180 90332
rect 35018 90278 35020 90330
rect 35082 90278 35094 90330
rect 35156 90278 35158 90330
rect 34996 90276 35020 90278
rect 35076 90276 35100 90278
rect 35156 90276 35180 90278
rect 34940 90256 35236 90276
rect 35164 90160 35216 90166
rect 35164 90102 35216 90108
rect 34888 90092 34940 90098
rect 34888 90034 34940 90040
rect 34796 89888 34848 89894
rect 34796 89830 34848 89836
rect 34900 89714 34928 90034
rect 34808 89686 34928 89714
rect 35176 89714 35204 90102
rect 35268 89962 35296 94454
rect 35256 89956 35308 89962
rect 35256 89898 35308 89904
rect 35176 89686 35296 89714
rect 34704 87304 34756 87310
rect 34808 87281 34836 89686
rect 34940 89244 35236 89264
rect 34996 89242 35020 89244
rect 35076 89242 35100 89244
rect 35156 89242 35180 89244
rect 35018 89190 35020 89242
rect 35082 89190 35094 89242
rect 35156 89190 35158 89242
rect 34996 89188 35020 89190
rect 35076 89188 35100 89190
rect 35156 89188 35180 89190
rect 34940 89168 35236 89188
rect 34940 88156 35236 88176
rect 34996 88154 35020 88156
rect 35076 88154 35100 88156
rect 35156 88154 35180 88156
rect 35018 88102 35020 88154
rect 35082 88102 35094 88154
rect 35156 88102 35158 88154
rect 34996 88100 35020 88102
rect 35076 88100 35100 88102
rect 35156 88100 35180 88102
rect 34940 88080 35236 88100
rect 35268 87854 35296 89686
rect 35256 87848 35308 87854
rect 35256 87790 35308 87796
rect 35256 87712 35308 87718
rect 35256 87654 35308 87660
rect 34704 87246 34756 87252
rect 34794 87272 34850 87281
rect 34794 87207 34850 87216
rect 34704 87168 34756 87174
rect 34704 87110 34756 87116
rect 34612 65068 34664 65074
rect 34612 65010 34664 65016
rect 34612 64864 34664 64870
rect 34612 64806 34664 64812
rect 34624 64025 34652 64806
rect 34610 64016 34666 64025
rect 34610 63951 34666 63960
rect 34612 63776 34664 63782
rect 34612 63718 34664 63724
rect 34624 62898 34652 63718
rect 34612 62892 34664 62898
rect 34612 62834 34664 62840
rect 34520 60240 34572 60246
rect 34520 60182 34572 60188
rect 34520 60036 34572 60042
rect 34520 59978 34572 59984
rect 34428 54800 34480 54806
rect 34428 54742 34480 54748
rect 34532 50386 34560 59978
rect 34612 51264 34664 51270
rect 34612 51206 34664 51212
rect 34520 50380 34572 50386
rect 34520 50322 34572 50328
rect 34532 49774 34560 50322
rect 34520 49768 34572 49774
rect 34520 49710 34572 49716
rect 34520 49088 34572 49094
rect 34520 49030 34572 49036
rect 34428 46980 34480 46986
rect 34428 46922 34480 46928
rect 34440 46374 34468 46922
rect 34532 46510 34560 49030
rect 34624 48142 34652 51206
rect 34612 48136 34664 48142
rect 34612 48078 34664 48084
rect 34612 48000 34664 48006
rect 34612 47942 34664 47948
rect 34520 46504 34572 46510
rect 34520 46446 34572 46452
rect 34428 46368 34480 46374
rect 34428 46310 34480 46316
rect 34520 46368 34572 46374
rect 34520 46310 34572 46316
rect 34336 46164 34388 46170
rect 34336 46106 34388 46112
rect 34440 46050 34468 46310
rect 34348 46034 34468 46050
rect 34244 46028 34296 46034
rect 34244 45970 34296 45976
rect 34336 46028 34468 46034
rect 34388 46022 34468 46028
rect 34336 45970 34388 45976
rect 34256 45354 34284 45970
rect 34348 45354 34376 45970
rect 34244 45348 34296 45354
rect 34244 45290 34296 45296
rect 34336 45348 34388 45354
rect 34336 45290 34388 45296
rect 34256 44402 34284 45290
rect 34348 44470 34376 45290
rect 34336 44464 34388 44470
rect 34336 44406 34388 44412
rect 34244 44396 34296 44402
rect 34244 44338 34296 44344
rect 34244 43988 34296 43994
rect 34244 43930 34296 43936
rect 34072 28966 34192 28994
rect 34072 22710 34100 28966
rect 34152 27872 34204 27878
rect 34152 27814 34204 27820
rect 34164 26314 34192 27814
rect 34256 27470 34284 43930
rect 34428 42560 34480 42566
rect 34428 42502 34480 42508
rect 34336 42016 34388 42022
rect 34336 41958 34388 41964
rect 34348 38554 34376 41958
rect 34440 41682 34468 42502
rect 34428 41676 34480 41682
rect 34428 41618 34480 41624
rect 34428 39296 34480 39302
rect 34428 39238 34480 39244
rect 34336 38548 34388 38554
rect 34336 38490 34388 38496
rect 34336 38412 34388 38418
rect 34336 38354 34388 38360
rect 34348 36650 34376 38354
rect 34440 37346 34468 39238
rect 34532 38418 34560 46310
rect 34624 46034 34652 47942
rect 34612 46028 34664 46034
rect 34612 45970 34664 45976
rect 34612 45348 34664 45354
rect 34612 45290 34664 45296
rect 34520 38412 34572 38418
rect 34520 38354 34572 38360
rect 34532 37466 34560 38354
rect 34520 37460 34572 37466
rect 34520 37402 34572 37408
rect 34440 37318 34560 37346
rect 34428 37256 34480 37262
rect 34428 37198 34480 37204
rect 34336 36644 34388 36650
rect 34336 36586 34388 36592
rect 34348 35494 34376 36586
rect 34440 35562 34468 37198
rect 34428 35556 34480 35562
rect 34428 35498 34480 35504
rect 34336 35488 34388 35494
rect 34336 35430 34388 35436
rect 34244 27464 34296 27470
rect 34244 27406 34296 27412
rect 34244 27328 34296 27334
rect 34244 27270 34296 27276
rect 34256 26450 34284 27270
rect 34244 26444 34296 26450
rect 34244 26386 34296 26392
rect 34348 26382 34376 35430
rect 34440 35222 34468 35498
rect 34428 35216 34480 35222
rect 34428 35158 34480 35164
rect 34428 34944 34480 34950
rect 34428 34886 34480 34892
rect 34440 32434 34468 34886
rect 34428 32428 34480 32434
rect 34428 32370 34480 32376
rect 34428 30592 34480 30598
rect 34428 30534 34480 30540
rect 34440 29238 34468 30534
rect 34428 29232 34480 29238
rect 34428 29174 34480 29180
rect 34428 27464 34480 27470
rect 34428 27406 34480 27412
rect 34336 26376 34388 26382
rect 34336 26318 34388 26324
rect 34152 26308 34204 26314
rect 34152 26250 34204 26256
rect 34164 25362 34192 26250
rect 34440 26234 34468 27406
rect 34348 26206 34468 26234
rect 34242 25528 34298 25537
rect 34242 25463 34298 25472
rect 34256 25430 34284 25463
rect 34244 25424 34296 25430
rect 34244 25366 34296 25372
rect 34152 25356 34204 25362
rect 34152 25298 34204 25304
rect 34164 24818 34192 25298
rect 34244 25152 34296 25158
rect 34244 25094 34296 25100
rect 34152 24812 34204 24818
rect 34152 24754 34204 24760
rect 34152 24608 34204 24614
rect 34152 24550 34204 24556
rect 34164 23254 34192 24550
rect 34256 24410 34284 25094
rect 34348 24585 34376 26206
rect 34428 25900 34480 25906
rect 34428 25842 34480 25848
rect 34440 25362 34468 25842
rect 34428 25356 34480 25362
rect 34428 25298 34480 25304
rect 34440 25226 34468 25298
rect 34532 25265 34560 37318
rect 34624 31754 34652 45290
rect 34716 36417 34744 87110
rect 34940 87068 35236 87088
rect 34996 87066 35020 87068
rect 35076 87066 35100 87068
rect 35156 87066 35180 87068
rect 35018 87014 35020 87066
rect 35082 87014 35094 87066
rect 35156 87014 35158 87066
rect 34996 87012 35020 87014
rect 35076 87012 35100 87014
rect 35156 87012 35180 87014
rect 34794 87000 34850 87009
rect 34940 86992 35236 87012
rect 34794 86935 34850 86944
rect 34808 86834 34836 86935
rect 34796 86828 34848 86834
rect 34796 86770 34848 86776
rect 34796 86692 34848 86698
rect 34796 86634 34848 86640
rect 34808 83910 34836 86634
rect 34940 85980 35236 86000
rect 34996 85978 35020 85980
rect 35076 85978 35100 85980
rect 35156 85978 35180 85980
rect 35018 85926 35020 85978
rect 35082 85926 35094 85978
rect 35156 85926 35158 85978
rect 34996 85924 35020 85926
rect 35076 85924 35100 85926
rect 35156 85924 35180 85926
rect 34940 85904 35236 85924
rect 34940 84892 35236 84912
rect 34996 84890 35020 84892
rect 35076 84890 35100 84892
rect 35156 84890 35180 84892
rect 35018 84838 35020 84890
rect 35082 84838 35094 84890
rect 35156 84838 35158 84890
rect 34996 84836 35020 84838
rect 35076 84836 35100 84838
rect 35156 84836 35180 84838
rect 34940 84816 35236 84836
rect 34796 83904 34848 83910
rect 34796 83846 34848 83852
rect 34940 83804 35236 83824
rect 34996 83802 35020 83804
rect 35076 83802 35100 83804
rect 35156 83802 35180 83804
rect 35018 83750 35020 83802
rect 35082 83750 35094 83802
rect 35156 83750 35158 83802
rect 34996 83748 35020 83750
rect 35076 83748 35100 83750
rect 35156 83748 35180 83750
rect 34940 83728 35236 83748
rect 34940 82716 35236 82736
rect 34996 82714 35020 82716
rect 35076 82714 35100 82716
rect 35156 82714 35180 82716
rect 35018 82662 35020 82714
rect 35082 82662 35094 82714
rect 35156 82662 35158 82714
rect 34996 82660 35020 82662
rect 35076 82660 35100 82662
rect 35156 82660 35180 82662
rect 34940 82640 35236 82660
rect 34940 81628 35236 81648
rect 34996 81626 35020 81628
rect 35076 81626 35100 81628
rect 35156 81626 35180 81628
rect 35018 81574 35020 81626
rect 35082 81574 35094 81626
rect 35156 81574 35158 81626
rect 34996 81572 35020 81574
rect 35076 81572 35100 81574
rect 35156 81572 35180 81574
rect 34940 81552 35236 81572
rect 34940 80540 35236 80560
rect 34996 80538 35020 80540
rect 35076 80538 35100 80540
rect 35156 80538 35180 80540
rect 35018 80486 35020 80538
rect 35082 80486 35094 80538
rect 35156 80486 35158 80538
rect 34996 80484 35020 80486
rect 35076 80484 35100 80486
rect 35156 80484 35180 80486
rect 34940 80464 35236 80484
rect 35268 80054 35296 87654
rect 34808 80026 35296 80054
rect 34808 73166 34836 80026
rect 34940 79452 35236 79472
rect 34996 79450 35020 79452
rect 35076 79450 35100 79452
rect 35156 79450 35180 79452
rect 35018 79398 35020 79450
rect 35082 79398 35094 79450
rect 35156 79398 35158 79450
rect 34996 79396 35020 79398
rect 35076 79396 35100 79398
rect 35156 79396 35180 79398
rect 34940 79376 35236 79396
rect 34940 78364 35236 78384
rect 34996 78362 35020 78364
rect 35076 78362 35100 78364
rect 35156 78362 35180 78364
rect 35018 78310 35020 78362
rect 35082 78310 35094 78362
rect 35156 78310 35158 78362
rect 34996 78308 35020 78310
rect 35076 78308 35100 78310
rect 35156 78308 35180 78310
rect 34940 78288 35236 78308
rect 34940 77276 35236 77296
rect 34996 77274 35020 77276
rect 35076 77274 35100 77276
rect 35156 77274 35180 77276
rect 35018 77222 35020 77274
rect 35082 77222 35094 77274
rect 35156 77222 35158 77274
rect 34996 77220 35020 77222
rect 35076 77220 35100 77222
rect 35156 77220 35180 77222
rect 34940 77200 35236 77220
rect 34940 76188 35236 76208
rect 34996 76186 35020 76188
rect 35076 76186 35100 76188
rect 35156 76186 35180 76188
rect 35018 76134 35020 76186
rect 35082 76134 35094 76186
rect 35156 76134 35158 76186
rect 34996 76132 35020 76134
rect 35076 76132 35100 76134
rect 35156 76132 35180 76134
rect 34940 76112 35236 76132
rect 35256 75948 35308 75954
rect 35256 75890 35308 75896
rect 34940 75100 35236 75120
rect 34996 75098 35020 75100
rect 35076 75098 35100 75100
rect 35156 75098 35180 75100
rect 35018 75046 35020 75098
rect 35082 75046 35094 75098
rect 35156 75046 35158 75098
rect 34996 75044 35020 75046
rect 35076 75044 35100 75046
rect 35156 75044 35180 75046
rect 34940 75024 35236 75044
rect 34940 74012 35236 74032
rect 34996 74010 35020 74012
rect 35076 74010 35100 74012
rect 35156 74010 35180 74012
rect 35018 73958 35020 74010
rect 35082 73958 35094 74010
rect 35156 73958 35158 74010
rect 34996 73956 35020 73958
rect 35076 73956 35100 73958
rect 35156 73956 35180 73958
rect 34940 73936 35236 73956
rect 34796 73160 34848 73166
rect 34796 73102 34848 73108
rect 34940 72924 35236 72944
rect 34996 72922 35020 72924
rect 35076 72922 35100 72924
rect 35156 72922 35180 72924
rect 35018 72870 35020 72922
rect 35082 72870 35094 72922
rect 35156 72870 35158 72922
rect 34996 72868 35020 72870
rect 35076 72868 35100 72870
rect 35156 72868 35180 72870
rect 34940 72848 35236 72868
rect 34940 71836 35236 71856
rect 34996 71834 35020 71836
rect 35076 71834 35100 71836
rect 35156 71834 35180 71836
rect 35018 71782 35020 71834
rect 35082 71782 35094 71834
rect 35156 71782 35158 71834
rect 34996 71780 35020 71782
rect 35076 71780 35100 71782
rect 35156 71780 35180 71782
rect 34940 71760 35236 71780
rect 34940 70748 35236 70768
rect 34996 70746 35020 70748
rect 35076 70746 35100 70748
rect 35156 70746 35180 70748
rect 35018 70694 35020 70746
rect 35082 70694 35094 70746
rect 35156 70694 35158 70746
rect 34996 70692 35020 70694
rect 35076 70692 35100 70694
rect 35156 70692 35180 70694
rect 34940 70672 35236 70692
rect 34940 69660 35236 69680
rect 34996 69658 35020 69660
rect 35076 69658 35100 69660
rect 35156 69658 35180 69660
rect 35018 69606 35020 69658
rect 35082 69606 35094 69658
rect 35156 69606 35158 69658
rect 34996 69604 35020 69606
rect 35076 69604 35100 69606
rect 35156 69604 35180 69606
rect 34940 69584 35236 69604
rect 34940 68572 35236 68592
rect 34996 68570 35020 68572
rect 35076 68570 35100 68572
rect 35156 68570 35180 68572
rect 35018 68518 35020 68570
rect 35082 68518 35094 68570
rect 35156 68518 35158 68570
rect 34996 68516 35020 68518
rect 35076 68516 35100 68518
rect 35156 68516 35180 68518
rect 34940 68496 35236 68516
rect 34940 67484 35236 67504
rect 34996 67482 35020 67484
rect 35076 67482 35100 67484
rect 35156 67482 35180 67484
rect 35018 67430 35020 67482
rect 35082 67430 35094 67482
rect 35156 67430 35158 67482
rect 34996 67428 35020 67430
rect 35076 67428 35100 67430
rect 35156 67428 35180 67430
rect 34940 67408 35236 67428
rect 34794 66872 34850 66881
rect 34794 66807 34850 66816
rect 34808 66706 34836 66807
rect 34796 66700 34848 66706
rect 34796 66642 34848 66648
rect 34940 66396 35236 66416
rect 34996 66394 35020 66396
rect 35076 66394 35100 66396
rect 35156 66394 35180 66396
rect 35018 66342 35020 66394
rect 35082 66342 35094 66394
rect 35156 66342 35158 66394
rect 34996 66340 35020 66342
rect 35076 66340 35100 66342
rect 35156 66340 35180 66342
rect 34940 66320 35236 66340
rect 35072 65612 35124 65618
rect 35072 65554 35124 65560
rect 35084 65521 35112 65554
rect 35070 65512 35126 65521
rect 35070 65447 35126 65456
rect 34796 65408 34848 65414
rect 34796 65350 34848 65356
rect 34808 65192 34836 65350
rect 34940 65308 35236 65328
rect 34996 65306 35020 65308
rect 35076 65306 35100 65308
rect 35156 65306 35180 65308
rect 35018 65254 35020 65306
rect 35082 65254 35094 65306
rect 35156 65254 35158 65306
rect 34996 65252 35020 65254
rect 35076 65252 35100 65254
rect 35156 65252 35180 65254
rect 34940 65232 35236 65252
rect 34808 65164 34928 65192
rect 34794 65104 34850 65113
rect 34794 65039 34850 65048
rect 34808 65006 34836 65039
rect 34796 65000 34848 65006
rect 34796 64942 34848 64948
rect 34796 64864 34848 64870
rect 34796 64806 34848 64812
rect 34808 64002 34836 64806
rect 34900 64530 34928 65164
rect 35164 65068 35216 65074
rect 35164 65010 35216 65016
rect 35070 64968 35126 64977
rect 35070 64903 35126 64912
rect 35084 64598 35112 64903
rect 35176 64648 35204 65010
rect 35268 64841 35296 75890
rect 35360 69222 35388 98602
rect 35440 98592 35492 98598
rect 35440 98534 35492 98540
rect 35452 94790 35480 98534
rect 35440 94784 35492 94790
rect 35440 94726 35492 94732
rect 35440 94376 35492 94382
rect 35440 94318 35492 94324
rect 35452 90098 35480 94318
rect 35440 90092 35492 90098
rect 35440 90034 35492 90040
rect 35440 89888 35492 89894
rect 35440 89830 35492 89836
rect 35452 87378 35480 89830
rect 35440 87372 35492 87378
rect 35440 87314 35492 87320
rect 35440 86828 35492 86834
rect 35440 86770 35492 86776
rect 35348 69216 35400 69222
rect 35348 69158 35400 69164
rect 35346 68504 35402 68513
rect 35346 68439 35402 68448
rect 35360 67930 35388 68439
rect 35348 67924 35400 67930
rect 35348 67866 35400 67872
rect 35348 66700 35400 66706
rect 35348 66642 35400 66648
rect 35360 66473 35388 66642
rect 35346 66464 35402 66473
rect 35346 66399 35402 66408
rect 35452 66254 35480 86770
rect 35544 83978 35572 106694
rect 35636 94518 35664 107306
rect 35624 94512 35676 94518
rect 35624 94454 35676 94460
rect 35624 93152 35676 93158
rect 35624 93094 35676 93100
rect 35636 91594 35664 93094
rect 35624 91588 35676 91594
rect 35624 91530 35676 91536
rect 35624 88392 35676 88398
rect 35624 88334 35676 88340
rect 35636 86834 35664 88334
rect 35624 86828 35676 86834
rect 35624 86770 35676 86776
rect 35624 86624 35676 86630
rect 35624 86566 35676 86572
rect 35636 85610 35664 86566
rect 35624 85604 35676 85610
rect 35624 85546 35676 85552
rect 35532 83972 35584 83978
rect 35532 83914 35584 83920
rect 35532 82272 35584 82278
rect 35532 82214 35584 82220
rect 35360 66226 35480 66254
rect 35360 64870 35388 66226
rect 35544 65550 35572 82214
rect 35728 80084 35756 113426
rect 35808 113416 35860 113422
rect 35808 113358 35860 113364
rect 35820 110129 35848 113358
rect 35900 112192 35952 112198
rect 35900 112134 35952 112140
rect 35806 110120 35862 110129
rect 35806 110055 35862 110064
rect 35808 110016 35860 110022
rect 35808 109958 35860 109964
rect 35820 109818 35848 109958
rect 35808 109812 35860 109818
rect 35808 109754 35860 109760
rect 35912 109682 35940 112134
rect 36004 111450 36032 115602
rect 36084 115048 36136 115054
rect 36084 114990 36136 114996
rect 36096 114442 36124 114990
rect 36280 114714 36308 116622
rect 36360 116272 36412 116278
rect 36360 116214 36412 116220
rect 36372 115734 36400 116214
rect 36360 115728 36412 115734
rect 36360 115670 36412 115676
rect 36360 115524 36412 115530
rect 36360 115466 36412 115472
rect 36268 114708 36320 114714
rect 36268 114650 36320 114656
rect 36176 114572 36228 114578
rect 36176 114514 36228 114520
rect 36084 114436 36136 114442
rect 36084 114378 36136 114384
rect 36084 113960 36136 113966
rect 36188 113914 36216 114514
rect 36268 114436 36320 114442
rect 36268 114378 36320 114384
rect 36280 113966 36308 114378
rect 36136 113908 36216 113914
rect 36084 113902 36216 113908
rect 36268 113960 36320 113966
rect 36268 113902 36320 113908
rect 36096 113886 36216 113902
rect 36084 112396 36136 112402
rect 36084 112338 36136 112344
rect 35992 111444 36044 111450
rect 35992 111386 36044 111392
rect 36096 110634 36124 112338
rect 36188 111722 36216 113886
rect 36280 113082 36308 113902
rect 36268 113076 36320 113082
rect 36268 113018 36320 113024
rect 36268 112804 36320 112810
rect 36268 112746 36320 112752
rect 36176 111716 36228 111722
rect 36176 111658 36228 111664
rect 36084 110628 36136 110634
rect 36084 110570 36136 110576
rect 35900 109676 35952 109682
rect 35900 109618 35952 109624
rect 35992 104576 36044 104582
rect 35992 104518 36044 104524
rect 35808 101448 35860 101454
rect 35808 101390 35860 101396
rect 35820 94382 35848 101390
rect 35900 94784 35952 94790
rect 35900 94726 35952 94732
rect 35808 94376 35860 94382
rect 35808 94318 35860 94324
rect 35808 94240 35860 94246
rect 35808 94182 35860 94188
rect 35820 82278 35848 94182
rect 35912 90166 35940 94726
rect 35900 90160 35952 90166
rect 35900 90102 35952 90108
rect 35900 89956 35952 89962
rect 35900 89898 35952 89904
rect 35912 87446 35940 89898
rect 35900 87440 35952 87446
rect 35900 87382 35952 87388
rect 35900 87168 35952 87174
rect 35900 87110 35952 87116
rect 35808 82272 35860 82278
rect 35808 82214 35860 82220
rect 35912 80850 35940 87110
rect 36004 83094 36032 104518
rect 36176 104032 36228 104038
rect 36176 103974 36228 103980
rect 36084 90160 36136 90166
rect 36084 90102 36136 90108
rect 35992 83088 36044 83094
rect 35992 83030 36044 83036
rect 36096 81938 36124 90102
rect 36188 86154 36216 103974
rect 36280 103514 36308 112746
rect 36372 111654 36400 115466
rect 36360 111648 36412 111654
rect 36360 111590 36412 111596
rect 36280 103486 36400 103514
rect 36268 100768 36320 100774
rect 36268 100710 36320 100716
rect 36176 86148 36228 86154
rect 36176 86090 36228 86096
rect 36176 85876 36228 85882
rect 36176 85818 36228 85824
rect 36084 81932 36136 81938
rect 36084 81874 36136 81880
rect 35900 80844 35952 80850
rect 35900 80786 35952 80792
rect 35636 80056 35756 80084
rect 35636 77294 35664 80056
rect 36188 80054 36216 85818
rect 36280 81802 36308 100710
rect 36268 81796 36320 81802
rect 36268 81738 36320 81744
rect 36268 81524 36320 81530
rect 36268 81466 36320 81472
rect 36096 80026 36216 80054
rect 35636 77266 35756 77294
rect 35624 74656 35676 74662
rect 35624 74598 35676 74604
rect 35532 65544 35584 65550
rect 35532 65486 35584 65492
rect 35440 65408 35492 65414
rect 35440 65350 35492 65356
rect 35532 65408 35584 65414
rect 35532 65350 35584 65356
rect 35348 64864 35400 64870
rect 35254 64832 35310 64841
rect 35348 64806 35400 64812
rect 35254 64767 35310 64776
rect 35452 64705 35480 65350
rect 35438 64696 35494 64705
rect 35176 64620 35388 64648
rect 35438 64631 35494 64640
rect 35072 64592 35124 64598
rect 35072 64534 35124 64540
rect 35254 64560 35310 64569
rect 34888 64524 34940 64530
rect 35360 64546 35388 64620
rect 35360 64518 35480 64546
rect 35254 64495 35310 64504
rect 34888 64466 34940 64472
rect 34900 64433 34928 64466
rect 34886 64424 34942 64433
rect 34886 64359 34942 64368
rect 34940 64220 35236 64240
rect 34996 64218 35020 64220
rect 35076 64218 35100 64220
rect 35156 64218 35180 64220
rect 35018 64166 35020 64218
rect 35082 64166 35094 64218
rect 35156 64166 35158 64218
rect 34996 64164 35020 64166
rect 35076 64164 35100 64166
rect 35156 64164 35180 64166
rect 34940 64144 35236 64164
rect 34808 63974 34928 64002
rect 34796 63912 34848 63918
rect 34796 63854 34848 63860
rect 34808 63345 34836 63854
rect 34794 63336 34850 63345
rect 34794 63271 34850 63280
rect 34900 63220 34928 63974
rect 34980 63912 35032 63918
rect 34980 63854 35032 63860
rect 35162 63880 35218 63889
rect 34992 63442 35020 63854
rect 35162 63815 35218 63824
rect 35176 63442 35204 63815
rect 34980 63436 35032 63442
rect 34980 63378 35032 63384
rect 35164 63436 35216 63442
rect 35164 63378 35216 63384
rect 34808 63192 34928 63220
rect 34808 59752 34836 63192
rect 34940 63132 35236 63152
rect 34996 63130 35020 63132
rect 35076 63130 35100 63132
rect 35156 63130 35180 63132
rect 35018 63078 35020 63130
rect 35082 63078 35094 63130
rect 35156 63078 35158 63130
rect 34996 63076 35020 63078
rect 35076 63076 35100 63078
rect 35156 63076 35180 63078
rect 34940 63056 35236 63076
rect 34940 62044 35236 62064
rect 34996 62042 35020 62044
rect 35076 62042 35100 62044
rect 35156 62042 35180 62044
rect 35018 61990 35020 62042
rect 35082 61990 35094 62042
rect 35156 61990 35158 62042
rect 34996 61988 35020 61990
rect 35076 61988 35100 61990
rect 35156 61988 35180 61990
rect 34940 61968 35236 61988
rect 34886 61432 34942 61441
rect 34886 61367 34942 61376
rect 34900 61266 34928 61367
rect 34888 61260 34940 61266
rect 34888 61202 34940 61208
rect 34940 60956 35236 60976
rect 34996 60954 35020 60956
rect 35076 60954 35100 60956
rect 35156 60954 35180 60956
rect 35018 60902 35020 60954
rect 35082 60902 35094 60954
rect 35156 60902 35158 60954
rect 34996 60900 35020 60902
rect 35076 60900 35100 60902
rect 35156 60900 35180 60902
rect 34940 60880 35236 60900
rect 34888 60784 34940 60790
rect 34888 60726 34940 60732
rect 35164 60784 35216 60790
rect 35164 60726 35216 60732
rect 34900 60042 34928 60726
rect 35176 60625 35204 60726
rect 35268 60654 35296 64495
rect 35348 64456 35400 64462
rect 35348 64398 35400 64404
rect 35360 64161 35388 64398
rect 35346 64152 35402 64161
rect 35346 64087 35402 64096
rect 35348 63912 35400 63918
rect 35348 63854 35400 63860
rect 35360 61146 35388 63854
rect 35452 61402 35480 64518
rect 35544 63889 35572 65350
rect 35530 63880 35586 63889
rect 35530 63815 35586 63824
rect 35532 63436 35584 63442
rect 35532 63378 35584 63384
rect 35544 61674 35572 63378
rect 35532 61668 35584 61674
rect 35532 61610 35584 61616
rect 35440 61396 35492 61402
rect 35440 61338 35492 61344
rect 35532 61260 35584 61266
rect 35532 61202 35584 61208
rect 35360 61118 35480 61146
rect 35348 61056 35400 61062
rect 35348 60998 35400 61004
rect 35256 60648 35308 60654
rect 35162 60616 35218 60625
rect 35256 60590 35308 60596
rect 35162 60551 35218 60560
rect 35360 60314 35388 60998
rect 35452 60586 35480 61118
rect 35544 60790 35572 61202
rect 35532 60784 35584 60790
rect 35532 60726 35584 60732
rect 35532 60648 35584 60654
rect 35532 60590 35584 60596
rect 35440 60580 35492 60586
rect 35440 60522 35492 60528
rect 35348 60308 35400 60314
rect 35348 60250 35400 60256
rect 35162 60208 35218 60217
rect 35162 60143 35164 60152
rect 35216 60143 35218 60152
rect 35164 60114 35216 60120
rect 34888 60036 34940 60042
rect 34888 59978 34940 59984
rect 35348 60036 35400 60042
rect 35348 59978 35400 59984
rect 34940 59868 35236 59888
rect 34996 59866 35020 59868
rect 35076 59866 35100 59868
rect 35156 59866 35180 59868
rect 35018 59814 35020 59866
rect 35082 59814 35094 59866
rect 35156 59814 35158 59866
rect 34996 59812 35020 59814
rect 35076 59812 35100 59814
rect 35156 59812 35180 59814
rect 34940 59792 35236 59812
rect 34808 59724 34928 59752
rect 34794 59664 34850 59673
rect 34794 59599 34850 59608
rect 34808 59566 34836 59599
rect 34796 59560 34848 59566
rect 34796 59502 34848 59508
rect 34900 59412 34928 59724
rect 35254 59528 35310 59537
rect 35254 59463 35310 59472
rect 34808 59384 34928 59412
rect 34808 58478 34836 59384
rect 34940 58780 35236 58800
rect 34996 58778 35020 58780
rect 35076 58778 35100 58780
rect 35156 58778 35180 58780
rect 35018 58726 35020 58778
rect 35082 58726 35094 58778
rect 35156 58726 35158 58778
rect 34996 58724 35020 58726
rect 35076 58724 35100 58726
rect 35156 58724 35180 58726
rect 34940 58704 35236 58724
rect 34796 58472 34848 58478
rect 34796 58414 34848 58420
rect 34940 57692 35236 57712
rect 34996 57690 35020 57692
rect 35076 57690 35100 57692
rect 35156 57690 35180 57692
rect 35018 57638 35020 57690
rect 35082 57638 35094 57690
rect 35156 57638 35158 57690
rect 34996 57636 35020 57638
rect 35076 57636 35100 57638
rect 35156 57636 35180 57638
rect 34940 57616 35236 57636
rect 34940 56604 35236 56624
rect 34996 56602 35020 56604
rect 35076 56602 35100 56604
rect 35156 56602 35180 56604
rect 35018 56550 35020 56602
rect 35082 56550 35094 56602
rect 35156 56550 35158 56602
rect 34996 56548 35020 56550
rect 35076 56548 35100 56550
rect 35156 56548 35180 56550
rect 34940 56528 35236 56548
rect 35268 55894 35296 59463
rect 35256 55888 35308 55894
rect 35256 55830 35308 55836
rect 35256 55752 35308 55758
rect 35256 55694 35308 55700
rect 34940 55516 35236 55536
rect 34996 55514 35020 55516
rect 35076 55514 35100 55516
rect 35156 55514 35180 55516
rect 35018 55462 35020 55514
rect 35082 55462 35094 55514
rect 35156 55462 35158 55514
rect 34996 55460 35020 55462
rect 35076 55460 35100 55462
rect 35156 55460 35180 55462
rect 34940 55440 35236 55460
rect 34940 54428 35236 54448
rect 34996 54426 35020 54428
rect 35076 54426 35100 54428
rect 35156 54426 35180 54428
rect 35018 54374 35020 54426
rect 35082 54374 35094 54426
rect 35156 54374 35158 54426
rect 34996 54372 35020 54374
rect 35076 54372 35100 54374
rect 35156 54372 35180 54374
rect 34940 54352 35236 54372
rect 34940 53340 35236 53360
rect 34996 53338 35020 53340
rect 35076 53338 35100 53340
rect 35156 53338 35180 53340
rect 35018 53286 35020 53338
rect 35082 53286 35094 53338
rect 35156 53286 35158 53338
rect 34996 53284 35020 53286
rect 35076 53284 35100 53286
rect 35156 53284 35180 53286
rect 34940 53264 35236 53284
rect 34940 52252 35236 52272
rect 34996 52250 35020 52252
rect 35076 52250 35100 52252
rect 35156 52250 35180 52252
rect 35018 52198 35020 52250
rect 35082 52198 35094 52250
rect 35156 52198 35158 52250
rect 34996 52196 35020 52198
rect 35076 52196 35100 52198
rect 35156 52196 35180 52198
rect 34940 52176 35236 52196
rect 34940 51164 35236 51184
rect 34996 51162 35020 51164
rect 35076 51162 35100 51164
rect 35156 51162 35180 51164
rect 35018 51110 35020 51162
rect 35082 51110 35094 51162
rect 35156 51110 35158 51162
rect 34996 51108 35020 51110
rect 35076 51108 35100 51110
rect 35156 51108 35180 51110
rect 34940 51088 35236 51108
rect 34940 50076 35236 50096
rect 34996 50074 35020 50076
rect 35076 50074 35100 50076
rect 35156 50074 35180 50076
rect 35018 50022 35020 50074
rect 35082 50022 35094 50074
rect 35156 50022 35158 50074
rect 34996 50020 35020 50022
rect 35076 50020 35100 50022
rect 35156 50020 35180 50022
rect 34940 50000 35236 50020
rect 34796 49768 34848 49774
rect 34796 49710 34848 49716
rect 34808 46510 34836 49710
rect 34940 48988 35236 49008
rect 34996 48986 35020 48988
rect 35076 48986 35100 48988
rect 35156 48986 35180 48988
rect 35018 48934 35020 48986
rect 35082 48934 35094 48986
rect 35156 48934 35158 48986
rect 34996 48932 35020 48934
rect 35076 48932 35100 48934
rect 35156 48932 35180 48934
rect 34940 48912 35236 48932
rect 34940 47900 35236 47920
rect 34996 47898 35020 47900
rect 35076 47898 35100 47900
rect 35156 47898 35180 47900
rect 35018 47846 35020 47898
rect 35082 47846 35094 47898
rect 35156 47846 35158 47898
rect 34996 47844 35020 47846
rect 35076 47844 35100 47846
rect 35156 47844 35180 47846
rect 34940 47824 35236 47844
rect 34940 46812 35236 46832
rect 34996 46810 35020 46812
rect 35076 46810 35100 46812
rect 35156 46810 35180 46812
rect 35018 46758 35020 46810
rect 35082 46758 35094 46810
rect 35156 46758 35158 46810
rect 34996 46756 35020 46758
rect 35076 46756 35100 46758
rect 35156 46756 35180 46758
rect 34940 46736 35236 46756
rect 34796 46504 34848 46510
rect 34796 46446 34848 46452
rect 34796 46368 34848 46374
rect 34796 46310 34848 46316
rect 34808 45422 34836 46310
rect 34940 45724 35236 45744
rect 34996 45722 35020 45724
rect 35076 45722 35100 45724
rect 35156 45722 35180 45724
rect 35018 45670 35020 45722
rect 35082 45670 35094 45722
rect 35156 45670 35158 45722
rect 34996 45668 35020 45670
rect 35076 45668 35100 45670
rect 35156 45668 35180 45670
rect 34940 45648 35236 45668
rect 34796 45416 34848 45422
rect 34796 45358 34848 45364
rect 34796 45280 34848 45286
rect 34796 45222 34848 45228
rect 34808 44334 34836 45222
rect 34940 44636 35236 44656
rect 34996 44634 35020 44636
rect 35076 44634 35100 44636
rect 35156 44634 35180 44636
rect 35018 44582 35020 44634
rect 35082 44582 35094 44634
rect 35156 44582 35158 44634
rect 34996 44580 35020 44582
rect 35076 44580 35100 44582
rect 35156 44580 35180 44582
rect 34940 44560 35236 44580
rect 34796 44328 34848 44334
rect 34796 44270 34848 44276
rect 35268 44146 35296 55694
rect 35360 46753 35388 59978
rect 35452 59498 35480 60522
rect 35440 59492 35492 59498
rect 35440 59434 35492 59440
rect 35452 59090 35480 59434
rect 35440 59084 35492 59090
rect 35440 59026 35492 59032
rect 35544 54738 35572 60590
rect 35636 60178 35664 74598
rect 35728 67658 35756 77266
rect 35900 75336 35952 75342
rect 35900 75278 35952 75284
rect 35912 71738 35940 75278
rect 35900 71732 35952 71738
rect 35900 71674 35952 71680
rect 35912 69290 35940 71674
rect 35992 71528 36044 71534
rect 35992 71470 36044 71476
rect 35900 69284 35952 69290
rect 35900 69226 35952 69232
rect 35808 68876 35860 68882
rect 35808 68818 35860 68824
rect 35820 68241 35848 68818
rect 35806 68232 35862 68241
rect 35806 68167 35862 68176
rect 35900 67788 35952 67794
rect 35900 67730 35952 67736
rect 35716 67652 35768 67658
rect 35716 67594 35768 67600
rect 35808 66020 35860 66026
rect 35808 65962 35860 65968
rect 35716 65612 35768 65618
rect 35716 65554 35768 65560
rect 35728 64569 35756 65554
rect 35714 64560 35770 64569
rect 35714 64495 35770 64504
rect 35716 64388 35768 64394
rect 35716 64330 35768 64336
rect 35728 63782 35756 64330
rect 35820 63918 35848 65962
rect 35808 63912 35860 63918
rect 35808 63854 35860 63860
rect 35716 63776 35768 63782
rect 35716 63718 35768 63724
rect 35728 63374 35756 63718
rect 35806 63608 35862 63617
rect 35806 63543 35808 63552
rect 35860 63543 35862 63552
rect 35808 63514 35860 63520
rect 35806 63472 35862 63481
rect 35806 63407 35808 63416
rect 35860 63407 35862 63416
rect 35808 63378 35860 63384
rect 35716 63368 35768 63374
rect 35716 63310 35768 63316
rect 35808 63232 35860 63238
rect 35808 63174 35860 63180
rect 35714 62792 35770 62801
rect 35714 62727 35770 62736
rect 35728 62354 35756 62727
rect 35716 62348 35768 62354
rect 35716 62290 35768 62296
rect 35820 61962 35848 63174
rect 35728 61934 35848 61962
rect 35624 60172 35676 60178
rect 35624 60114 35676 60120
rect 35624 59696 35676 59702
rect 35624 59638 35676 59644
rect 35532 54732 35584 54738
rect 35532 54674 35584 54680
rect 35532 52080 35584 52086
rect 35532 52022 35584 52028
rect 35440 51808 35492 51814
rect 35440 51750 35492 51756
rect 35452 50454 35480 51750
rect 35440 50448 35492 50454
rect 35440 50390 35492 50396
rect 35440 48136 35492 48142
rect 35440 48078 35492 48084
rect 35346 46744 35402 46753
rect 35346 46679 35402 46688
rect 35348 46640 35400 46646
rect 35348 46582 35400 46588
rect 34808 44118 35296 44146
rect 34808 38706 34836 44118
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 35256 41540 35308 41546
rect 35256 41482 35308 41488
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 35268 41070 35296 41482
rect 35256 41064 35308 41070
rect 35256 41006 35308 41012
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 34808 38678 35296 38706
rect 34796 38548 34848 38554
rect 34796 38490 34848 38496
rect 34702 36408 34758 36417
rect 34702 36343 34758 36352
rect 34704 36304 34756 36310
rect 34704 36246 34756 36252
rect 34716 32978 34744 36246
rect 34704 32972 34756 32978
rect 34704 32914 34756 32920
rect 34624 31726 34744 31754
rect 34612 31136 34664 31142
rect 34612 31078 34664 31084
rect 34624 26489 34652 31078
rect 34610 26480 34666 26489
rect 34610 26415 34666 26424
rect 34612 26308 34664 26314
rect 34612 26250 34664 26256
rect 34518 25256 34574 25265
rect 34428 25220 34480 25226
rect 34518 25191 34574 25200
rect 34428 25162 34480 25168
rect 34520 25152 34572 25158
rect 34520 25094 34572 25100
rect 34532 24800 34560 25094
rect 34440 24772 34560 24800
rect 34334 24576 34390 24585
rect 34334 24511 34390 24520
rect 34244 24404 34296 24410
rect 34244 24346 34296 24352
rect 34336 24132 34388 24138
rect 34336 24074 34388 24080
rect 34244 23724 34296 23730
rect 34244 23666 34296 23672
rect 34152 23248 34204 23254
rect 34152 23190 34204 23196
rect 34060 22704 34112 22710
rect 34060 22646 34112 22652
rect 34152 22704 34204 22710
rect 34152 22646 34204 22652
rect 34164 22386 34192 22646
rect 34072 22358 34192 22386
rect 34072 21962 34100 22358
rect 34150 22264 34206 22273
rect 34150 22199 34206 22208
rect 34060 21956 34112 21962
rect 34060 21898 34112 21904
rect 34058 21856 34114 21865
rect 34058 21791 34114 21800
rect 34072 21418 34100 21791
rect 34060 21412 34112 21418
rect 34060 21354 34112 21360
rect 34164 21298 34192 22199
rect 34072 21270 34192 21298
rect 34072 19666 34100 21270
rect 34150 21176 34206 21185
rect 34150 21111 34206 21120
rect 34164 19802 34192 21111
rect 34256 20806 34284 23666
rect 34348 22438 34376 24074
rect 34440 23866 34468 24772
rect 34520 24676 34572 24682
rect 34520 24618 34572 24624
rect 34428 23860 34480 23866
rect 34428 23802 34480 23808
rect 34426 22944 34482 22953
rect 34426 22879 34482 22888
rect 34440 22574 34468 22879
rect 34428 22568 34480 22574
rect 34428 22510 34480 22516
rect 34336 22432 34388 22438
rect 34336 22374 34388 22380
rect 34440 22166 34468 22510
rect 34428 22160 34480 22166
rect 34334 22128 34390 22137
rect 34428 22102 34480 22108
rect 34334 22063 34390 22072
rect 34348 21457 34376 22063
rect 34426 21992 34482 22001
rect 34426 21927 34482 21936
rect 34334 21448 34390 21457
rect 34334 21383 34390 21392
rect 34336 21344 34388 21350
rect 34336 21286 34388 21292
rect 34244 20800 34296 20806
rect 34244 20742 34296 20748
rect 34256 20466 34284 20742
rect 34244 20460 34296 20466
rect 34244 20402 34296 20408
rect 34244 20256 34296 20262
rect 34244 20198 34296 20204
rect 34256 19990 34284 20198
rect 34244 19984 34296 19990
rect 34244 19926 34296 19932
rect 34164 19774 34284 19802
rect 34072 19638 34192 19666
rect 34058 19544 34114 19553
rect 34058 19479 34114 19488
rect 34072 18834 34100 19479
rect 34164 18970 34192 19638
rect 34152 18964 34204 18970
rect 34152 18906 34204 18912
rect 34060 18828 34112 18834
rect 34060 18770 34112 18776
rect 34060 18692 34112 18698
rect 34060 18634 34112 18640
rect 34072 17882 34100 18634
rect 34060 17876 34112 17882
rect 34060 17818 34112 17824
rect 34164 17218 34192 18906
rect 34072 17190 34192 17218
rect 33966 17096 34022 17105
rect 33966 17031 34022 17040
rect 33966 16960 34022 16969
rect 33966 16895 34022 16904
rect 33980 15978 34008 16895
rect 34072 16436 34100 17190
rect 34152 17128 34204 17134
rect 34152 17070 34204 17076
rect 34164 16726 34192 17070
rect 34152 16720 34204 16726
rect 34152 16662 34204 16668
rect 34152 16584 34204 16590
rect 34150 16552 34152 16561
rect 34204 16552 34206 16561
rect 34150 16487 34206 16496
rect 34072 16408 34192 16436
rect 33968 15972 34020 15978
rect 33968 15914 34020 15920
rect 33980 15609 34008 15914
rect 34060 15632 34112 15638
rect 33966 15600 34022 15609
rect 34060 15574 34112 15580
rect 33966 15535 34022 15544
rect 33968 15360 34020 15366
rect 33966 15328 33968 15337
rect 34020 15328 34022 15337
rect 33966 15263 34022 15272
rect 34072 14362 34100 15574
rect 33980 14334 34100 14362
rect 33980 14074 34008 14334
rect 34060 14272 34112 14278
rect 34060 14214 34112 14220
rect 33968 14068 34020 14074
rect 33968 14010 34020 14016
rect 33968 13864 34020 13870
rect 33968 13806 34020 13812
rect 33876 11756 33928 11762
rect 33876 11698 33928 11704
rect 33784 5296 33836 5302
rect 33784 5238 33836 5244
rect 33600 4684 33652 4690
rect 33600 4626 33652 4632
rect 33508 3936 33560 3942
rect 33508 3878 33560 3884
rect 33416 2644 33468 2650
rect 33416 2586 33468 2592
rect 33612 800 33640 4626
rect 33692 3392 33744 3398
rect 33692 3334 33744 3340
rect 33704 3194 33732 3334
rect 33692 3188 33744 3194
rect 33692 3130 33744 3136
rect 33876 2508 33928 2514
rect 33876 2450 33928 2456
rect 33888 800 33916 2450
rect 33980 2446 34008 13806
rect 34072 12918 34100 14214
rect 34060 12912 34112 12918
rect 34060 12854 34112 12860
rect 34164 2990 34192 16408
rect 34256 15638 34284 19774
rect 34348 17134 34376 21286
rect 34440 17882 34468 21927
rect 34532 21468 34560 24618
rect 34624 23497 34652 26250
rect 34716 25362 34744 31726
rect 34808 26382 34836 38490
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34888 36236 34940 36242
rect 34888 36178 34940 36184
rect 34900 36145 34928 36178
rect 34886 36136 34942 36145
rect 34886 36071 34942 36080
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 35268 35766 35296 38678
rect 35360 36174 35388 46582
rect 35452 41414 35480 48078
rect 35544 45354 35572 52022
rect 35636 50998 35664 59638
rect 35728 55758 35756 61934
rect 35808 61736 35860 61742
rect 35808 61678 35860 61684
rect 35820 61033 35848 61678
rect 35806 61024 35862 61033
rect 35806 60959 35862 60968
rect 35808 59968 35860 59974
rect 35808 59910 35860 59916
rect 35820 59634 35848 59910
rect 35808 59628 35860 59634
rect 35808 59570 35860 59576
rect 35806 59256 35862 59265
rect 35806 59191 35862 59200
rect 35820 58478 35848 59191
rect 35808 58472 35860 58478
rect 35808 58414 35860 58420
rect 35808 55888 35860 55894
rect 35808 55830 35860 55836
rect 35716 55752 35768 55758
rect 35716 55694 35768 55700
rect 35820 51074 35848 55830
rect 35728 51046 35848 51074
rect 35912 51074 35940 67730
rect 36004 67182 36032 71470
rect 36096 68950 36124 80026
rect 36280 77382 36308 81466
rect 36268 77376 36320 77382
rect 36268 77318 36320 77324
rect 36268 75200 36320 75206
rect 36268 75142 36320 75148
rect 36176 73568 36228 73574
rect 36176 73510 36228 73516
rect 36084 68944 36136 68950
rect 36084 68886 36136 68892
rect 36188 68338 36216 73510
rect 36280 68474 36308 75142
rect 36372 75002 36400 103486
rect 36360 74996 36412 75002
rect 36360 74938 36412 74944
rect 36360 72480 36412 72486
rect 36360 72422 36412 72428
rect 36268 68468 36320 68474
rect 36268 68410 36320 68416
rect 36176 68332 36228 68338
rect 36176 68274 36228 68280
rect 36268 68264 36320 68270
rect 36268 68206 36320 68212
rect 36176 68128 36228 68134
rect 36176 68070 36228 68076
rect 36084 67584 36136 67590
rect 36084 67526 36136 67532
rect 36096 67386 36124 67526
rect 36084 67380 36136 67386
rect 36084 67322 36136 67328
rect 35992 67176 36044 67182
rect 35992 67118 36044 67124
rect 36004 66094 36032 67118
rect 36084 67040 36136 67046
rect 36084 66982 36136 66988
rect 35992 66088 36044 66094
rect 35992 66030 36044 66036
rect 36004 65006 36032 66030
rect 35992 65000 36044 65006
rect 35992 64942 36044 64948
rect 35992 64524 36044 64530
rect 36096 64512 36124 66982
rect 36188 66706 36216 68070
rect 36280 67697 36308 68206
rect 36266 67688 36322 67697
rect 36266 67623 36322 67632
rect 36176 66700 36228 66706
rect 36176 66642 36228 66648
rect 36268 66632 36320 66638
rect 36268 66574 36320 66580
rect 36176 65408 36228 65414
rect 36176 65350 36228 65356
rect 36044 64484 36124 64512
rect 35992 64466 36044 64472
rect 36004 63850 36032 64466
rect 36082 64424 36138 64433
rect 36082 64359 36138 64368
rect 35992 63844 36044 63850
rect 35992 63786 36044 63792
rect 36004 63578 36032 63786
rect 35992 63572 36044 63578
rect 35992 63514 36044 63520
rect 36096 63356 36124 64359
rect 36188 63442 36216 65350
rect 36280 64666 36308 66574
rect 36268 64660 36320 64666
rect 36268 64602 36320 64608
rect 36268 64456 36320 64462
rect 36372 64433 36400 72422
rect 36464 71534 36492 117030
rect 36556 116890 36584 117030
rect 36648 116890 36676 119200
rect 36544 116884 36596 116890
rect 36544 116826 36596 116832
rect 36636 116884 36688 116890
rect 36636 116826 36688 116832
rect 36542 116784 36598 116793
rect 36542 116719 36544 116728
rect 36596 116719 36598 116728
rect 36544 116690 36596 116696
rect 36832 116618 36860 119200
rect 36910 117872 36966 117881
rect 36910 117807 36966 117816
rect 36820 116612 36872 116618
rect 36820 116554 36872 116560
rect 36728 116544 36780 116550
rect 36728 116486 36780 116492
rect 36544 115456 36596 115462
rect 36544 115398 36596 115404
rect 36556 114753 36584 115398
rect 36542 114744 36598 114753
rect 36542 114679 36598 114688
rect 36544 113484 36596 113490
rect 36544 113426 36596 113432
rect 36556 108730 36584 113426
rect 36544 108724 36596 108730
rect 36544 108666 36596 108672
rect 36740 102202 36768 116486
rect 36820 115660 36872 115666
rect 36820 115602 36872 115608
rect 36832 103154 36860 115602
rect 36924 113558 36952 117807
rect 37108 117230 37136 119200
rect 37278 119200 37334 120800
rect 37554 119200 37610 120800
rect 37738 119200 37794 120800
rect 38014 119200 38070 120800
rect 38198 119200 38254 120800
rect 38474 119200 38530 120800
rect 38658 119200 38714 120800
rect 38934 119200 38990 120800
rect 39118 119200 39174 120800
rect 39394 119200 39450 120800
rect 39578 119200 39634 120800
rect 39854 119200 39910 120800
rect 37186 119167 37242 119176
rect 37096 117224 37148 117230
rect 37096 117166 37148 117172
rect 37004 116068 37056 116074
rect 37004 116010 37056 116016
rect 36912 113552 36964 113558
rect 36912 113494 36964 113500
rect 37016 113354 37044 116010
rect 37200 113626 37228 119167
rect 37292 115598 37320 119200
rect 37568 116142 37596 119200
rect 37752 117094 37780 119200
rect 37740 117088 37792 117094
rect 37740 117030 37792 117036
rect 38028 116278 38056 119200
rect 38212 116822 38240 119200
rect 38200 116816 38252 116822
rect 38200 116758 38252 116764
rect 38016 116272 38068 116278
rect 38016 116214 38068 116220
rect 37556 116136 37608 116142
rect 37556 116078 37608 116084
rect 37280 115592 37332 115598
rect 37280 115534 37332 115540
rect 37372 115524 37424 115530
rect 37372 115466 37424 115472
rect 37384 115161 37412 115466
rect 37370 115152 37426 115161
rect 37370 115087 37426 115096
rect 37924 114980 37976 114986
rect 37924 114922 37976 114928
rect 37740 114912 37792 114918
rect 37740 114854 37792 114860
rect 37372 113824 37424 113830
rect 37372 113766 37424 113772
rect 37188 113620 37240 113626
rect 37188 113562 37240 113568
rect 37188 113484 37240 113490
rect 37188 113426 37240 113432
rect 37200 113393 37228 113426
rect 37186 113384 37242 113393
rect 37004 113348 37056 113354
rect 37186 113319 37242 113328
rect 37004 113290 37056 113296
rect 37280 113280 37332 113286
rect 37280 113222 37332 113228
rect 37188 112804 37240 112810
rect 37188 112746 37240 112752
rect 37094 112568 37150 112577
rect 37094 112503 37150 112512
rect 37108 112402 37136 112503
rect 37200 112470 37228 112746
rect 37188 112464 37240 112470
rect 37188 112406 37240 112412
rect 37096 112396 37148 112402
rect 37096 112338 37148 112344
rect 37094 112024 37150 112033
rect 37094 111959 37150 111968
rect 37108 111790 37136 111959
rect 37096 111784 37148 111790
rect 37096 111726 37148 111732
rect 37096 111308 37148 111314
rect 37096 111250 37148 111256
rect 37108 111217 37136 111250
rect 37094 111208 37150 111217
rect 37094 111143 37150 111152
rect 37094 110256 37150 110265
rect 37094 110191 37096 110200
rect 37148 110191 37150 110200
rect 37096 110162 37148 110168
rect 37094 109848 37150 109857
rect 37094 109783 37150 109792
rect 37108 109614 37136 109783
rect 37096 109608 37148 109614
rect 37096 109550 37148 109556
rect 36912 109268 36964 109274
rect 36912 109210 36964 109216
rect 36820 103148 36872 103154
rect 36820 103090 36872 103096
rect 36728 102196 36780 102202
rect 36728 102138 36780 102144
rect 36728 101856 36780 101862
rect 36728 101798 36780 101804
rect 36544 100020 36596 100026
rect 36544 99962 36596 99968
rect 36556 86222 36584 99962
rect 36636 93832 36688 93838
rect 36636 93774 36688 93780
rect 36648 87514 36676 93774
rect 36636 87508 36688 87514
rect 36636 87450 36688 87456
rect 36636 87236 36688 87242
rect 36636 87178 36688 87184
rect 36544 86216 36596 86222
rect 36544 86158 36596 86164
rect 36648 85898 36676 87178
rect 36740 87145 36768 101798
rect 36820 99680 36872 99686
rect 36820 99622 36872 99628
rect 36832 87281 36860 99622
rect 36818 87272 36874 87281
rect 36924 87242 36952 109210
rect 37096 109132 37148 109138
rect 37096 109074 37148 109080
rect 37108 108905 37136 109074
rect 37094 108896 37150 108905
rect 37094 108831 37150 108840
rect 37186 108080 37242 108089
rect 37186 108015 37188 108024
rect 37240 108015 37242 108024
rect 37188 107986 37240 107992
rect 37186 107536 37242 107545
rect 37186 107471 37242 107480
rect 37200 107438 37228 107471
rect 37188 107432 37240 107438
rect 37188 107374 37240 107380
rect 37188 106956 37240 106962
rect 37188 106898 37240 106904
rect 37200 106729 37228 106898
rect 37186 106720 37242 106729
rect 37186 106655 37242 106664
rect 37188 105868 37240 105874
rect 37188 105810 37240 105816
rect 37200 105777 37228 105810
rect 37186 105768 37242 105777
rect 37186 105703 37242 105712
rect 37186 104952 37242 104961
rect 37186 104887 37242 104896
rect 37200 104854 37228 104887
rect 37188 104848 37240 104854
rect 37188 104790 37240 104796
rect 37186 104408 37242 104417
rect 37186 104343 37242 104352
rect 37200 104174 37228 104343
rect 37188 104168 37240 104174
rect 37188 104110 37240 104116
rect 37188 103692 37240 103698
rect 37188 103634 37240 103640
rect 37200 103601 37228 103634
rect 37186 103592 37242 103601
rect 37186 103527 37242 103536
rect 37186 102640 37242 102649
rect 37186 102575 37188 102584
rect 37240 102575 37242 102584
rect 37188 102546 37240 102552
rect 37004 102400 37056 102406
rect 37004 102342 37056 102348
rect 37016 96234 37044 102342
rect 37186 102232 37242 102241
rect 37186 102167 37242 102176
rect 37200 101998 37228 102167
rect 37188 101992 37240 101998
rect 37188 101934 37240 101940
rect 37188 101516 37240 101522
rect 37188 101458 37240 101464
rect 37200 101289 37228 101458
rect 37186 101280 37242 101289
rect 37186 101215 37242 101224
rect 37186 100464 37242 100473
rect 37186 100399 37188 100408
rect 37240 100399 37242 100408
rect 37188 100370 37240 100376
rect 37292 100026 37320 113222
rect 37280 100020 37332 100026
rect 37280 99962 37332 99968
rect 37278 99920 37334 99929
rect 37278 99855 37334 99864
rect 37292 99822 37320 99855
rect 37280 99816 37332 99822
rect 37280 99758 37332 99764
rect 37186 99512 37242 99521
rect 37186 99447 37242 99456
rect 37200 99346 37228 99447
rect 37188 99340 37240 99346
rect 37188 99282 37240 99288
rect 37096 98252 37148 98258
rect 37096 98194 37148 98200
rect 37108 98161 37136 98194
rect 37094 98152 37150 98161
rect 37094 98087 37150 98096
rect 37094 97336 37150 97345
rect 37094 97271 37150 97280
rect 37108 97170 37136 97271
rect 37096 97164 37148 97170
rect 37096 97106 37148 97112
rect 37094 96792 37150 96801
rect 37094 96727 37150 96736
rect 37108 96558 37136 96727
rect 37096 96552 37148 96558
rect 37096 96494 37148 96500
rect 37016 96206 37136 96234
rect 37004 94784 37056 94790
rect 37004 94726 37056 94732
rect 36818 87207 36874 87216
rect 36912 87236 36964 87242
rect 36912 87178 36964 87184
rect 36726 87136 36782 87145
rect 36726 87071 36782 87080
rect 36910 87136 36966 87145
rect 36910 87071 36966 87080
rect 36818 87000 36874 87009
rect 36818 86935 36874 86944
rect 36728 86896 36780 86902
rect 36728 86838 36780 86844
rect 36556 85870 36676 85898
rect 36556 84794 36584 85870
rect 36636 85808 36688 85814
rect 36636 85750 36688 85756
rect 36544 84788 36596 84794
rect 36544 84730 36596 84736
rect 36544 83360 36596 83366
rect 36544 83302 36596 83308
rect 36452 71528 36504 71534
rect 36452 71470 36504 71476
rect 36452 68468 36504 68474
rect 36452 68410 36504 68416
rect 36464 66994 36492 68410
rect 36556 67182 36584 83302
rect 36648 69358 36676 85750
rect 36740 81530 36768 86838
rect 36832 86766 36860 86935
rect 36820 86760 36872 86766
rect 36820 86702 36872 86708
rect 36820 84448 36872 84454
rect 36820 84390 36872 84396
rect 36728 81524 36780 81530
rect 36728 81466 36780 81472
rect 36726 70000 36782 70009
rect 36726 69935 36728 69944
rect 36780 69935 36782 69944
rect 36728 69906 36780 69912
rect 36636 69352 36688 69358
rect 36636 69294 36688 69300
rect 36728 69284 36780 69290
rect 36728 69226 36780 69232
rect 36740 69018 36768 69226
rect 36728 69012 36780 69018
rect 36728 68954 36780 68960
rect 36740 68406 36768 68954
rect 36728 68400 36780 68406
rect 36728 68342 36780 68348
rect 36636 68332 36688 68338
rect 36636 68274 36688 68280
rect 36648 67674 36676 68274
rect 36740 67930 36768 68342
rect 36832 68270 36860 84390
rect 36924 80782 36952 87071
rect 36912 80776 36964 80782
rect 36912 80718 36964 80724
rect 37016 73098 37044 94726
rect 37108 86306 37136 96206
rect 37188 96076 37240 96082
rect 37188 96018 37240 96024
rect 37200 95985 37228 96018
rect 37186 95976 37242 95985
rect 37186 95911 37242 95920
rect 37186 95024 37242 95033
rect 37186 94959 37188 94968
rect 37240 94959 37242 94968
rect 37188 94930 37240 94936
rect 37186 94616 37242 94625
rect 37186 94551 37242 94560
rect 37200 94382 37228 94551
rect 37188 94376 37240 94382
rect 37188 94318 37240 94324
rect 37188 93900 37240 93906
rect 37188 93842 37240 93848
rect 37200 93673 37228 93842
rect 37384 93838 37412 113766
rect 37648 112736 37700 112742
rect 37648 112678 37700 112684
rect 37660 100502 37688 112678
rect 37752 101454 37780 114854
rect 37936 114345 37964 114922
rect 37922 114336 37978 114345
rect 37922 114271 37978 114280
rect 37924 113892 37976 113898
rect 37924 113834 37976 113840
rect 37936 113801 37964 113834
rect 37922 113792 37978 113801
rect 37922 113727 37978 113736
rect 37922 112976 37978 112985
rect 38488 112946 38516 119200
rect 38568 117156 38620 117162
rect 38568 117098 38620 117104
rect 37922 112911 37978 112920
rect 38476 112940 38528 112946
rect 37936 112878 37964 112911
rect 38476 112882 38528 112888
rect 37924 112872 37976 112878
rect 37924 112814 37976 112820
rect 37832 111784 37884 111790
rect 37832 111726 37884 111732
rect 37844 111625 37872 111726
rect 38476 111716 38528 111722
rect 38476 111658 38528 111664
rect 37830 111616 37886 111625
rect 37830 111551 37886 111560
rect 37832 110696 37884 110702
rect 37830 110664 37832 110673
rect 37884 110664 37886 110673
rect 37830 110599 37886 110608
rect 37832 109608 37884 109614
rect 37832 109550 37884 109556
rect 37844 109449 37872 109550
rect 37830 109440 37886 109449
rect 37830 109375 37886 109384
rect 37832 108520 37884 108526
rect 37830 108488 37832 108497
rect 37884 108488 37886 108497
rect 37830 108423 37886 108432
rect 37924 107364 37976 107370
rect 37924 107306 37976 107312
rect 37936 107137 37964 107306
rect 37922 107128 37978 107137
rect 37922 107063 37978 107072
rect 37924 106344 37976 106350
rect 37924 106286 37976 106292
rect 37936 106185 37964 106286
rect 37922 106176 37978 106185
rect 37922 106111 37978 106120
rect 37922 105360 37978 105369
rect 37922 105295 37978 105304
rect 37936 105262 37964 105295
rect 37924 105256 37976 105262
rect 37924 105198 37976 105204
rect 37924 104100 37976 104106
rect 37924 104042 37976 104048
rect 37936 104009 37964 104042
rect 37922 104000 37978 104009
rect 37922 103935 37978 103944
rect 38200 103556 38252 103562
rect 38200 103498 38252 103504
rect 37922 103048 37978 103057
rect 37922 102983 37924 102992
rect 37976 102983 37978 102992
rect 37924 102954 37976 102960
rect 37924 101924 37976 101930
rect 37924 101866 37976 101872
rect 37936 101833 37964 101866
rect 37922 101824 37978 101833
rect 37922 101759 37978 101768
rect 37740 101448 37792 101454
rect 37740 101390 37792 101396
rect 37922 100872 37978 100881
rect 37922 100807 37924 100816
rect 37976 100807 37978 100816
rect 37924 100778 37976 100784
rect 37648 100496 37700 100502
rect 37648 100438 37700 100444
rect 37924 99816 37976 99822
rect 37924 99758 37976 99764
rect 37936 99113 37964 99758
rect 37922 99104 37978 99113
rect 37922 99039 37978 99048
rect 37924 98728 37976 98734
rect 37922 98696 37924 98705
rect 37976 98696 37978 98705
rect 37922 98631 37978 98640
rect 37830 97744 37886 97753
rect 37830 97679 37886 97688
rect 37844 97646 37872 97679
rect 37832 97640 37884 97646
rect 37832 97582 37884 97588
rect 37924 96484 37976 96490
rect 37924 96426 37976 96432
rect 37936 96393 37964 96426
rect 37922 96384 37978 96393
rect 37922 96319 37978 96328
rect 37922 95432 37978 95441
rect 37922 95367 37924 95376
rect 37976 95367 37978 95376
rect 37924 95338 37976 95344
rect 37924 94308 37976 94314
rect 37924 94250 37976 94256
rect 37556 94240 37608 94246
rect 37936 94217 37964 94250
rect 37556 94182 37608 94188
rect 37922 94208 37978 94217
rect 37372 93832 37424 93838
rect 37372 93774 37424 93780
rect 37186 93664 37242 93673
rect 37186 93599 37242 93608
rect 37280 93288 37332 93294
rect 37278 93256 37280 93265
rect 37332 93256 37334 93265
rect 37278 93191 37334 93200
rect 37278 92304 37334 92313
rect 37278 92239 37334 92248
rect 37292 92206 37320 92239
rect 37280 92200 37332 92206
rect 37280 92142 37332 92148
rect 37372 92064 37424 92070
rect 37372 92006 37424 92012
rect 37186 91896 37242 91905
rect 37186 91831 37242 91840
rect 37200 91730 37228 91831
rect 37188 91724 37240 91730
rect 37188 91666 37240 91672
rect 37280 91520 37332 91526
rect 37280 91462 37332 91468
rect 37188 91112 37240 91118
rect 37186 91080 37188 91089
rect 37240 91080 37242 91089
rect 37186 91015 37242 91024
rect 37292 90250 37320 91462
rect 37200 90222 37320 90250
rect 37200 89842 37228 90222
rect 37278 90128 37334 90137
rect 37278 90063 37334 90072
rect 37292 90030 37320 90063
rect 37280 90024 37332 90030
rect 37280 89966 37332 89972
rect 37200 89814 37320 89842
rect 37186 89720 37242 89729
rect 37186 89655 37242 89664
rect 37200 89554 37228 89655
rect 37188 89548 37240 89554
rect 37188 89490 37240 89496
rect 37292 89026 37320 89814
rect 37200 88998 37320 89026
rect 37200 87514 37228 88998
rect 37280 88936 37332 88942
rect 37280 88878 37332 88884
rect 37292 88777 37320 88878
rect 37278 88768 37334 88777
rect 37278 88703 37334 88712
rect 37278 87952 37334 87961
rect 37278 87887 37334 87896
rect 37292 87854 37320 87887
rect 37280 87848 37332 87854
rect 37280 87790 37332 87796
rect 37188 87508 37240 87514
rect 37188 87450 37240 87456
rect 37186 87408 37242 87417
rect 37186 87343 37188 87352
rect 37240 87343 37242 87352
rect 37188 87314 37240 87320
rect 37188 87236 37240 87242
rect 37188 87178 37240 87184
rect 37200 86698 37228 87178
rect 37280 86760 37332 86766
rect 37280 86702 37332 86708
rect 37188 86692 37240 86698
rect 37188 86634 37240 86640
rect 37292 86601 37320 86702
rect 37278 86592 37334 86601
rect 37278 86527 37334 86536
rect 37108 86278 37228 86306
rect 37096 86148 37148 86154
rect 37096 86090 37148 86096
rect 37108 82822 37136 86090
rect 37200 84402 37228 86278
rect 37280 85672 37332 85678
rect 37278 85640 37280 85649
rect 37332 85640 37334 85649
rect 37278 85575 37334 85584
rect 37278 84824 37334 84833
rect 37278 84759 37334 84768
rect 37292 84590 37320 84759
rect 37280 84584 37332 84590
rect 37280 84526 37332 84532
rect 37200 84374 37320 84402
rect 37186 84280 37242 84289
rect 37186 84215 37242 84224
rect 37200 84114 37228 84215
rect 37188 84108 37240 84114
rect 37188 84050 37240 84056
rect 37292 83994 37320 84374
rect 37384 84182 37412 92006
rect 37464 90976 37516 90982
rect 37464 90918 37516 90924
rect 37476 90030 37504 90918
rect 37464 90024 37516 90030
rect 37464 89966 37516 89972
rect 37464 89888 37516 89894
rect 37464 89830 37516 89836
rect 37476 87802 37504 89830
rect 37568 88398 37596 94182
rect 37922 94143 37978 94152
rect 37924 93288 37976 93294
rect 37924 93230 37976 93236
rect 37936 92857 37964 93230
rect 38108 93152 38160 93158
rect 38108 93094 38160 93100
rect 37922 92848 37978 92857
rect 37922 92783 37978 92792
rect 37924 92200 37976 92206
rect 37924 92142 37976 92148
rect 37832 92064 37884 92070
rect 37832 92006 37884 92012
rect 37740 91248 37792 91254
rect 37740 91190 37792 91196
rect 37648 89344 37700 89350
rect 37648 89286 37700 89292
rect 37556 88392 37608 88398
rect 37556 88334 37608 88340
rect 37476 87774 37596 87802
rect 37464 87712 37516 87718
rect 37464 87654 37516 87660
rect 37372 84176 37424 84182
rect 37372 84118 37424 84124
rect 37200 83966 37320 83994
rect 37096 82816 37148 82822
rect 37096 82758 37148 82764
rect 37200 82226 37228 83966
rect 37372 83904 37424 83910
rect 37372 83846 37424 83852
rect 37280 83496 37332 83502
rect 37278 83464 37280 83473
rect 37332 83464 37334 83473
rect 37278 83399 37334 83408
rect 37278 82512 37334 82521
rect 37278 82447 37334 82456
rect 37292 82414 37320 82447
rect 37280 82408 37332 82414
rect 37280 82350 37332 82356
rect 37108 82198 37228 82226
rect 37108 80102 37136 82198
rect 37186 82104 37242 82113
rect 37186 82039 37242 82048
rect 37200 81938 37228 82039
rect 37188 81932 37240 81938
rect 37188 81874 37240 81880
rect 37188 81796 37240 81802
rect 37188 81738 37240 81744
rect 37096 80096 37148 80102
rect 37096 80038 37148 80044
rect 37200 79898 37228 81738
rect 37280 81320 37332 81326
rect 37280 81262 37332 81268
rect 37292 81161 37320 81262
rect 37278 81152 37334 81161
rect 37278 81087 37334 81096
rect 37278 80336 37334 80345
rect 37278 80271 37334 80280
rect 37292 80238 37320 80271
rect 37280 80232 37332 80238
rect 37280 80174 37332 80180
rect 37188 79892 37240 79898
rect 37188 79834 37240 79840
rect 37186 79792 37242 79801
rect 37186 79727 37188 79736
rect 37240 79727 37242 79736
rect 37188 79698 37240 79704
rect 37280 79144 37332 79150
rect 37280 79086 37332 79092
rect 37292 78985 37320 79086
rect 37278 78976 37334 78985
rect 37278 78911 37334 78920
rect 37280 78056 37332 78062
rect 37278 78024 37280 78033
rect 37332 78024 37334 78033
rect 37278 77959 37334 77968
rect 37278 77208 37334 77217
rect 37278 77143 37334 77152
rect 37292 76974 37320 77143
rect 37280 76968 37332 76974
rect 37280 76910 37332 76916
rect 37280 75880 37332 75886
rect 37278 75848 37280 75857
rect 37332 75848 37334 75857
rect 37278 75783 37334 75792
rect 37188 75404 37240 75410
rect 37188 75346 37240 75352
rect 37200 75313 37228 75346
rect 37186 75304 37242 75313
rect 37186 75239 37242 75248
rect 37278 74896 37334 74905
rect 37278 74831 37334 74840
rect 37292 74798 37320 74831
rect 37280 74792 37332 74798
rect 37280 74734 37332 74740
rect 37186 74488 37242 74497
rect 37186 74423 37242 74432
rect 37200 74322 37228 74423
rect 37188 74316 37240 74322
rect 37188 74258 37240 74264
rect 37096 73840 37148 73846
rect 37096 73782 37148 73788
rect 37004 73092 37056 73098
rect 37004 73034 37056 73040
rect 37108 72026 37136 73782
rect 37280 73704 37332 73710
rect 37280 73646 37332 73652
rect 37292 73545 37320 73646
rect 37278 73536 37334 73545
rect 37278 73471 37334 73480
rect 37278 72720 37334 72729
rect 37278 72655 37334 72664
rect 37292 72622 37320 72655
rect 37280 72616 37332 72622
rect 37280 72558 37332 72564
rect 37186 72176 37242 72185
rect 37186 72111 37188 72120
rect 37240 72111 37242 72120
rect 37188 72082 37240 72088
rect 37108 71998 37228 72026
rect 36912 71936 36964 71942
rect 36912 71878 36964 71884
rect 36924 69873 36952 71878
rect 37096 70848 37148 70854
rect 37096 70790 37148 70796
rect 36910 69864 36966 69873
rect 36910 69799 36966 69808
rect 37004 69828 37056 69834
rect 37004 69770 37056 69776
rect 36912 69760 36964 69766
rect 36912 69702 36964 69708
rect 36820 68264 36872 68270
rect 36820 68206 36872 68212
rect 36728 67924 36780 67930
rect 36728 67866 36780 67872
rect 36820 67924 36872 67930
rect 36820 67866 36872 67872
rect 36728 67788 36780 67794
rect 36832 67776 36860 67866
rect 36780 67748 36860 67776
rect 36728 67730 36780 67736
rect 36648 67646 36860 67674
rect 36636 67584 36688 67590
rect 36636 67526 36688 67532
rect 36544 67176 36596 67182
rect 36544 67118 36596 67124
rect 36464 66966 36584 66994
rect 36452 65612 36504 65618
rect 36452 65554 36504 65560
rect 36268 64398 36320 64404
rect 36358 64424 36414 64433
rect 36176 63436 36228 63442
rect 36176 63378 36228 63384
rect 36004 63328 36124 63356
rect 36004 60654 36032 63328
rect 36082 63064 36138 63073
rect 36082 62999 36138 63008
rect 36096 62830 36124 62999
rect 36084 62824 36136 62830
rect 36084 62766 36136 62772
rect 36280 62506 36308 64398
rect 36358 64359 36414 64368
rect 36360 64320 36412 64326
rect 36360 64262 36412 64268
rect 36096 62478 36308 62506
rect 35992 60648 36044 60654
rect 35992 60590 36044 60596
rect 35992 60172 36044 60178
rect 35992 60114 36044 60120
rect 36004 59770 36032 60114
rect 35992 59764 36044 59770
rect 35992 59706 36044 59712
rect 36096 59566 36124 62478
rect 36266 62384 36322 62393
rect 36266 62319 36268 62328
rect 36320 62319 36322 62328
rect 36268 62290 36320 62296
rect 36176 62144 36228 62150
rect 36176 62086 36228 62092
rect 36084 59560 36136 59566
rect 36084 59502 36136 59508
rect 36188 59242 36216 62086
rect 36268 61260 36320 61266
rect 36268 61202 36320 61208
rect 36096 59214 36216 59242
rect 35992 59084 36044 59090
rect 35992 59026 36044 59032
rect 36004 58070 36032 59026
rect 35992 58064 36044 58070
rect 35992 58006 36044 58012
rect 36096 55894 36124 59214
rect 36176 58880 36228 58886
rect 36176 58822 36228 58828
rect 36084 55888 36136 55894
rect 36084 55830 36136 55836
rect 35912 51046 36032 51074
rect 35624 50992 35676 50998
rect 35624 50934 35676 50940
rect 35624 50176 35676 50182
rect 35624 50118 35676 50124
rect 35532 45348 35584 45354
rect 35532 45290 35584 45296
rect 35452 41386 35572 41414
rect 35440 40928 35492 40934
rect 35440 40870 35492 40876
rect 35348 36168 35400 36174
rect 35348 36110 35400 36116
rect 35348 36032 35400 36038
rect 35348 35974 35400 35980
rect 35256 35760 35308 35766
rect 35256 35702 35308 35708
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 35360 32314 35388 35974
rect 35268 32286 35388 32314
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34888 29232 34940 29238
rect 34888 29174 34940 29180
rect 34900 28490 34928 29174
rect 34888 28484 34940 28490
rect 34888 28426 34940 28432
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34796 26376 34848 26382
rect 34796 26318 34848 26324
rect 34796 26240 34848 26246
rect 34796 26182 34848 26188
rect 34704 25356 34756 25362
rect 34704 25298 34756 25304
rect 34702 25256 34758 25265
rect 34702 25191 34758 25200
rect 34610 23488 34666 23497
rect 34610 23423 34666 23432
rect 34612 23180 34664 23186
rect 34612 23122 34664 23128
rect 34624 23089 34652 23122
rect 34610 23080 34666 23089
rect 34610 23015 34666 23024
rect 34612 22976 34664 22982
rect 34612 22918 34664 22924
rect 34624 22098 34652 22918
rect 34716 22522 34744 25191
rect 34808 22624 34836 26182
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 34886 25936 34942 25945
rect 34886 25871 34942 25880
rect 34900 25265 34928 25871
rect 34980 25832 35032 25838
rect 34980 25774 35032 25780
rect 34992 25401 35020 25774
rect 35164 25764 35216 25770
rect 35164 25706 35216 25712
rect 35176 25430 35204 25706
rect 35164 25424 35216 25430
rect 34978 25392 35034 25401
rect 35164 25366 35216 25372
rect 34978 25327 35034 25336
rect 34886 25256 34942 25265
rect 34886 25191 34942 25200
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 35162 24882 35218 24891
rect 35162 24817 35218 24826
rect 35176 24138 35204 24817
rect 35268 24682 35296 32286
rect 35348 32224 35400 32230
rect 35348 32166 35400 32172
rect 35256 24676 35308 24682
rect 35256 24618 35308 24624
rect 35256 24404 35308 24410
rect 35256 24346 35308 24352
rect 35164 24132 35216 24138
rect 35164 24074 35216 24080
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34980 23724 35032 23730
rect 34980 23666 35032 23672
rect 34992 23254 35020 23666
rect 35268 23662 35296 24346
rect 35256 23656 35308 23662
rect 35256 23598 35308 23604
rect 34980 23248 35032 23254
rect 35360 23236 35388 32166
rect 34980 23190 35032 23196
rect 35268 23208 35388 23236
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 35072 22704 35124 22710
rect 35072 22646 35124 22652
rect 34808 22596 35020 22624
rect 34716 22494 34836 22522
rect 34704 22432 34756 22438
rect 34704 22374 34756 22380
rect 34612 22092 34664 22098
rect 34612 22034 34664 22040
rect 34612 21956 34664 21962
rect 34612 21898 34664 21904
rect 34624 21622 34652 21898
rect 34612 21616 34664 21622
rect 34612 21558 34664 21564
rect 34532 21440 34652 21468
rect 34520 20800 34572 20806
rect 34520 20742 34572 20748
rect 34532 20602 34560 20742
rect 34520 20596 34572 20602
rect 34520 20538 34572 20544
rect 34518 20496 34574 20505
rect 34518 20431 34574 20440
rect 34532 19990 34560 20431
rect 34520 19984 34572 19990
rect 34518 19952 34520 19961
rect 34572 19952 34574 19961
rect 34518 19887 34574 19896
rect 34520 19848 34572 19854
rect 34520 19790 34572 19796
rect 34532 19310 34560 19790
rect 34520 19304 34572 19310
rect 34520 19246 34572 19252
rect 34532 18902 34560 19246
rect 34520 18896 34572 18902
rect 34520 18838 34572 18844
rect 34520 18216 34572 18222
rect 34624 18204 34652 21440
rect 34716 19310 34744 22374
rect 34808 20398 34836 22494
rect 34888 22432 34940 22438
rect 34992 22420 35020 22596
rect 35084 22545 35112 22646
rect 35268 22574 35296 23208
rect 35348 23044 35400 23050
rect 35348 22986 35400 22992
rect 35256 22568 35308 22574
rect 35070 22536 35126 22545
rect 35256 22510 35308 22516
rect 35070 22471 35126 22480
rect 34992 22392 35296 22420
rect 34888 22374 34940 22380
rect 34900 22001 34928 22374
rect 35070 22128 35126 22137
rect 35070 22063 35072 22072
rect 35124 22063 35126 22072
rect 35072 22034 35124 22040
rect 34886 21992 34942 22001
rect 34886 21927 34942 21936
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 35268 21672 35296 22392
rect 35176 21644 35296 21672
rect 35176 20913 35204 21644
rect 35256 21548 35308 21554
rect 35256 21490 35308 21496
rect 35162 20904 35218 20913
rect 35162 20839 35218 20848
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 34796 20392 34848 20398
rect 34796 20334 34848 20340
rect 34886 20360 34942 20369
rect 34886 20295 34942 20304
rect 34796 20256 34848 20262
rect 34796 20198 34848 20204
rect 34704 19304 34756 19310
rect 34704 19246 34756 19252
rect 34704 18896 34756 18902
rect 34704 18838 34756 18844
rect 34716 18358 34744 18838
rect 34704 18352 34756 18358
rect 34704 18294 34756 18300
rect 34704 18216 34756 18222
rect 34624 18176 34704 18204
rect 34520 18158 34572 18164
rect 34704 18158 34756 18164
rect 34428 17876 34480 17882
rect 34428 17818 34480 17824
rect 34336 17128 34388 17134
rect 34336 17070 34388 17076
rect 34334 16960 34390 16969
rect 34334 16895 34390 16904
rect 34348 16658 34376 16895
rect 34336 16652 34388 16658
rect 34336 16594 34388 16600
rect 34334 16008 34390 16017
rect 34334 15943 34390 15952
rect 34244 15632 34296 15638
rect 34244 15574 34296 15580
rect 34348 15570 34376 15943
rect 34336 15564 34388 15570
rect 34336 15506 34388 15512
rect 34244 15428 34296 15434
rect 34244 15370 34296 15376
rect 34256 14958 34284 15370
rect 34334 15192 34390 15201
rect 34334 15127 34390 15136
rect 34244 14952 34296 14958
rect 34244 14894 34296 14900
rect 34348 14822 34376 15127
rect 34336 14816 34388 14822
rect 34336 14758 34388 14764
rect 34348 14634 34376 14758
rect 34256 14606 34376 14634
rect 34256 13870 34284 14606
rect 34334 14512 34390 14521
rect 34334 14447 34336 14456
rect 34388 14447 34390 14456
rect 34336 14418 34388 14424
rect 34348 14074 34376 14418
rect 34336 14068 34388 14074
rect 34336 14010 34388 14016
rect 34348 13938 34376 14010
rect 34336 13932 34388 13938
rect 34336 13874 34388 13880
rect 34244 13864 34296 13870
rect 34244 13806 34296 13812
rect 34440 4758 34468 17818
rect 34532 17678 34560 18158
rect 34704 18080 34756 18086
rect 34704 18022 34756 18028
rect 34612 17808 34664 17814
rect 34612 17750 34664 17756
rect 34520 17672 34572 17678
rect 34520 17614 34572 17620
rect 34532 17202 34560 17614
rect 34520 17196 34572 17202
rect 34520 17138 34572 17144
rect 34624 16794 34652 17750
rect 34716 17066 34744 18022
rect 34704 17060 34756 17066
rect 34704 17002 34756 17008
rect 34612 16788 34664 16794
rect 34612 16730 34664 16736
rect 34612 16652 34664 16658
rect 34532 16612 34612 16640
rect 34532 11694 34560 16612
rect 34612 16594 34664 16600
rect 34612 16448 34664 16454
rect 34612 16390 34664 16396
rect 34624 15910 34652 16390
rect 34716 16182 34744 17002
rect 34704 16176 34756 16182
rect 34704 16118 34756 16124
rect 34612 15904 34664 15910
rect 34612 15846 34664 15852
rect 34612 15564 34664 15570
rect 34612 15506 34664 15512
rect 34624 14890 34652 15506
rect 34612 14884 34664 14890
rect 34612 14826 34664 14832
rect 34624 14618 34652 14826
rect 34612 14612 34664 14618
rect 34612 14554 34664 14560
rect 34624 14006 34652 14554
rect 34612 14000 34664 14006
rect 34612 13942 34664 13948
rect 34808 12434 34836 20198
rect 34900 19825 34928 20295
rect 34886 19816 34942 19825
rect 34886 19751 34942 19760
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 35072 19440 35124 19446
rect 34886 19408 34942 19417
rect 35072 19382 35124 19388
rect 34886 19343 34942 19352
rect 34900 18970 34928 19343
rect 34888 18964 34940 18970
rect 34888 18906 34940 18912
rect 35084 18737 35112 19382
rect 35164 19304 35216 19310
rect 35164 19246 35216 19252
rect 35070 18728 35126 18737
rect 35176 18698 35204 19246
rect 35070 18663 35126 18672
rect 35164 18692 35216 18698
rect 35164 18634 35216 18640
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 34886 18320 34942 18329
rect 34886 18255 34942 18264
rect 34900 18222 34928 18255
rect 34888 18216 34940 18222
rect 34888 18158 34940 18164
rect 34900 17746 34928 18158
rect 34888 17740 34940 17746
rect 34888 17682 34940 17688
rect 35072 17740 35124 17746
rect 35072 17682 35124 17688
rect 35084 17610 35112 17682
rect 35072 17604 35124 17610
rect 35072 17546 35124 17552
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 35268 16658 35296 21490
rect 35360 21185 35388 22986
rect 35346 21176 35402 21185
rect 35346 21111 35402 21120
rect 35452 21010 35480 40870
rect 35544 36530 35572 41386
rect 35636 36700 35664 50118
rect 35728 45490 35756 51046
rect 35808 50720 35860 50726
rect 35808 50662 35860 50668
rect 35820 46866 35848 50662
rect 35820 46838 35940 46866
rect 35806 46744 35862 46753
rect 35806 46679 35862 46688
rect 35716 45484 35768 45490
rect 35716 45426 35768 45432
rect 35716 45348 35768 45354
rect 35716 45290 35768 45296
rect 35728 36825 35756 45290
rect 35820 38758 35848 46679
rect 35912 45354 35940 46838
rect 35900 45348 35952 45354
rect 35900 45290 35952 45296
rect 35900 41472 35952 41478
rect 35900 41414 35952 41420
rect 35808 38752 35860 38758
rect 35808 38694 35860 38700
rect 35714 36816 35770 36825
rect 35714 36751 35770 36760
rect 35636 36672 35848 36700
rect 35714 36544 35770 36553
rect 35544 36502 35664 36530
rect 35530 36408 35586 36417
rect 35530 36343 35586 36352
rect 35544 31754 35572 36343
rect 35532 31748 35584 31754
rect 35532 31690 35584 31696
rect 35532 31476 35584 31482
rect 35532 31418 35584 31424
rect 35348 21004 35400 21010
rect 35348 20946 35400 20952
rect 35440 21004 35492 21010
rect 35440 20946 35492 20952
rect 35360 20330 35388 20946
rect 35438 20904 35494 20913
rect 35438 20839 35494 20848
rect 35348 20324 35400 20330
rect 35348 20266 35400 20272
rect 35360 19922 35388 20266
rect 35348 19916 35400 19922
rect 35348 19858 35400 19864
rect 35360 19174 35388 19858
rect 35348 19168 35400 19174
rect 35348 19110 35400 19116
rect 35348 18828 35400 18834
rect 35348 18770 35400 18776
rect 35360 18290 35388 18770
rect 35452 18714 35480 20839
rect 35544 18834 35572 31418
rect 35636 27606 35664 36502
rect 35714 36479 35770 36488
rect 35624 27600 35676 27606
rect 35624 27542 35676 27548
rect 35624 25696 35676 25702
rect 35624 25638 35676 25644
rect 35636 23594 35664 25638
rect 35728 25362 35756 36479
rect 35820 33862 35848 36672
rect 35808 33856 35860 33862
rect 35808 33798 35860 33804
rect 35808 32972 35860 32978
rect 35808 32914 35860 32920
rect 35716 25356 35768 25362
rect 35716 25298 35768 25304
rect 35716 25220 35768 25226
rect 35716 25162 35768 25168
rect 35728 24886 35756 25162
rect 35716 24880 35768 24886
rect 35716 24822 35768 24828
rect 35728 24274 35756 24822
rect 35716 24268 35768 24274
rect 35716 24210 35768 24216
rect 35728 23866 35756 24210
rect 35716 23860 35768 23866
rect 35716 23802 35768 23808
rect 35624 23588 35676 23594
rect 35624 23530 35676 23536
rect 35716 23520 35768 23526
rect 35622 23488 35678 23497
rect 35716 23462 35768 23468
rect 35622 23423 35678 23432
rect 35636 22098 35664 23423
rect 35728 22710 35756 23462
rect 35716 22704 35768 22710
rect 35716 22646 35768 22652
rect 35716 22568 35768 22574
rect 35716 22510 35768 22516
rect 35624 22092 35676 22098
rect 35624 22034 35676 22040
rect 35622 21992 35678 22001
rect 35622 21927 35678 21936
rect 35532 18828 35584 18834
rect 35532 18770 35584 18776
rect 35452 18686 35572 18714
rect 35440 18624 35492 18630
rect 35440 18566 35492 18572
rect 35348 18284 35400 18290
rect 35348 18226 35400 18232
rect 35348 17604 35400 17610
rect 35348 17546 35400 17552
rect 35256 16652 35308 16658
rect 35256 16594 35308 16600
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34624 12406 34836 12434
rect 34520 11688 34572 11694
rect 34520 11630 34572 11636
rect 34624 8634 34652 12406
rect 35360 12374 35388 17546
rect 35452 15609 35480 18566
rect 35438 15600 35494 15609
rect 35438 15535 35494 15544
rect 35440 15496 35492 15502
rect 35440 15438 35492 15444
rect 34704 12368 34756 12374
rect 34704 12310 34756 12316
rect 35348 12368 35400 12374
rect 35348 12310 35400 12316
rect 34612 8628 34664 8634
rect 34612 8570 34664 8576
rect 34520 5772 34572 5778
rect 34520 5714 34572 5720
rect 34428 4752 34480 4758
rect 34428 4694 34480 4700
rect 34336 4140 34388 4146
rect 34336 4082 34388 4088
rect 34348 3602 34376 4082
rect 34336 3596 34388 3602
rect 34336 3538 34388 3544
rect 34244 3392 34296 3398
rect 34244 3334 34296 3340
rect 34152 2984 34204 2990
rect 34152 2926 34204 2932
rect 33968 2440 34020 2446
rect 33968 2382 34020 2388
rect 34256 800 34284 3334
rect 34532 800 34560 5714
rect 34716 5642 34744 12310
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 34796 11688 34848 11694
rect 35452 11642 35480 15438
rect 35544 14958 35572 18686
rect 35636 15570 35664 21927
rect 35728 17746 35756 22510
rect 35820 19922 35848 32914
rect 35912 25294 35940 41414
rect 35900 25288 35952 25294
rect 35900 25230 35952 25236
rect 35900 25152 35952 25158
rect 35900 25094 35952 25100
rect 35912 23798 35940 25094
rect 35900 23792 35952 23798
rect 35900 23734 35952 23740
rect 35900 23520 35952 23526
rect 35900 23462 35952 23468
rect 35912 22001 35940 23462
rect 35898 21992 35954 22001
rect 35898 21927 35954 21936
rect 35900 21888 35952 21894
rect 35900 21830 35952 21836
rect 35912 21146 35940 21830
rect 35900 21140 35952 21146
rect 35900 21082 35952 21088
rect 35900 20868 35952 20874
rect 35900 20810 35952 20816
rect 35912 20097 35940 20810
rect 35898 20088 35954 20097
rect 35898 20023 35954 20032
rect 35808 19916 35860 19922
rect 35808 19858 35860 19864
rect 35900 19916 35952 19922
rect 35900 19858 35952 19864
rect 35912 18902 35940 19858
rect 35900 18896 35952 18902
rect 35900 18838 35952 18844
rect 35808 18624 35860 18630
rect 35808 18566 35860 18572
rect 35716 17740 35768 17746
rect 35716 17682 35768 17688
rect 35716 16788 35768 16794
rect 35716 16730 35768 16736
rect 35624 15564 35676 15570
rect 35624 15506 35676 15512
rect 35622 15464 35678 15473
rect 35622 15399 35678 15408
rect 35532 14952 35584 14958
rect 35532 14894 35584 14900
rect 35530 14376 35586 14385
rect 35636 14362 35664 15399
rect 35728 14482 35756 16730
rect 35716 14476 35768 14482
rect 35716 14418 35768 14424
rect 35636 14334 35756 14362
rect 35530 14311 35586 14320
rect 34796 11630 34848 11636
rect 34704 5636 34756 5642
rect 34704 5578 34756 5584
rect 34808 5370 34836 11630
rect 35360 11614 35480 11642
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 35360 5370 35388 11614
rect 35544 6914 35572 14311
rect 35624 12300 35676 12306
rect 35624 12242 35676 12248
rect 35452 6886 35572 6914
rect 35636 6914 35664 12242
rect 35728 8566 35756 14334
rect 35820 10742 35848 18566
rect 35912 15434 35940 18838
rect 35900 15428 35952 15434
rect 35900 15370 35952 15376
rect 35912 15162 35940 15370
rect 35900 15156 35952 15162
rect 35900 15098 35952 15104
rect 35900 15020 35952 15026
rect 35900 14962 35952 14968
rect 35808 10736 35860 10742
rect 35808 10678 35860 10684
rect 35716 8560 35768 8566
rect 35716 8502 35768 8508
rect 35636 6886 35756 6914
rect 35452 5914 35480 6886
rect 35440 5908 35492 5914
rect 35440 5850 35492 5856
rect 35532 5772 35584 5778
rect 35532 5714 35584 5720
rect 34796 5364 34848 5370
rect 34796 5306 34848 5312
rect 35348 5364 35400 5370
rect 35348 5306 35400 5312
rect 34612 5160 34664 5166
rect 34612 5102 34664 5108
rect 34624 4185 34652 5102
rect 34704 5092 34756 5098
rect 34704 5034 34756 5040
rect 34610 4176 34666 4185
rect 34610 4111 34666 4120
rect 34612 4004 34664 4010
rect 34612 3946 34664 3952
rect 34624 3466 34652 3946
rect 34716 3942 34744 5034
rect 34796 4548 34848 4554
rect 34796 4490 34848 4496
rect 34808 4078 34836 4490
rect 35256 4480 35308 4486
rect 35256 4422 35308 4428
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34796 4072 34848 4078
rect 34796 4014 34848 4020
rect 34704 3936 34756 3942
rect 34704 3878 34756 3884
rect 34612 3460 34664 3466
rect 34612 3402 34664 3408
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 34796 2984 34848 2990
rect 34796 2926 34848 2932
rect 34612 2644 34664 2650
rect 34612 2586 34664 2592
rect 34624 2417 34652 2586
rect 34610 2408 34666 2417
rect 34610 2343 34666 2352
rect 34808 1578 34836 2926
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 35268 1986 35296 4422
rect 35544 3777 35572 5714
rect 35728 4826 35756 6886
rect 35912 5914 35940 14962
rect 35900 5908 35952 5914
rect 35900 5850 35952 5856
rect 35900 5772 35952 5778
rect 35900 5714 35952 5720
rect 35808 5704 35860 5710
rect 35808 5646 35860 5652
rect 35716 4820 35768 4826
rect 35716 4762 35768 4768
rect 35624 4684 35676 4690
rect 35624 4626 35676 4632
rect 35530 3768 35586 3777
rect 35530 3703 35586 3712
rect 35532 2372 35584 2378
rect 35532 2314 35584 2320
rect 35176 1958 35296 1986
rect 34808 1550 34928 1578
rect 34900 800 34928 1550
rect 35176 800 35204 1958
rect 35544 800 35572 2314
rect 35636 2009 35664 4626
rect 35622 2000 35678 2009
rect 35622 1935 35678 1944
rect 35820 1057 35848 5646
rect 35912 3369 35940 5714
rect 35898 3360 35954 3369
rect 35898 3295 35954 3304
rect 36004 2582 36032 51046
rect 36084 46980 36136 46986
rect 36084 46922 36136 46928
rect 36096 24274 36124 46922
rect 36188 40390 36216 58822
rect 36280 58585 36308 61202
rect 36266 58576 36322 58585
rect 36266 58511 36322 58520
rect 36268 58472 36320 58478
rect 36268 58414 36320 58420
rect 36280 52426 36308 58414
rect 36268 52420 36320 52426
rect 36268 52362 36320 52368
rect 36176 40384 36228 40390
rect 36176 40326 36228 40332
rect 36176 40112 36228 40118
rect 36176 40054 36228 40060
rect 36188 35834 36216 40054
rect 36372 38486 36400 64262
rect 36464 63753 36492 65554
rect 36450 63744 36506 63753
rect 36450 63679 36506 63688
rect 36452 63572 36504 63578
rect 36452 63514 36504 63520
rect 36464 62694 36492 63514
rect 36556 63034 36584 66966
rect 36648 66842 36676 67526
rect 36728 67108 36780 67114
rect 36728 67050 36780 67056
rect 36636 66836 36688 66842
rect 36636 66778 36688 66784
rect 36740 66774 36768 67050
rect 36728 66768 36780 66774
rect 36728 66710 36780 66716
rect 36636 65952 36688 65958
rect 36636 65894 36688 65900
rect 36544 63028 36596 63034
rect 36544 62970 36596 62976
rect 36648 62898 36676 65894
rect 36728 65544 36780 65550
rect 36728 65486 36780 65492
rect 36740 64938 36768 65486
rect 36728 64932 36780 64938
rect 36728 64874 36780 64880
rect 36740 64598 36768 64874
rect 36728 64592 36780 64598
rect 36728 64534 36780 64540
rect 36740 63617 36768 64534
rect 36726 63608 36782 63617
rect 36726 63543 36782 63552
rect 36728 63504 36780 63510
rect 36728 63446 36780 63452
rect 36636 62892 36688 62898
rect 36556 62852 36636 62880
rect 36452 62688 36504 62694
rect 36452 62630 36504 62636
rect 36556 62422 36584 62852
rect 36636 62834 36688 62840
rect 36740 62762 36768 63446
rect 36728 62756 36780 62762
rect 36728 62698 36780 62704
rect 36636 62688 36688 62694
rect 36636 62630 36688 62636
rect 36544 62416 36596 62422
rect 36544 62358 36596 62364
rect 36544 61668 36596 61674
rect 36544 61610 36596 61616
rect 36556 60722 36584 61610
rect 36544 60716 36596 60722
rect 36544 60658 36596 60664
rect 36452 60648 36504 60654
rect 36452 60590 36504 60596
rect 36464 58682 36492 60590
rect 36544 60512 36596 60518
rect 36544 60454 36596 60460
rect 36452 58676 36504 58682
rect 36452 58618 36504 58624
rect 36450 58576 36506 58585
rect 36450 58511 36506 58520
rect 36464 55962 36492 58511
rect 36452 55956 36504 55962
rect 36452 55898 36504 55904
rect 36452 45552 36504 45558
rect 36452 45494 36504 45500
rect 36360 38480 36412 38486
rect 36360 38422 36412 38428
rect 36360 36916 36412 36922
rect 36360 36858 36412 36864
rect 36268 36168 36320 36174
rect 36268 36110 36320 36116
rect 36176 35828 36228 35834
rect 36176 35770 36228 35776
rect 36176 35624 36228 35630
rect 36176 35566 36228 35572
rect 36188 33658 36216 35566
rect 36176 33652 36228 33658
rect 36176 33594 36228 33600
rect 36176 33516 36228 33522
rect 36176 33458 36228 33464
rect 36188 26518 36216 33458
rect 36176 26512 36228 26518
rect 36176 26454 36228 26460
rect 36176 25832 36228 25838
rect 36176 25774 36228 25780
rect 36188 24886 36216 25774
rect 36176 24880 36228 24886
rect 36176 24822 36228 24828
rect 36280 24750 36308 36110
rect 36372 33522 36400 36858
rect 36360 33516 36412 33522
rect 36360 33458 36412 33464
rect 36360 31680 36412 31686
rect 36360 31622 36412 31628
rect 36372 29034 36400 31622
rect 36360 29028 36412 29034
rect 36360 28970 36412 28976
rect 36360 27600 36412 27606
rect 36360 27542 36412 27548
rect 36372 25838 36400 27542
rect 36360 25832 36412 25838
rect 36360 25774 36412 25780
rect 36360 25356 36412 25362
rect 36360 25298 36412 25304
rect 36268 24744 36320 24750
rect 36268 24686 36320 24692
rect 36176 24608 36228 24614
rect 36176 24550 36228 24556
rect 36268 24608 36320 24614
rect 36268 24550 36320 24556
rect 36084 24268 36136 24274
rect 36084 24210 36136 24216
rect 36084 24132 36136 24138
rect 36188 24120 36216 24550
rect 36136 24092 36216 24120
rect 36084 24074 36136 24080
rect 36096 23730 36124 24074
rect 36084 23724 36136 23730
rect 36084 23666 36136 23672
rect 36096 23050 36124 23666
rect 36176 23656 36228 23662
rect 36176 23598 36228 23604
rect 36188 23118 36216 23598
rect 36176 23112 36228 23118
rect 36176 23054 36228 23060
rect 36084 23044 36136 23050
rect 36084 22986 36136 22992
rect 36096 22642 36124 22986
rect 36084 22636 36136 22642
rect 36084 22578 36136 22584
rect 36188 22574 36216 23054
rect 36176 22568 36228 22574
rect 36176 22510 36228 22516
rect 36084 22228 36136 22234
rect 36188 22216 36216 22510
rect 36136 22188 36216 22216
rect 36084 22170 36136 22176
rect 36096 20534 36124 22170
rect 36176 21956 36228 21962
rect 36176 21898 36228 21904
rect 36188 21010 36216 21898
rect 36176 21004 36228 21010
rect 36176 20946 36228 20952
rect 36188 20874 36216 20946
rect 36176 20868 36228 20874
rect 36176 20810 36228 20816
rect 36084 20528 36136 20534
rect 36084 20470 36136 20476
rect 36188 20466 36216 20810
rect 36176 20460 36228 20466
rect 36176 20402 36228 20408
rect 36084 20392 36136 20398
rect 36084 20334 36136 20340
rect 36096 19446 36124 20334
rect 36084 19440 36136 19446
rect 36084 19382 36136 19388
rect 36084 18964 36136 18970
rect 36084 18906 36136 18912
rect 36096 16794 36124 18906
rect 36188 18902 36216 20402
rect 36176 18896 36228 18902
rect 36176 18838 36228 18844
rect 36084 16788 36136 16794
rect 36084 16730 36136 16736
rect 36174 16552 36230 16561
rect 36174 16487 36230 16496
rect 36084 15088 36136 15094
rect 36084 15030 36136 15036
rect 36096 5914 36124 15030
rect 36188 6390 36216 16487
rect 36176 6384 36228 6390
rect 36176 6326 36228 6332
rect 36084 5908 36136 5914
rect 36084 5850 36136 5856
rect 36084 5160 36136 5166
rect 36084 5102 36136 5108
rect 35992 2576 36044 2582
rect 35992 2518 36044 2524
rect 35900 2508 35952 2514
rect 35900 2450 35952 2456
rect 35806 1048 35862 1057
rect 35806 983 35862 992
rect 35912 800 35940 2450
rect 36096 1465 36124 5102
rect 36280 3670 36308 24550
rect 36372 12986 36400 25298
rect 36464 23662 36492 45494
rect 36556 36922 36584 60454
rect 36648 40118 36676 62630
rect 36726 62248 36782 62257
rect 36726 62183 36728 62192
rect 36780 62183 36782 62192
rect 36728 62154 36780 62160
rect 36726 61976 36782 61985
rect 36726 61911 36782 61920
rect 36740 61742 36768 61911
rect 36728 61736 36780 61742
rect 36728 61678 36780 61684
rect 36728 61260 36780 61266
rect 36728 61202 36780 61208
rect 36740 61062 36768 61202
rect 36728 61056 36780 61062
rect 36728 60998 36780 61004
rect 36728 60716 36780 60722
rect 36728 60658 36780 60664
rect 36740 59566 36768 60658
rect 36728 59560 36780 59566
rect 36728 59502 36780 59508
rect 36740 59226 36768 59502
rect 36728 59220 36780 59226
rect 36728 59162 36780 59168
rect 36832 59090 36860 67646
rect 36924 67182 36952 69702
rect 37016 68762 37044 69770
rect 37108 68882 37136 70790
rect 37200 68921 37228 71998
rect 37280 71392 37332 71398
rect 37280 71334 37332 71340
rect 37292 69358 37320 71334
rect 37384 71176 37412 83846
rect 37476 81394 37504 87654
rect 37568 82890 37596 87774
rect 37556 82884 37608 82890
rect 37556 82826 37608 82832
rect 37556 82272 37608 82278
rect 37556 82214 37608 82220
rect 37464 81388 37516 81394
rect 37464 81330 37516 81336
rect 37568 71602 37596 82214
rect 37660 82074 37688 89286
rect 37752 83026 37780 91190
rect 37844 89026 37872 92006
rect 37936 91497 37964 92142
rect 37922 91488 37978 91497
rect 37922 91423 37978 91432
rect 37924 91112 37976 91118
rect 37924 91054 37976 91060
rect 37936 90545 37964 91054
rect 37922 90536 37978 90545
rect 37922 90471 37978 90480
rect 37924 90024 37976 90030
rect 37924 89966 37976 89972
rect 37936 89185 37964 89966
rect 37922 89176 37978 89185
rect 37922 89111 37978 89120
rect 37844 88998 38056 89026
rect 37924 88936 37976 88942
rect 37924 88878 37976 88884
rect 37832 88800 37884 88806
rect 37832 88742 37884 88748
rect 37740 83020 37792 83026
rect 37740 82962 37792 82968
rect 37740 82884 37792 82890
rect 37740 82826 37792 82832
rect 37648 82068 37700 82074
rect 37648 82010 37700 82016
rect 37648 81388 37700 81394
rect 37648 81330 37700 81336
rect 37660 80054 37688 81330
rect 37752 81326 37780 82826
rect 37740 81320 37792 81326
rect 37740 81262 37792 81268
rect 37844 80646 37872 88742
rect 37936 88369 37964 88878
rect 37922 88360 37978 88369
rect 37922 88295 37978 88304
rect 37924 87848 37976 87854
rect 37924 87790 37976 87796
rect 37936 87009 37964 87790
rect 37922 87000 37978 87009
rect 37922 86935 37978 86944
rect 37924 86760 37976 86766
rect 37924 86702 37976 86708
rect 37936 86057 37964 86702
rect 37922 86048 37978 86057
rect 37922 85983 37978 85992
rect 37924 85672 37976 85678
rect 37924 85614 37976 85620
rect 37936 85241 37964 85614
rect 37922 85232 37978 85241
rect 37922 85167 37978 85176
rect 37924 84584 37976 84590
rect 37924 84526 37976 84532
rect 37936 83881 37964 84526
rect 37922 83872 37978 83881
rect 37922 83807 37978 83816
rect 37924 83496 37976 83502
rect 37924 83438 37976 83444
rect 37936 82929 37964 83438
rect 37922 82920 37978 82929
rect 37922 82855 37978 82864
rect 38028 82482 38056 88998
rect 38120 83570 38148 93094
rect 38108 83564 38160 83570
rect 38108 83506 38160 83512
rect 38016 82476 38068 82482
rect 38016 82418 38068 82424
rect 37924 82408 37976 82414
rect 37924 82350 37976 82356
rect 37936 81569 37964 82350
rect 38212 82006 38240 103498
rect 38384 95940 38436 95946
rect 38384 95882 38436 95888
rect 38292 88800 38344 88806
rect 38292 88742 38344 88748
rect 38200 82000 38252 82006
rect 38200 81942 38252 81948
rect 37922 81560 37978 81569
rect 37922 81495 37978 81504
rect 37924 81320 37976 81326
rect 38304 81274 38332 88742
rect 37924 81262 37976 81268
rect 37936 80753 37964 81262
rect 38212 81246 38332 81274
rect 37922 80744 37978 80753
rect 37922 80679 37978 80688
rect 37832 80640 37884 80646
rect 37832 80582 37884 80588
rect 38212 80306 38240 81246
rect 38292 81184 38344 81190
rect 38292 81126 38344 81132
rect 38200 80300 38252 80306
rect 38200 80242 38252 80248
rect 37924 80232 37976 80238
rect 37924 80174 37976 80180
rect 37660 80026 37780 80054
rect 37648 76832 37700 76838
rect 37648 76774 37700 76780
rect 37556 71596 37608 71602
rect 37556 71538 37608 71544
rect 37464 71528 37516 71534
rect 37464 71470 37516 71476
rect 37476 71369 37504 71470
rect 37556 71392 37608 71398
rect 37462 71360 37518 71369
rect 37556 71334 37608 71340
rect 37462 71295 37518 71304
rect 37384 71148 37504 71176
rect 37372 71052 37424 71058
rect 37372 70994 37424 71000
rect 37384 70825 37412 70994
rect 37370 70816 37426 70825
rect 37370 70751 37426 70760
rect 37476 70530 37504 71148
rect 37384 70502 37504 70530
rect 37384 70106 37412 70502
rect 37464 70440 37516 70446
rect 37464 70382 37516 70388
rect 37372 70100 37424 70106
rect 37372 70042 37424 70048
rect 37372 69964 37424 69970
rect 37372 69906 37424 69912
rect 37280 69352 37332 69358
rect 37280 69294 37332 69300
rect 37280 69216 37332 69222
rect 37280 69158 37332 69164
rect 37292 68950 37320 69158
rect 37384 69057 37412 69906
rect 37476 69601 37504 70382
rect 37462 69592 37518 69601
rect 37462 69527 37518 69536
rect 37462 69456 37518 69465
rect 37462 69391 37518 69400
rect 37370 69048 37426 69057
rect 37370 68983 37426 68992
rect 37280 68944 37332 68950
rect 37186 68912 37242 68921
rect 37096 68876 37148 68882
rect 37280 68886 37332 68892
rect 37186 68847 37242 68856
rect 37096 68818 37148 68824
rect 37016 68734 37136 68762
rect 37002 68640 37058 68649
rect 37002 68575 37058 68584
rect 36912 67176 36964 67182
rect 36912 67118 36964 67124
rect 36912 66836 36964 66842
rect 36912 66778 36964 66784
rect 36924 66706 36952 66778
rect 36912 66700 36964 66706
rect 36912 66642 36964 66648
rect 36912 66496 36964 66502
rect 36912 66438 36964 66444
rect 36924 65006 36952 66438
rect 36912 65000 36964 65006
rect 36912 64942 36964 64948
rect 36910 64832 36966 64841
rect 36910 64767 36966 64776
rect 36924 64530 36952 64767
rect 36912 64524 36964 64530
rect 36912 64466 36964 64472
rect 36910 64016 36966 64025
rect 36910 63951 36966 63960
rect 36924 63918 36952 63951
rect 36912 63912 36964 63918
rect 36912 63854 36964 63860
rect 36912 63028 36964 63034
rect 36912 62970 36964 62976
rect 36924 60654 36952 62970
rect 36912 60648 36964 60654
rect 36912 60590 36964 60596
rect 36912 59492 36964 59498
rect 36912 59434 36964 59440
rect 36820 59084 36872 59090
rect 36820 59026 36872 59032
rect 36728 58880 36780 58886
rect 36728 58822 36780 58828
rect 36818 58848 36874 58857
rect 36740 58614 36768 58822
rect 36818 58783 36874 58792
rect 36728 58608 36780 58614
rect 36728 58550 36780 58556
rect 36728 58472 36780 58478
rect 36728 58414 36780 58420
rect 36740 58313 36768 58414
rect 36726 58304 36782 58313
rect 36726 58239 36782 58248
rect 36832 58002 36860 58783
rect 36924 58002 36952 59434
rect 37016 58478 37044 68575
rect 37108 67794 37136 68734
rect 37188 68740 37240 68746
rect 37188 68682 37240 68688
rect 37096 67788 37148 67794
rect 37096 67730 37148 67736
rect 37096 67108 37148 67114
rect 37096 67050 37148 67056
rect 37108 66706 37136 67050
rect 37200 66706 37228 68682
rect 37292 68202 37320 68886
rect 37370 68504 37426 68513
rect 37370 68439 37372 68448
rect 37424 68439 37426 68448
rect 37372 68410 37424 68416
rect 37372 68332 37424 68338
rect 37372 68274 37424 68280
rect 37280 68196 37332 68202
rect 37280 68138 37332 68144
rect 37292 67862 37320 68138
rect 37280 67856 37332 67862
rect 37280 67798 37332 67804
rect 37280 66768 37332 66774
rect 37280 66710 37332 66716
rect 37096 66700 37148 66706
rect 37096 66642 37148 66648
rect 37188 66700 37240 66706
rect 37188 66642 37240 66648
rect 37108 65958 37136 66642
rect 37292 66026 37320 66710
rect 37280 66020 37332 66026
rect 37280 65962 37332 65968
rect 37096 65952 37148 65958
rect 37096 65894 37148 65900
rect 37096 65612 37148 65618
rect 37096 65554 37148 65560
rect 37108 64938 37136 65554
rect 37188 65204 37240 65210
rect 37188 65146 37240 65152
rect 37096 64932 37148 64938
rect 37096 64874 37148 64880
rect 37108 64598 37136 64874
rect 37096 64592 37148 64598
rect 37096 64534 37148 64540
rect 37096 63776 37148 63782
rect 37096 63718 37148 63724
rect 37004 58472 37056 58478
rect 37004 58414 37056 58420
rect 36820 57996 36872 58002
rect 36820 57938 36872 57944
rect 36912 57996 36964 58002
rect 36912 57938 36964 57944
rect 37004 55956 37056 55962
rect 37004 55898 37056 55904
rect 36820 55888 36872 55894
rect 36820 55830 36872 55836
rect 36728 53644 36780 53650
rect 36728 53586 36780 53592
rect 36740 53417 36768 53586
rect 36726 53408 36782 53417
rect 36726 53343 36782 53352
rect 36728 44192 36780 44198
rect 36728 44134 36780 44140
rect 36636 40112 36688 40118
rect 36636 40054 36688 40060
rect 36636 39840 36688 39846
rect 36636 39782 36688 39788
rect 36544 36916 36596 36922
rect 36544 36858 36596 36864
rect 36544 33856 36596 33862
rect 36544 33798 36596 33804
rect 36556 25430 36584 33798
rect 36648 31822 36676 39782
rect 36740 32858 36768 44134
rect 36832 42770 36860 55830
rect 36820 42764 36872 42770
rect 36820 42706 36872 42712
rect 36820 40384 36872 40390
rect 36820 40326 36872 40332
rect 36832 33046 36860 40326
rect 36820 33040 36872 33046
rect 36820 32982 36872 32988
rect 36740 32830 36952 32858
rect 36820 31884 36872 31890
rect 36820 31826 36872 31832
rect 36636 31816 36688 31822
rect 36636 31758 36688 31764
rect 36728 31408 36780 31414
rect 36728 31350 36780 31356
rect 36636 30796 36688 30802
rect 36636 30738 36688 30744
rect 36648 26586 36676 30738
rect 36636 26580 36688 26586
rect 36636 26522 36688 26528
rect 36636 25764 36688 25770
rect 36636 25706 36688 25712
rect 36544 25424 36596 25430
rect 36544 25366 36596 25372
rect 36544 25288 36596 25294
rect 36544 25230 36596 25236
rect 36452 23656 36504 23662
rect 36452 23598 36504 23604
rect 36556 22778 36584 25230
rect 36544 22772 36596 22778
rect 36544 22714 36596 22720
rect 36544 22636 36596 22642
rect 36544 22578 36596 22584
rect 36452 22500 36504 22506
rect 36452 22442 36504 22448
rect 36360 12980 36412 12986
rect 36360 12922 36412 12928
rect 36464 10810 36492 22442
rect 36556 19990 36584 22578
rect 36544 19984 36596 19990
rect 36544 19926 36596 19932
rect 36648 17320 36676 25706
rect 36740 22574 36768 31350
rect 36832 29306 36860 31826
rect 36924 31414 36952 32830
rect 36912 31408 36964 31414
rect 36912 31350 36964 31356
rect 36912 31272 36964 31278
rect 36912 31214 36964 31220
rect 36820 29300 36872 29306
rect 36820 29242 36872 29248
rect 36820 29028 36872 29034
rect 36820 28970 36872 28976
rect 36832 24614 36860 28970
rect 36924 28218 36952 31214
rect 36912 28212 36964 28218
rect 36912 28154 36964 28160
rect 36912 28008 36964 28014
rect 36912 27950 36964 27956
rect 36924 27062 36952 27950
rect 36912 27056 36964 27062
rect 36912 26998 36964 27004
rect 36912 25764 36964 25770
rect 36912 25706 36964 25712
rect 36820 24608 36872 24614
rect 36820 24550 36872 24556
rect 36820 23588 36872 23594
rect 36820 23530 36872 23536
rect 36728 22568 36780 22574
rect 36728 22510 36780 22516
rect 36728 22432 36780 22438
rect 36728 22374 36780 22380
rect 36740 22098 36768 22374
rect 36728 22092 36780 22098
rect 36728 22034 36780 22040
rect 36728 21412 36780 21418
rect 36728 21354 36780 21360
rect 36740 20398 36768 21354
rect 36728 20392 36780 20398
rect 36728 20334 36780 20340
rect 36648 17292 36768 17320
rect 36544 17264 36596 17270
rect 36544 17206 36596 17212
rect 36556 11898 36584 17206
rect 36636 17196 36688 17202
rect 36636 17138 36688 17144
rect 36544 11892 36596 11898
rect 36544 11834 36596 11840
rect 36648 11830 36676 17138
rect 36740 13530 36768 17292
rect 36832 17202 36860 23530
rect 36924 21010 36952 25706
rect 36912 21004 36964 21010
rect 36912 20946 36964 20952
rect 36912 18760 36964 18766
rect 36912 18702 36964 18708
rect 36820 17196 36872 17202
rect 36820 17138 36872 17144
rect 36728 13524 36780 13530
rect 36728 13466 36780 13472
rect 36820 12096 36872 12102
rect 36820 12038 36872 12044
rect 36636 11824 36688 11830
rect 36636 11766 36688 11772
rect 36452 10804 36504 10810
rect 36452 10746 36504 10752
rect 36832 6458 36860 12038
rect 36924 7478 36952 18702
rect 36912 7472 36964 7478
rect 36912 7414 36964 7420
rect 36820 6452 36872 6458
rect 36820 6394 36872 6400
rect 36912 6248 36964 6254
rect 36912 6190 36964 6196
rect 36728 5160 36780 5166
rect 36728 5102 36780 5108
rect 36360 4752 36412 4758
rect 36360 4694 36412 4700
rect 36372 3942 36400 4694
rect 36452 4684 36504 4690
rect 36452 4626 36504 4632
rect 36464 4593 36492 4626
rect 36450 4584 36506 4593
rect 36450 4519 36506 4528
rect 36636 4004 36688 4010
rect 36636 3946 36688 3952
rect 36360 3936 36412 3942
rect 36360 3878 36412 3884
rect 36268 3664 36320 3670
rect 36268 3606 36320 3612
rect 36648 3602 36676 3946
rect 36636 3596 36688 3602
rect 36636 3538 36688 3544
rect 36176 3392 36228 3398
rect 36176 3334 36228 3340
rect 36082 1456 36138 1465
rect 36082 1391 36138 1400
rect 36188 800 36216 3334
rect 36544 2848 36596 2854
rect 36544 2790 36596 2796
rect 36556 800 36584 2790
rect 2870 368 2926 377
rect 2870 303 2926 312
rect 2962 -800 3018 800
rect 3330 -800 3386 800
rect 3606 -800 3662 800
rect 3974 -800 4030 800
rect 4250 -800 4306 800
rect 4618 -800 4674 800
rect 4986 -800 5042 800
rect 5262 -800 5318 800
rect 5630 -800 5686 800
rect 5906 -800 5962 800
rect 6274 -800 6330 800
rect 6550 -800 6606 800
rect 6918 -800 6974 800
rect 7194 -800 7250 800
rect 7562 -800 7618 800
rect 7838 -800 7894 800
rect 8206 -800 8262 800
rect 8482 -800 8538 800
rect 8850 -800 8906 800
rect 9218 -800 9274 800
rect 9494 -800 9550 800
rect 9862 -800 9918 800
rect 10138 -800 10194 800
rect 10506 -800 10562 800
rect 10782 -800 10838 800
rect 11150 -800 11206 800
rect 11426 -800 11482 800
rect 11794 -800 11850 800
rect 12070 -800 12126 800
rect 12438 -800 12494 800
rect 12714 -800 12770 800
rect 13082 -800 13138 800
rect 13450 -800 13506 800
rect 13726 -800 13782 800
rect 14094 -800 14150 800
rect 14370 -800 14426 800
rect 14738 -800 14794 800
rect 15014 -800 15070 800
rect 15382 -800 15438 800
rect 15658 -800 15714 800
rect 16026 -800 16082 800
rect 16302 -800 16358 800
rect 16670 -800 16726 800
rect 16946 -800 17002 800
rect 17314 -800 17370 800
rect 17590 -800 17646 800
rect 17958 -800 18014 800
rect 18326 -800 18382 800
rect 18602 -800 18658 800
rect 18970 -800 19026 800
rect 19246 -800 19302 800
rect 19614 -800 19670 800
rect 19890 -800 19946 800
rect 20258 -800 20314 800
rect 20534 -800 20590 800
rect 20902 -800 20958 800
rect 21178 -800 21234 800
rect 21546 -800 21602 800
rect 21822 -800 21878 800
rect 22190 -800 22246 800
rect 22558 -800 22614 800
rect 22834 -800 22890 800
rect 23202 -800 23258 800
rect 23478 -800 23534 800
rect 23846 -800 23902 800
rect 24122 -800 24178 800
rect 24490 -800 24546 800
rect 24766 -800 24822 800
rect 25134 -800 25190 800
rect 25410 -800 25466 800
rect 25778 -800 25834 800
rect 26054 -800 26110 800
rect 26422 -800 26478 800
rect 26790 -800 26846 800
rect 27066 -800 27122 800
rect 27434 -800 27490 800
rect 27710 -800 27766 800
rect 28078 -800 28134 800
rect 28354 -800 28410 800
rect 28722 -800 28778 800
rect 28998 -800 29054 800
rect 29366 -800 29422 800
rect 29642 -800 29698 800
rect 30010 -800 30066 800
rect 30286 -800 30342 800
rect 30654 -800 30710 800
rect 30930 -800 30986 800
rect 31298 -800 31354 800
rect 31666 -800 31722 800
rect 31942 -800 31998 800
rect 32310 -800 32366 800
rect 32586 -800 32642 800
rect 32954 -800 33010 800
rect 33230 -800 33286 800
rect 33598 -800 33654 800
rect 33874 -800 33930 800
rect 34242 -800 34298 800
rect 34518 -800 34574 800
rect 34886 -800 34942 800
rect 35162 -800 35218 800
rect 35530 -800 35586 800
rect 35898 -800 35954 800
rect 36174 -800 36230 800
rect 36542 -800 36598 800
rect 36740 649 36768 5102
rect 36820 3460 36872 3466
rect 36820 3402 36872 3408
rect 36832 800 36860 3402
rect 36924 2825 36952 6190
rect 36910 2816 36966 2825
rect 36910 2751 36966 2760
rect 37016 2310 37044 55898
rect 37108 37874 37136 63718
rect 37200 60092 37228 65146
rect 37292 64122 37320 65962
rect 37280 64116 37332 64122
rect 37280 64058 37332 64064
rect 37278 63880 37334 63889
rect 37278 63815 37334 63824
rect 37292 63442 37320 63815
rect 37280 63436 37332 63442
rect 37280 63378 37332 63384
rect 37280 62960 37332 62966
rect 37278 62928 37280 62937
rect 37332 62928 37334 62937
rect 37278 62863 37334 62872
rect 37280 62416 37332 62422
rect 37280 62358 37332 62364
rect 37292 61674 37320 62358
rect 37384 61810 37412 68274
rect 37476 67634 37504 69391
rect 37568 68270 37596 71334
rect 37660 70258 37688 76774
rect 37752 73030 37780 80026
rect 37936 79393 37964 80174
rect 37922 79384 37978 79393
rect 37922 79319 37978 79328
rect 37924 79144 37976 79150
rect 37924 79086 37976 79092
rect 37936 78441 37964 79086
rect 37922 78432 37978 78441
rect 37922 78367 37978 78376
rect 37924 78056 37976 78062
rect 37924 77998 37976 78004
rect 37936 77625 37964 77998
rect 38200 77920 38252 77926
rect 38200 77862 38252 77868
rect 37922 77616 37978 77625
rect 37922 77551 37978 77560
rect 38016 76968 38068 76974
rect 38016 76910 38068 76916
rect 37832 76832 37884 76838
rect 37832 76774 37884 76780
rect 37740 73024 37792 73030
rect 37740 72966 37792 72972
rect 37844 72842 37872 76774
rect 37922 76664 37978 76673
rect 37922 76599 37978 76608
rect 37936 75886 37964 76599
rect 38028 76265 38056 76910
rect 38014 76256 38070 76265
rect 38014 76191 38070 76200
rect 37924 75880 37976 75886
rect 37924 75822 37976 75828
rect 37924 74792 37976 74798
rect 37924 74734 37976 74740
rect 37936 74089 37964 74734
rect 37922 74080 37978 74089
rect 37922 74015 37978 74024
rect 37924 73704 37976 73710
rect 37924 73646 37976 73652
rect 37936 73137 37964 73646
rect 37922 73128 37978 73137
rect 37922 73063 37978 73072
rect 37924 73024 37976 73030
rect 37924 72966 37976 72972
rect 37752 72814 37872 72842
rect 37752 70378 37780 72814
rect 37832 70576 37884 70582
rect 37832 70518 37884 70524
rect 37740 70372 37792 70378
rect 37740 70314 37792 70320
rect 37660 70230 37780 70258
rect 37648 70100 37700 70106
rect 37648 70042 37700 70048
rect 37556 68264 37608 68270
rect 37556 68206 37608 68212
rect 37660 67930 37688 70042
rect 37648 67924 37700 67930
rect 37648 67866 37700 67872
rect 37476 67606 37596 67634
rect 37464 64864 37516 64870
rect 37464 64806 37516 64812
rect 37568 64818 37596 67606
rect 37648 67108 37700 67114
rect 37648 67050 37700 67056
rect 37660 66774 37688 67050
rect 37648 66768 37700 66774
rect 37648 66710 37700 66716
rect 37648 65680 37700 65686
rect 37648 65622 37700 65628
rect 37660 64977 37688 65622
rect 37646 64968 37702 64977
rect 37646 64903 37702 64912
rect 37476 64598 37504 64806
rect 37568 64790 37688 64818
rect 37554 64696 37610 64705
rect 37554 64631 37610 64640
rect 37464 64592 37516 64598
rect 37464 64534 37516 64540
rect 37476 63850 37504 64534
rect 37568 64530 37596 64631
rect 37556 64524 37608 64530
rect 37556 64466 37608 64472
rect 37660 64462 37688 64790
rect 37648 64456 37700 64462
rect 37648 64398 37700 64404
rect 37556 64116 37608 64122
rect 37556 64058 37608 64064
rect 37568 63918 37596 64058
rect 37556 63912 37608 63918
rect 37556 63854 37608 63860
rect 37648 63912 37700 63918
rect 37648 63854 37700 63860
rect 37464 63844 37516 63850
rect 37464 63786 37516 63792
rect 37476 63306 37504 63786
rect 37660 63617 37688 63854
rect 37646 63608 37702 63617
rect 37646 63543 37702 63552
rect 37556 63504 37608 63510
rect 37554 63472 37556 63481
rect 37608 63472 37610 63481
rect 37554 63407 37610 63416
rect 37464 63300 37516 63306
rect 37464 63242 37516 63248
rect 37752 63050 37780 70230
rect 37844 67250 37872 70518
rect 37936 70417 37964 72966
rect 38108 71528 38160 71534
rect 38108 71470 38160 71476
rect 38016 70576 38068 70582
rect 38016 70518 38068 70524
rect 37922 70408 37978 70417
rect 37922 70343 37978 70352
rect 37924 70304 37976 70310
rect 37924 70246 37976 70252
rect 37936 68338 37964 70246
rect 38028 69306 38056 70518
rect 38120 70417 38148 71470
rect 38106 70408 38162 70417
rect 38106 70343 38162 70352
rect 38212 69562 38240 77862
rect 38304 75002 38332 81126
rect 38396 76022 38424 95882
rect 38384 76016 38436 76022
rect 38384 75958 38436 75964
rect 38292 74996 38344 75002
rect 38292 74938 38344 74944
rect 38384 72480 38436 72486
rect 38384 72422 38436 72428
rect 38292 70440 38344 70446
rect 38292 70382 38344 70388
rect 38200 69556 38252 69562
rect 38200 69498 38252 69504
rect 38200 69420 38252 69426
rect 38200 69362 38252 69368
rect 38028 69278 38148 69306
rect 38016 69216 38068 69222
rect 38016 69158 38068 69164
rect 37924 68332 37976 68338
rect 37924 68274 37976 68280
rect 37924 68128 37976 68134
rect 37924 68070 37976 68076
rect 37832 67244 37884 67250
rect 37832 67186 37884 67192
rect 37832 66496 37884 66502
rect 37832 66438 37884 66444
rect 37660 63022 37780 63050
rect 37556 62960 37608 62966
rect 37556 62902 37608 62908
rect 37464 62824 37516 62830
rect 37464 62766 37516 62772
rect 37476 62490 37504 62766
rect 37464 62484 37516 62490
rect 37464 62426 37516 62432
rect 37464 62348 37516 62354
rect 37464 62290 37516 62296
rect 37476 62257 37504 62290
rect 37568 62286 37596 62902
rect 37660 62694 37688 63022
rect 37648 62688 37700 62694
rect 37648 62630 37700 62636
rect 37556 62280 37608 62286
rect 37462 62248 37518 62257
rect 37556 62222 37608 62228
rect 37462 62183 37518 62192
rect 37464 61872 37516 61878
rect 37464 61814 37516 61820
rect 37372 61804 37424 61810
rect 37372 61746 37424 61752
rect 37280 61668 37332 61674
rect 37280 61610 37332 61616
rect 37292 61334 37320 61610
rect 37280 61328 37332 61334
rect 37280 61270 37332 61276
rect 37292 60654 37320 61270
rect 37476 60654 37504 61814
rect 37568 61674 37596 62222
rect 37740 61872 37792 61878
rect 37740 61814 37792 61820
rect 37556 61668 37608 61674
rect 37556 61610 37608 61616
rect 37568 61402 37596 61610
rect 37556 61396 37608 61402
rect 37556 61338 37608 61344
rect 37280 60648 37332 60654
rect 37280 60590 37332 60596
rect 37464 60648 37516 60654
rect 37464 60590 37516 60596
rect 37568 60586 37596 61338
rect 37556 60580 37608 60586
rect 37556 60522 37608 60528
rect 37372 60240 37424 60246
rect 37372 60182 37424 60188
rect 37280 60104 37332 60110
rect 37200 60064 37280 60092
rect 37200 59974 37228 60064
rect 37280 60046 37332 60052
rect 37188 59968 37240 59974
rect 37188 59910 37240 59916
rect 37200 59498 37228 59910
rect 37384 59498 37412 60182
rect 37188 59492 37240 59498
rect 37188 59434 37240 59440
rect 37372 59492 37424 59498
rect 37372 59434 37424 59440
rect 37200 59226 37228 59434
rect 37188 59220 37240 59226
rect 37188 59162 37240 59168
rect 37200 58562 37228 59162
rect 37384 59158 37412 59434
rect 37372 59152 37424 59158
rect 37372 59094 37424 59100
rect 37280 59084 37332 59090
rect 37280 59026 37332 59032
rect 37292 58682 37320 59026
rect 37280 58676 37332 58682
rect 37280 58618 37332 58624
rect 37200 58534 37320 58562
rect 37188 58472 37240 58478
rect 37188 58414 37240 58420
rect 37200 58138 37228 58414
rect 37292 58410 37320 58534
rect 37384 58410 37412 59094
rect 37280 58404 37332 58410
rect 37280 58346 37332 58352
rect 37372 58404 37424 58410
rect 37372 58346 37424 58352
rect 37188 58132 37240 58138
rect 37188 58074 37240 58080
rect 37280 58064 37332 58070
rect 37280 58006 37332 58012
rect 37188 57996 37240 58002
rect 37188 57938 37240 57944
rect 37200 57905 37228 57938
rect 37186 57896 37242 57905
rect 37186 57831 37242 57840
rect 37292 57594 37320 58006
rect 37280 57588 37332 57594
rect 37280 57530 37332 57536
rect 37462 57488 37518 57497
rect 37462 57423 37518 57432
rect 37476 57390 37504 57423
rect 37464 57384 37516 57390
rect 37464 57326 37516 57332
rect 37648 56704 37700 56710
rect 37648 56646 37700 56652
rect 37464 56296 37516 56302
rect 37464 56238 37516 56244
rect 37476 56137 37504 56238
rect 37556 56160 37608 56166
rect 37462 56128 37518 56137
rect 37556 56102 37608 56108
rect 37462 56063 37518 56072
rect 37188 55820 37240 55826
rect 37188 55762 37240 55768
rect 37200 55729 37228 55762
rect 37186 55720 37242 55729
rect 37186 55655 37242 55664
rect 37464 55208 37516 55214
rect 37464 55150 37516 55156
rect 37372 55072 37424 55078
rect 37372 55014 37424 55020
rect 37188 54732 37240 54738
rect 37188 54674 37240 54680
rect 37200 54369 37228 54674
rect 37186 54360 37242 54369
rect 37186 54295 37242 54304
rect 37186 53816 37242 53825
rect 37186 53751 37242 53760
rect 37200 53650 37228 53751
rect 37188 53644 37240 53650
rect 37188 53586 37240 53592
rect 37280 53032 37332 53038
rect 37278 53000 37280 53009
rect 37332 53000 37334 53009
rect 37278 52935 37334 52944
rect 37186 51640 37242 51649
rect 37186 51575 37242 51584
rect 37200 51474 37228 51575
rect 37384 51542 37412 55014
rect 37476 54777 37504 55150
rect 37462 54768 37518 54777
rect 37462 54703 37518 54712
rect 37462 52048 37518 52057
rect 37568 52018 37596 56102
rect 37462 51983 37518 51992
rect 37556 52012 37608 52018
rect 37476 51950 37504 51983
rect 37556 51954 37608 51960
rect 37464 51944 37516 51950
rect 37464 51886 37516 51892
rect 37372 51536 37424 51542
rect 37372 51478 37424 51484
rect 37188 51468 37240 51474
rect 37188 51410 37240 51416
rect 37464 50856 37516 50862
rect 37464 50798 37516 50804
rect 37476 50697 37504 50798
rect 37556 50720 37608 50726
rect 37462 50688 37518 50697
rect 37556 50662 37608 50668
rect 37462 50623 37518 50632
rect 37370 49464 37426 49473
rect 37370 49399 37426 49408
rect 37384 49298 37412 49399
rect 37372 49292 37424 49298
rect 37372 49234 37424 49240
rect 37278 48920 37334 48929
rect 37278 48855 37334 48864
rect 37292 48686 37320 48855
rect 37280 48680 37332 48686
rect 37280 48622 37332 48628
rect 37372 48204 37424 48210
rect 37372 48146 37424 48152
rect 37384 48113 37412 48146
rect 37370 48104 37426 48113
rect 37370 48039 37426 48048
rect 37280 47592 37332 47598
rect 37278 47560 37280 47569
rect 37332 47560 37334 47569
rect 37278 47495 37334 47504
rect 37568 47122 37596 50662
rect 37556 47116 37608 47122
rect 37556 47058 37608 47064
rect 37462 46744 37518 46753
rect 37462 46679 37518 46688
rect 37476 46510 37504 46679
rect 37464 46504 37516 46510
rect 37464 46446 37516 46452
rect 37186 46200 37242 46209
rect 37186 46135 37242 46144
rect 37200 46034 37228 46135
rect 37188 46028 37240 46034
rect 37188 45970 37240 45976
rect 37464 45416 37516 45422
rect 37462 45384 37464 45393
rect 37516 45384 37518 45393
rect 37462 45319 37518 45328
rect 37188 44328 37240 44334
rect 37188 44270 37240 44276
rect 37200 44033 37228 44270
rect 37280 44192 37332 44198
rect 37280 44134 37332 44140
rect 37186 44024 37242 44033
rect 37186 43959 37242 43968
rect 37188 43852 37240 43858
rect 37188 43794 37240 43800
rect 37200 43625 37228 43794
rect 37186 43616 37242 43625
rect 37186 43551 37242 43560
rect 37292 42362 37320 44134
rect 37372 42764 37424 42770
rect 37372 42706 37424 42712
rect 37384 42673 37412 42706
rect 37370 42664 37426 42673
rect 37370 42599 37426 42608
rect 37280 42356 37332 42362
rect 37280 42298 37332 42304
rect 37278 42256 37334 42265
rect 37278 42191 37334 42200
rect 37292 42158 37320 42191
rect 37280 42152 37332 42158
rect 37280 42094 37332 42100
rect 37188 41676 37240 41682
rect 37188 41618 37240 41624
rect 37200 41313 37228 41618
rect 37186 41304 37242 41313
rect 37186 41239 37242 41248
rect 37280 41064 37332 41070
rect 37280 41006 37332 41012
rect 37292 40905 37320 41006
rect 37278 40896 37334 40905
rect 37278 40831 37334 40840
rect 37464 39976 37516 39982
rect 37462 39944 37464 39953
rect 37516 39944 37518 39953
rect 37462 39879 37518 39888
rect 37280 39500 37332 39506
rect 37280 39442 37332 39448
rect 37292 39098 37320 39442
rect 37280 39092 37332 39098
rect 37280 39034 37332 39040
rect 37464 38888 37516 38894
rect 37464 38830 37516 38836
rect 37476 38729 37504 38830
rect 37462 38720 37518 38729
rect 37462 38655 37518 38664
rect 37188 38412 37240 38418
rect 37188 38354 37240 38360
rect 37200 38185 37228 38354
rect 37186 38176 37242 38185
rect 37186 38111 37242 38120
rect 37096 37868 37148 37874
rect 37096 37810 37148 37816
rect 37188 37800 37240 37806
rect 37188 37742 37240 37748
rect 37200 37466 37228 37742
rect 37188 37460 37240 37466
rect 37188 37402 37240 37408
rect 37370 37360 37426 37369
rect 37370 37295 37372 37304
rect 37424 37295 37426 37304
rect 37372 37266 37424 37272
rect 37278 36816 37334 36825
rect 37278 36751 37334 36760
rect 37292 36718 37320 36751
rect 37096 36712 37148 36718
rect 37096 36654 37148 36660
rect 37280 36712 37332 36718
rect 37280 36654 37332 36660
rect 37108 36378 37136 36654
rect 37096 36372 37148 36378
rect 37096 36314 37148 36320
rect 37372 36236 37424 36242
rect 37372 36178 37424 36184
rect 37384 36009 37412 36178
rect 37370 36000 37426 36009
rect 37370 35935 37426 35944
rect 37280 35624 37332 35630
rect 37280 35566 37332 35572
rect 37292 35465 37320 35566
rect 37278 35456 37334 35465
rect 37278 35391 37334 35400
rect 37096 35080 37148 35086
rect 37096 35022 37148 35028
rect 37108 32026 37136 35022
rect 37462 34640 37518 34649
rect 37462 34575 37518 34584
rect 37476 34542 37504 34575
rect 37464 34536 37516 34542
rect 37464 34478 37516 34484
rect 37464 33448 37516 33454
rect 37464 33390 37516 33396
rect 37476 33289 37504 33390
rect 37462 33280 37518 33289
rect 37462 33215 37518 33224
rect 37188 32972 37240 32978
rect 37188 32914 37240 32920
rect 37200 32881 37228 32914
rect 37186 32872 37242 32881
rect 37186 32807 37242 32816
rect 37188 32360 37240 32366
rect 37188 32302 37240 32308
rect 37096 32020 37148 32026
rect 37096 31962 37148 31968
rect 37096 31816 37148 31822
rect 37096 31758 37148 31764
rect 37108 25770 37136 31758
rect 37200 30938 37228 32302
rect 37370 31920 37426 31929
rect 37370 31855 37372 31864
rect 37424 31855 37426 31864
rect 37372 31826 37424 31832
rect 37278 31512 37334 31521
rect 37278 31447 37334 31456
rect 37292 31278 37320 31447
rect 37280 31272 37332 31278
rect 37280 31214 37332 31220
rect 37188 30932 37240 30938
rect 37188 30874 37240 30880
rect 37372 30796 37424 30802
rect 37372 30738 37424 30744
rect 37384 30569 37412 30738
rect 37370 30560 37426 30569
rect 37370 30495 37426 30504
rect 37280 30184 37332 30190
rect 37278 30152 37280 30161
rect 37332 30152 37334 30161
rect 37278 30087 37334 30096
rect 37280 30048 37332 30054
rect 37280 29990 37332 29996
rect 37188 27532 37240 27538
rect 37188 27474 37240 27480
rect 37200 27441 37228 27474
rect 37186 27432 37242 27441
rect 37186 27367 37242 27376
rect 37188 27056 37240 27062
rect 37188 26998 37240 27004
rect 37096 25764 37148 25770
rect 37096 25706 37148 25712
rect 37200 25514 37228 26998
rect 37292 26330 37320 29990
rect 37462 29200 37518 29209
rect 37462 29135 37518 29144
rect 37476 29102 37504 29135
rect 37464 29096 37516 29102
rect 37464 29038 37516 29044
rect 37464 28008 37516 28014
rect 37462 27976 37464 27985
rect 37516 27976 37518 27985
rect 37462 27911 37518 27920
rect 37464 27600 37516 27606
rect 37464 27542 37516 27548
rect 37370 26616 37426 26625
rect 37370 26551 37426 26560
rect 37384 26450 37412 26551
rect 37372 26444 37424 26450
rect 37372 26386 37424 26392
rect 37292 26302 37412 26330
rect 37278 26072 37334 26081
rect 37278 26007 37334 26016
rect 37292 25838 37320 26007
rect 37280 25832 37332 25838
rect 37280 25774 37332 25780
rect 37108 25486 37228 25514
rect 37384 25498 37412 26302
rect 37372 25492 37424 25498
rect 37108 25106 37136 25486
rect 37372 25434 37424 25440
rect 37188 25356 37240 25362
rect 37188 25298 37240 25304
rect 37200 25265 37228 25298
rect 37186 25256 37242 25265
rect 37186 25191 37242 25200
rect 37108 25078 37228 25106
rect 37096 24676 37148 24682
rect 37096 24618 37148 24624
rect 37108 17270 37136 24618
rect 37200 24410 37228 25078
rect 37278 24848 37334 24857
rect 37278 24783 37334 24792
rect 37292 24750 37320 24783
rect 37280 24744 37332 24750
rect 37280 24686 37332 24692
rect 37188 24404 37240 24410
rect 37188 24346 37240 24352
rect 37372 24268 37424 24274
rect 37372 24210 37424 24216
rect 37384 23905 37412 24210
rect 37370 23896 37426 23905
rect 37188 23860 37240 23866
rect 37370 23831 37426 23840
rect 37188 23802 37240 23808
rect 37200 21622 37228 23802
rect 37280 23656 37332 23662
rect 37280 23598 37332 23604
rect 37292 23497 37320 23598
rect 37278 23488 37334 23497
rect 37278 23423 37334 23432
rect 37372 22976 37424 22982
rect 37372 22918 37424 22924
rect 37280 22568 37332 22574
rect 37278 22536 37280 22545
rect 37332 22536 37334 22545
rect 37278 22471 37334 22480
rect 37188 21616 37240 21622
rect 37188 21558 37240 21564
rect 37280 21480 37332 21486
rect 37280 21422 37332 21428
rect 37292 21185 37320 21422
rect 37278 21176 37334 21185
rect 37278 21111 37334 21120
rect 37188 21004 37240 21010
rect 37188 20946 37240 20952
rect 37200 20777 37228 20946
rect 37186 20768 37242 20777
rect 37186 20703 37242 20712
rect 37188 19916 37240 19922
rect 37188 19858 37240 19864
rect 37200 19825 37228 19858
rect 37186 19816 37242 19825
rect 37186 19751 37242 19760
rect 37384 19700 37412 22918
rect 37476 22778 37504 27542
rect 37556 26920 37608 26926
rect 37556 26862 37608 26868
rect 37464 22772 37516 22778
rect 37464 22714 37516 22720
rect 37462 22128 37518 22137
rect 37462 22063 37518 22072
rect 37476 20890 37504 22063
rect 37568 21690 37596 26862
rect 37556 21684 37608 21690
rect 37556 21626 37608 21632
rect 37476 20862 37596 20890
rect 37464 20800 37516 20806
rect 37464 20742 37516 20748
rect 37200 19672 37412 19700
rect 37200 18986 37228 19672
rect 37278 19408 37334 19417
rect 37278 19343 37334 19352
rect 37292 19310 37320 19343
rect 37280 19304 37332 19310
rect 37280 19246 37332 19252
rect 37200 18958 37320 18986
rect 37188 18828 37240 18834
rect 37188 18770 37240 18776
rect 37200 18465 37228 18770
rect 37186 18456 37242 18465
rect 37186 18391 37242 18400
rect 37292 18306 37320 18958
rect 37200 18278 37320 18306
rect 37096 17264 37148 17270
rect 37096 17206 37148 17212
rect 37200 17082 37228 18278
rect 37280 18216 37332 18222
rect 37280 18158 37332 18164
rect 37292 18057 37320 18158
rect 37278 18048 37334 18057
rect 37278 17983 37334 17992
rect 37278 17232 37334 17241
rect 37278 17167 37334 17176
rect 37292 17134 37320 17167
rect 37108 17054 37228 17082
rect 37280 17128 37332 17134
rect 37280 17070 37332 17076
rect 37108 11354 37136 17054
rect 37476 16674 37504 20742
rect 37568 18630 37596 20862
rect 37556 18624 37608 18630
rect 37556 18566 37608 18572
rect 37556 16992 37608 16998
rect 37556 16934 37608 16940
rect 37384 16646 37504 16674
rect 37280 16040 37332 16046
rect 37280 15982 37332 15988
rect 37292 15881 37320 15982
rect 37278 15872 37334 15881
rect 37278 15807 37334 15816
rect 37188 15564 37240 15570
rect 37188 15506 37240 15512
rect 37200 15337 37228 15506
rect 37186 15328 37242 15337
rect 37186 15263 37242 15272
rect 37186 14512 37242 14521
rect 37186 14447 37188 14456
rect 37240 14447 37242 14456
rect 37188 14418 37240 14424
rect 37278 14104 37334 14113
rect 37278 14039 37334 14048
rect 37292 13870 37320 14039
rect 37280 13864 37332 13870
rect 37280 13806 37332 13812
rect 37186 13560 37242 13569
rect 37186 13495 37242 13504
rect 37200 13394 37228 13495
rect 37188 13388 37240 13394
rect 37188 13330 37240 13336
rect 37280 12776 37332 12782
rect 37278 12744 37280 12753
rect 37332 12744 37334 12753
rect 37278 12679 37334 12688
rect 37278 11792 37334 11801
rect 37278 11727 37334 11736
rect 37292 11694 37320 11727
rect 37280 11688 37332 11694
rect 37280 11630 37332 11636
rect 37186 11384 37242 11393
rect 37096 11348 37148 11354
rect 37186 11319 37242 11328
rect 37096 11290 37148 11296
rect 37200 11218 37228 11319
rect 37188 11212 37240 11218
rect 37188 11154 37240 11160
rect 37280 10600 37332 10606
rect 37280 10542 37332 10548
rect 37292 10441 37320 10542
rect 37278 10432 37334 10441
rect 37278 10367 37334 10376
rect 37278 9616 37334 9625
rect 37278 9551 37334 9560
rect 37292 9518 37320 9551
rect 37280 9512 37332 9518
rect 37280 9454 37332 9460
rect 37384 9178 37412 16646
rect 37568 12434 37596 16934
rect 37476 12406 37596 12434
rect 37372 9172 37424 9178
rect 37372 9114 37424 9120
rect 37186 9072 37242 9081
rect 37186 9007 37188 9016
rect 37240 9007 37242 9016
rect 37188 8978 37240 8984
rect 37188 8424 37240 8430
rect 37188 8366 37240 8372
rect 37200 8265 37228 8366
rect 37186 8256 37242 8265
rect 37186 8191 37242 8200
rect 37280 7336 37332 7342
rect 37278 7304 37280 7313
rect 37332 7304 37334 7313
rect 37278 7239 37334 7248
rect 37186 6896 37242 6905
rect 37186 6831 37188 6840
rect 37240 6831 37242 6840
rect 37188 6802 37240 6808
rect 37476 6458 37504 12406
rect 37464 6452 37516 6458
rect 37464 6394 37516 6400
rect 37280 6248 37332 6254
rect 37280 6190 37332 6196
rect 37292 5953 37320 6190
rect 37278 5944 37334 5953
rect 37278 5879 37334 5888
rect 37188 5772 37240 5778
rect 37188 5714 37240 5720
rect 37200 5545 37228 5714
rect 37186 5536 37242 5545
rect 37186 5471 37242 5480
rect 37096 5160 37148 5166
rect 37096 5102 37148 5108
rect 37004 2304 37056 2310
rect 37004 2246 37056 2252
rect 36726 640 36782 649
rect 36726 575 36782 584
rect 36818 -800 36874 800
rect 37108 241 37136 5102
rect 37188 3120 37240 3126
rect 37188 3062 37240 3068
rect 37200 800 37228 3062
rect 37660 2582 37688 56646
rect 37752 31482 37780 61814
rect 37844 59537 37872 66438
rect 37936 63918 37964 68070
rect 38028 65006 38056 69158
rect 38120 66094 38148 69278
rect 38212 68354 38240 69362
rect 38304 68649 38332 70382
rect 38396 69494 38424 72422
rect 38384 69488 38436 69494
rect 38384 69430 38436 69436
rect 38384 69352 38436 69358
rect 38384 69294 38436 69300
rect 38290 68640 38346 68649
rect 38290 68575 38346 68584
rect 38212 68326 38332 68354
rect 38200 68264 38252 68270
rect 38200 68206 38252 68212
rect 38108 66088 38160 66094
rect 38108 66030 38160 66036
rect 38212 65929 38240 68206
rect 38198 65920 38254 65929
rect 38198 65855 38254 65864
rect 38016 65000 38068 65006
rect 38016 64942 38068 64948
rect 37924 63912 37976 63918
rect 38304 63866 38332 68326
rect 38396 67289 38424 69294
rect 38382 67280 38438 67289
rect 38382 67215 38438 67224
rect 38384 67176 38436 67182
rect 38384 67118 38436 67124
rect 37924 63854 37976 63860
rect 38028 63838 38332 63866
rect 38028 60734 38056 63838
rect 38108 63776 38160 63782
rect 38108 63718 38160 63724
rect 37936 60706 38056 60734
rect 37830 59528 37886 59537
rect 37830 59463 37886 59472
rect 37936 58954 37964 60706
rect 37924 58948 37976 58954
rect 37924 58890 37976 58896
rect 37832 58608 37884 58614
rect 37832 58550 37884 58556
rect 37740 31476 37792 31482
rect 37740 31418 37792 31424
rect 37844 28762 37872 58550
rect 37924 57384 37976 57390
rect 37924 57326 37976 57332
rect 37936 56953 37964 57326
rect 37922 56944 37978 56953
rect 37922 56879 37978 56888
rect 37922 56536 37978 56545
rect 37922 56471 37978 56480
rect 37936 56302 37964 56471
rect 37924 56296 37976 56302
rect 37924 56238 37976 56244
rect 37924 55208 37976 55214
rect 37922 55176 37924 55185
rect 37976 55176 37978 55185
rect 37922 55111 37978 55120
rect 37924 53032 37976 53038
rect 37924 52974 37976 52980
rect 37936 52601 37964 52974
rect 37922 52592 37978 52601
rect 37922 52527 37978 52536
rect 37924 51944 37976 51950
rect 37924 51886 37976 51892
rect 37936 51241 37964 51886
rect 37922 51232 37978 51241
rect 37922 51167 37978 51176
rect 37924 50856 37976 50862
rect 37924 50798 37976 50804
rect 37936 50289 37964 50798
rect 37922 50280 37978 50289
rect 37922 50215 37978 50224
rect 37922 49872 37978 49881
rect 37922 49807 37978 49816
rect 37936 49774 37964 49807
rect 37924 49768 37976 49774
rect 37924 49710 37976 49716
rect 37924 48680 37976 48686
rect 37924 48622 37976 48628
rect 37936 48521 37964 48622
rect 37922 48512 37978 48521
rect 37922 48447 37978 48456
rect 37924 47592 37976 47598
rect 37924 47534 37976 47540
rect 37936 47161 37964 47534
rect 37922 47152 37978 47161
rect 37922 47087 37978 47096
rect 37924 46504 37976 46510
rect 37924 46446 37976 46452
rect 37936 45801 37964 46446
rect 37922 45792 37978 45801
rect 37922 45727 37978 45736
rect 37924 45416 37976 45422
rect 37924 45358 37976 45364
rect 37936 44985 37964 45358
rect 37922 44976 37978 44985
rect 37922 44911 37978 44920
rect 37922 44432 37978 44441
rect 37922 44367 37978 44376
rect 37936 44334 37964 44367
rect 37924 44328 37976 44334
rect 37924 44270 37976 44276
rect 37924 43240 37976 43246
rect 37924 43182 37976 43188
rect 37936 43081 37964 43182
rect 37922 43072 37978 43081
rect 37922 43007 37978 43016
rect 37924 42152 37976 42158
rect 37924 42094 37976 42100
rect 37936 41857 37964 42094
rect 37922 41848 37978 41857
rect 37922 41783 37978 41792
rect 37924 41064 37976 41070
rect 37924 41006 37976 41012
rect 37936 40497 37964 41006
rect 37922 40488 37978 40497
rect 37922 40423 37978 40432
rect 38120 40050 38148 63718
rect 38396 63510 38424 67118
rect 38384 63504 38436 63510
rect 38384 63446 38436 63452
rect 38292 63232 38344 63238
rect 38292 63174 38344 63180
rect 38200 54052 38252 54058
rect 38200 53994 38252 54000
rect 38108 40044 38160 40050
rect 38108 39986 38160 39992
rect 37924 39976 37976 39982
rect 37924 39918 37976 39924
rect 37936 39545 37964 39918
rect 37922 39536 37978 39545
rect 37922 39471 37978 39480
rect 37922 39128 37978 39137
rect 37922 39063 37978 39072
rect 37936 38894 37964 39063
rect 37924 38888 37976 38894
rect 37924 38830 37976 38836
rect 37924 37800 37976 37806
rect 37922 37768 37924 37777
rect 37976 37768 37978 37777
rect 37922 37703 37978 37712
rect 37924 36712 37976 36718
rect 37924 36654 37976 36660
rect 37936 36417 37964 36654
rect 37922 36408 37978 36417
rect 37922 36343 37978 36352
rect 37924 35624 37976 35630
rect 37924 35566 37976 35572
rect 37936 35057 37964 35566
rect 37922 35048 37978 35057
rect 37922 34983 37978 34992
rect 37924 34536 37976 34542
rect 37924 34478 37976 34484
rect 37936 34241 37964 34478
rect 37922 34232 37978 34241
rect 37922 34167 37978 34176
rect 37922 33688 37978 33697
rect 37922 33623 37978 33632
rect 37936 33454 37964 33623
rect 37924 33448 37976 33454
rect 37924 33390 37976 33396
rect 37924 32360 37976 32366
rect 37922 32328 37924 32337
rect 37976 32328 37978 32337
rect 37922 32263 37978 32272
rect 37924 31272 37976 31278
rect 37924 31214 37976 31220
rect 37936 31113 37964 31214
rect 37922 31104 37978 31113
rect 37922 31039 37978 31048
rect 37924 30184 37976 30190
rect 37924 30126 37976 30132
rect 37936 29753 37964 30126
rect 37922 29744 37978 29753
rect 37922 29679 37978 29688
rect 37924 29096 37976 29102
rect 37924 29038 37976 29044
rect 37832 28756 37884 28762
rect 37832 28698 37884 28704
rect 37936 28393 37964 29038
rect 38014 28792 38070 28801
rect 38014 28727 38070 28736
rect 37922 28384 37978 28393
rect 37922 28319 37978 28328
rect 38028 28014 38056 28727
rect 38016 28008 38068 28014
rect 38016 27950 38068 27956
rect 37922 27024 37978 27033
rect 37922 26959 37978 26968
rect 37936 26926 37964 26959
rect 37924 26920 37976 26926
rect 37924 26862 37976 26868
rect 37832 26512 37884 26518
rect 37832 26454 37884 26460
rect 37738 25392 37794 25401
rect 37738 25327 37794 25336
rect 37752 18970 37780 25327
rect 37844 20058 37872 26454
rect 37924 25832 37976 25838
rect 37924 25774 37976 25780
rect 37936 25673 37964 25774
rect 37922 25664 37978 25673
rect 37922 25599 37978 25608
rect 38106 25528 38162 25537
rect 38106 25463 38162 25472
rect 37924 24744 37976 24750
rect 37924 24686 37976 24692
rect 37936 24313 37964 24686
rect 37922 24304 37978 24313
rect 37922 24239 37978 24248
rect 38016 24064 38068 24070
rect 38016 24006 38068 24012
rect 37924 23656 37976 23662
rect 37924 23598 37976 23604
rect 37936 22953 37964 23598
rect 37922 22944 37978 22953
rect 37922 22879 37978 22888
rect 37924 22568 37976 22574
rect 37924 22510 37976 22516
rect 37936 22137 37964 22510
rect 37922 22128 37978 22137
rect 37922 22063 37978 22072
rect 37922 21584 37978 21593
rect 37922 21519 37978 21528
rect 37936 21486 37964 21519
rect 37924 21480 37976 21486
rect 37924 21422 37976 21428
rect 37924 20392 37976 20398
rect 37922 20360 37924 20369
rect 37976 20360 37978 20369
rect 37922 20295 37978 20304
rect 37832 20052 37884 20058
rect 37832 19994 37884 20000
rect 37832 19848 37884 19854
rect 37832 19790 37884 19796
rect 37740 18964 37792 18970
rect 37740 18906 37792 18912
rect 37844 12850 37872 19790
rect 37924 19304 37976 19310
rect 37924 19246 37976 19252
rect 37936 19009 37964 19246
rect 37922 19000 37978 19009
rect 37922 18935 37978 18944
rect 37924 18216 37976 18222
rect 37924 18158 37976 18164
rect 37936 17649 37964 18158
rect 37922 17640 37978 17649
rect 37922 17575 37978 17584
rect 37924 17128 37976 17134
rect 37924 17070 37976 17076
rect 37936 16697 37964 17070
rect 37922 16688 37978 16697
rect 37922 16623 37978 16632
rect 37922 16280 37978 16289
rect 37922 16215 37978 16224
rect 37936 16046 37964 16215
rect 37924 16040 37976 16046
rect 37924 15982 37976 15988
rect 37924 14952 37976 14958
rect 37922 14920 37924 14929
rect 37976 14920 37978 14929
rect 37922 14855 37978 14864
rect 38028 14618 38056 24006
rect 38120 16250 38148 25463
rect 38108 16244 38160 16250
rect 38108 16186 38160 16192
rect 38016 14612 38068 14618
rect 38016 14554 38068 14560
rect 37924 13864 37976 13870
rect 37924 13806 37976 13812
rect 37936 13161 37964 13806
rect 37922 13152 37978 13161
rect 37922 13087 37978 13096
rect 37832 12844 37884 12850
rect 37832 12786 37884 12792
rect 37924 12776 37976 12782
rect 37924 12718 37976 12724
rect 37936 12209 37964 12718
rect 37922 12200 37978 12209
rect 37922 12135 37978 12144
rect 37924 10600 37976 10606
rect 37924 10542 37976 10548
rect 37936 10033 37964 10542
rect 37922 10024 37978 10033
rect 37922 9959 37978 9968
rect 37924 9512 37976 9518
rect 37924 9454 37976 9460
rect 37936 8673 37964 9454
rect 37922 8664 37978 8673
rect 37922 8599 37978 8608
rect 37924 8424 37976 8430
rect 37924 8366 37976 8372
rect 37936 7721 37964 8366
rect 37922 7712 37978 7721
rect 37922 7647 37978 7656
rect 37924 7336 37976 7342
rect 37924 7278 37976 7284
rect 37936 6497 37964 7278
rect 37922 6488 37978 6497
rect 37922 6423 37978 6432
rect 37832 3460 37884 3466
rect 37832 3402 37884 3408
rect 37648 2576 37700 2582
rect 37648 2518 37700 2524
rect 37464 2508 37516 2514
rect 37464 2450 37516 2456
rect 37476 800 37504 2450
rect 37844 800 37872 3402
rect 38212 3194 38240 53994
rect 38304 36854 38332 63174
rect 38384 59696 38436 59702
rect 38384 59638 38436 59644
rect 38292 36848 38344 36854
rect 38292 36790 38344 36796
rect 38396 28422 38424 59638
rect 38488 55894 38516 111658
rect 38580 96014 38608 117098
rect 38672 115802 38700 119200
rect 38660 115796 38712 115802
rect 38660 115738 38712 115744
rect 38948 113014 38976 119200
rect 39132 113082 39160 119200
rect 39408 113966 39436 119200
rect 39592 115734 39620 119200
rect 39580 115728 39632 115734
rect 39580 115670 39632 115676
rect 39868 115122 39896 119200
rect 39856 115116 39908 115122
rect 39856 115058 39908 115064
rect 39396 113960 39448 113966
rect 39396 113902 39448 113908
rect 39120 113076 39172 113082
rect 39120 113018 39172 113024
rect 38936 113008 38988 113014
rect 38936 112950 38988 112956
rect 39120 111648 39172 111654
rect 39120 111590 39172 111596
rect 38660 110016 38712 110022
rect 38660 109958 38712 109964
rect 38568 96008 38620 96014
rect 38568 95950 38620 95956
rect 38672 80054 38700 109958
rect 38844 109472 38896 109478
rect 38844 109414 38896 109420
rect 38752 101992 38804 101998
rect 38752 101934 38804 101940
rect 38764 80986 38792 101934
rect 38856 89714 38884 109414
rect 39132 89714 39160 111590
rect 38856 89686 38976 89714
rect 39132 89686 39252 89714
rect 38752 80980 38804 80986
rect 38752 80922 38804 80928
rect 38672 80026 38792 80054
rect 38568 79552 38620 79558
rect 38568 79494 38620 79500
rect 38580 70258 38608 79494
rect 38764 79370 38792 80026
rect 38764 79342 38884 79370
rect 38752 79280 38804 79286
rect 38752 79222 38804 79228
rect 38660 75744 38712 75750
rect 38660 75686 38712 75692
rect 38672 70378 38700 75686
rect 38660 70372 38712 70378
rect 38660 70314 38712 70320
rect 38580 70230 38700 70258
rect 38566 70136 38622 70145
rect 38566 70071 38622 70080
rect 38580 65482 38608 70071
rect 38568 65476 38620 65482
rect 38568 65418 38620 65424
rect 38672 64841 38700 70230
rect 38658 64832 38714 64841
rect 38658 64767 38714 64776
rect 38568 64320 38620 64326
rect 38568 64262 38620 64268
rect 38476 55888 38528 55894
rect 38476 55830 38528 55836
rect 38580 39438 38608 64262
rect 38764 63374 38792 79222
rect 38856 74458 38884 79342
rect 38948 75274 38976 89686
rect 39028 83360 39080 83366
rect 39028 83302 39080 83308
rect 38936 75268 38988 75274
rect 38936 75210 38988 75216
rect 38844 74452 38896 74458
rect 38844 74394 38896 74400
rect 38844 74112 38896 74118
rect 38844 74054 38896 74060
rect 38856 71618 38884 74054
rect 38936 71800 38988 71806
rect 38934 71768 38936 71777
rect 38988 71768 38990 71777
rect 38934 71703 38990 71712
rect 38856 71590 38976 71618
rect 38844 71528 38896 71534
rect 38844 71470 38896 71476
rect 38856 66842 38884 71470
rect 38844 66836 38896 66842
rect 38844 66778 38896 66784
rect 38844 65748 38896 65754
rect 38844 65690 38896 65696
rect 38856 63850 38884 65690
rect 38844 63844 38896 63850
rect 38844 63786 38896 63792
rect 38948 63730 38976 71590
rect 39040 66162 39068 83302
rect 39120 79008 39172 79014
rect 39120 78950 39172 78956
rect 39132 72468 39160 78950
rect 39224 75954 39252 89686
rect 39396 84448 39448 84454
rect 39396 84390 39448 84396
rect 39304 78192 39356 78198
rect 39304 78134 39356 78140
rect 39212 75948 39264 75954
rect 39212 75890 39264 75896
rect 39316 75070 39344 78134
rect 39408 75274 39436 84390
rect 39948 82272 40000 82278
rect 39948 82214 40000 82220
rect 39672 81728 39724 81734
rect 39672 81670 39724 81676
rect 39488 80096 39540 80102
rect 39488 80038 39540 80044
rect 39396 75268 39448 75274
rect 39396 75210 39448 75216
rect 39304 75064 39356 75070
rect 39304 75006 39356 75012
rect 39132 72440 39436 72468
rect 39304 70372 39356 70378
rect 39304 70314 39356 70320
rect 39120 70168 39172 70174
rect 39120 70110 39172 70116
rect 39028 66156 39080 66162
rect 39028 66098 39080 66104
rect 39028 65408 39080 65414
rect 39028 65350 39080 65356
rect 38856 63702 38976 63730
rect 38752 63368 38804 63374
rect 38752 63310 38804 63316
rect 38752 62960 38804 62966
rect 38752 62902 38804 62908
rect 38660 59968 38712 59974
rect 38660 59910 38712 59916
rect 38672 53174 38700 59910
rect 38660 53168 38712 53174
rect 38660 53110 38712 53116
rect 38764 51882 38792 62902
rect 38856 59430 38884 63702
rect 38936 63640 38988 63646
rect 38936 63582 38988 63588
rect 38844 59424 38896 59430
rect 38844 59366 38896 59372
rect 38948 54330 38976 63582
rect 38936 54324 38988 54330
rect 38936 54266 38988 54272
rect 38936 53168 38988 53174
rect 38936 53110 38988 53116
rect 38752 51876 38804 51882
rect 38752 51818 38804 51824
rect 38752 51604 38804 51610
rect 38752 51546 38804 51552
rect 38568 39432 38620 39438
rect 38568 39374 38620 39380
rect 38764 32298 38792 51546
rect 38752 32292 38804 32298
rect 38752 32234 38804 32240
rect 38476 28484 38528 28490
rect 38476 28426 38528 28432
rect 38384 28416 38436 28422
rect 38384 28358 38436 28364
rect 38384 25696 38436 25702
rect 38384 25638 38436 25644
rect 38292 24336 38344 24342
rect 38292 24278 38344 24284
rect 38304 12986 38332 24278
rect 38396 14006 38424 25638
rect 38488 21554 38516 28426
rect 38948 27946 38976 53110
rect 39040 41614 39068 65350
rect 39132 62218 39160 70110
rect 39212 69216 39264 69222
rect 39212 69158 39264 69164
rect 39224 67590 39252 69158
rect 39212 67584 39264 67590
rect 39212 67526 39264 67532
rect 39120 62212 39172 62218
rect 39120 62154 39172 62160
rect 39316 60042 39344 70314
rect 39408 65686 39436 72440
rect 39396 65680 39448 65686
rect 39396 65622 39448 65628
rect 39396 65136 39448 65142
rect 39396 65078 39448 65084
rect 39304 60036 39356 60042
rect 39304 59978 39356 59984
rect 39408 45082 39436 65078
rect 39500 63986 39528 80038
rect 39580 75268 39632 75274
rect 39580 75210 39632 75216
rect 39592 67318 39620 75210
rect 39684 75138 39712 81670
rect 39856 80368 39908 80374
rect 39856 80310 39908 80316
rect 39764 75812 39816 75818
rect 39764 75754 39816 75760
rect 39672 75132 39724 75138
rect 39672 75074 39724 75080
rect 39672 74996 39724 75002
rect 39672 74938 39724 74944
rect 39580 67312 39632 67318
rect 39580 67254 39632 67260
rect 39580 67176 39632 67182
rect 39580 67118 39632 67124
rect 39488 63980 39540 63986
rect 39488 63922 39540 63928
rect 39592 61062 39620 67118
rect 39684 65210 39712 74938
rect 39776 69698 39804 75754
rect 39764 69692 39816 69698
rect 39764 69634 39816 69640
rect 39764 69556 39816 69562
rect 39764 69498 39816 69504
rect 39672 65204 39724 65210
rect 39672 65146 39724 65152
rect 39776 63073 39804 69498
rect 39868 64122 39896 80310
rect 39960 65074 39988 82214
rect 39948 65068 40000 65074
rect 39948 65010 40000 65016
rect 39856 64116 39908 64122
rect 39856 64058 39908 64064
rect 39762 63064 39818 63073
rect 39762 62999 39818 63008
rect 39580 61056 39632 61062
rect 39580 60998 39632 61004
rect 39396 45076 39448 45082
rect 39396 45018 39448 45024
rect 39028 41608 39080 41614
rect 39028 41550 39080 41556
rect 38936 27940 38988 27946
rect 38936 27882 38988 27888
rect 38660 26376 38712 26382
rect 38660 26318 38712 26324
rect 38568 22024 38620 22030
rect 38568 21966 38620 21972
rect 38476 21548 38528 21554
rect 38476 21490 38528 21496
rect 38476 20936 38528 20942
rect 38476 20878 38528 20884
rect 38384 14000 38436 14006
rect 38384 13942 38436 13948
rect 38292 12980 38344 12986
rect 38292 12922 38344 12928
rect 38292 12844 38344 12850
rect 38292 12786 38344 12792
rect 38304 7546 38332 12786
rect 38488 9654 38516 20878
rect 38476 9648 38528 9654
rect 38476 9590 38528 9596
rect 38580 9382 38608 21966
rect 38672 17338 38700 26318
rect 38752 25424 38804 25430
rect 38752 25366 38804 25372
rect 38660 17332 38712 17338
rect 38660 17274 38712 17280
rect 38764 14074 38792 25366
rect 38752 14068 38804 14074
rect 38752 14010 38804 14016
rect 38936 11076 38988 11082
rect 38936 11018 38988 11024
rect 38948 10849 38976 11018
rect 38934 10840 38990 10849
rect 38934 10775 38990 10784
rect 38568 9376 38620 9382
rect 38568 9318 38620 9324
rect 38292 7540 38344 7546
rect 38292 7482 38344 7488
rect 38936 5568 38988 5574
rect 38936 5510 38988 5516
rect 38948 5137 38976 5510
rect 38934 5128 38990 5137
rect 38934 5063 38990 5072
rect 39396 5092 39448 5098
rect 39396 5034 39448 5040
rect 39120 4072 39172 4078
rect 39120 4014 39172 4020
rect 38476 4004 38528 4010
rect 38476 3946 38528 3952
rect 38200 3188 38252 3194
rect 38200 3130 38252 3136
rect 37922 3088 37978 3097
rect 37922 3023 37978 3032
rect 37936 2990 37964 3023
rect 37924 2984 37976 2990
rect 37924 2926 37976 2932
rect 38108 2916 38160 2922
rect 38108 2858 38160 2864
rect 38120 800 38148 2858
rect 38488 800 38516 3946
rect 38752 3936 38804 3942
rect 38752 3878 38804 3884
rect 38764 800 38792 3878
rect 39132 800 39160 4014
rect 39408 800 39436 5034
rect 39764 4548 39816 4554
rect 39764 4490 39816 4496
rect 39776 800 39804 4490
rect 37094 232 37150 241
rect 37094 167 37150 176
rect 37186 -800 37242 800
rect 37462 -800 37518 800
rect 37830 -800 37886 800
rect 38106 -800 38162 800
rect 38474 -800 38530 800
rect 38750 -800 38806 800
rect 39118 -800 39174 800
rect 39394 -800 39450 800
rect 39762 -800 39818 800
<< via2 >>
rect 3422 119448 3478 119504
rect 1398 117816 1454 117872
rect 2042 116204 2098 116240
rect 2042 116184 2044 116204
rect 2044 116184 2096 116204
rect 2096 116184 2098 116204
rect 1398 105868 1454 105904
rect 1398 105848 1400 105868
rect 1400 105848 1452 105868
rect 1452 105848 1454 105868
rect 1490 104216 1546 104272
rect 1398 101768 1454 101824
rect 1398 100952 1454 101008
rect 1398 100272 1454 100328
rect 1398 99456 1454 99512
rect 1398 98676 1400 98696
rect 1400 98676 1452 98696
rect 1452 98676 1454 98696
rect 1398 98640 1454 98676
rect 1398 97824 1454 97880
rect 1398 97008 1454 97064
rect 1398 96192 1454 96248
rect 1398 95412 1400 95432
rect 1400 95412 1452 95432
rect 1452 95412 1454 95432
rect 1398 95376 1454 95412
rect 1398 94560 1454 94616
rect 1398 93744 1454 93800
rect 1398 93064 1454 93120
rect 1398 92248 1454 92304
rect 1398 91432 1454 91488
rect 1398 89800 1454 89856
rect 1398 88984 1454 89040
rect 1398 88168 1454 88224
rect 1398 87372 1454 87408
rect 1398 87352 1400 87372
rect 1400 87352 1452 87372
rect 1452 87352 1454 87372
rect 1398 86708 1400 86728
rect 1400 86708 1452 86728
rect 1452 86708 1454 86728
rect 1398 86672 1454 86708
rect 1398 85856 1454 85912
rect 1398 85040 1454 85096
rect 1398 84224 1454 84280
rect 1398 83444 1400 83464
rect 1400 83444 1452 83464
rect 1452 83444 1454 83464
rect 1398 83408 1454 83444
rect 1398 82592 1454 82648
rect 1398 81776 1454 81832
rect 1398 80960 1454 81016
rect 1398 80280 1454 80336
rect 1398 79464 1454 79520
rect 1398 78668 1454 78704
rect 1398 78648 1400 78668
rect 1400 78648 1452 78668
rect 1452 78648 1454 78668
rect 1398 77832 1454 77888
rect 1398 77016 1454 77072
rect 1398 76200 1454 76256
rect 1398 75404 1454 75440
rect 1398 75384 1400 75404
rect 1400 75384 1452 75404
rect 1452 75384 1454 75404
rect 1398 74568 1454 74624
rect 1398 73752 1454 73808
rect 1398 73072 1454 73128
rect 1398 72256 1454 72312
rect 1398 71476 1400 71496
rect 1400 71476 1452 71496
rect 1452 71476 1454 71496
rect 1398 71440 1454 71476
rect 1398 70624 1454 70680
rect 1398 69808 1454 69864
rect 1398 68992 1454 69048
rect 1398 68212 1400 68232
rect 1400 68212 1452 68232
rect 1452 68212 1454 68232
rect 1398 68176 1454 68212
rect 1398 67360 1454 67416
rect 1398 66700 1454 66736
rect 1398 66680 1400 66700
rect 1400 66680 1452 66700
rect 1452 66680 1454 66700
rect 1398 65864 1454 65920
rect 1398 65048 1454 65104
rect 1398 64232 1454 64288
rect 1398 63436 1454 63472
rect 1398 63416 1400 63436
rect 1400 63416 1452 63436
rect 1452 63416 1454 63436
rect 1398 62600 1454 62656
rect 1398 61784 1454 61840
rect 1398 60968 1454 61024
rect 1398 60288 1454 60344
rect 1398 59508 1400 59528
rect 1400 59508 1452 59528
rect 1452 59508 1454 59528
rect 1398 59472 1454 59508
rect 1398 58656 1454 58712
rect 1398 57840 1454 57896
rect 1398 57024 1454 57080
rect 1398 56244 1400 56264
rect 1400 56244 1452 56264
rect 1452 56244 1454 56264
rect 1398 56208 1454 56244
rect 1398 55392 1454 55448
rect 1398 54576 1454 54632
rect 1398 53760 1454 53816
rect 1398 53080 1454 53136
rect 1398 52264 1454 52320
rect 1398 51468 1454 51504
rect 1398 51448 1400 51468
rect 1400 51448 1452 51468
rect 1452 51448 1454 51468
rect 1950 115404 1952 115424
rect 1952 115404 2004 115424
rect 2004 115404 2006 115424
rect 1950 115368 2006 115404
rect 2042 114552 2098 114608
rect 1858 113736 1914 113792
rect 2870 118632 2926 118688
rect 2778 117000 2834 117056
rect 1950 113076 2006 113112
rect 1950 113056 1952 113076
rect 1952 113056 2004 113076
rect 2004 113056 2006 113076
rect 2042 112276 2044 112296
rect 2044 112276 2096 112296
rect 2096 112276 2098 112296
rect 2042 112240 2098 112276
rect 1950 111444 2006 111480
rect 1950 111424 1952 111444
rect 1952 111424 2004 111444
rect 2004 111424 2006 111444
rect 2042 110628 2098 110664
rect 2042 110608 2044 110628
rect 2044 110608 2096 110628
rect 2096 110608 2098 110628
rect 1950 109812 2006 109848
rect 1950 109792 1952 109812
rect 1952 109792 2004 109812
rect 2004 109792 2006 109812
rect 1858 108976 1914 109032
rect 1950 108180 2006 108216
rect 1950 108160 1952 108180
rect 1952 108160 2004 108180
rect 2004 108160 2006 108180
rect 2042 107364 2098 107400
rect 2042 107344 2044 107364
rect 2044 107344 2096 107364
rect 2096 107344 2098 107364
rect 1950 106700 1952 106720
rect 1952 106700 2004 106720
rect 2004 106700 2006 106720
rect 1950 106664 2006 106700
rect 1950 105068 1952 105088
rect 1952 105068 2004 105088
rect 2004 105068 2006 105088
rect 1950 105032 2006 105068
rect 2042 103400 2098 103456
rect 2042 102604 2098 102640
rect 2042 102584 2044 102604
rect 2044 102584 2096 102604
rect 2096 102584 2098 102604
rect 2042 90636 2098 90672
rect 2042 90616 2044 90636
rect 2044 90616 2096 90636
rect 2096 90616 2098 90636
rect 36082 119584 36138 119640
rect 1858 50632 1914 50688
rect 1858 49816 1914 49872
rect 1858 49000 1914 49056
rect 1858 48204 1914 48240
rect 1858 48184 1860 48204
rect 1860 48184 1912 48204
rect 1912 48184 1914 48204
rect 1858 47368 1914 47424
rect 1858 46688 1914 46744
rect 1858 45872 1914 45928
rect 1858 45056 1914 45112
rect 1858 44260 1914 44296
rect 1858 44240 1860 44260
rect 1860 44240 1912 44260
rect 1912 44240 1914 44260
rect 1858 43424 1914 43480
rect 1858 42608 1914 42664
rect 1858 41792 1914 41848
rect 1858 40996 1914 41032
rect 1858 40976 1860 40996
rect 1860 40976 1912 40996
rect 1912 40976 1914 40996
rect 1858 40296 1914 40352
rect 1858 39500 1914 39536
rect 1858 39480 1860 39500
rect 1860 39480 1912 39500
rect 1912 39480 1914 39500
rect 1858 38664 1914 38720
rect 1858 37848 1914 37904
rect 1858 37032 1914 37088
rect 1858 36236 1914 36272
rect 1858 36216 1860 36236
rect 1860 36216 1912 36236
rect 1912 36216 1914 36236
rect 1858 35400 1914 35456
rect 1858 34584 1914 34640
rect 1858 33768 1914 33824
rect 1858 33088 1914 33144
rect 1858 32292 1914 32328
rect 1858 32272 1860 32292
rect 1860 32272 1912 32292
rect 1912 32272 1914 32292
rect 1858 31456 1914 31512
rect 1858 30640 1914 30696
rect 1858 29824 1914 29880
rect 1858 29044 1860 29064
rect 1860 29044 1912 29064
rect 1912 29044 1914 29064
rect 1858 29008 1914 29044
rect 1858 28192 1914 28248
rect 1858 27376 1914 27432
rect 1858 26696 1914 26752
rect 1858 25880 1914 25936
rect 1858 25064 1914 25120
rect 1858 24268 1914 24304
rect 1858 24248 1860 24268
rect 1860 24248 1912 24268
rect 1912 24248 1914 24268
rect 1858 23432 1914 23488
rect 1858 22616 1914 22672
rect 1858 21800 1914 21856
rect 1858 21004 1914 21040
rect 1858 20984 1860 21004
rect 1860 20984 1912 21004
rect 1912 20984 1914 21004
rect 1858 20324 1914 20360
rect 1858 20304 1860 20324
rect 1860 20304 1912 20324
rect 1912 20304 1914 20324
rect 1858 19488 1914 19544
rect 1858 18672 1914 18728
rect 1858 17856 1914 17912
rect 1858 17060 1914 17096
rect 1858 17040 1860 17060
rect 1860 17040 1912 17060
rect 1912 17040 1914 17060
rect 1398 2624 1454 2680
rect 1858 16224 1914 16280
rect 1858 15408 1914 15464
rect 1858 14592 1914 14648
rect 1858 13812 1860 13832
rect 1860 13812 1912 13832
rect 1912 13812 1914 13832
rect 1858 13776 1914 13812
rect 1858 13096 1914 13152
rect 1858 12300 1914 12336
rect 1858 12280 1860 12300
rect 1860 12280 1912 12300
rect 1912 12280 1914 12300
rect 1858 11464 1914 11520
rect 1858 10648 1914 10704
rect 1858 9832 1914 9888
rect 1858 9036 1914 9072
rect 1858 9016 1860 9036
rect 1860 9016 1912 9036
rect 1912 9016 1914 9036
rect 1858 8200 1914 8256
rect 1858 7384 1914 7440
rect 1858 6704 1914 6760
rect 1858 5888 1914 5944
rect 1858 5092 1914 5128
rect 1858 5072 1860 5092
rect 1860 5072 1912 5092
rect 1912 5072 1914 5092
rect 1858 4256 1914 4312
rect 1858 3440 1914 3496
rect 1858 992 1914 1048
rect 4220 117530 4276 117532
rect 4300 117530 4356 117532
rect 4380 117530 4436 117532
rect 4460 117530 4516 117532
rect 4220 117478 4246 117530
rect 4246 117478 4276 117530
rect 4300 117478 4310 117530
rect 4310 117478 4356 117530
rect 4380 117478 4426 117530
rect 4426 117478 4436 117530
rect 4460 117478 4490 117530
rect 4490 117478 4516 117530
rect 4220 117476 4276 117478
rect 4300 117476 4356 117478
rect 4380 117476 4436 117478
rect 4460 117476 4516 117478
rect 4220 116442 4276 116444
rect 4300 116442 4356 116444
rect 4380 116442 4436 116444
rect 4460 116442 4516 116444
rect 4220 116390 4246 116442
rect 4246 116390 4276 116442
rect 4300 116390 4310 116442
rect 4310 116390 4356 116442
rect 4380 116390 4426 116442
rect 4426 116390 4436 116442
rect 4460 116390 4490 116442
rect 4490 116390 4516 116442
rect 4220 116388 4276 116390
rect 4300 116388 4356 116390
rect 4380 116388 4436 116390
rect 4460 116388 4516 116390
rect 4220 115354 4276 115356
rect 4300 115354 4356 115356
rect 4380 115354 4436 115356
rect 4460 115354 4516 115356
rect 4220 115302 4246 115354
rect 4246 115302 4276 115354
rect 4300 115302 4310 115354
rect 4310 115302 4356 115354
rect 4380 115302 4426 115354
rect 4426 115302 4436 115354
rect 4460 115302 4490 115354
rect 4490 115302 4516 115354
rect 4220 115300 4276 115302
rect 4300 115300 4356 115302
rect 4380 115300 4436 115302
rect 4460 115300 4516 115302
rect 4220 114266 4276 114268
rect 4300 114266 4356 114268
rect 4380 114266 4436 114268
rect 4460 114266 4516 114268
rect 4220 114214 4246 114266
rect 4246 114214 4276 114266
rect 4300 114214 4310 114266
rect 4310 114214 4356 114266
rect 4380 114214 4426 114266
rect 4426 114214 4436 114266
rect 4460 114214 4490 114266
rect 4490 114214 4516 114266
rect 4220 114212 4276 114214
rect 4300 114212 4356 114214
rect 4380 114212 4436 114214
rect 4460 114212 4516 114214
rect 4220 113178 4276 113180
rect 4300 113178 4356 113180
rect 4380 113178 4436 113180
rect 4460 113178 4516 113180
rect 4220 113126 4246 113178
rect 4246 113126 4276 113178
rect 4300 113126 4310 113178
rect 4310 113126 4356 113178
rect 4380 113126 4426 113178
rect 4426 113126 4436 113178
rect 4460 113126 4490 113178
rect 4490 113126 4516 113178
rect 4220 113124 4276 113126
rect 4300 113124 4356 113126
rect 4380 113124 4436 113126
rect 4460 113124 4516 113126
rect 4220 112090 4276 112092
rect 4300 112090 4356 112092
rect 4380 112090 4436 112092
rect 4460 112090 4516 112092
rect 4220 112038 4246 112090
rect 4246 112038 4276 112090
rect 4300 112038 4310 112090
rect 4310 112038 4356 112090
rect 4380 112038 4426 112090
rect 4426 112038 4436 112090
rect 4460 112038 4490 112090
rect 4490 112038 4516 112090
rect 4220 112036 4276 112038
rect 4300 112036 4356 112038
rect 4380 112036 4436 112038
rect 4460 112036 4516 112038
rect 4220 111002 4276 111004
rect 4300 111002 4356 111004
rect 4380 111002 4436 111004
rect 4460 111002 4516 111004
rect 4220 110950 4246 111002
rect 4246 110950 4276 111002
rect 4300 110950 4310 111002
rect 4310 110950 4356 111002
rect 4380 110950 4426 111002
rect 4426 110950 4436 111002
rect 4460 110950 4490 111002
rect 4490 110950 4516 111002
rect 4220 110948 4276 110950
rect 4300 110948 4356 110950
rect 4380 110948 4436 110950
rect 4460 110948 4516 110950
rect 4220 109914 4276 109916
rect 4300 109914 4356 109916
rect 4380 109914 4436 109916
rect 4460 109914 4516 109916
rect 4220 109862 4246 109914
rect 4246 109862 4276 109914
rect 4300 109862 4310 109914
rect 4310 109862 4356 109914
rect 4380 109862 4426 109914
rect 4426 109862 4436 109914
rect 4460 109862 4490 109914
rect 4490 109862 4516 109914
rect 4220 109860 4276 109862
rect 4300 109860 4356 109862
rect 4380 109860 4436 109862
rect 4460 109860 4516 109862
rect 4220 108826 4276 108828
rect 4300 108826 4356 108828
rect 4380 108826 4436 108828
rect 4460 108826 4516 108828
rect 4220 108774 4246 108826
rect 4246 108774 4276 108826
rect 4300 108774 4310 108826
rect 4310 108774 4356 108826
rect 4380 108774 4426 108826
rect 4426 108774 4436 108826
rect 4460 108774 4490 108826
rect 4490 108774 4516 108826
rect 4220 108772 4276 108774
rect 4300 108772 4356 108774
rect 4380 108772 4436 108774
rect 4460 108772 4516 108774
rect 4220 107738 4276 107740
rect 4300 107738 4356 107740
rect 4380 107738 4436 107740
rect 4460 107738 4516 107740
rect 4220 107686 4246 107738
rect 4246 107686 4276 107738
rect 4300 107686 4310 107738
rect 4310 107686 4356 107738
rect 4380 107686 4426 107738
rect 4426 107686 4436 107738
rect 4460 107686 4490 107738
rect 4490 107686 4516 107738
rect 4220 107684 4276 107686
rect 4300 107684 4356 107686
rect 4380 107684 4436 107686
rect 4460 107684 4516 107686
rect 4220 106650 4276 106652
rect 4300 106650 4356 106652
rect 4380 106650 4436 106652
rect 4460 106650 4516 106652
rect 4220 106598 4246 106650
rect 4246 106598 4276 106650
rect 4300 106598 4310 106650
rect 4310 106598 4356 106650
rect 4380 106598 4426 106650
rect 4426 106598 4436 106650
rect 4460 106598 4490 106650
rect 4490 106598 4516 106650
rect 4220 106596 4276 106598
rect 4300 106596 4356 106598
rect 4380 106596 4436 106598
rect 4460 106596 4516 106598
rect 4220 105562 4276 105564
rect 4300 105562 4356 105564
rect 4380 105562 4436 105564
rect 4460 105562 4516 105564
rect 4220 105510 4246 105562
rect 4246 105510 4276 105562
rect 4300 105510 4310 105562
rect 4310 105510 4356 105562
rect 4380 105510 4426 105562
rect 4426 105510 4436 105562
rect 4460 105510 4490 105562
rect 4490 105510 4516 105562
rect 4220 105508 4276 105510
rect 4300 105508 4356 105510
rect 4380 105508 4436 105510
rect 4460 105508 4516 105510
rect 4220 104474 4276 104476
rect 4300 104474 4356 104476
rect 4380 104474 4436 104476
rect 4460 104474 4516 104476
rect 4220 104422 4246 104474
rect 4246 104422 4276 104474
rect 4300 104422 4310 104474
rect 4310 104422 4356 104474
rect 4380 104422 4426 104474
rect 4426 104422 4436 104474
rect 4460 104422 4490 104474
rect 4490 104422 4516 104474
rect 4220 104420 4276 104422
rect 4300 104420 4356 104422
rect 4380 104420 4436 104422
rect 4460 104420 4516 104422
rect 4220 103386 4276 103388
rect 4300 103386 4356 103388
rect 4380 103386 4436 103388
rect 4460 103386 4516 103388
rect 4220 103334 4246 103386
rect 4246 103334 4276 103386
rect 4300 103334 4310 103386
rect 4310 103334 4356 103386
rect 4380 103334 4426 103386
rect 4426 103334 4436 103386
rect 4460 103334 4490 103386
rect 4490 103334 4516 103386
rect 4220 103332 4276 103334
rect 4300 103332 4356 103334
rect 4380 103332 4436 103334
rect 4460 103332 4516 103334
rect 4220 102298 4276 102300
rect 4300 102298 4356 102300
rect 4380 102298 4436 102300
rect 4460 102298 4516 102300
rect 4220 102246 4246 102298
rect 4246 102246 4276 102298
rect 4300 102246 4310 102298
rect 4310 102246 4356 102298
rect 4380 102246 4426 102298
rect 4426 102246 4436 102298
rect 4460 102246 4490 102298
rect 4490 102246 4516 102298
rect 4220 102244 4276 102246
rect 4300 102244 4356 102246
rect 4380 102244 4436 102246
rect 4460 102244 4516 102246
rect 4220 101210 4276 101212
rect 4300 101210 4356 101212
rect 4380 101210 4436 101212
rect 4460 101210 4516 101212
rect 4220 101158 4246 101210
rect 4246 101158 4276 101210
rect 4300 101158 4310 101210
rect 4310 101158 4356 101210
rect 4380 101158 4426 101210
rect 4426 101158 4436 101210
rect 4460 101158 4490 101210
rect 4490 101158 4516 101210
rect 4220 101156 4276 101158
rect 4300 101156 4356 101158
rect 4380 101156 4436 101158
rect 4460 101156 4516 101158
rect 4220 100122 4276 100124
rect 4300 100122 4356 100124
rect 4380 100122 4436 100124
rect 4460 100122 4516 100124
rect 4220 100070 4246 100122
rect 4246 100070 4276 100122
rect 4300 100070 4310 100122
rect 4310 100070 4356 100122
rect 4380 100070 4426 100122
rect 4426 100070 4436 100122
rect 4460 100070 4490 100122
rect 4490 100070 4516 100122
rect 4220 100068 4276 100070
rect 4300 100068 4356 100070
rect 4380 100068 4436 100070
rect 4460 100068 4516 100070
rect 4220 99034 4276 99036
rect 4300 99034 4356 99036
rect 4380 99034 4436 99036
rect 4460 99034 4516 99036
rect 4220 98982 4246 99034
rect 4246 98982 4276 99034
rect 4300 98982 4310 99034
rect 4310 98982 4356 99034
rect 4380 98982 4426 99034
rect 4426 98982 4436 99034
rect 4460 98982 4490 99034
rect 4490 98982 4516 99034
rect 4220 98980 4276 98982
rect 4300 98980 4356 98982
rect 4380 98980 4436 98982
rect 4460 98980 4516 98982
rect 4220 97946 4276 97948
rect 4300 97946 4356 97948
rect 4380 97946 4436 97948
rect 4460 97946 4516 97948
rect 4220 97894 4246 97946
rect 4246 97894 4276 97946
rect 4300 97894 4310 97946
rect 4310 97894 4356 97946
rect 4380 97894 4426 97946
rect 4426 97894 4436 97946
rect 4460 97894 4490 97946
rect 4490 97894 4516 97946
rect 4220 97892 4276 97894
rect 4300 97892 4356 97894
rect 4380 97892 4436 97894
rect 4460 97892 4516 97894
rect 4220 96858 4276 96860
rect 4300 96858 4356 96860
rect 4380 96858 4436 96860
rect 4460 96858 4516 96860
rect 4220 96806 4246 96858
rect 4246 96806 4276 96858
rect 4300 96806 4310 96858
rect 4310 96806 4356 96858
rect 4380 96806 4426 96858
rect 4426 96806 4436 96858
rect 4460 96806 4490 96858
rect 4490 96806 4516 96858
rect 4220 96804 4276 96806
rect 4300 96804 4356 96806
rect 4380 96804 4436 96806
rect 4460 96804 4516 96806
rect 4220 95770 4276 95772
rect 4300 95770 4356 95772
rect 4380 95770 4436 95772
rect 4460 95770 4516 95772
rect 4220 95718 4246 95770
rect 4246 95718 4276 95770
rect 4300 95718 4310 95770
rect 4310 95718 4356 95770
rect 4380 95718 4426 95770
rect 4426 95718 4436 95770
rect 4460 95718 4490 95770
rect 4490 95718 4516 95770
rect 4220 95716 4276 95718
rect 4300 95716 4356 95718
rect 4380 95716 4436 95718
rect 4460 95716 4516 95718
rect 4220 94682 4276 94684
rect 4300 94682 4356 94684
rect 4380 94682 4436 94684
rect 4460 94682 4516 94684
rect 4220 94630 4246 94682
rect 4246 94630 4276 94682
rect 4300 94630 4310 94682
rect 4310 94630 4356 94682
rect 4380 94630 4426 94682
rect 4426 94630 4436 94682
rect 4460 94630 4490 94682
rect 4490 94630 4516 94682
rect 4220 94628 4276 94630
rect 4300 94628 4356 94630
rect 4380 94628 4436 94630
rect 4460 94628 4516 94630
rect 4220 93594 4276 93596
rect 4300 93594 4356 93596
rect 4380 93594 4436 93596
rect 4460 93594 4516 93596
rect 4220 93542 4246 93594
rect 4246 93542 4276 93594
rect 4300 93542 4310 93594
rect 4310 93542 4356 93594
rect 4380 93542 4426 93594
rect 4426 93542 4436 93594
rect 4460 93542 4490 93594
rect 4490 93542 4516 93594
rect 4220 93540 4276 93542
rect 4300 93540 4356 93542
rect 4380 93540 4436 93542
rect 4460 93540 4516 93542
rect 4220 92506 4276 92508
rect 4300 92506 4356 92508
rect 4380 92506 4436 92508
rect 4460 92506 4516 92508
rect 4220 92454 4246 92506
rect 4246 92454 4276 92506
rect 4300 92454 4310 92506
rect 4310 92454 4356 92506
rect 4380 92454 4426 92506
rect 4426 92454 4436 92506
rect 4460 92454 4490 92506
rect 4490 92454 4516 92506
rect 4220 92452 4276 92454
rect 4300 92452 4356 92454
rect 4380 92452 4436 92454
rect 4460 92452 4516 92454
rect 4220 91418 4276 91420
rect 4300 91418 4356 91420
rect 4380 91418 4436 91420
rect 4460 91418 4516 91420
rect 4220 91366 4246 91418
rect 4246 91366 4276 91418
rect 4300 91366 4310 91418
rect 4310 91366 4356 91418
rect 4380 91366 4426 91418
rect 4426 91366 4436 91418
rect 4460 91366 4490 91418
rect 4490 91366 4516 91418
rect 4220 91364 4276 91366
rect 4300 91364 4356 91366
rect 4380 91364 4436 91366
rect 4460 91364 4516 91366
rect 4220 90330 4276 90332
rect 4300 90330 4356 90332
rect 4380 90330 4436 90332
rect 4460 90330 4516 90332
rect 4220 90278 4246 90330
rect 4246 90278 4276 90330
rect 4300 90278 4310 90330
rect 4310 90278 4356 90330
rect 4380 90278 4426 90330
rect 4426 90278 4436 90330
rect 4460 90278 4490 90330
rect 4490 90278 4516 90330
rect 4220 90276 4276 90278
rect 4300 90276 4356 90278
rect 4380 90276 4436 90278
rect 4460 90276 4516 90278
rect 4220 89242 4276 89244
rect 4300 89242 4356 89244
rect 4380 89242 4436 89244
rect 4460 89242 4516 89244
rect 4220 89190 4246 89242
rect 4246 89190 4276 89242
rect 4300 89190 4310 89242
rect 4310 89190 4356 89242
rect 4380 89190 4426 89242
rect 4426 89190 4436 89242
rect 4460 89190 4490 89242
rect 4490 89190 4516 89242
rect 4220 89188 4276 89190
rect 4300 89188 4356 89190
rect 4380 89188 4436 89190
rect 4460 89188 4516 89190
rect 4220 88154 4276 88156
rect 4300 88154 4356 88156
rect 4380 88154 4436 88156
rect 4460 88154 4516 88156
rect 4220 88102 4246 88154
rect 4246 88102 4276 88154
rect 4300 88102 4310 88154
rect 4310 88102 4356 88154
rect 4380 88102 4426 88154
rect 4426 88102 4436 88154
rect 4460 88102 4490 88154
rect 4490 88102 4516 88154
rect 4220 88100 4276 88102
rect 4300 88100 4356 88102
rect 4380 88100 4436 88102
rect 4460 88100 4516 88102
rect 4220 87066 4276 87068
rect 4300 87066 4356 87068
rect 4380 87066 4436 87068
rect 4460 87066 4516 87068
rect 4220 87014 4246 87066
rect 4246 87014 4276 87066
rect 4300 87014 4310 87066
rect 4310 87014 4356 87066
rect 4380 87014 4426 87066
rect 4426 87014 4436 87066
rect 4460 87014 4490 87066
rect 4490 87014 4516 87066
rect 4220 87012 4276 87014
rect 4300 87012 4356 87014
rect 4380 87012 4436 87014
rect 4460 87012 4516 87014
rect 4220 85978 4276 85980
rect 4300 85978 4356 85980
rect 4380 85978 4436 85980
rect 4460 85978 4516 85980
rect 4220 85926 4246 85978
rect 4246 85926 4276 85978
rect 4300 85926 4310 85978
rect 4310 85926 4356 85978
rect 4380 85926 4426 85978
rect 4426 85926 4436 85978
rect 4460 85926 4490 85978
rect 4490 85926 4516 85978
rect 4220 85924 4276 85926
rect 4300 85924 4356 85926
rect 4380 85924 4436 85926
rect 4460 85924 4516 85926
rect 4220 84890 4276 84892
rect 4300 84890 4356 84892
rect 4380 84890 4436 84892
rect 4460 84890 4516 84892
rect 4220 84838 4246 84890
rect 4246 84838 4276 84890
rect 4300 84838 4310 84890
rect 4310 84838 4356 84890
rect 4380 84838 4426 84890
rect 4426 84838 4436 84890
rect 4460 84838 4490 84890
rect 4490 84838 4516 84890
rect 4220 84836 4276 84838
rect 4300 84836 4356 84838
rect 4380 84836 4436 84838
rect 4460 84836 4516 84838
rect 4220 83802 4276 83804
rect 4300 83802 4356 83804
rect 4380 83802 4436 83804
rect 4460 83802 4516 83804
rect 4220 83750 4246 83802
rect 4246 83750 4276 83802
rect 4300 83750 4310 83802
rect 4310 83750 4356 83802
rect 4380 83750 4426 83802
rect 4426 83750 4436 83802
rect 4460 83750 4490 83802
rect 4490 83750 4516 83802
rect 4220 83748 4276 83750
rect 4300 83748 4356 83750
rect 4380 83748 4436 83750
rect 4460 83748 4516 83750
rect 4220 82714 4276 82716
rect 4300 82714 4356 82716
rect 4380 82714 4436 82716
rect 4460 82714 4516 82716
rect 4220 82662 4246 82714
rect 4246 82662 4276 82714
rect 4300 82662 4310 82714
rect 4310 82662 4356 82714
rect 4380 82662 4426 82714
rect 4426 82662 4436 82714
rect 4460 82662 4490 82714
rect 4490 82662 4516 82714
rect 4220 82660 4276 82662
rect 4300 82660 4356 82662
rect 4380 82660 4436 82662
rect 4460 82660 4516 82662
rect 4220 81626 4276 81628
rect 4300 81626 4356 81628
rect 4380 81626 4436 81628
rect 4460 81626 4516 81628
rect 4220 81574 4246 81626
rect 4246 81574 4276 81626
rect 4300 81574 4310 81626
rect 4310 81574 4356 81626
rect 4380 81574 4426 81626
rect 4426 81574 4436 81626
rect 4460 81574 4490 81626
rect 4490 81574 4516 81626
rect 4220 81572 4276 81574
rect 4300 81572 4356 81574
rect 4380 81572 4436 81574
rect 4460 81572 4516 81574
rect 4220 80538 4276 80540
rect 4300 80538 4356 80540
rect 4380 80538 4436 80540
rect 4460 80538 4516 80540
rect 4220 80486 4246 80538
rect 4246 80486 4276 80538
rect 4300 80486 4310 80538
rect 4310 80486 4356 80538
rect 4380 80486 4426 80538
rect 4426 80486 4436 80538
rect 4460 80486 4490 80538
rect 4490 80486 4516 80538
rect 4220 80484 4276 80486
rect 4300 80484 4356 80486
rect 4380 80484 4436 80486
rect 4460 80484 4516 80486
rect 4220 79450 4276 79452
rect 4300 79450 4356 79452
rect 4380 79450 4436 79452
rect 4460 79450 4516 79452
rect 4220 79398 4246 79450
rect 4246 79398 4276 79450
rect 4300 79398 4310 79450
rect 4310 79398 4356 79450
rect 4380 79398 4426 79450
rect 4426 79398 4436 79450
rect 4460 79398 4490 79450
rect 4490 79398 4516 79450
rect 4220 79396 4276 79398
rect 4300 79396 4356 79398
rect 4380 79396 4436 79398
rect 4460 79396 4516 79398
rect 4220 78362 4276 78364
rect 4300 78362 4356 78364
rect 4380 78362 4436 78364
rect 4460 78362 4516 78364
rect 4220 78310 4246 78362
rect 4246 78310 4276 78362
rect 4300 78310 4310 78362
rect 4310 78310 4356 78362
rect 4380 78310 4426 78362
rect 4426 78310 4436 78362
rect 4460 78310 4490 78362
rect 4490 78310 4516 78362
rect 4220 78308 4276 78310
rect 4300 78308 4356 78310
rect 4380 78308 4436 78310
rect 4460 78308 4516 78310
rect 4220 77274 4276 77276
rect 4300 77274 4356 77276
rect 4380 77274 4436 77276
rect 4460 77274 4516 77276
rect 4220 77222 4246 77274
rect 4246 77222 4276 77274
rect 4300 77222 4310 77274
rect 4310 77222 4356 77274
rect 4380 77222 4426 77274
rect 4426 77222 4436 77274
rect 4460 77222 4490 77274
rect 4490 77222 4516 77274
rect 4220 77220 4276 77222
rect 4300 77220 4356 77222
rect 4380 77220 4436 77222
rect 4460 77220 4516 77222
rect 4220 76186 4276 76188
rect 4300 76186 4356 76188
rect 4380 76186 4436 76188
rect 4460 76186 4516 76188
rect 4220 76134 4246 76186
rect 4246 76134 4276 76186
rect 4300 76134 4310 76186
rect 4310 76134 4356 76186
rect 4380 76134 4426 76186
rect 4426 76134 4436 76186
rect 4460 76134 4490 76186
rect 4490 76134 4516 76186
rect 4220 76132 4276 76134
rect 4300 76132 4356 76134
rect 4380 76132 4436 76134
rect 4460 76132 4516 76134
rect 4220 75098 4276 75100
rect 4300 75098 4356 75100
rect 4380 75098 4436 75100
rect 4460 75098 4516 75100
rect 4220 75046 4246 75098
rect 4246 75046 4276 75098
rect 4300 75046 4310 75098
rect 4310 75046 4356 75098
rect 4380 75046 4426 75098
rect 4426 75046 4436 75098
rect 4460 75046 4490 75098
rect 4490 75046 4516 75098
rect 4220 75044 4276 75046
rect 4300 75044 4356 75046
rect 4380 75044 4436 75046
rect 4460 75044 4516 75046
rect 4220 74010 4276 74012
rect 4300 74010 4356 74012
rect 4380 74010 4436 74012
rect 4460 74010 4516 74012
rect 4220 73958 4246 74010
rect 4246 73958 4276 74010
rect 4300 73958 4310 74010
rect 4310 73958 4356 74010
rect 4380 73958 4426 74010
rect 4426 73958 4436 74010
rect 4460 73958 4490 74010
rect 4490 73958 4516 74010
rect 4220 73956 4276 73958
rect 4300 73956 4356 73958
rect 4380 73956 4436 73958
rect 4460 73956 4516 73958
rect 4220 72922 4276 72924
rect 4300 72922 4356 72924
rect 4380 72922 4436 72924
rect 4460 72922 4516 72924
rect 4220 72870 4246 72922
rect 4246 72870 4276 72922
rect 4300 72870 4310 72922
rect 4310 72870 4356 72922
rect 4380 72870 4426 72922
rect 4426 72870 4436 72922
rect 4460 72870 4490 72922
rect 4490 72870 4516 72922
rect 4220 72868 4276 72870
rect 4300 72868 4356 72870
rect 4380 72868 4436 72870
rect 4460 72868 4516 72870
rect 4220 71834 4276 71836
rect 4300 71834 4356 71836
rect 4380 71834 4436 71836
rect 4460 71834 4516 71836
rect 4220 71782 4246 71834
rect 4246 71782 4276 71834
rect 4300 71782 4310 71834
rect 4310 71782 4356 71834
rect 4380 71782 4426 71834
rect 4426 71782 4436 71834
rect 4460 71782 4490 71834
rect 4490 71782 4516 71834
rect 4220 71780 4276 71782
rect 4300 71780 4356 71782
rect 4380 71780 4436 71782
rect 4460 71780 4516 71782
rect 4220 70746 4276 70748
rect 4300 70746 4356 70748
rect 4380 70746 4436 70748
rect 4460 70746 4516 70748
rect 4220 70694 4246 70746
rect 4246 70694 4276 70746
rect 4300 70694 4310 70746
rect 4310 70694 4356 70746
rect 4380 70694 4426 70746
rect 4426 70694 4436 70746
rect 4460 70694 4490 70746
rect 4490 70694 4516 70746
rect 4220 70692 4276 70694
rect 4300 70692 4356 70694
rect 4380 70692 4436 70694
rect 4460 70692 4516 70694
rect 4220 69658 4276 69660
rect 4300 69658 4356 69660
rect 4380 69658 4436 69660
rect 4460 69658 4516 69660
rect 4220 69606 4246 69658
rect 4246 69606 4276 69658
rect 4300 69606 4310 69658
rect 4310 69606 4356 69658
rect 4380 69606 4426 69658
rect 4426 69606 4436 69658
rect 4460 69606 4490 69658
rect 4490 69606 4516 69658
rect 4220 69604 4276 69606
rect 4300 69604 4356 69606
rect 4380 69604 4436 69606
rect 4460 69604 4516 69606
rect 4220 68570 4276 68572
rect 4300 68570 4356 68572
rect 4380 68570 4436 68572
rect 4460 68570 4516 68572
rect 4220 68518 4246 68570
rect 4246 68518 4276 68570
rect 4300 68518 4310 68570
rect 4310 68518 4356 68570
rect 4380 68518 4426 68570
rect 4426 68518 4436 68570
rect 4460 68518 4490 68570
rect 4490 68518 4516 68570
rect 4220 68516 4276 68518
rect 4300 68516 4356 68518
rect 4380 68516 4436 68518
rect 4460 68516 4516 68518
rect 4220 67482 4276 67484
rect 4300 67482 4356 67484
rect 4380 67482 4436 67484
rect 4460 67482 4516 67484
rect 4220 67430 4246 67482
rect 4246 67430 4276 67482
rect 4300 67430 4310 67482
rect 4310 67430 4356 67482
rect 4380 67430 4426 67482
rect 4426 67430 4436 67482
rect 4460 67430 4490 67482
rect 4490 67430 4516 67482
rect 4220 67428 4276 67430
rect 4300 67428 4356 67430
rect 4380 67428 4436 67430
rect 4460 67428 4516 67430
rect 4220 66394 4276 66396
rect 4300 66394 4356 66396
rect 4380 66394 4436 66396
rect 4460 66394 4516 66396
rect 4220 66342 4246 66394
rect 4246 66342 4276 66394
rect 4300 66342 4310 66394
rect 4310 66342 4356 66394
rect 4380 66342 4426 66394
rect 4426 66342 4436 66394
rect 4460 66342 4490 66394
rect 4490 66342 4516 66394
rect 4220 66340 4276 66342
rect 4300 66340 4356 66342
rect 4380 66340 4436 66342
rect 4460 66340 4516 66342
rect 4220 65306 4276 65308
rect 4300 65306 4356 65308
rect 4380 65306 4436 65308
rect 4460 65306 4516 65308
rect 4220 65254 4246 65306
rect 4246 65254 4276 65306
rect 4300 65254 4310 65306
rect 4310 65254 4356 65306
rect 4380 65254 4426 65306
rect 4426 65254 4436 65306
rect 4460 65254 4490 65306
rect 4490 65254 4516 65306
rect 4220 65252 4276 65254
rect 4300 65252 4356 65254
rect 4380 65252 4436 65254
rect 4460 65252 4516 65254
rect 4220 64218 4276 64220
rect 4300 64218 4356 64220
rect 4380 64218 4436 64220
rect 4460 64218 4516 64220
rect 4220 64166 4246 64218
rect 4246 64166 4276 64218
rect 4300 64166 4310 64218
rect 4310 64166 4356 64218
rect 4380 64166 4426 64218
rect 4426 64166 4436 64218
rect 4460 64166 4490 64218
rect 4490 64166 4516 64218
rect 4220 64164 4276 64166
rect 4300 64164 4356 64166
rect 4380 64164 4436 64166
rect 4460 64164 4516 64166
rect 4220 63130 4276 63132
rect 4300 63130 4356 63132
rect 4380 63130 4436 63132
rect 4460 63130 4516 63132
rect 4220 63078 4246 63130
rect 4246 63078 4276 63130
rect 4300 63078 4310 63130
rect 4310 63078 4356 63130
rect 4380 63078 4426 63130
rect 4426 63078 4436 63130
rect 4460 63078 4490 63130
rect 4490 63078 4516 63130
rect 4220 63076 4276 63078
rect 4300 63076 4356 63078
rect 4380 63076 4436 63078
rect 4460 63076 4516 63078
rect 4220 62042 4276 62044
rect 4300 62042 4356 62044
rect 4380 62042 4436 62044
rect 4460 62042 4516 62044
rect 4220 61990 4246 62042
rect 4246 61990 4276 62042
rect 4300 61990 4310 62042
rect 4310 61990 4356 62042
rect 4380 61990 4426 62042
rect 4426 61990 4436 62042
rect 4460 61990 4490 62042
rect 4490 61990 4516 62042
rect 4220 61988 4276 61990
rect 4300 61988 4356 61990
rect 4380 61988 4436 61990
rect 4460 61988 4516 61990
rect 4220 60954 4276 60956
rect 4300 60954 4356 60956
rect 4380 60954 4436 60956
rect 4460 60954 4516 60956
rect 4220 60902 4246 60954
rect 4246 60902 4276 60954
rect 4300 60902 4310 60954
rect 4310 60902 4356 60954
rect 4380 60902 4426 60954
rect 4426 60902 4436 60954
rect 4460 60902 4490 60954
rect 4490 60902 4516 60954
rect 4220 60900 4276 60902
rect 4300 60900 4356 60902
rect 4380 60900 4436 60902
rect 4460 60900 4516 60902
rect 4220 59866 4276 59868
rect 4300 59866 4356 59868
rect 4380 59866 4436 59868
rect 4460 59866 4516 59868
rect 4220 59814 4246 59866
rect 4246 59814 4276 59866
rect 4300 59814 4310 59866
rect 4310 59814 4356 59866
rect 4380 59814 4426 59866
rect 4426 59814 4436 59866
rect 4460 59814 4490 59866
rect 4490 59814 4516 59866
rect 4220 59812 4276 59814
rect 4300 59812 4356 59814
rect 4380 59812 4436 59814
rect 4460 59812 4516 59814
rect 4220 58778 4276 58780
rect 4300 58778 4356 58780
rect 4380 58778 4436 58780
rect 4460 58778 4516 58780
rect 4220 58726 4246 58778
rect 4246 58726 4276 58778
rect 4300 58726 4310 58778
rect 4310 58726 4356 58778
rect 4380 58726 4426 58778
rect 4426 58726 4436 58778
rect 4460 58726 4490 58778
rect 4490 58726 4516 58778
rect 4220 58724 4276 58726
rect 4300 58724 4356 58726
rect 4380 58724 4436 58726
rect 4460 58724 4516 58726
rect 4220 57690 4276 57692
rect 4300 57690 4356 57692
rect 4380 57690 4436 57692
rect 4460 57690 4516 57692
rect 4220 57638 4246 57690
rect 4246 57638 4276 57690
rect 4300 57638 4310 57690
rect 4310 57638 4356 57690
rect 4380 57638 4426 57690
rect 4426 57638 4436 57690
rect 4460 57638 4490 57690
rect 4490 57638 4516 57690
rect 4220 57636 4276 57638
rect 4300 57636 4356 57638
rect 4380 57636 4436 57638
rect 4460 57636 4516 57638
rect 4220 56602 4276 56604
rect 4300 56602 4356 56604
rect 4380 56602 4436 56604
rect 4460 56602 4516 56604
rect 4220 56550 4246 56602
rect 4246 56550 4276 56602
rect 4300 56550 4310 56602
rect 4310 56550 4356 56602
rect 4380 56550 4426 56602
rect 4426 56550 4436 56602
rect 4460 56550 4490 56602
rect 4490 56550 4516 56602
rect 4220 56548 4276 56550
rect 4300 56548 4356 56550
rect 4380 56548 4436 56550
rect 4460 56548 4516 56550
rect 4220 55514 4276 55516
rect 4300 55514 4356 55516
rect 4380 55514 4436 55516
rect 4460 55514 4516 55516
rect 4220 55462 4246 55514
rect 4246 55462 4276 55514
rect 4300 55462 4310 55514
rect 4310 55462 4356 55514
rect 4380 55462 4426 55514
rect 4426 55462 4436 55514
rect 4460 55462 4490 55514
rect 4490 55462 4516 55514
rect 4220 55460 4276 55462
rect 4300 55460 4356 55462
rect 4380 55460 4436 55462
rect 4460 55460 4516 55462
rect 4220 54426 4276 54428
rect 4300 54426 4356 54428
rect 4380 54426 4436 54428
rect 4460 54426 4516 54428
rect 4220 54374 4246 54426
rect 4246 54374 4276 54426
rect 4300 54374 4310 54426
rect 4310 54374 4356 54426
rect 4380 54374 4426 54426
rect 4426 54374 4436 54426
rect 4460 54374 4490 54426
rect 4490 54374 4516 54426
rect 4220 54372 4276 54374
rect 4300 54372 4356 54374
rect 4380 54372 4436 54374
rect 4460 54372 4516 54374
rect 4220 53338 4276 53340
rect 4300 53338 4356 53340
rect 4380 53338 4436 53340
rect 4460 53338 4516 53340
rect 4220 53286 4246 53338
rect 4246 53286 4276 53338
rect 4300 53286 4310 53338
rect 4310 53286 4356 53338
rect 4380 53286 4426 53338
rect 4426 53286 4436 53338
rect 4460 53286 4490 53338
rect 4490 53286 4516 53338
rect 4220 53284 4276 53286
rect 4300 53284 4356 53286
rect 4380 53284 4436 53286
rect 4460 53284 4516 53286
rect 4220 52250 4276 52252
rect 4300 52250 4356 52252
rect 4380 52250 4436 52252
rect 4460 52250 4516 52252
rect 4220 52198 4246 52250
rect 4246 52198 4276 52250
rect 4300 52198 4310 52250
rect 4310 52198 4356 52250
rect 4380 52198 4426 52250
rect 4426 52198 4436 52250
rect 4460 52198 4490 52250
rect 4490 52198 4516 52250
rect 4220 52196 4276 52198
rect 4300 52196 4356 52198
rect 4380 52196 4436 52198
rect 4460 52196 4516 52198
rect 4220 51162 4276 51164
rect 4300 51162 4356 51164
rect 4380 51162 4436 51164
rect 4460 51162 4516 51164
rect 4220 51110 4246 51162
rect 4246 51110 4276 51162
rect 4300 51110 4310 51162
rect 4310 51110 4356 51162
rect 4380 51110 4426 51162
rect 4426 51110 4436 51162
rect 4460 51110 4490 51162
rect 4490 51110 4516 51162
rect 4220 51108 4276 51110
rect 4300 51108 4356 51110
rect 4380 51108 4436 51110
rect 4460 51108 4516 51110
rect 4220 50074 4276 50076
rect 4300 50074 4356 50076
rect 4380 50074 4436 50076
rect 4460 50074 4516 50076
rect 4220 50022 4246 50074
rect 4246 50022 4276 50074
rect 4300 50022 4310 50074
rect 4310 50022 4356 50074
rect 4380 50022 4426 50074
rect 4426 50022 4436 50074
rect 4460 50022 4490 50074
rect 4490 50022 4516 50074
rect 4220 50020 4276 50022
rect 4300 50020 4356 50022
rect 4380 50020 4436 50022
rect 4460 50020 4516 50022
rect 4220 48986 4276 48988
rect 4300 48986 4356 48988
rect 4380 48986 4436 48988
rect 4460 48986 4516 48988
rect 4220 48934 4246 48986
rect 4246 48934 4276 48986
rect 4300 48934 4310 48986
rect 4310 48934 4356 48986
rect 4380 48934 4426 48986
rect 4426 48934 4436 48986
rect 4460 48934 4490 48986
rect 4490 48934 4516 48986
rect 4220 48932 4276 48934
rect 4300 48932 4356 48934
rect 4380 48932 4436 48934
rect 4460 48932 4516 48934
rect 4220 47898 4276 47900
rect 4300 47898 4356 47900
rect 4380 47898 4436 47900
rect 4460 47898 4516 47900
rect 4220 47846 4246 47898
rect 4246 47846 4276 47898
rect 4300 47846 4310 47898
rect 4310 47846 4356 47898
rect 4380 47846 4426 47898
rect 4426 47846 4436 47898
rect 4460 47846 4490 47898
rect 4490 47846 4516 47898
rect 4220 47844 4276 47846
rect 4300 47844 4356 47846
rect 4380 47844 4436 47846
rect 4460 47844 4516 47846
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 2778 1808 2834 1864
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 19580 116986 19636 116988
rect 19660 116986 19716 116988
rect 19740 116986 19796 116988
rect 19820 116986 19876 116988
rect 19580 116934 19606 116986
rect 19606 116934 19636 116986
rect 19660 116934 19670 116986
rect 19670 116934 19716 116986
rect 19740 116934 19786 116986
rect 19786 116934 19796 116986
rect 19820 116934 19850 116986
rect 19850 116934 19876 116986
rect 19580 116932 19636 116934
rect 19660 116932 19716 116934
rect 19740 116932 19796 116934
rect 19820 116932 19876 116934
rect 19580 115898 19636 115900
rect 19660 115898 19716 115900
rect 19740 115898 19796 115900
rect 19820 115898 19876 115900
rect 19580 115846 19606 115898
rect 19606 115846 19636 115898
rect 19660 115846 19670 115898
rect 19670 115846 19716 115898
rect 19740 115846 19786 115898
rect 19786 115846 19796 115898
rect 19820 115846 19850 115898
rect 19850 115846 19876 115898
rect 19580 115844 19636 115846
rect 19660 115844 19716 115846
rect 19740 115844 19796 115846
rect 19820 115844 19876 115846
rect 19580 114810 19636 114812
rect 19660 114810 19716 114812
rect 19740 114810 19796 114812
rect 19820 114810 19876 114812
rect 19580 114758 19606 114810
rect 19606 114758 19636 114810
rect 19660 114758 19670 114810
rect 19670 114758 19716 114810
rect 19740 114758 19786 114810
rect 19786 114758 19796 114810
rect 19820 114758 19850 114810
rect 19850 114758 19876 114810
rect 19580 114756 19636 114758
rect 19660 114756 19716 114758
rect 19740 114756 19796 114758
rect 19820 114756 19876 114758
rect 21454 115132 21456 115152
rect 21456 115132 21508 115152
rect 21508 115132 21510 115152
rect 21454 115096 21510 115132
rect 22650 116320 22706 116376
rect 22466 116204 22522 116240
rect 22466 116184 22468 116204
rect 22468 116184 22520 116204
rect 22520 116184 22522 116204
rect 23110 116728 23166 116784
rect 23018 115096 23074 115152
rect 19580 113722 19636 113724
rect 19660 113722 19716 113724
rect 19740 113722 19796 113724
rect 19820 113722 19876 113724
rect 19580 113670 19606 113722
rect 19606 113670 19636 113722
rect 19660 113670 19670 113722
rect 19670 113670 19716 113722
rect 19740 113670 19786 113722
rect 19786 113670 19796 113722
rect 19820 113670 19850 113722
rect 19850 113670 19876 113722
rect 19580 113668 19636 113670
rect 19660 113668 19716 113670
rect 19740 113668 19796 113670
rect 19820 113668 19876 113670
rect 19580 112634 19636 112636
rect 19660 112634 19716 112636
rect 19740 112634 19796 112636
rect 19820 112634 19876 112636
rect 19580 112582 19606 112634
rect 19606 112582 19636 112634
rect 19660 112582 19670 112634
rect 19670 112582 19716 112634
rect 19740 112582 19786 112634
rect 19786 112582 19796 112634
rect 19820 112582 19850 112634
rect 19850 112582 19876 112634
rect 19580 112580 19636 112582
rect 19660 112580 19716 112582
rect 19740 112580 19796 112582
rect 19820 112580 19876 112582
rect 19580 111546 19636 111548
rect 19660 111546 19716 111548
rect 19740 111546 19796 111548
rect 19820 111546 19876 111548
rect 19580 111494 19606 111546
rect 19606 111494 19636 111546
rect 19660 111494 19670 111546
rect 19670 111494 19716 111546
rect 19740 111494 19786 111546
rect 19786 111494 19796 111546
rect 19820 111494 19850 111546
rect 19850 111494 19876 111546
rect 19580 111492 19636 111494
rect 19660 111492 19716 111494
rect 19740 111492 19796 111494
rect 19820 111492 19876 111494
rect 19580 110458 19636 110460
rect 19660 110458 19716 110460
rect 19740 110458 19796 110460
rect 19820 110458 19876 110460
rect 19580 110406 19606 110458
rect 19606 110406 19636 110458
rect 19660 110406 19670 110458
rect 19670 110406 19716 110458
rect 19740 110406 19786 110458
rect 19786 110406 19796 110458
rect 19820 110406 19850 110458
rect 19850 110406 19876 110458
rect 19580 110404 19636 110406
rect 19660 110404 19716 110406
rect 19740 110404 19796 110406
rect 19820 110404 19876 110406
rect 19580 109370 19636 109372
rect 19660 109370 19716 109372
rect 19740 109370 19796 109372
rect 19820 109370 19876 109372
rect 19580 109318 19606 109370
rect 19606 109318 19636 109370
rect 19660 109318 19670 109370
rect 19670 109318 19716 109370
rect 19740 109318 19786 109370
rect 19786 109318 19796 109370
rect 19820 109318 19850 109370
rect 19850 109318 19876 109370
rect 19580 109316 19636 109318
rect 19660 109316 19716 109318
rect 19740 109316 19796 109318
rect 19820 109316 19876 109318
rect 24030 115132 24032 115152
rect 24032 115132 24084 115152
rect 24084 115132 24086 115152
rect 24030 115096 24086 115132
rect 24766 116048 24822 116104
rect 24950 117000 25006 117056
rect 25410 116320 25466 116376
rect 25778 117272 25834 117328
rect 26422 116184 26478 116240
rect 26422 114996 26424 115016
rect 26424 114996 26476 115016
rect 26476 114996 26478 115016
rect 26422 114960 26478 114996
rect 26974 117272 27030 117328
rect 28630 117000 28686 117056
rect 28354 116048 28410 116104
rect 19580 108282 19636 108284
rect 19660 108282 19716 108284
rect 19740 108282 19796 108284
rect 19820 108282 19876 108284
rect 19580 108230 19606 108282
rect 19606 108230 19636 108282
rect 19660 108230 19670 108282
rect 19670 108230 19716 108282
rect 19740 108230 19786 108282
rect 19786 108230 19796 108282
rect 19820 108230 19850 108282
rect 19850 108230 19876 108282
rect 19580 108228 19636 108230
rect 19660 108228 19716 108230
rect 19740 108228 19796 108230
rect 19820 108228 19876 108230
rect 19580 107194 19636 107196
rect 19660 107194 19716 107196
rect 19740 107194 19796 107196
rect 19820 107194 19876 107196
rect 19580 107142 19606 107194
rect 19606 107142 19636 107194
rect 19660 107142 19670 107194
rect 19670 107142 19716 107194
rect 19740 107142 19786 107194
rect 19786 107142 19796 107194
rect 19820 107142 19850 107194
rect 19850 107142 19876 107194
rect 19580 107140 19636 107142
rect 19660 107140 19716 107142
rect 19740 107140 19796 107142
rect 19820 107140 19876 107142
rect 19580 106106 19636 106108
rect 19660 106106 19716 106108
rect 19740 106106 19796 106108
rect 19820 106106 19876 106108
rect 19580 106054 19606 106106
rect 19606 106054 19636 106106
rect 19660 106054 19670 106106
rect 19670 106054 19716 106106
rect 19740 106054 19786 106106
rect 19786 106054 19796 106106
rect 19820 106054 19850 106106
rect 19850 106054 19876 106106
rect 19580 106052 19636 106054
rect 19660 106052 19716 106054
rect 19740 106052 19796 106054
rect 19820 106052 19876 106054
rect 19580 105018 19636 105020
rect 19660 105018 19716 105020
rect 19740 105018 19796 105020
rect 19820 105018 19876 105020
rect 19580 104966 19606 105018
rect 19606 104966 19636 105018
rect 19660 104966 19670 105018
rect 19670 104966 19716 105018
rect 19740 104966 19786 105018
rect 19786 104966 19796 105018
rect 19820 104966 19850 105018
rect 19850 104966 19876 105018
rect 19580 104964 19636 104966
rect 19660 104964 19716 104966
rect 19740 104964 19796 104966
rect 19820 104964 19876 104966
rect 19580 103930 19636 103932
rect 19660 103930 19716 103932
rect 19740 103930 19796 103932
rect 19820 103930 19876 103932
rect 19580 103878 19606 103930
rect 19606 103878 19636 103930
rect 19660 103878 19670 103930
rect 19670 103878 19716 103930
rect 19740 103878 19786 103930
rect 19786 103878 19796 103930
rect 19820 103878 19850 103930
rect 19850 103878 19876 103930
rect 19580 103876 19636 103878
rect 19660 103876 19716 103878
rect 19740 103876 19796 103878
rect 19820 103876 19876 103878
rect 19580 102842 19636 102844
rect 19660 102842 19716 102844
rect 19740 102842 19796 102844
rect 19820 102842 19876 102844
rect 19580 102790 19606 102842
rect 19606 102790 19636 102842
rect 19660 102790 19670 102842
rect 19670 102790 19716 102842
rect 19740 102790 19786 102842
rect 19786 102790 19796 102842
rect 19820 102790 19850 102842
rect 19850 102790 19876 102842
rect 19580 102788 19636 102790
rect 19660 102788 19716 102790
rect 19740 102788 19796 102790
rect 19820 102788 19876 102790
rect 19580 101754 19636 101756
rect 19660 101754 19716 101756
rect 19740 101754 19796 101756
rect 19820 101754 19876 101756
rect 19580 101702 19606 101754
rect 19606 101702 19636 101754
rect 19660 101702 19670 101754
rect 19670 101702 19716 101754
rect 19740 101702 19786 101754
rect 19786 101702 19796 101754
rect 19820 101702 19850 101754
rect 19850 101702 19876 101754
rect 19580 101700 19636 101702
rect 19660 101700 19716 101702
rect 19740 101700 19796 101702
rect 19820 101700 19876 101702
rect 19580 100666 19636 100668
rect 19660 100666 19716 100668
rect 19740 100666 19796 100668
rect 19820 100666 19876 100668
rect 19580 100614 19606 100666
rect 19606 100614 19636 100666
rect 19660 100614 19670 100666
rect 19670 100614 19716 100666
rect 19740 100614 19786 100666
rect 19786 100614 19796 100666
rect 19820 100614 19850 100666
rect 19850 100614 19876 100666
rect 19580 100612 19636 100614
rect 19660 100612 19716 100614
rect 19740 100612 19796 100614
rect 19820 100612 19876 100614
rect 19580 99578 19636 99580
rect 19660 99578 19716 99580
rect 19740 99578 19796 99580
rect 19820 99578 19876 99580
rect 19580 99526 19606 99578
rect 19606 99526 19636 99578
rect 19660 99526 19670 99578
rect 19670 99526 19716 99578
rect 19740 99526 19786 99578
rect 19786 99526 19796 99578
rect 19820 99526 19850 99578
rect 19850 99526 19876 99578
rect 19580 99524 19636 99526
rect 19660 99524 19716 99526
rect 19740 99524 19796 99526
rect 19820 99524 19876 99526
rect 19580 98490 19636 98492
rect 19660 98490 19716 98492
rect 19740 98490 19796 98492
rect 19820 98490 19876 98492
rect 19580 98438 19606 98490
rect 19606 98438 19636 98490
rect 19660 98438 19670 98490
rect 19670 98438 19716 98490
rect 19740 98438 19786 98490
rect 19786 98438 19796 98490
rect 19820 98438 19850 98490
rect 19850 98438 19876 98490
rect 19580 98436 19636 98438
rect 19660 98436 19716 98438
rect 19740 98436 19796 98438
rect 19820 98436 19876 98438
rect 19580 97402 19636 97404
rect 19660 97402 19716 97404
rect 19740 97402 19796 97404
rect 19820 97402 19876 97404
rect 19580 97350 19606 97402
rect 19606 97350 19636 97402
rect 19660 97350 19670 97402
rect 19670 97350 19716 97402
rect 19740 97350 19786 97402
rect 19786 97350 19796 97402
rect 19820 97350 19850 97402
rect 19850 97350 19876 97402
rect 19580 97348 19636 97350
rect 19660 97348 19716 97350
rect 19740 97348 19796 97350
rect 19820 97348 19876 97350
rect 19580 96314 19636 96316
rect 19660 96314 19716 96316
rect 19740 96314 19796 96316
rect 19820 96314 19876 96316
rect 19580 96262 19606 96314
rect 19606 96262 19636 96314
rect 19660 96262 19670 96314
rect 19670 96262 19716 96314
rect 19740 96262 19786 96314
rect 19786 96262 19796 96314
rect 19820 96262 19850 96314
rect 19850 96262 19876 96314
rect 19580 96260 19636 96262
rect 19660 96260 19716 96262
rect 19740 96260 19796 96262
rect 19820 96260 19876 96262
rect 19580 95226 19636 95228
rect 19660 95226 19716 95228
rect 19740 95226 19796 95228
rect 19820 95226 19876 95228
rect 19580 95174 19606 95226
rect 19606 95174 19636 95226
rect 19660 95174 19670 95226
rect 19670 95174 19716 95226
rect 19740 95174 19786 95226
rect 19786 95174 19796 95226
rect 19820 95174 19850 95226
rect 19850 95174 19876 95226
rect 19580 95172 19636 95174
rect 19660 95172 19716 95174
rect 19740 95172 19796 95174
rect 19820 95172 19876 95174
rect 19580 94138 19636 94140
rect 19660 94138 19716 94140
rect 19740 94138 19796 94140
rect 19820 94138 19876 94140
rect 19580 94086 19606 94138
rect 19606 94086 19636 94138
rect 19660 94086 19670 94138
rect 19670 94086 19716 94138
rect 19740 94086 19786 94138
rect 19786 94086 19796 94138
rect 19820 94086 19850 94138
rect 19850 94086 19876 94138
rect 19580 94084 19636 94086
rect 19660 94084 19716 94086
rect 19740 94084 19796 94086
rect 19820 94084 19876 94086
rect 19580 93050 19636 93052
rect 19660 93050 19716 93052
rect 19740 93050 19796 93052
rect 19820 93050 19876 93052
rect 19580 92998 19606 93050
rect 19606 92998 19636 93050
rect 19660 92998 19670 93050
rect 19670 92998 19716 93050
rect 19740 92998 19786 93050
rect 19786 92998 19796 93050
rect 19820 92998 19850 93050
rect 19850 92998 19876 93050
rect 19580 92996 19636 92998
rect 19660 92996 19716 92998
rect 19740 92996 19796 92998
rect 19820 92996 19876 92998
rect 19580 91962 19636 91964
rect 19660 91962 19716 91964
rect 19740 91962 19796 91964
rect 19820 91962 19876 91964
rect 19580 91910 19606 91962
rect 19606 91910 19636 91962
rect 19660 91910 19670 91962
rect 19670 91910 19716 91962
rect 19740 91910 19786 91962
rect 19786 91910 19796 91962
rect 19820 91910 19850 91962
rect 19850 91910 19876 91962
rect 19580 91908 19636 91910
rect 19660 91908 19716 91910
rect 19740 91908 19796 91910
rect 19820 91908 19876 91910
rect 19580 90874 19636 90876
rect 19660 90874 19716 90876
rect 19740 90874 19796 90876
rect 19820 90874 19876 90876
rect 19580 90822 19606 90874
rect 19606 90822 19636 90874
rect 19660 90822 19670 90874
rect 19670 90822 19716 90874
rect 19740 90822 19786 90874
rect 19786 90822 19796 90874
rect 19820 90822 19850 90874
rect 19850 90822 19876 90874
rect 19580 90820 19636 90822
rect 19660 90820 19716 90822
rect 19740 90820 19796 90822
rect 19820 90820 19876 90822
rect 19580 89786 19636 89788
rect 19660 89786 19716 89788
rect 19740 89786 19796 89788
rect 19820 89786 19876 89788
rect 19580 89734 19606 89786
rect 19606 89734 19636 89786
rect 19660 89734 19670 89786
rect 19670 89734 19716 89786
rect 19740 89734 19786 89786
rect 19786 89734 19796 89786
rect 19820 89734 19850 89786
rect 19850 89734 19876 89786
rect 19580 89732 19636 89734
rect 19660 89732 19716 89734
rect 19740 89732 19796 89734
rect 19820 89732 19876 89734
rect 19580 88698 19636 88700
rect 19660 88698 19716 88700
rect 19740 88698 19796 88700
rect 19820 88698 19876 88700
rect 19580 88646 19606 88698
rect 19606 88646 19636 88698
rect 19660 88646 19670 88698
rect 19670 88646 19716 88698
rect 19740 88646 19786 88698
rect 19786 88646 19796 88698
rect 19820 88646 19850 88698
rect 19850 88646 19876 88698
rect 19580 88644 19636 88646
rect 19660 88644 19716 88646
rect 19740 88644 19796 88646
rect 19820 88644 19876 88646
rect 19580 87610 19636 87612
rect 19660 87610 19716 87612
rect 19740 87610 19796 87612
rect 19820 87610 19876 87612
rect 19580 87558 19606 87610
rect 19606 87558 19636 87610
rect 19660 87558 19670 87610
rect 19670 87558 19716 87610
rect 19740 87558 19786 87610
rect 19786 87558 19796 87610
rect 19820 87558 19850 87610
rect 19850 87558 19876 87610
rect 19580 87556 19636 87558
rect 19660 87556 19716 87558
rect 19740 87556 19796 87558
rect 19820 87556 19876 87558
rect 19580 86522 19636 86524
rect 19660 86522 19716 86524
rect 19740 86522 19796 86524
rect 19820 86522 19876 86524
rect 19580 86470 19606 86522
rect 19606 86470 19636 86522
rect 19660 86470 19670 86522
rect 19670 86470 19716 86522
rect 19740 86470 19786 86522
rect 19786 86470 19796 86522
rect 19820 86470 19850 86522
rect 19850 86470 19876 86522
rect 19580 86468 19636 86470
rect 19660 86468 19716 86470
rect 19740 86468 19796 86470
rect 19820 86468 19876 86470
rect 19580 85434 19636 85436
rect 19660 85434 19716 85436
rect 19740 85434 19796 85436
rect 19820 85434 19876 85436
rect 19580 85382 19606 85434
rect 19606 85382 19636 85434
rect 19660 85382 19670 85434
rect 19670 85382 19716 85434
rect 19740 85382 19786 85434
rect 19786 85382 19796 85434
rect 19820 85382 19850 85434
rect 19850 85382 19876 85434
rect 19580 85380 19636 85382
rect 19660 85380 19716 85382
rect 19740 85380 19796 85382
rect 19820 85380 19876 85382
rect 19580 84346 19636 84348
rect 19660 84346 19716 84348
rect 19740 84346 19796 84348
rect 19820 84346 19876 84348
rect 19580 84294 19606 84346
rect 19606 84294 19636 84346
rect 19660 84294 19670 84346
rect 19670 84294 19716 84346
rect 19740 84294 19786 84346
rect 19786 84294 19796 84346
rect 19820 84294 19850 84346
rect 19850 84294 19876 84346
rect 19580 84292 19636 84294
rect 19660 84292 19716 84294
rect 19740 84292 19796 84294
rect 19820 84292 19876 84294
rect 19580 83258 19636 83260
rect 19660 83258 19716 83260
rect 19740 83258 19796 83260
rect 19820 83258 19876 83260
rect 19580 83206 19606 83258
rect 19606 83206 19636 83258
rect 19660 83206 19670 83258
rect 19670 83206 19716 83258
rect 19740 83206 19786 83258
rect 19786 83206 19796 83258
rect 19820 83206 19850 83258
rect 19850 83206 19876 83258
rect 19580 83204 19636 83206
rect 19660 83204 19716 83206
rect 19740 83204 19796 83206
rect 19820 83204 19876 83206
rect 19580 82170 19636 82172
rect 19660 82170 19716 82172
rect 19740 82170 19796 82172
rect 19820 82170 19876 82172
rect 19580 82118 19606 82170
rect 19606 82118 19636 82170
rect 19660 82118 19670 82170
rect 19670 82118 19716 82170
rect 19740 82118 19786 82170
rect 19786 82118 19796 82170
rect 19820 82118 19850 82170
rect 19850 82118 19876 82170
rect 19580 82116 19636 82118
rect 19660 82116 19716 82118
rect 19740 82116 19796 82118
rect 19820 82116 19876 82118
rect 19580 81082 19636 81084
rect 19660 81082 19716 81084
rect 19740 81082 19796 81084
rect 19820 81082 19876 81084
rect 19580 81030 19606 81082
rect 19606 81030 19636 81082
rect 19660 81030 19670 81082
rect 19670 81030 19716 81082
rect 19740 81030 19786 81082
rect 19786 81030 19796 81082
rect 19820 81030 19850 81082
rect 19850 81030 19876 81082
rect 19580 81028 19636 81030
rect 19660 81028 19716 81030
rect 19740 81028 19796 81030
rect 19820 81028 19876 81030
rect 19580 79994 19636 79996
rect 19660 79994 19716 79996
rect 19740 79994 19796 79996
rect 19820 79994 19876 79996
rect 19580 79942 19606 79994
rect 19606 79942 19636 79994
rect 19660 79942 19670 79994
rect 19670 79942 19716 79994
rect 19740 79942 19786 79994
rect 19786 79942 19796 79994
rect 19820 79942 19850 79994
rect 19850 79942 19876 79994
rect 19580 79940 19636 79942
rect 19660 79940 19716 79942
rect 19740 79940 19796 79942
rect 19820 79940 19876 79942
rect 19580 78906 19636 78908
rect 19660 78906 19716 78908
rect 19740 78906 19796 78908
rect 19820 78906 19876 78908
rect 19580 78854 19606 78906
rect 19606 78854 19636 78906
rect 19660 78854 19670 78906
rect 19670 78854 19716 78906
rect 19740 78854 19786 78906
rect 19786 78854 19796 78906
rect 19820 78854 19850 78906
rect 19850 78854 19876 78906
rect 19580 78852 19636 78854
rect 19660 78852 19716 78854
rect 19740 78852 19796 78854
rect 19820 78852 19876 78854
rect 19580 77818 19636 77820
rect 19660 77818 19716 77820
rect 19740 77818 19796 77820
rect 19820 77818 19876 77820
rect 19580 77766 19606 77818
rect 19606 77766 19636 77818
rect 19660 77766 19670 77818
rect 19670 77766 19716 77818
rect 19740 77766 19786 77818
rect 19786 77766 19796 77818
rect 19820 77766 19850 77818
rect 19850 77766 19876 77818
rect 19580 77764 19636 77766
rect 19660 77764 19716 77766
rect 19740 77764 19796 77766
rect 19820 77764 19876 77766
rect 19580 76730 19636 76732
rect 19660 76730 19716 76732
rect 19740 76730 19796 76732
rect 19820 76730 19876 76732
rect 19580 76678 19606 76730
rect 19606 76678 19636 76730
rect 19660 76678 19670 76730
rect 19670 76678 19716 76730
rect 19740 76678 19786 76730
rect 19786 76678 19796 76730
rect 19820 76678 19850 76730
rect 19850 76678 19876 76730
rect 19580 76676 19636 76678
rect 19660 76676 19716 76678
rect 19740 76676 19796 76678
rect 19820 76676 19876 76678
rect 19580 75642 19636 75644
rect 19660 75642 19716 75644
rect 19740 75642 19796 75644
rect 19820 75642 19876 75644
rect 19580 75590 19606 75642
rect 19606 75590 19636 75642
rect 19660 75590 19670 75642
rect 19670 75590 19716 75642
rect 19740 75590 19786 75642
rect 19786 75590 19796 75642
rect 19820 75590 19850 75642
rect 19850 75590 19876 75642
rect 19580 75588 19636 75590
rect 19660 75588 19716 75590
rect 19740 75588 19796 75590
rect 19820 75588 19876 75590
rect 19580 74554 19636 74556
rect 19660 74554 19716 74556
rect 19740 74554 19796 74556
rect 19820 74554 19876 74556
rect 19580 74502 19606 74554
rect 19606 74502 19636 74554
rect 19660 74502 19670 74554
rect 19670 74502 19716 74554
rect 19740 74502 19786 74554
rect 19786 74502 19796 74554
rect 19820 74502 19850 74554
rect 19850 74502 19876 74554
rect 19580 74500 19636 74502
rect 19660 74500 19716 74502
rect 19740 74500 19796 74502
rect 19820 74500 19876 74502
rect 19580 73466 19636 73468
rect 19660 73466 19716 73468
rect 19740 73466 19796 73468
rect 19820 73466 19876 73468
rect 19580 73414 19606 73466
rect 19606 73414 19636 73466
rect 19660 73414 19670 73466
rect 19670 73414 19716 73466
rect 19740 73414 19786 73466
rect 19786 73414 19796 73466
rect 19820 73414 19850 73466
rect 19850 73414 19876 73466
rect 19580 73412 19636 73414
rect 19660 73412 19716 73414
rect 19740 73412 19796 73414
rect 19820 73412 19876 73414
rect 19580 72378 19636 72380
rect 19660 72378 19716 72380
rect 19740 72378 19796 72380
rect 19820 72378 19876 72380
rect 19580 72326 19606 72378
rect 19606 72326 19636 72378
rect 19660 72326 19670 72378
rect 19670 72326 19716 72378
rect 19740 72326 19786 72378
rect 19786 72326 19796 72378
rect 19820 72326 19850 72378
rect 19850 72326 19876 72378
rect 19580 72324 19636 72326
rect 19660 72324 19716 72326
rect 19740 72324 19796 72326
rect 19820 72324 19876 72326
rect 19580 71290 19636 71292
rect 19660 71290 19716 71292
rect 19740 71290 19796 71292
rect 19820 71290 19876 71292
rect 19580 71238 19606 71290
rect 19606 71238 19636 71290
rect 19660 71238 19670 71290
rect 19670 71238 19716 71290
rect 19740 71238 19786 71290
rect 19786 71238 19796 71290
rect 19820 71238 19850 71290
rect 19850 71238 19876 71290
rect 19580 71236 19636 71238
rect 19660 71236 19716 71238
rect 19740 71236 19796 71238
rect 19820 71236 19876 71238
rect 19580 70202 19636 70204
rect 19660 70202 19716 70204
rect 19740 70202 19796 70204
rect 19820 70202 19876 70204
rect 19580 70150 19606 70202
rect 19606 70150 19636 70202
rect 19660 70150 19670 70202
rect 19670 70150 19716 70202
rect 19740 70150 19786 70202
rect 19786 70150 19796 70202
rect 19820 70150 19850 70202
rect 19850 70150 19876 70202
rect 19580 70148 19636 70150
rect 19660 70148 19716 70150
rect 19740 70148 19796 70150
rect 19820 70148 19876 70150
rect 19580 69114 19636 69116
rect 19660 69114 19716 69116
rect 19740 69114 19796 69116
rect 19820 69114 19876 69116
rect 19580 69062 19606 69114
rect 19606 69062 19636 69114
rect 19660 69062 19670 69114
rect 19670 69062 19716 69114
rect 19740 69062 19786 69114
rect 19786 69062 19796 69114
rect 19820 69062 19850 69114
rect 19850 69062 19876 69114
rect 19580 69060 19636 69062
rect 19660 69060 19716 69062
rect 19740 69060 19796 69062
rect 19820 69060 19876 69062
rect 19580 68026 19636 68028
rect 19660 68026 19716 68028
rect 19740 68026 19796 68028
rect 19820 68026 19876 68028
rect 19580 67974 19606 68026
rect 19606 67974 19636 68026
rect 19660 67974 19670 68026
rect 19670 67974 19716 68026
rect 19740 67974 19786 68026
rect 19786 67974 19796 68026
rect 19820 67974 19850 68026
rect 19850 67974 19876 68026
rect 19580 67972 19636 67974
rect 19660 67972 19716 67974
rect 19740 67972 19796 67974
rect 19820 67972 19876 67974
rect 19580 66938 19636 66940
rect 19660 66938 19716 66940
rect 19740 66938 19796 66940
rect 19820 66938 19876 66940
rect 19580 66886 19606 66938
rect 19606 66886 19636 66938
rect 19660 66886 19670 66938
rect 19670 66886 19716 66938
rect 19740 66886 19786 66938
rect 19786 66886 19796 66938
rect 19820 66886 19850 66938
rect 19850 66886 19876 66938
rect 19580 66884 19636 66886
rect 19660 66884 19716 66886
rect 19740 66884 19796 66886
rect 19820 66884 19876 66886
rect 19580 65850 19636 65852
rect 19660 65850 19716 65852
rect 19740 65850 19796 65852
rect 19820 65850 19876 65852
rect 19580 65798 19606 65850
rect 19606 65798 19636 65850
rect 19660 65798 19670 65850
rect 19670 65798 19716 65850
rect 19740 65798 19786 65850
rect 19786 65798 19796 65850
rect 19820 65798 19850 65850
rect 19850 65798 19876 65850
rect 19580 65796 19636 65798
rect 19660 65796 19716 65798
rect 19740 65796 19796 65798
rect 19820 65796 19876 65798
rect 19580 64762 19636 64764
rect 19660 64762 19716 64764
rect 19740 64762 19796 64764
rect 19820 64762 19876 64764
rect 19580 64710 19606 64762
rect 19606 64710 19636 64762
rect 19660 64710 19670 64762
rect 19670 64710 19716 64762
rect 19740 64710 19786 64762
rect 19786 64710 19796 64762
rect 19820 64710 19850 64762
rect 19850 64710 19876 64762
rect 19580 64708 19636 64710
rect 19660 64708 19716 64710
rect 19740 64708 19796 64710
rect 19820 64708 19876 64710
rect 19580 63674 19636 63676
rect 19660 63674 19716 63676
rect 19740 63674 19796 63676
rect 19820 63674 19876 63676
rect 19580 63622 19606 63674
rect 19606 63622 19636 63674
rect 19660 63622 19670 63674
rect 19670 63622 19716 63674
rect 19740 63622 19786 63674
rect 19786 63622 19796 63674
rect 19820 63622 19850 63674
rect 19850 63622 19876 63674
rect 19580 63620 19636 63622
rect 19660 63620 19716 63622
rect 19740 63620 19796 63622
rect 19820 63620 19876 63622
rect 19580 62586 19636 62588
rect 19660 62586 19716 62588
rect 19740 62586 19796 62588
rect 19820 62586 19876 62588
rect 19580 62534 19606 62586
rect 19606 62534 19636 62586
rect 19660 62534 19670 62586
rect 19670 62534 19716 62586
rect 19740 62534 19786 62586
rect 19786 62534 19796 62586
rect 19820 62534 19850 62586
rect 19850 62534 19876 62586
rect 19580 62532 19636 62534
rect 19660 62532 19716 62534
rect 19740 62532 19796 62534
rect 19820 62532 19876 62534
rect 19580 61498 19636 61500
rect 19660 61498 19716 61500
rect 19740 61498 19796 61500
rect 19820 61498 19876 61500
rect 19580 61446 19606 61498
rect 19606 61446 19636 61498
rect 19660 61446 19670 61498
rect 19670 61446 19716 61498
rect 19740 61446 19786 61498
rect 19786 61446 19796 61498
rect 19820 61446 19850 61498
rect 19850 61446 19876 61498
rect 19580 61444 19636 61446
rect 19660 61444 19716 61446
rect 19740 61444 19796 61446
rect 19820 61444 19876 61446
rect 19580 60410 19636 60412
rect 19660 60410 19716 60412
rect 19740 60410 19796 60412
rect 19820 60410 19876 60412
rect 19580 60358 19606 60410
rect 19606 60358 19636 60410
rect 19660 60358 19670 60410
rect 19670 60358 19716 60410
rect 19740 60358 19786 60410
rect 19786 60358 19796 60410
rect 19820 60358 19850 60410
rect 19850 60358 19876 60410
rect 19580 60356 19636 60358
rect 19660 60356 19716 60358
rect 19740 60356 19796 60358
rect 19820 60356 19876 60358
rect 19580 59322 19636 59324
rect 19660 59322 19716 59324
rect 19740 59322 19796 59324
rect 19820 59322 19876 59324
rect 19580 59270 19606 59322
rect 19606 59270 19636 59322
rect 19660 59270 19670 59322
rect 19670 59270 19716 59322
rect 19740 59270 19786 59322
rect 19786 59270 19796 59322
rect 19820 59270 19850 59322
rect 19850 59270 19876 59322
rect 19580 59268 19636 59270
rect 19660 59268 19716 59270
rect 19740 59268 19796 59270
rect 19820 59268 19876 59270
rect 19580 58234 19636 58236
rect 19660 58234 19716 58236
rect 19740 58234 19796 58236
rect 19820 58234 19876 58236
rect 19580 58182 19606 58234
rect 19606 58182 19636 58234
rect 19660 58182 19670 58234
rect 19670 58182 19716 58234
rect 19740 58182 19786 58234
rect 19786 58182 19796 58234
rect 19820 58182 19850 58234
rect 19850 58182 19876 58234
rect 19580 58180 19636 58182
rect 19660 58180 19716 58182
rect 19740 58180 19796 58182
rect 19820 58180 19876 58182
rect 19580 57146 19636 57148
rect 19660 57146 19716 57148
rect 19740 57146 19796 57148
rect 19820 57146 19876 57148
rect 19580 57094 19606 57146
rect 19606 57094 19636 57146
rect 19660 57094 19670 57146
rect 19670 57094 19716 57146
rect 19740 57094 19786 57146
rect 19786 57094 19796 57146
rect 19820 57094 19850 57146
rect 19850 57094 19876 57146
rect 19580 57092 19636 57094
rect 19660 57092 19716 57094
rect 19740 57092 19796 57094
rect 19820 57092 19876 57094
rect 19580 56058 19636 56060
rect 19660 56058 19716 56060
rect 19740 56058 19796 56060
rect 19820 56058 19876 56060
rect 19580 56006 19606 56058
rect 19606 56006 19636 56058
rect 19660 56006 19670 56058
rect 19670 56006 19716 56058
rect 19740 56006 19786 56058
rect 19786 56006 19796 56058
rect 19820 56006 19850 56058
rect 19850 56006 19876 56058
rect 19580 56004 19636 56006
rect 19660 56004 19716 56006
rect 19740 56004 19796 56006
rect 19820 56004 19876 56006
rect 19580 54970 19636 54972
rect 19660 54970 19716 54972
rect 19740 54970 19796 54972
rect 19820 54970 19876 54972
rect 19580 54918 19606 54970
rect 19606 54918 19636 54970
rect 19660 54918 19670 54970
rect 19670 54918 19716 54970
rect 19740 54918 19786 54970
rect 19786 54918 19796 54970
rect 19820 54918 19850 54970
rect 19850 54918 19876 54970
rect 19580 54916 19636 54918
rect 19660 54916 19716 54918
rect 19740 54916 19796 54918
rect 19820 54916 19876 54918
rect 19580 53882 19636 53884
rect 19660 53882 19716 53884
rect 19740 53882 19796 53884
rect 19820 53882 19876 53884
rect 19580 53830 19606 53882
rect 19606 53830 19636 53882
rect 19660 53830 19670 53882
rect 19670 53830 19716 53882
rect 19740 53830 19786 53882
rect 19786 53830 19796 53882
rect 19820 53830 19850 53882
rect 19850 53830 19876 53882
rect 19580 53828 19636 53830
rect 19660 53828 19716 53830
rect 19740 53828 19796 53830
rect 19820 53828 19876 53830
rect 19580 52794 19636 52796
rect 19660 52794 19716 52796
rect 19740 52794 19796 52796
rect 19820 52794 19876 52796
rect 19580 52742 19606 52794
rect 19606 52742 19636 52794
rect 19660 52742 19670 52794
rect 19670 52742 19716 52794
rect 19740 52742 19786 52794
rect 19786 52742 19796 52794
rect 19820 52742 19850 52794
rect 19850 52742 19876 52794
rect 19580 52740 19636 52742
rect 19660 52740 19716 52742
rect 19740 52740 19796 52742
rect 19820 52740 19876 52742
rect 19580 51706 19636 51708
rect 19660 51706 19716 51708
rect 19740 51706 19796 51708
rect 19820 51706 19876 51708
rect 19580 51654 19606 51706
rect 19606 51654 19636 51706
rect 19660 51654 19670 51706
rect 19670 51654 19716 51706
rect 19740 51654 19786 51706
rect 19786 51654 19796 51706
rect 19820 51654 19850 51706
rect 19850 51654 19876 51706
rect 19580 51652 19636 51654
rect 19660 51652 19716 51654
rect 19740 51652 19796 51654
rect 19820 51652 19876 51654
rect 19580 50618 19636 50620
rect 19660 50618 19716 50620
rect 19740 50618 19796 50620
rect 19820 50618 19876 50620
rect 19580 50566 19606 50618
rect 19606 50566 19636 50618
rect 19660 50566 19670 50618
rect 19670 50566 19716 50618
rect 19740 50566 19786 50618
rect 19786 50566 19796 50618
rect 19820 50566 19850 50618
rect 19850 50566 19876 50618
rect 19580 50564 19636 50566
rect 19660 50564 19716 50566
rect 19740 50564 19796 50566
rect 19820 50564 19876 50566
rect 19580 49530 19636 49532
rect 19660 49530 19716 49532
rect 19740 49530 19796 49532
rect 19820 49530 19876 49532
rect 19580 49478 19606 49530
rect 19606 49478 19636 49530
rect 19660 49478 19670 49530
rect 19670 49478 19716 49530
rect 19740 49478 19786 49530
rect 19786 49478 19796 49530
rect 19820 49478 19850 49530
rect 19850 49478 19876 49530
rect 19580 49476 19636 49478
rect 19660 49476 19716 49478
rect 19740 49476 19796 49478
rect 19820 49476 19876 49478
rect 19580 48442 19636 48444
rect 19660 48442 19716 48444
rect 19740 48442 19796 48444
rect 19820 48442 19876 48444
rect 19580 48390 19606 48442
rect 19606 48390 19636 48442
rect 19660 48390 19670 48442
rect 19670 48390 19716 48442
rect 19740 48390 19786 48442
rect 19786 48390 19796 48442
rect 19820 48390 19850 48442
rect 19850 48390 19876 48442
rect 19580 48388 19636 48390
rect 19660 48388 19716 48390
rect 19740 48388 19796 48390
rect 19820 48388 19876 48390
rect 19580 47354 19636 47356
rect 19660 47354 19716 47356
rect 19740 47354 19796 47356
rect 19820 47354 19876 47356
rect 19580 47302 19606 47354
rect 19606 47302 19636 47354
rect 19660 47302 19670 47354
rect 19670 47302 19716 47354
rect 19740 47302 19786 47354
rect 19786 47302 19796 47354
rect 19820 47302 19850 47354
rect 19850 47302 19876 47354
rect 19580 47300 19636 47302
rect 19660 47300 19716 47302
rect 19740 47300 19796 47302
rect 19820 47300 19876 47302
rect 19580 46266 19636 46268
rect 19660 46266 19716 46268
rect 19740 46266 19796 46268
rect 19820 46266 19876 46268
rect 19580 46214 19606 46266
rect 19606 46214 19636 46266
rect 19660 46214 19670 46266
rect 19670 46214 19716 46266
rect 19740 46214 19786 46266
rect 19786 46214 19796 46266
rect 19820 46214 19850 46266
rect 19850 46214 19876 46266
rect 19580 46212 19636 46214
rect 19660 46212 19716 46214
rect 19740 46212 19796 46214
rect 19820 46212 19876 46214
rect 19580 45178 19636 45180
rect 19660 45178 19716 45180
rect 19740 45178 19796 45180
rect 19820 45178 19876 45180
rect 19580 45126 19606 45178
rect 19606 45126 19636 45178
rect 19660 45126 19670 45178
rect 19670 45126 19716 45178
rect 19740 45126 19786 45178
rect 19786 45126 19796 45178
rect 19820 45126 19850 45178
rect 19850 45126 19876 45178
rect 19580 45124 19636 45126
rect 19660 45124 19716 45126
rect 19740 45124 19796 45126
rect 19820 45124 19876 45126
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 23570 14728 23626 14784
rect 23478 14476 23534 14512
rect 23478 14456 23480 14476
rect 23480 14456 23532 14476
rect 23532 14456 23534 14476
rect 23662 14356 23664 14376
rect 23664 14356 23716 14376
rect 23716 14356 23718 14376
rect 23662 14320 23718 14356
rect 24214 13504 24270 13560
rect 25134 18672 25190 18728
rect 25134 14728 25190 14784
rect 26054 14456 26110 14512
rect 26606 18672 26662 18728
rect 28998 115892 29054 115948
rect 29182 115776 29238 115832
rect 29182 115232 29238 115288
rect 28814 114996 28816 115016
rect 28816 114996 28868 115016
rect 28868 114996 28870 115016
rect 28814 114960 28870 114996
rect 29550 115796 29606 115832
rect 29550 115776 29552 115796
rect 29552 115776 29604 115796
rect 29604 115776 29606 115796
rect 29550 115640 29606 115696
rect 29366 115096 29422 115152
rect 30378 115912 30434 115968
rect 30286 115232 30342 115288
rect 25042 3460 25098 3496
rect 25042 3440 25044 3460
rect 25044 3440 25096 3460
rect 25096 3440 25098 3460
rect 26330 3712 26386 3768
rect 26606 3168 26662 3224
rect 26330 2896 26386 2952
rect 27434 14728 27490 14784
rect 27618 13504 27674 13560
rect 27894 15408 27950 15464
rect 27802 14456 27858 14512
rect 28262 18672 28318 18728
rect 28998 17584 29054 17640
rect 28906 14900 28908 14920
rect 28908 14900 28960 14920
rect 28960 14900 28962 14920
rect 28906 14864 28962 14900
rect 28906 14728 28962 14784
rect 29642 86264 29698 86320
rect 29550 18400 29606 18456
rect 29182 14356 29184 14376
rect 29184 14356 29236 14376
rect 29236 14356 29238 14376
rect 29182 14320 29238 14356
rect 29734 14728 29790 14784
rect 28630 3188 28686 3224
rect 28630 3168 28632 3188
rect 28632 3168 28684 3188
rect 28684 3168 28686 3188
rect 28998 3068 29000 3088
rect 29000 3068 29052 3088
rect 29052 3068 29054 3088
rect 28998 3032 29054 3068
rect 30930 116068 30986 116104
rect 30930 116048 30932 116068
rect 30932 116048 30984 116068
rect 30984 116048 30986 116068
rect 30194 17584 30250 17640
rect 30562 19760 30618 19816
rect 30286 16496 30342 16552
rect 31758 116084 31760 116104
rect 31760 116084 31812 116104
rect 31812 116084 31814 116104
rect 31758 116048 31814 116084
rect 32402 115912 32458 115968
rect 30746 19760 30802 19816
rect 30378 14864 30434 14920
rect 29366 3848 29422 3904
rect 29182 2896 29238 2952
rect 30930 20032 30986 20088
rect 30010 3576 30066 3632
rect 30470 3032 30526 3088
rect 30654 3032 30710 3088
rect 31022 3848 31078 3904
rect 31114 3596 31170 3632
rect 31114 3576 31116 3596
rect 31116 3576 31168 3596
rect 31168 3576 31170 3596
rect 31482 23044 31538 23080
rect 31482 23024 31484 23044
rect 31484 23024 31536 23044
rect 31536 23024 31538 23044
rect 31390 15428 31446 15464
rect 31390 15408 31392 15428
rect 31392 15408 31444 15428
rect 31444 15408 31446 15428
rect 32402 36080 32458 36136
rect 32770 81504 32826 81560
rect 33046 81912 33102 81968
rect 34610 118768 34666 118824
rect 34940 117530 34996 117532
rect 35020 117530 35076 117532
rect 35100 117530 35156 117532
rect 35180 117530 35236 117532
rect 34940 117478 34966 117530
rect 34966 117478 34996 117530
rect 35020 117478 35030 117530
rect 35030 117478 35076 117530
rect 35100 117478 35146 117530
rect 35146 117478 35156 117530
rect 35180 117478 35210 117530
rect 35210 117478 35236 117530
rect 34940 117476 34996 117478
rect 35020 117476 35076 117478
rect 35100 117476 35156 117478
rect 35180 117476 35236 117478
rect 33598 62872 33654 62928
rect 34518 115676 34520 115696
rect 34520 115676 34572 115696
rect 34572 115676 34574 115696
rect 34518 115640 34574 115676
rect 32034 21664 32090 21720
rect 32310 22208 32366 22264
rect 32218 21528 32274 21584
rect 32310 19352 32366 19408
rect 31758 16496 31814 16552
rect 31666 15272 31722 15328
rect 32494 21528 32550 21584
rect 32954 24520 33010 24576
rect 32862 22480 32918 22536
rect 32770 20848 32826 20904
rect 33046 22072 33102 22128
rect 32862 20304 32918 20360
rect 32770 19488 32826 19544
rect 31850 4020 31852 4040
rect 31852 4020 31904 4040
rect 31904 4020 31906 4040
rect 31390 3712 31446 3768
rect 31850 3984 31906 4020
rect 31666 3848 31722 3904
rect 31574 3440 31630 3496
rect 32310 15952 32366 16008
rect 34334 86284 34390 86320
rect 34334 86264 34336 86284
rect 34336 86264 34388 86284
rect 34388 86264 34390 86284
rect 33782 36080 33838 36136
rect 33322 22344 33378 22400
rect 33230 21936 33286 21992
rect 33138 20712 33194 20768
rect 33322 21120 33378 21176
rect 33322 20304 33378 20360
rect 33322 19896 33378 19952
rect 32954 14320 33010 14376
rect 33322 16904 33378 16960
rect 33322 14476 33378 14512
rect 33322 14456 33324 14476
rect 33324 14456 33376 14476
rect 33376 14456 33378 14476
rect 33690 23024 33746 23080
rect 33690 21936 33746 21992
rect 33874 23024 33930 23080
rect 33874 19760 33930 19816
rect 35346 118224 35402 118280
rect 35622 117408 35678 117464
rect 35530 116864 35586 116920
rect 34940 116442 34996 116444
rect 35020 116442 35076 116444
rect 35100 116442 35156 116444
rect 35180 116442 35236 116444
rect 34940 116390 34966 116442
rect 34966 116390 34996 116442
rect 35020 116390 35030 116442
rect 35030 116390 35076 116442
rect 35100 116390 35146 116442
rect 35146 116390 35156 116442
rect 35180 116390 35210 116442
rect 35210 116390 35236 116442
rect 34940 116388 34996 116390
rect 35020 116388 35076 116390
rect 35100 116388 35156 116390
rect 35180 116388 35236 116390
rect 35162 116048 35218 116104
rect 35346 116456 35402 116512
rect 35162 115504 35218 115560
rect 34940 115354 34996 115356
rect 35020 115354 35076 115356
rect 35100 115354 35156 115356
rect 35180 115354 35236 115356
rect 34940 115302 34966 115354
rect 34966 115302 34996 115354
rect 35020 115302 35030 115354
rect 35030 115302 35076 115354
rect 35100 115302 35146 115354
rect 35146 115302 35156 115354
rect 35180 115302 35210 115354
rect 35210 115302 35236 115354
rect 34940 115300 34996 115302
rect 35020 115300 35076 115302
rect 35100 115300 35156 115302
rect 35180 115300 35236 115302
rect 35346 115096 35402 115152
rect 34940 114266 34996 114268
rect 35020 114266 35076 114268
rect 35100 114266 35156 114268
rect 35180 114266 35236 114268
rect 34940 114214 34966 114266
rect 34966 114214 34996 114266
rect 35020 114214 35030 114266
rect 35030 114214 35076 114266
rect 35100 114214 35146 114266
rect 35146 114214 35156 114266
rect 35180 114214 35210 114266
rect 35210 114214 35236 114266
rect 34940 114212 34996 114214
rect 35020 114212 35076 114214
rect 35100 114212 35156 114214
rect 35180 114212 35236 114214
rect 34940 113178 34996 113180
rect 35020 113178 35076 113180
rect 35100 113178 35156 113180
rect 35180 113178 35236 113180
rect 34940 113126 34966 113178
rect 34966 113126 34996 113178
rect 35020 113126 35030 113178
rect 35030 113126 35076 113178
rect 35100 113126 35146 113178
rect 35146 113126 35156 113178
rect 35180 113126 35210 113178
rect 35210 113126 35236 113178
rect 34940 113124 34996 113126
rect 35020 113124 35076 113126
rect 35100 113124 35156 113126
rect 35180 113124 35236 113126
rect 34940 112090 34996 112092
rect 35020 112090 35076 112092
rect 35100 112090 35156 112092
rect 35180 112090 35236 112092
rect 34940 112038 34966 112090
rect 34966 112038 34996 112090
rect 35020 112038 35030 112090
rect 35030 112038 35076 112090
rect 35100 112038 35146 112090
rect 35146 112038 35156 112090
rect 35180 112038 35210 112090
rect 35210 112038 35236 112090
rect 34940 112036 34996 112038
rect 35020 112036 35076 112038
rect 35100 112036 35156 112038
rect 35180 112036 35236 112038
rect 34940 111002 34996 111004
rect 35020 111002 35076 111004
rect 35100 111002 35156 111004
rect 35180 111002 35236 111004
rect 34940 110950 34966 111002
rect 34966 110950 34996 111002
rect 35020 110950 35030 111002
rect 35030 110950 35076 111002
rect 35100 110950 35146 111002
rect 35146 110950 35156 111002
rect 35180 110950 35210 111002
rect 35210 110950 35236 111002
rect 34940 110948 34996 110950
rect 35020 110948 35076 110950
rect 35100 110948 35156 110950
rect 35180 110948 35236 110950
rect 34940 109914 34996 109916
rect 35020 109914 35076 109916
rect 35100 109914 35156 109916
rect 35180 109914 35236 109916
rect 34940 109862 34966 109914
rect 34966 109862 34996 109914
rect 35020 109862 35030 109914
rect 35030 109862 35076 109914
rect 35100 109862 35146 109914
rect 35146 109862 35156 109914
rect 35180 109862 35210 109914
rect 35210 109862 35236 109914
rect 34940 109860 34996 109862
rect 35020 109860 35076 109862
rect 35100 109860 35156 109862
rect 35180 109860 35236 109862
rect 34940 108826 34996 108828
rect 35020 108826 35076 108828
rect 35100 108826 35156 108828
rect 35180 108826 35236 108828
rect 34940 108774 34966 108826
rect 34966 108774 34996 108826
rect 35020 108774 35030 108826
rect 35030 108774 35076 108826
rect 35100 108774 35146 108826
rect 35146 108774 35156 108826
rect 35180 108774 35210 108826
rect 35210 108774 35236 108826
rect 34940 108772 34996 108774
rect 35020 108772 35076 108774
rect 35100 108772 35156 108774
rect 35180 108772 35236 108774
rect 34940 107738 34996 107740
rect 35020 107738 35076 107740
rect 35100 107738 35156 107740
rect 35180 107738 35236 107740
rect 34940 107686 34966 107738
rect 34966 107686 34996 107738
rect 35020 107686 35030 107738
rect 35030 107686 35076 107738
rect 35100 107686 35146 107738
rect 35146 107686 35156 107738
rect 35180 107686 35210 107738
rect 35210 107686 35236 107738
rect 34940 107684 34996 107686
rect 35020 107684 35076 107686
rect 35100 107684 35156 107686
rect 35180 107684 35236 107686
rect 34940 106650 34996 106652
rect 35020 106650 35076 106652
rect 35100 106650 35156 106652
rect 35180 106650 35236 106652
rect 34940 106598 34966 106650
rect 34966 106598 34996 106650
rect 35020 106598 35030 106650
rect 35030 106598 35076 106650
rect 35100 106598 35146 106650
rect 35146 106598 35156 106650
rect 35180 106598 35210 106650
rect 35210 106598 35236 106650
rect 34940 106596 34996 106598
rect 35020 106596 35076 106598
rect 35100 106596 35156 106598
rect 35180 106596 35236 106598
rect 34940 105562 34996 105564
rect 35020 105562 35076 105564
rect 35100 105562 35156 105564
rect 35180 105562 35236 105564
rect 34940 105510 34966 105562
rect 34966 105510 34996 105562
rect 35020 105510 35030 105562
rect 35030 105510 35076 105562
rect 35100 105510 35146 105562
rect 35146 105510 35156 105562
rect 35180 105510 35210 105562
rect 35210 105510 35236 105562
rect 34940 105508 34996 105510
rect 35020 105508 35076 105510
rect 35100 105508 35156 105510
rect 35180 105508 35236 105510
rect 34940 104474 34996 104476
rect 35020 104474 35076 104476
rect 35100 104474 35156 104476
rect 35180 104474 35236 104476
rect 34940 104422 34966 104474
rect 34966 104422 34996 104474
rect 35020 104422 35030 104474
rect 35030 104422 35076 104474
rect 35100 104422 35146 104474
rect 35146 104422 35156 104474
rect 35180 104422 35210 104474
rect 35210 104422 35236 104474
rect 34940 104420 34996 104422
rect 35020 104420 35076 104422
rect 35100 104420 35156 104422
rect 35180 104420 35236 104422
rect 34940 103386 34996 103388
rect 35020 103386 35076 103388
rect 35100 103386 35156 103388
rect 35180 103386 35236 103388
rect 34940 103334 34966 103386
rect 34966 103334 34996 103386
rect 35020 103334 35030 103386
rect 35030 103334 35076 103386
rect 35100 103334 35146 103386
rect 35146 103334 35156 103386
rect 35180 103334 35210 103386
rect 35210 103334 35236 103386
rect 34940 103332 34996 103334
rect 35020 103332 35076 103334
rect 35100 103332 35156 103334
rect 35180 103332 35236 103334
rect 34940 102298 34996 102300
rect 35020 102298 35076 102300
rect 35100 102298 35156 102300
rect 35180 102298 35236 102300
rect 34940 102246 34966 102298
rect 34966 102246 34996 102298
rect 35020 102246 35030 102298
rect 35030 102246 35076 102298
rect 35100 102246 35146 102298
rect 35146 102246 35156 102298
rect 35180 102246 35210 102298
rect 35210 102246 35236 102298
rect 34940 102244 34996 102246
rect 35020 102244 35076 102246
rect 35100 102244 35156 102246
rect 35180 102244 35236 102246
rect 34940 101210 34996 101212
rect 35020 101210 35076 101212
rect 35100 101210 35156 101212
rect 35180 101210 35236 101212
rect 34940 101158 34966 101210
rect 34966 101158 34996 101210
rect 35020 101158 35030 101210
rect 35030 101158 35076 101210
rect 35100 101158 35146 101210
rect 35146 101158 35156 101210
rect 35180 101158 35210 101210
rect 35210 101158 35236 101210
rect 34940 101156 34996 101158
rect 35020 101156 35076 101158
rect 35100 101156 35156 101158
rect 35180 101156 35236 101158
rect 34940 100122 34996 100124
rect 35020 100122 35076 100124
rect 35100 100122 35156 100124
rect 35180 100122 35236 100124
rect 34940 100070 34966 100122
rect 34966 100070 34996 100122
rect 35020 100070 35030 100122
rect 35030 100070 35076 100122
rect 35100 100070 35146 100122
rect 35146 100070 35156 100122
rect 35180 100070 35210 100122
rect 35210 100070 35236 100122
rect 34940 100068 34996 100070
rect 35020 100068 35076 100070
rect 35100 100068 35156 100070
rect 35180 100068 35236 100070
rect 34940 99034 34996 99036
rect 35020 99034 35076 99036
rect 35100 99034 35156 99036
rect 35180 99034 35236 99036
rect 34940 98982 34966 99034
rect 34966 98982 34996 99034
rect 35020 98982 35030 99034
rect 35030 98982 35076 99034
rect 35100 98982 35146 99034
rect 35146 98982 35156 99034
rect 35180 98982 35210 99034
rect 35210 98982 35236 99034
rect 34940 98980 34996 98982
rect 35020 98980 35076 98982
rect 35100 98980 35156 98982
rect 35180 98980 35236 98982
rect 35438 109656 35494 109712
rect 34940 97946 34996 97948
rect 35020 97946 35076 97948
rect 35100 97946 35156 97948
rect 35180 97946 35236 97948
rect 34940 97894 34966 97946
rect 34966 97894 34996 97946
rect 35020 97894 35030 97946
rect 35030 97894 35076 97946
rect 35100 97894 35146 97946
rect 35146 97894 35156 97946
rect 35180 97894 35210 97946
rect 35210 97894 35236 97946
rect 34940 97892 34996 97894
rect 35020 97892 35076 97894
rect 35100 97892 35156 97894
rect 35180 97892 35236 97894
rect 34940 96858 34996 96860
rect 35020 96858 35076 96860
rect 35100 96858 35156 96860
rect 35180 96858 35236 96860
rect 34940 96806 34966 96858
rect 34966 96806 34996 96858
rect 35020 96806 35030 96858
rect 35030 96806 35076 96858
rect 35100 96806 35146 96858
rect 35146 96806 35156 96858
rect 35180 96806 35210 96858
rect 35210 96806 35236 96858
rect 34940 96804 34996 96806
rect 35020 96804 35076 96806
rect 35100 96804 35156 96806
rect 35180 96804 35236 96806
rect 34940 95770 34996 95772
rect 35020 95770 35076 95772
rect 35100 95770 35156 95772
rect 35180 95770 35236 95772
rect 34940 95718 34966 95770
rect 34966 95718 34996 95770
rect 35020 95718 35030 95770
rect 35030 95718 35076 95770
rect 35100 95718 35146 95770
rect 35146 95718 35156 95770
rect 35180 95718 35210 95770
rect 35210 95718 35236 95770
rect 34940 95716 34996 95718
rect 35020 95716 35076 95718
rect 35100 95716 35156 95718
rect 35180 95716 35236 95718
rect 34940 94682 34996 94684
rect 35020 94682 35076 94684
rect 35100 94682 35156 94684
rect 35180 94682 35236 94684
rect 34940 94630 34966 94682
rect 34966 94630 34996 94682
rect 35020 94630 35030 94682
rect 35030 94630 35076 94682
rect 35100 94630 35146 94682
rect 35146 94630 35156 94682
rect 35180 94630 35210 94682
rect 35210 94630 35236 94682
rect 34940 94628 34996 94630
rect 35020 94628 35076 94630
rect 35100 94628 35156 94630
rect 35180 94628 35236 94630
rect 34940 93594 34996 93596
rect 35020 93594 35076 93596
rect 35100 93594 35156 93596
rect 35180 93594 35236 93596
rect 34940 93542 34966 93594
rect 34966 93542 34996 93594
rect 35020 93542 35030 93594
rect 35030 93542 35076 93594
rect 35100 93542 35146 93594
rect 35146 93542 35156 93594
rect 35180 93542 35210 93594
rect 35210 93542 35236 93594
rect 34940 93540 34996 93542
rect 35020 93540 35076 93542
rect 35100 93540 35156 93542
rect 35180 93540 35236 93542
rect 34940 92506 34996 92508
rect 35020 92506 35076 92508
rect 35100 92506 35156 92508
rect 35180 92506 35236 92508
rect 34940 92454 34966 92506
rect 34966 92454 34996 92506
rect 35020 92454 35030 92506
rect 35030 92454 35076 92506
rect 35100 92454 35146 92506
rect 35146 92454 35156 92506
rect 35180 92454 35210 92506
rect 35210 92454 35236 92506
rect 34940 92452 34996 92454
rect 35020 92452 35076 92454
rect 35100 92452 35156 92454
rect 35180 92452 35236 92454
rect 34940 91418 34996 91420
rect 35020 91418 35076 91420
rect 35100 91418 35156 91420
rect 35180 91418 35236 91420
rect 34940 91366 34966 91418
rect 34966 91366 34996 91418
rect 35020 91366 35030 91418
rect 35030 91366 35076 91418
rect 35100 91366 35146 91418
rect 35146 91366 35156 91418
rect 35180 91366 35210 91418
rect 35210 91366 35236 91418
rect 34940 91364 34996 91366
rect 35020 91364 35076 91366
rect 35100 91364 35156 91366
rect 35180 91364 35236 91366
rect 34940 90330 34996 90332
rect 35020 90330 35076 90332
rect 35100 90330 35156 90332
rect 35180 90330 35236 90332
rect 34940 90278 34966 90330
rect 34966 90278 34996 90330
rect 35020 90278 35030 90330
rect 35030 90278 35076 90330
rect 35100 90278 35146 90330
rect 35146 90278 35156 90330
rect 35180 90278 35210 90330
rect 35210 90278 35236 90330
rect 34940 90276 34996 90278
rect 35020 90276 35076 90278
rect 35100 90276 35156 90278
rect 35180 90276 35236 90278
rect 34940 89242 34996 89244
rect 35020 89242 35076 89244
rect 35100 89242 35156 89244
rect 35180 89242 35236 89244
rect 34940 89190 34966 89242
rect 34966 89190 34996 89242
rect 35020 89190 35030 89242
rect 35030 89190 35076 89242
rect 35100 89190 35146 89242
rect 35146 89190 35156 89242
rect 35180 89190 35210 89242
rect 35210 89190 35236 89242
rect 34940 89188 34996 89190
rect 35020 89188 35076 89190
rect 35100 89188 35156 89190
rect 35180 89188 35236 89190
rect 34940 88154 34996 88156
rect 35020 88154 35076 88156
rect 35100 88154 35156 88156
rect 35180 88154 35236 88156
rect 34940 88102 34966 88154
rect 34966 88102 34996 88154
rect 35020 88102 35030 88154
rect 35030 88102 35076 88154
rect 35100 88102 35146 88154
rect 35146 88102 35156 88154
rect 35180 88102 35210 88154
rect 35210 88102 35236 88154
rect 34940 88100 34996 88102
rect 35020 88100 35076 88102
rect 35100 88100 35156 88102
rect 35180 88100 35236 88102
rect 34794 87216 34850 87272
rect 34610 63960 34666 64016
rect 34242 25472 34298 25528
rect 34940 87066 34996 87068
rect 35020 87066 35076 87068
rect 35100 87066 35156 87068
rect 35180 87066 35236 87068
rect 34940 87014 34966 87066
rect 34966 87014 34996 87066
rect 35020 87014 35030 87066
rect 35030 87014 35076 87066
rect 35100 87014 35146 87066
rect 35146 87014 35156 87066
rect 35180 87014 35210 87066
rect 35210 87014 35236 87066
rect 34940 87012 34996 87014
rect 35020 87012 35076 87014
rect 35100 87012 35156 87014
rect 35180 87012 35236 87014
rect 34794 86944 34850 87000
rect 34940 85978 34996 85980
rect 35020 85978 35076 85980
rect 35100 85978 35156 85980
rect 35180 85978 35236 85980
rect 34940 85926 34966 85978
rect 34966 85926 34996 85978
rect 35020 85926 35030 85978
rect 35030 85926 35076 85978
rect 35100 85926 35146 85978
rect 35146 85926 35156 85978
rect 35180 85926 35210 85978
rect 35210 85926 35236 85978
rect 34940 85924 34996 85926
rect 35020 85924 35076 85926
rect 35100 85924 35156 85926
rect 35180 85924 35236 85926
rect 34940 84890 34996 84892
rect 35020 84890 35076 84892
rect 35100 84890 35156 84892
rect 35180 84890 35236 84892
rect 34940 84838 34966 84890
rect 34966 84838 34996 84890
rect 35020 84838 35030 84890
rect 35030 84838 35076 84890
rect 35100 84838 35146 84890
rect 35146 84838 35156 84890
rect 35180 84838 35210 84890
rect 35210 84838 35236 84890
rect 34940 84836 34996 84838
rect 35020 84836 35076 84838
rect 35100 84836 35156 84838
rect 35180 84836 35236 84838
rect 34940 83802 34996 83804
rect 35020 83802 35076 83804
rect 35100 83802 35156 83804
rect 35180 83802 35236 83804
rect 34940 83750 34966 83802
rect 34966 83750 34996 83802
rect 35020 83750 35030 83802
rect 35030 83750 35076 83802
rect 35100 83750 35146 83802
rect 35146 83750 35156 83802
rect 35180 83750 35210 83802
rect 35210 83750 35236 83802
rect 34940 83748 34996 83750
rect 35020 83748 35076 83750
rect 35100 83748 35156 83750
rect 35180 83748 35236 83750
rect 34940 82714 34996 82716
rect 35020 82714 35076 82716
rect 35100 82714 35156 82716
rect 35180 82714 35236 82716
rect 34940 82662 34966 82714
rect 34966 82662 34996 82714
rect 35020 82662 35030 82714
rect 35030 82662 35076 82714
rect 35100 82662 35146 82714
rect 35146 82662 35156 82714
rect 35180 82662 35210 82714
rect 35210 82662 35236 82714
rect 34940 82660 34996 82662
rect 35020 82660 35076 82662
rect 35100 82660 35156 82662
rect 35180 82660 35236 82662
rect 34940 81626 34996 81628
rect 35020 81626 35076 81628
rect 35100 81626 35156 81628
rect 35180 81626 35236 81628
rect 34940 81574 34966 81626
rect 34966 81574 34996 81626
rect 35020 81574 35030 81626
rect 35030 81574 35076 81626
rect 35100 81574 35146 81626
rect 35146 81574 35156 81626
rect 35180 81574 35210 81626
rect 35210 81574 35236 81626
rect 34940 81572 34996 81574
rect 35020 81572 35076 81574
rect 35100 81572 35156 81574
rect 35180 81572 35236 81574
rect 34940 80538 34996 80540
rect 35020 80538 35076 80540
rect 35100 80538 35156 80540
rect 35180 80538 35236 80540
rect 34940 80486 34966 80538
rect 34966 80486 34996 80538
rect 35020 80486 35030 80538
rect 35030 80486 35076 80538
rect 35100 80486 35146 80538
rect 35146 80486 35156 80538
rect 35180 80486 35210 80538
rect 35210 80486 35236 80538
rect 34940 80484 34996 80486
rect 35020 80484 35076 80486
rect 35100 80484 35156 80486
rect 35180 80484 35236 80486
rect 34940 79450 34996 79452
rect 35020 79450 35076 79452
rect 35100 79450 35156 79452
rect 35180 79450 35236 79452
rect 34940 79398 34966 79450
rect 34966 79398 34996 79450
rect 35020 79398 35030 79450
rect 35030 79398 35076 79450
rect 35100 79398 35146 79450
rect 35146 79398 35156 79450
rect 35180 79398 35210 79450
rect 35210 79398 35236 79450
rect 34940 79396 34996 79398
rect 35020 79396 35076 79398
rect 35100 79396 35156 79398
rect 35180 79396 35236 79398
rect 34940 78362 34996 78364
rect 35020 78362 35076 78364
rect 35100 78362 35156 78364
rect 35180 78362 35236 78364
rect 34940 78310 34966 78362
rect 34966 78310 34996 78362
rect 35020 78310 35030 78362
rect 35030 78310 35076 78362
rect 35100 78310 35146 78362
rect 35146 78310 35156 78362
rect 35180 78310 35210 78362
rect 35210 78310 35236 78362
rect 34940 78308 34996 78310
rect 35020 78308 35076 78310
rect 35100 78308 35156 78310
rect 35180 78308 35236 78310
rect 34940 77274 34996 77276
rect 35020 77274 35076 77276
rect 35100 77274 35156 77276
rect 35180 77274 35236 77276
rect 34940 77222 34966 77274
rect 34966 77222 34996 77274
rect 35020 77222 35030 77274
rect 35030 77222 35076 77274
rect 35100 77222 35146 77274
rect 35146 77222 35156 77274
rect 35180 77222 35210 77274
rect 35210 77222 35236 77274
rect 34940 77220 34996 77222
rect 35020 77220 35076 77222
rect 35100 77220 35156 77222
rect 35180 77220 35236 77222
rect 34940 76186 34996 76188
rect 35020 76186 35076 76188
rect 35100 76186 35156 76188
rect 35180 76186 35236 76188
rect 34940 76134 34966 76186
rect 34966 76134 34996 76186
rect 35020 76134 35030 76186
rect 35030 76134 35076 76186
rect 35100 76134 35146 76186
rect 35146 76134 35156 76186
rect 35180 76134 35210 76186
rect 35210 76134 35236 76186
rect 34940 76132 34996 76134
rect 35020 76132 35076 76134
rect 35100 76132 35156 76134
rect 35180 76132 35236 76134
rect 34940 75098 34996 75100
rect 35020 75098 35076 75100
rect 35100 75098 35156 75100
rect 35180 75098 35236 75100
rect 34940 75046 34966 75098
rect 34966 75046 34996 75098
rect 35020 75046 35030 75098
rect 35030 75046 35076 75098
rect 35100 75046 35146 75098
rect 35146 75046 35156 75098
rect 35180 75046 35210 75098
rect 35210 75046 35236 75098
rect 34940 75044 34996 75046
rect 35020 75044 35076 75046
rect 35100 75044 35156 75046
rect 35180 75044 35236 75046
rect 34940 74010 34996 74012
rect 35020 74010 35076 74012
rect 35100 74010 35156 74012
rect 35180 74010 35236 74012
rect 34940 73958 34966 74010
rect 34966 73958 34996 74010
rect 35020 73958 35030 74010
rect 35030 73958 35076 74010
rect 35100 73958 35146 74010
rect 35146 73958 35156 74010
rect 35180 73958 35210 74010
rect 35210 73958 35236 74010
rect 34940 73956 34996 73958
rect 35020 73956 35076 73958
rect 35100 73956 35156 73958
rect 35180 73956 35236 73958
rect 34940 72922 34996 72924
rect 35020 72922 35076 72924
rect 35100 72922 35156 72924
rect 35180 72922 35236 72924
rect 34940 72870 34966 72922
rect 34966 72870 34996 72922
rect 35020 72870 35030 72922
rect 35030 72870 35076 72922
rect 35100 72870 35146 72922
rect 35146 72870 35156 72922
rect 35180 72870 35210 72922
rect 35210 72870 35236 72922
rect 34940 72868 34996 72870
rect 35020 72868 35076 72870
rect 35100 72868 35156 72870
rect 35180 72868 35236 72870
rect 34940 71834 34996 71836
rect 35020 71834 35076 71836
rect 35100 71834 35156 71836
rect 35180 71834 35236 71836
rect 34940 71782 34966 71834
rect 34966 71782 34996 71834
rect 35020 71782 35030 71834
rect 35030 71782 35076 71834
rect 35100 71782 35146 71834
rect 35146 71782 35156 71834
rect 35180 71782 35210 71834
rect 35210 71782 35236 71834
rect 34940 71780 34996 71782
rect 35020 71780 35076 71782
rect 35100 71780 35156 71782
rect 35180 71780 35236 71782
rect 34940 70746 34996 70748
rect 35020 70746 35076 70748
rect 35100 70746 35156 70748
rect 35180 70746 35236 70748
rect 34940 70694 34966 70746
rect 34966 70694 34996 70746
rect 35020 70694 35030 70746
rect 35030 70694 35076 70746
rect 35100 70694 35146 70746
rect 35146 70694 35156 70746
rect 35180 70694 35210 70746
rect 35210 70694 35236 70746
rect 34940 70692 34996 70694
rect 35020 70692 35076 70694
rect 35100 70692 35156 70694
rect 35180 70692 35236 70694
rect 34940 69658 34996 69660
rect 35020 69658 35076 69660
rect 35100 69658 35156 69660
rect 35180 69658 35236 69660
rect 34940 69606 34966 69658
rect 34966 69606 34996 69658
rect 35020 69606 35030 69658
rect 35030 69606 35076 69658
rect 35100 69606 35146 69658
rect 35146 69606 35156 69658
rect 35180 69606 35210 69658
rect 35210 69606 35236 69658
rect 34940 69604 34996 69606
rect 35020 69604 35076 69606
rect 35100 69604 35156 69606
rect 35180 69604 35236 69606
rect 34940 68570 34996 68572
rect 35020 68570 35076 68572
rect 35100 68570 35156 68572
rect 35180 68570 35236 68572
rect 34940 68518 34966 68570
rect 34966 68518 34996 68570
rect 35020 68518 35030 68570
rect 35030 68518 35076 68570
rect 35100 68518 35146 68570
rect 35146 68518 35156 68570
rect 35180 68518 35210 68570
rect 35210 68518 35236 68570
rect 34940 68516 34996 68518
rect 35020 68516 35076 68518
rect 35100 68516 35156 68518
rect 35180 68516 35236 68518
rect 34940 67482 34996 67484
rect 35020 67482 35076 67484
rect 35100 67482 35156 67484
rect 35180 67482 35236 67484
rect 34940 67430 34966 67482
rect 34966 67430 34996 67482
rect 35020 67430 35030 67482
rect 35030 67430 35076 67482
rect 35100 67430 35146 67482
rect 35146 67430 35156 67482
rect 35180 67430 35210 67482
rect 35210 67430 35236 67482
rect 34940 67428 34996 67430
rect 35020 67428 35076 67430
rect 35100 67428 35156 67430
rect 35180 67428 35236 67430
rect 34794 66816 34850 66872
rect 34940 66394 34996 66396
rect 35020 66394 35076 66396
rect 35100 66394 35156 66396
rect 35180 66394 35236 66396
rect 34940 66342 34966 66394
rect 34966 66342 34996 66394
rect 35020 66342 35030 66394
rect 35030 66342 35076 66394
rect 35100 66342 35146 66394
rect 35146 66342 35156 66394
rect 35180 66342 35210 66394
rect 35210 66342 35236 66394
rect 34940 66340 34996 66342
rect 35020 66340 35076 66342
rect 35100 66340 35156 66342
rect 35180 66340 35236 66342
rect 35070 65456 35126 65512
rect 34940 65306 34996 65308
rect 35020 65306 35076 65308
rect 35100 65306 35156 65308
rect 35180 65306 35236 65308
rect 34940 65254 34966 65306
rect 34966 65254 34996 65306
rect 35020 65254 35030 65306
rect 35030 65254 35076 65306
rect 35100 65254 35146 65306
rect 35146 65254 35156 65306
rect 35180 65254 35210 65306
rect 35210 65254 35236 65306
rect 34940 65252 34996 65254
rect 35020 65252 35076 65254
rect 35100 65252 35156 65254
rect 35180 65252 35236 65254
rect 34794 65048 34850 65104
rect 35070 64912 35126 64968
rect 35346 68448 35402 68504
rect 35346 66408 35402 66464
rect 35806 110064 35862 110120
rect 35254 64776 35310 64832
rect 35438 64640 35494 64696
rect 35254 64504 35310 64560
rect 34886 64368 34942 64424
rect 34940 64218 34996 64220
rect 35020 64218 35076 64220
rect 35100 64218 35156 64220
rect 35180 64218 35236 64220
rect 34940 64166 34966 64218
rect 34966 64166 34996 64218
rect 35020 64166 35030 64218
rect 35030 64166 35076 64218
rect 35100 64166 35146 64218
rect 35146 64166 35156 64218
rect 35180 64166 35210 64218
rect 35210 64166 35236 64218
rect 34940 64164 34996 64166
rect 35020 64164 35076 64166
rect 35100 64164 35156 64166
rect 35180 64164 35236 64166
rect 34794 63280 34850 63336
rect 35162 63824 35218 63880
rect 34940 63130 34996 63132
rect 35020 63130 35076 63132
rect 35100 63130 35156 63132
rect 35180 63130 35236 63132
rect 34940 63078 34966 63130
rect 34966 63078 34996 63130
rect 35020 63078 35030 63130
rect 35030 63078 35076 63130
rect 35100 63078 35146 63130
rect 35146 63078 35156 63130
rect 35180 63078 35210 63130
rect 35210 63078 35236 63130
rect 34940 63076 34996 63078
rect 35020 63076 35076 63078
rect 35100 63076 35156 63078
rect 35180 63076 35236 63078
rect 34940 62042 34996 62044
rect 35020 62042 35076 62044
rect 35100 62042 35156 62044
rect 35180 62042 35236 62044
rect 34940 61990 34966 62042
rect 34966 61990 34996 62042
rect 35020 61990 35030 62042
rect 35030 61990 35076 62042
rect 35100 61990 35146 62042
rect 35146 61990 35156 62042
rect 35180 61990 35210 62042
rect 35210 61990 35236 62042
rect 34940 61988 34996 61990
rect 35020 61988 35076 61990
rect 35100 61988 35156 61990
rect 35180 61988 35236 61990
rect 34886 61376 34942 61432
rect 34940 60954 34996 60956
rect 35020 60954 35076 60956
rect 35100 60954 35156 60956
rect 35180 60954 35236 60956
rect 34940 60902 34966 60954
rect 34966 60902 34996 60954
rect 35020 60902 35030 60954
rect 35030 60902 35076 60954
rect 35100 60902 35146 60954
rect 35146 60902 35156 60954
rect 35180 60902 35210 60954
rect 35210 60902 35236 60954
rect 34940 60900 34996 60902
rect 35020 60900 35076 60902
rect 35100 60900 35156 60902
rect 35180 60900 35236 60902
rect 35346 64096 35402 64152
rect 35530 63824 35586 63880
rect 35162 60560 35218 60616
rect 35162 60172 35218 60208
rect 35162 60152 35164 60172
rect 35164 60152 35216 60172
rect 35216 60152 35218 60172
rect 34940 59866 34996 59868
rect 35020 59866 35076 59868
rect 35100 59866 35156 59868
rect 35180 59866 35236 59868
rect 34940 59814 34966 59866
rect 34966 59814 34996 59866
rect 35020 59814 35030 59866
rect 35030 59814 35076 59866
rect 35100 59814 35146 59866
rect 35146 59814 35156 59866
rect 35180 59814 35210 59866
rect 35210 59814 35236 59866
rect 34940 59812 34996 59814
rect 35020 59812 35076 59814
rect 35100 59812 35156 59814
rect 35180 59812 35236 59814
rect 34794 59608 34850 59664
rect 35254 59472 35310 59528
rect 34940 58778 34996 58780
rect 35020 58778 35076 58780
rect 35100 58778 35156 58780
rect 35180 58778 35236 58780
rect 34940 58726 34966 58778
rect 34966 58726 34996 58778
rect 35020 58726 35030 58778
rect 35030 58726 35076 58778
rect 35100 58726 35146 58778
rect 35146 58726 35156 58778
rect 35180 58726 35210 58778
rect 35210 58726 35236 58778
rect 34940 58724 34996 58726
rect 35020 58724 35076 58726
rect 35100 58724 35156 58726
rect 35180 58724 35236 58726
rect 34940 57690 34996 57692
rect 35020 57690 35076 57692
rect 35100 57690 35156 57692
rect 35180 57690 35236 57692
rect 34940 57638 34966 57690
rect 34966 57638 34996 57690
rect 35020 57638 35030 57690
rect 35030 57638 35076 57690
rect 35100 57638 35146 57690
rect 35146 57638 35156 57690
rect 35180 57638 35210 57690
rect 35210 57638 35236 57690
rect 34940 57636 34996 57638
rect 35020 57636 35076 57638
rect 35100 57636 35156 57638
rect 35180 57636 35236 57638
rect 34940 56602 34996 56604
rect 35020 56602 35076 56604
rect 35100 56602 35156 56604
rect 35180 56602 35236 56604
rect 34940 56550 34966 56602
rect 34966 56550 34996 56602
rect 35020 56550 35030 56602
rect 35030 56550 35076 56602
rect 35100 56550 35146 56602
rect 35146 56550 35156 56602
rect 35180 56550 35210 56602
rect 35210 56550 35236 56602
rect 34940 56548 34996 56550
rect 35020 56548 35076 56550
rect 35100 56548 35156 56550
rect 35180 56548 35236 56550
rect 34940 55514 34996 55516
rect 35020 55514 35076 55516
rect 35100 55514 35156 55516
rect 35180 55514 35236 55516
rect 34940 55462 34966 55514
rect 34966 55462 34996 55514
rect 35020 55462 35030 55514
rect 35030 55462 35076 55514
rect 35100 55462 35146 55514
rect 35146 55462 35156 55514
rect 35180 55462 35210 55514
rect 35210 55462 35236 55514
rect 34940 55460 34996 55462
rect 35020 55460 35076 55462
rect 35100 55460 35156 55462
rect 35180 55460 35236 55462
rect 34940 54426 34996 54428
rect 35020 54426 35076 54428
rect 35100 54426 35156 54428
rect 35180 54426 35236 54428
rect 34940 54374 34966 54426
rect 34966 54374 34996 54426
rect 35020 54374 35030 54426
rect 35030 54374 35076 54426
rect 35100 54374 35146 54426
rect 35146 54374 35156 54426
rect 35180 54374 35210 54426
rect 35210 54374 35236 54426
rect 34940 54372 34996 54374
rect 35020 54372 35076 54374
rect 35100 54372 35156 54374
rect 35180 54372 35236 54374
rect 34940 53338 34996 53340
rect 35020 53338 35076 53340
rect 35100 53338 35156 53340
rect 35180 53338 35236 53340
rect 34940 53286 34966 53338
rect 34966 53286 34996 53338
rect 35020 53286 35030 53338
rect 35030 53286 35076 53338
rect 35100 53286 35146 53338
rect 35146 53286 35156 53338
rect 35180 53286 35210 53338
rect 35210 53286 35236 53338
rect 34940 53284 34996 53286
rect 35020 53284 35076 53286
rect 35100 53284 35156 53286
rect 35180 53284 35236 53286
rect 34940 52250 34996 52252
rect 35020 52250 35076 52252
rect 35100 52250 35156 52252
rect 35180 52250 35236 52252
rect 34940 52198 34966 52250
rect 34966 52198 34996 52250
rect 35020 52198 35030 52250
rect 35030 52198 35076 52250
rect 35100 52198 35146 52250
rect 35146 52198 35156 52250
rect 35180 52198 35210 52250
rect 35210 52198 35236 52250
rect 34940 52196 34996 52198
rect 35020 52196 35076 52198
rect 35100 52196 35156 52198
rect 35180 52196 35236 52198
rect 34940 51162 34996 51164
rect 35020 51162 35076 51164
rect 35100 51162 35156 51164
rect 35180 51162 35236 51164
rect 34940 51110 34966 51162
rect 34966 51110 34996 51162
rect 35020 51110 35030 51162
rect 35030 51110 35076 51162
rect 35100 51110 35146 51162
rect 35146 51110 35156 51162
rect 35180 51110 35210 51162
rect 35210 51110 35236 51162
rect 34940 51108 34996 51110
rect 35020 51108 35076 51110
rect 35100 51108 35156 51110
rect 35180 51108 35236 51110
rect 34940 50074 34996 50076
rect 35020 50074 35076 50076
rect 35100 50074 35156 50076
rect 35180 50074 35236 50076
rect 34940 50022 34966 50074
rect 34966 50022 34996 50074
rect 35020 50022 35030 50074
rect 35030 50022 35076 50074
rect 35100 50022 35146 50074
rect 35146 50022 35156 50074
rect 35180 50022 35210 50074
rect 35210 50022 35236 50074
rect 34940 50020 34996 50022
rect 35020 50020 35076 50022
rect 35100 50020 35156 50022
rect 35180 50020 35236 50022
rect 34940 48986 34996 48988
rect 35020 48986 35076 48988
rect 35100 48986 35156 48988
rect 35180 48986 35236 48988
rect 34940 48934 34966 48986
rect 34966 48934 34996 48986
rect 35020 48934 35030 48986
rect 35030 48934 35076 48986
rect 35100 48934 35146 48986
rect 35146 48934 35156 48986
rect 35180 48934 35210 48986
rect 35210 48934 35236 48986
rect 34940 48932 34996 48934
rect 35020 48932 35076 48934
rect 35100 48932 35156 48934
rect 35180 48932 35236 48934
rect 34940 47898 34996 47900
rect 35020 47898 35076 47900
rect 35100 47898 35156 47900
rect 35180 47898 35236 47900
rect 34940 47846 34966 47898
rect 34966 47846 34996 47898
rect 35020 47846 35030 47898
rect 35030 47846 35076 47898
rect 35100 47846 35146 47898
rect 35146 47846 35156 47898
rect 35180 47846 35210 47898
rect 35210 47846 35236 47898
rect 34940 47844 34996 47846
rect 35020 47844 35076 47846
rect 35100 47844 35156 47846
rect 35180 47844 35236 47846
rect 34940 46810 34996 46812
rect 35020 46810 35076 46812
rect 35100 46810 35156 46812
rect 35180 46810 35236 46812
rect 34940 46758 34966 46810
rect 34966 46758 34996 46810
rect 35020 46758 35030 46810
rect 35030 46758 35076 46810
rect 35100 46758 35146 46810
rect 35146 46758 35156 46810
rect 35180 46758 35210 46810
rect 35210 46758 35236 46810
rect 34940 46756 34996 46758
rect 35020 46756 35076 46758
rect 35100 46756 35156 46758
rect 35180 46756 35236 46758
rect 34940 45722 34996 45724
rect 35020 45722 35076 45724
rect 35100 45722 35156 45724
rect 35180 45722 35236 45724
rect 34940 45670 34966 45722
rect 34966 45670 34996 45722
rect 35020 45670 35030 45722
rect 35030 45670 35076 45722
rect 35100 45670 35146 45722
rect 35146 45670 35156 45722
rect 35180 45670 35210 45722
rect 35210 45670 35236 45722
rect 34940 45668 34996 45670
rect 35020 45668 35076 45670
rect 35100 45668 35156 45670
rect 35180 45668 35236 45670
rect 34940 44634 34996 44636
rect 35020 44634 35076 44636
rect 35100 44634 35156 44636
rect 35180 44634 35236 44636
rect 34940 44582 34966 44634
rect 34966 44582 34996 44634
rect 35020 44582 35030 44634
rect 35030 44582 35076 44634
rect 35100 44582 35146 44634
rect 35146 44582 35156 44634
rect 35180 44582 35210 44634
rect 35210 44582 35236 44634
rect 34940 44580 34996 44582
rect 35020 44580 35076 44582
rect 35100 44580 35156 44582
rect 35180 44580 35236 44582
rect 35806 68176 35862 68232
rect 35714 64504 35770 64560
rect 35806 63572 35862 63608
rect 35806 63552 35808 63572
rect 35808 63552 35860 63572
rect 35860 63552 35862 63572
rect 35806 63436 35862 63472
rect 35806 63416 35808 63436
rect 35808 63416 35860 63436
rect 35860 63416 35862 63436
rect 35714 62736 35770 62792
rect 35346 46688 35402 46744
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 34702 36352 34758 36408
rect 34610 26424 34666 26480
rect 34518 25200 34574 25256
rect 34334 24520 34390 24576
rect 34150 22208 34206 22264
rect 34058 21800 34114 21856
rect 34150 21120 34206 21176
rect 34426 22888 34482 22944
rect 34334 22072 34390 22128
rect 34426 21936 34482 21992
rect 34334 21392 34390 21448
rect 34058 19488 34114 19544
rect 33966 17040 34022 17096
rect 33966 16904 34022 16960
rect 34150 16532 34152 16552
rect 34152 16532 34204 16552
rect 34204 16532 34206 16552
rect 34150 16496 34206 16532
rect 33966 15544 34022 15600
rect 33966 15308 33968 15328
rect 33968 15308 34020 15328
rect 34020 15308 34022 15328
rect 33966 15272 34022 15308
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34886 36080 34942 36136
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 35806 60968 35862 61024
rect 35806 59200 35862 59256
rect 36266 67632 36322 67688
rect 36082 64368 36138 64424
rect 36542 116748 36598 116784
rect 36542 116728 36544 116748
rect 36544 116728 36596 116748
rect 36596 116728 36598 116748
rect 36910 117816 36966 117872
rect 36542 114688 36598 114744
rect 37186 119176 37242 119232
rect 37370 115096 37426 115152
rect 37186 113328 37242 113384
rect 37094 112512 37150 112568
rect 37094 111968 37150 112024
rect 37094 111152 37150 111208
rect 37094 110220 37150 110256
rect 37094 110200 37096 110220
rect 37096 110200 37148 110220
rect 37148 110200 37150 110220
rect 37094 109792 37150 109848
rect 36818 87216 36874 87272
rect 37094 108840 37150 108896
rect 37186 108044 37242 108080
rect 37186 108024 37188 108044
rect 37188 108024 37240 108044
rect 37240 108024 37242 108044
rect 37186 107480 37242 107536
rect 37186 106664 37242 106720
rect 37186 105712 37242 105768
rect 37186 104896 37242 104952
rect 37186 104352 37242 104408
rect 37186 103536 37242 103592
rect 37186 102604 37242 102640
rect 37186 102584 37188 102604
rect 37188 102584 37240 102604
rect 37240 102584 37242 102604
rect 37186 102176 37242 102232
rect 37186 101224 37242 101280
rect 37186 100428 37242 100464
rect 37186 100408 37188 100428
rect 37188 100408 37240 100428
rect 37240 100408 37242 100428
rect 37278 99864 37334 99920
rect 37186 99456 37242 99512
rect 37094 98096 37150 98152
rect 37094 97280 37150 97336
rect 37094 96736 37150 96792
rect 36726 87080 36782 87136
rect 36910 87080 36966 87136
rect 36818 86944 36874 87000
rect 36726 69964 36782 70000
rect 36726 69944 36728 69964
rect 36728 69944 36780 69964
rect 36780 69944 36782 69964
rect 37186 95920 37242 95976
rect 37186 94988 37242 95024
rect 37186 94968 37188 94988
rect 37188 94968 37240 94988
rect 37240 94968 37242 94988
rect 37186 94560 37242 94616
rect 37922 114280 37978 114336
rect 37922 113736 37978 113792
rect 37922 112920 37978 112976
rect 37830 111560 37886 111616
rect 37830 110644 37832 110664
rect 37832 110644 37884 110664
rect 37884 110644 37886 110664
rect 37830 110608 37886 110644
rect 37830 109384 37886 109440
rect 37830 108468 37832 108488
rect 37832 108468 37884 108488
rect 37884 108468 37886 108488
rect 37830 108432 37886 108468
rect 37922 107072 37978 107128
rect 37922 106120 37978 106176
rect 37922 105304 37978 105360
rect 37922 103944 37978 104000
rect 37922 103012 37978 103048
rect 37922 102992 37924 103012
rect 37924 102992 37976 103012
rect 37976 102992 37978 103012
rect 37922 101768 37978 101824
rect 37922 100836 37978 100872
rect 37922 100816 37924 100836
rect 37924 100816 37976 100836
rect 37976 100816 37978 100836
rect 37922 99048 37978 99104
rect 37922 98676 37924 98696
rect 37924 98676 37976 98696
rect 37976 98676 37978 98696
rect 37922 98640 37978 98676
rect 37830 97688 37886 97744
rect 37922 96328 37978 96384
rect 37922 95396 37978 95432
rect 37922 95376 37924 95396
rect 37924 95376 37976 95396
rect 37976 95376 37978 95396
rect 37186 93608 37242 93664
rect 37278 93236 37280 93256
rect 37280 93236 37332 93256
rect 37332 93236 37334 93256
rect 37278 93200 37334 93236
rect 37278 92248 37334 92304
rect 37186 91840 37242 91896
rect 37186 91060 37188 91080
rect 37188 91060 37240 91080
rect 37240 91060 37242 91080
rect 37186 91024 37242 91060
rect 37278 90072 37334 90128
rect 37186 89664 37242 89720
rect 37278 88712 37334 88768
rect 37278 87896 37334 87952
rect 37186 87372 37242 87408
rect 37186 87352 37188 87372
rect 37188 87352 37240 87372
rect 37240 87352 37242 87372
rect 37278 86536 37334 86592
rect 37278 85620 37280 85640
rect 37280 85620 37332 85640
rect 37332 85620 37334 85640
rect 37278 85584 37334 85620
rect 37278 84768 37334 84824
rect 37186 84224 37242 84280
rect 37922 94152 37978 94208
rect 37922 92792 37978 92848
rect 37278 83444 37280 83464
rect 37280 83444 37332 83464
rect 37332 83444 37334 83464
rect 37278 83408 37334 83444
rect 37278 82456 37334 82512
rect 37186 82048 37242 82104
rect 37278 81096 37334 81152
rect 37278 80280 37334 80336
rect 37186 79756 37242 79792
rect 37186 79736 37188 79756
rect 37188 79736 37240 79756
rect 37240 79736 37242 79756
rect 37278 78920 37334 78976
rect 37278 78004 37280 78024
rect 37280 78004 37332 78024
rect 37332 78004 37334 78024
rect 37278 77968 37334 78004
rect 37278 77152 37334 77208
rect 37278 75828 37280 75848
rect 37280 75828 37332 75848
rect 37332 75828 37334 75848
rect 37278 75792 37334 75828
rect 37186 75248 37242 75304
rect 37278 74840 37334 74896
rect 37186 74432 37242 74488
rect 37278 73480 37334 73536
rect 37278 72664 37334 72720
rect 37186 72140 37242 72176
rect 37186 72120 37188 72140
rect 37188 72120 37240 72140
rect 37240 72120 37242 72140
rect 36910 69808 36966 69864
rect 36082 63008 36138 63064
rect 36358 64368 36414 64424
rect 36266 62348 36322 62384
rect 36266 62328 36268 62348
rect 36268 62328 36320 62348
rect 36320 62328 36322 62348
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34702 25200 34758 25256
rect 34610 23432 34666 23488
rect 34610 23024 34666 23080
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34886 25880 34942 25936
rect 34978 25336 35034 25392
rect 34886 25200 34942 25256
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 35162 24826 35218 24882
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 34518 20440 34574 20496
rect 34518 19932 34520 19952
rect 34520 19932 34572 19952
rect 34572 19932 34574 19952
rect 34518 19896 34574 19932
rect 35070 22480 35126 22536
rect 35070 22092 35126 22128
rect 35070 22072 35072 22092
rect 35072 22072 35124 22092
rect 35124 22072 35126 22092
rect 34886 21936 34942 21992
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 35162 20848 35218 20904
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 34886 20304 34942 20360
rect 34334 16904 34390 16960
rect 34334 15952 34390 16008
rect 34334 15136 34390 15192
rect 34334 14476 34390 14512
rect 34334 14456 34336 14476
rect 34336 14456 34388 14476
rect 34388 14456 34390 14476
rect 34886 19760 34942 19816
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34886 19352 34942 19408
rect 35070 18672 35126 18728
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34886 18264 34942 18320
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 35346 21120 35402 21176
rect 35806 46688 35862 46744
rect 35714 36760 35770 36816
rect 35530 36352 35586 36408
rect 35438 20848 35494 20904
rect 35714 36488 35770 36544
rect 35622 23432 35678 23488
rect 35622 21936 35678 21992
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 35438 15544 35494 15600
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 35898 21936 35954 21992
rect 35898 20032 35954 20088
rect 35622 15408 35678 15464
rect 35530 14320 35586 14376
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34610 4120 34666 4176
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34610 2352 34666 2408
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 35530 3712 35586 3768
rect 35622 1944 35678 2000
rect 35898 3304 35954 3360
rect 36266 58520 36322 58576
rect 36450 63688 36506 63744
rect 36726 63552 36782 63608
rect 36450 58520 36506 58576
rect 36174 16496 36230 16552
rect 35806 992 35862 1048
rect 36726 62212 36782 62248
rect 36726 62192 36728 62212
rect 36728 62192 36780 62212
rect 36780 62192 36782 62212
rect 36726 61920 36782 61976
rect 37922 91432 37978 91488
rect 37922 90480 37978 90536
rect 37922 89120 37978 89176
rect 37922 88304 37978 88360
rect 37922 86944 37978 87000
rect 37922 85992 37978 86048
rect 37922 85176 37978 85232
rect 37922 83816 37978 83872
rect 37922 82864 37978 82920
rect 37922 81504 37978 81560
rect 37922 80688 37978 80744
rect 37462 71304 37518 71360
rect 37370 70760 37426 70816
rect 37462 69536 37518 69592
rect 37462 69400 37518 69456
rect 37370 68992 37426 69048
rect 37186 68856 37242 68912
rect 37002 68584 37058 68640
rect 36910 64776 36966 64832
rect 36910 63960 36966 64016
rect 36818 58792 36874 58848
rect 36726 58248 36782 58304
rect 37370 68468 37426 68504
rect 37370 68448 37372 68468
rect 37372 68448 37424 68468
rect 37424 68448 37426 68468
rect 36726 53352 36782 53408
rect 36450 4528 36506 4584
rect 36082 1400 36138 1456
rect 2870 312 2926 368
rect 36910 2760 36966 2816
rect 37278 63824 37334 63880
rect 37278 62908 37280 62928
rect 37280 62908 37332 62928
rect 37332 62908 37334 62928
rect 37278 62872 37334 62908
rect 37922 79328 37978 79384
rect 37922 78376 37978 78432
rect 37922 77560 37978 77616
rect 37922 76608 37978 76664
rect 38014 76200 38070 76256
rect 37922 74024 37978 74080
rect 37922 73072 37978 73128
rect 37646 64912 37702 64968
rect 37554 64640 37610 64696
rect 37646 63552 37702 63608
rect 37554 63452 37556 63472
rect 37556 63452 37608 63472
rect 37608 63452 37610 63472
rect 37554 63416 37610 63452
rect 37922 70352 37978 70408
rect 38106 70352 38162 70408
rect 37462 62192 37518 62248
rect 37186 57840 37242 57896
rect 37462 57432 37518 57488
rect 37462 56072 37518 56128
rect 37186 55664 37242 55720
rect 37186 54304 37242 54360
rect 37186 53760 37242 53816
rect 37278 52980 37280 53000
rect 37280 52980 37332 53000
rect 37332 52980 37334 53000
rect 37278 52944 37334 52980
rect 37186 51584 37242 51640
rect 37462 54712 37518 54768
rect 37462 51992 37518 52048
rect 37462 50632 37518 50688
rect 37370 49408 37426 49464
rect 37278 48864 37334 48920
rect 37370 48048 37426 48104
rect 37278 47540 37280 47560
rect 37280 47540 37332 47560
rect 37332 47540 37334 47560
rect 37278 47504 37334 47540
rect 37462 46688 37518 46744
rect 37186 46144 37242 46200
rect 37462 45364 37464 45384
rect 37464 45364 37516 45384
rect 37516 45364 37518 45384
rect 37462 45328 37518 45364
rect 37186 43968 37242 44024
rect 37186 43560 37242 43616
rect 37370 42608 37426 42664
rect 37278 42200 37334 42256
rect 37186 41248 37242 41304
rect 37278 40840 37334 40896
rect 37462 39924 37464 39944
rect 37464 39924 37516 39944
rect 37516 39924 37518 39944
rect 37462 39888 37518 39924
rect 37462 38664 37518 38720
rect 37186 38120 37242 38176
rect 37370 37324 37426 37360
rect 37370 37304 37372 37324
rect 37372 37304 37424 37324
rect 37424 37304 37426 37324
rect 37278 36760 37334 36816
rect 37370 35944 37426 36000
rect 37278 35400 37334 35456
rect 37462 34584 37518 34640
rect 37462 33224 37518 33280
rect 37186 32816 37242 32872
rect 37370 31884 37426 31920
rect 37370 31864 37372 31884
rect 37372 31864 37424 31884
rect 37424 31864 37426 31884
rect 37278 31456 37334 31512
rect 37370 30504 37426 30560
rect 37278 30132 37280 30152
rect 37280 30132 37332 30152
rect 37332 30132 37334 30152
rect 37278 30096 37334 30132
rect 37186 27376 37242 27432
rect 37462 29144 37518 29200
rect 37462 27956 37464 27976
rect 37464 27956 37516 27976
rect 37516 27956 37518 27976
rect 37462 27920 37518 27956
rect 37370 26560 37426 26616
rect 37278 26016 37334 26072
rect 37186 25200 37242 25256
rect 37278 24792 37334 24848
rect 37370 23840 37426 23896
rect 37278 23432 37334 23488
rect 37278 22516 37280 22536
rect 37280 22516 37332 22536
rect 37332 22516 37334 22536
rect 37278 22480 37334 22516
rect 37278 21120 37334 21176
rect 37186 20712 37242 20768
rect 37186 19760 37242 19816
rect 37462 22072 37518 22128
rect 37278 19352 37334 19408
rect 37186 18400 37242 18456
rect 37278 17992 37334 18048
rect 37278 17176 37334 17232
rect 37278 15816 37334 15872
rect 37186 15272 37242 15328
rect 37186 14476 37242 14512
rect 37186 14456 37188 14476
rect 37188 14456 37240 14476
rect 37240 14456 37242 14476
rect 37278 14048 37334 14104
rect 37186 13504 37242 13560
rect 37278 12724 37280 12744
rect 37280 12724 37332 12744
rect 37332 12724 37334 12744
rect 37278 12688 37334 12724
rect 37278 11736 37334 11792
rect 37186 11328 37242 11384
rect 37278 10376 37334 10432
rect 37278 9560 37334 9616
rect 37186 9036 37242 9072
rect 37186 9016 37188 9036
rect 37188 9016 37240 9036
rect 37240 9016 37242 9036
rect 37186 8200 37242 8256
rect 37278 7284 37280 7304
rect 37280 7284 37332 7304
rect 37332 7284 37334 7304
rect 37278 7248 37334 7284
rect 37186 6860 37242 6896
rect 37186 6840 37188 6860
rect 37188 6840 37240 6860
rect 37240 6840 37242 6860
rect 37278 5888 37334 5944
rect 37186 5480 37242 5536
rect 36726 584 36782 640
rect 38290 68584 38346 68640
rect 38198 65864 38254 65920
rect 38382 67224 38438 67280
rect 37830 59472 37886 59528
rect 37922 56888 37978 56944
rect 37922 56480 37978 56536
rect 37922 55156 37924 55176
rect 37924 55156 37976 55176
rect 37976 55156 37978 55176
rect 37922 55120 37978 55156
rect 37922 52536 37978 52592
rect 37922 51176 37978 51232
rect 37922 50224 37978 50280
rect 37922 49816 37978 49872
rect 37922 48456 37978 48512
rect 37922 47096 37978 47152
rect 37922 45736 37978 45792
rect 37922 44920 37978 44976
rect 37922 44376 37978 44432
rect 37922 43016 37978 43072
rect 37922 41792 37978 41848
rect 37922 40432 37978 40488
rect 37922 39480 37978 39536
rect 37922 39072 37978 39128
rect 37922 37748 37924 37768
rect 37924 37748 37976 37768
rect 37976 37748 37978 37768
rect 37922 37712 37978 37748
rect 37922 36352 37978 36408
rect 37922 34992 37978 35048
rect 37922 34176 37978 34232
rect 37922 33632 37978 33688
rect 37922 32308 37924 32328
rect 37924 32308 37976 32328
rect 37976 32308 37978 32328
rect 37922 32272 37978 32308
rect 37922 31048 37978 31104
rect 37922 29688 37978 29744
rect 38014 28736 38070 28792
rect 37922 28328 37978 28384
rect 37922 26968 37978 27024
rect 37738 25336 37794 25392
rect 37922 25608 37978 25664
rect 38106 25472 38162 25528
rect 37922 24248 37978 24304
rect 37922 22888 37978 22944
rect 37922 22072 37978 22128
rect 37922 21528 37978 21584
rect 37922 20340 37924 20360
rect 37924 20340 37976 20360
rect 37976 20340 37978 20360
rect 37922 20304 37978 20340
rect 37922 18944 37978 19000
rect 37922 17584 37978 17640
rect 37922 16632 37978 16688
rect 37922 16224 37978 16280
rect 37922 14900 37924 14920
rect 37924 14900 37976 14920
rect 37976 14900 37978 14920
rect 37922 14864 37978 14900
rect 37922 13096 37978 13152
rect 37922 12144 37978 12200
rect 37922 9968 37978 10024
rect 37922 8608 37978 8664
rect 37922 7656 37978 7712
rect 37922 6432 37978 6488
rect 38566 70080 38622 70136
rect 38658 64776 38714 64832
rect 38934 71748 38936 71768
rect 38936 71748 38988 71768
rect 38988 71748 38990 71768
rect 38934 71712 38990 71748
rect 39762 63008 39818 63064
rect 38934 10784 38990 10840
rect 38934 5072 38990 5128
rect 37922 3032 37978 3088
rect 37094 176 37150 232
<< metal3 >>
rect 36077 119642 36143 119645
rect 39200 119642 40800 119672
rect 36077 119640 40800 119642
rect 36077 119584 36082 119640
rect 36138 119584 40800 119640
rect 36077 119582 40800 119584
rect 36077 119579 36143 119582
rect 39200 119552 40800 119582
rect -800 119506 800 119536
rect 3417 119506 3483 119509
rect -800 119504 3483 119506
rect -800 119448 3422 119504
rect 3478 119448 3483 119504
rect -800 119446 3483 119448
rect -800 119416 800 119446
rect 3417 119443 3483 119446
rect 37181 119234 37247 119237
rect 39200 119234 40800 119264
rect 37181 119232 40800 119234
rect 37181 119176 37186 119232
rect 37242 119176 40800 119232
rect 37181 119174 40800 119176
rect 37181 119171 37247 119174
rect 39200 119144 40800 119174
rect 34605 118826 34671 118829
rect 39200 118826 40800 118856
rect 34605 118824 40800 118826
rect 34605 118768 34610 118824
rect 34666 118768 40800 118824
rect 34605 118766 40800 118768
rect 34605 118763 34671 118766
rect 39200 118736 40800 118766
rect -800 118690 800 118720
rect 2865 118690 2931 118693
rect -800 118688 2931 118690
rect -800 118632 2870 118688
rect 2926 118632 2931 118688
rect -800 118630 2931 118632
rect -800 118600 800 118630
rect 2865 118627 2931 118630
rect 35341 118282 35407 118285
rect 39200 118282 40800 118312
rect 35341 118280 40800 118282
rect 35341 118224 35346 118280
rect 35402 118224 40800 118280
rect 35341 118222 40800 118224
rect 35341 118219 35407 118222
rect 39200 118192 40800 118222
rect -800 117874 800 117904
rect 1393 117874 1459 117877
rect -800 117872 1459 117874
rect -800 117816 1398 117872
rect 1454 117816 1459 117872
rect -800 117814 1459 117816
rect -800 117784 800 117814
rect 1393 117811 1459 117814
rect 36905 117874 36971 117877
rect 39200 117874 40800 117904
rect 36905 117872 40800 117874
rect 36905 117816 36910 117872
rect 36966 117816 40800 117872
rect 36905 117814 40800 117816
rect 36905 117811 36971 117814
rect 39200 117784 40800 117814
rect 4208 117536 4528 117537
rect 4208 117472 4216 117536
rect 4280 117472 4296 117536
rect 4360 117472 4376 117536
rect 4440 117472 4456 117536
rect 4520 117472 4528 117536
rect 4208 117471 4528 117472
rect 34928 117536 35248 117537
rect 34928 117472 34936 117536
rect 35000 117472 35016 117536
rect 35080 117472 35096 117536
rect 35160 117472 35176 117536
rect 35240 117472 35248 117536
rect 34928 117471 35248 117472
rect 35617 117466 35683 117469
rect 39200 117466 40800 117496
rect 35617 117464 40800 117466
rect 35617 117408 35622 117464
rect 35678 117408 40800 117464
rect 35617 117406 40800 117408
rect 35617 117403 35683 117406
rect 39200 117376 40800 117406
rect 25773 117330 25839 117333
rect 26969 117330 27035 117333
rect 25773 117328 27035 117330
rect 25773 117272 25778 117328
rect 25834 117272 26974 117328
rect 27030 117272 27035 117328
rect 25773 117270 27035 117272
rect 25773 117267 25839 117270
rect 26969 117267 27035 117270
rect -800 117058 800 117088
rect 2773 117058 2839 117061
rect -800 117056 2839 117058
rect -800 117000 2778 117056
rect 2834 117000 2839 117056
rect -800 116998 2839 117000
rect -800 116968 800 116998
rect 2773 116995 2839 116998
rect 24945 117058 25011 117061
rect 28625 117058 28691 117061
rect 24945 117056 28691 117058
rect 24945 117000 24950 117056
rect 25006 117000 28630 117056
rect 28686 117000 28691 117056
rect 24945 116998 28691 117000
rect 24945 116995 25011 116998
rect 28625 116995 28691 116998
rect 19568 116992 19888 116993
rect 19568 116928 19576 116992
rect 19640 116928 19656 116992
rect 19720 116928 19736 116992
rect 19800 116928 19816 116992
rect 19880 116928 19888 116992
rect 19568 116927 19888 116928
rect 35525 116922 35591 116925
rect 39200 116922 40800 116952
rect 35525 116920 40800 116922
rect 35525 116864 35530 116920
rect 35586 116864 40800 116920
rect 35525 116862 40800 116864
rect 35525 116859 35591 116862
rect 39200 116832 40800 116862
rect 23105 116786 23171 116789
rect 36537 116786 36603 116789
rect 23105 116784 36603 116786
rect 23105 116728 23110 116784
rect 23166 116728 36542 116784
rect 36598 116728 36603 116784
rect 23105 116726 36603 116728
rect 23105 116723 23171 116726
rect 36537 116723 36603 116726
rect 35341 116514 35407 116517
rect 39200 116514 40800 116544
rect 35341 116512 40800 116514
rect 35341 116456 35346 116512
rect 35402 116456 40800 116512
rect 35341 116454 40800 116456
rect 35341 116451 35407 116454
rect 4208 116448 4528 116449
rect 4208 116384 4216 116448
rect 4280 116384 4296 116448
rect 4360 116384 4376 116448
rect 4440 116384 4456 116448
rect 4520 116384 4528 116448
rect 4208 116383 4528 116384
rect 34928 116448 35248 116449
rect 34928 116384 34936 116448
rect 35000 116384 35016 116448
rect 35080 116384 35096 116448
rect 35160 116384 35176 116448
rect 35240 116384 35248 116448
rect 39200 116424 40800 116454
rect 34928 116383 35248 116384
rect 22645 116378 22711 116381
rect 25405 116378 25471 116381
rect 22645 116376 25471 116378
rect 22645 116320 22650 116376
rect 22706 116320 25410 116376
rect 25466 116320 25471 116376
rect 22645 116318 25471 116320
rect 22645 116315 22711 116318
rect 25405 116315 25471 116318
rect -800 116242 800 116272
rect 2037 116242 2103 116245
rect -800 116240 2103 116242
rect -800 116184 2042 116240
rect 2098 116184 2103 116240
rect -800 116182 2103 116184
rect -800 116152 800 116182
rect 2037 116179 2103 116182
rect 22461 116242 22527 116245
rect 26417 116242 26483 116245
rect 22461 116240 26483 116242
rect 22461 116184 22466 116240
rect 22522 116184 26422 116240
rect 26478 116184 26483 116240
rect 22461 116182 26483 116184
rect 22461 116179 22527 116182
rect 26417 116179 26483 116182
rect 24761 116106 24827 116109
rect 28349 116106 28415 116109
rect 24761 116104 28415 116106
rect 24761 116048 24766 116104
rect 24822 116048 28354 116104
rect 28410 116048 28415 116104
rect 24761 116046 28415 116048
rect 24761 116043 24827 116046
rect 28349 116043 28415 116046
rect 30925 116106 30991 116109
rect 31753 116106 31819 116109
rect 30925 116104 31819 116106
rect 30925 116048 30930 116104
rect 30986 116048 31758 116104
rect 31814 116048 31819 116104
rect 30925 116046 31819 116048
rect 30925 116043 30991 116046
rect 31753 116043 31819 116046
rect 35157 116106 35223 116109
rect 39200 116106 40800 116136
rect 35157 116104 40800 116106
rect 35157 116048 35162 116104
rect 35218 116048 40800 116104
rect 35157 116046 40800 116048
rect 35157 116043 35223 116046
rect 39200 116016 40800 116046
rect 30373 115970 30439 115973
rect 32397 115970 32463 115973
rect 30373 115968 32463 115970
rect 28993 115950 29059 115953
rect 28950 115948 29059 115950
rect 19568 115904 19888 115905
rect 19568 115840 19576 115904
rect 19640 115840 19656 115904
rect 19720 115840 19736 115904
rect 19800 115840 19816 115904
rect 19880 115840 19888 115904
rect 19568 115839 19888 115840
rect 28950 115892 28998 115948
rect 29054 115892 29059 115948
rect 30373 115912 30378 115968
rect 30434 115912 32402 115968
rect 32458 115912 32463 115968
rect 30373 115910 32463 115912
rect 30373 115907 30439 115910
rect 32397 115907 32463 115910
rect 28950 115887 29059 115892
rect 28950 115698 29010 115887
rect 29177 115834 29243 115837
rect 29545 115834 29611 115837
rect 29177 115832 29611 115834
rect 29177 115776 29182 115832
rect 29238 115776 29550 115832
rect 29606 115776 29611 115832
rect 29177 115774 29611 115776
rect 29177 115771 29243 115774
rect 29545 115771 29611 115774
rect 29545 115698 29611 115701
rect 28950 115696 29611 115698
rect 28950 115640 29550 115696
rect 29606 115640 29611 115696
rect 28950 115638 29611 115640
rect 29545 115635 29611 115638
rect 34513 115698 34579 115701
rect 39200 115698 40800 115728
rect 34513 115696 40800 115698
rect 34513 115640 34518 115696
rect 34574 115640 40800 115696
rect 34513 115638 40800 115640
rect 34513 115635 34579 115638
rect 39200 115608 40800 115638
rect 35157 115562 35223 115565
rect 35157 115560 35450 115562
rect 35157 115504 35162 115560
rect 35218 115504 35450 115560
rect 35157 115502 35450 115504
rect 35157 115499 35223 115502
rect -800 115426 800 115456
rect 1945 115426 2011 115429
rect -800 115424 2011 115426
rect -800 115368 1950 115424
rect 2006 115368 2011 115424
rect -800 115366 2011 115368
rect -800 115336 800 115366
rect 1945 115363 2011 115366
rect 4208 115360 4528 115361
rect 4208 115296 4216 115360
rect 4280 115296 4296 115360
rect 4360 115296 4376 115360
rect 4440 115296 4456 115360
rect 4520 115296 4528 115360
rect 4208 115295 4528 115296
rect 34928 115360 35248 115361
rect 34928 115296 34936 115360
rect 35000 115296 35016 115360
rect 35080 115296 35096 115360
rect 35160 115296 35176 115360
rect 35240 115296 35248 115360
rect 34928 115295 35248 115296
rect 29177 115290 29243 115293
rect 30281 115290 30347 115293
rect 29177 115288 30347 115290
rect 29177 115232 29182 115288
rect 29238 115232 30286 115288
rect 30342 115232 30347 115288
rect 29177 115230 30347 115232
rect 29177 115227 29243 115230
rect 30281 115227 30347 115230
rect 35390 115157 35450 115502
rect 21449 115154 21515 115157
rect 23013 115154 23079 115157
rect 21449 115152 23079 115154
rect 21449 115096 21454 115152
rect 21510 115096 23018 115152
rect 23074 115096 23079 115152
rect 21449 115094 23079 115096
rect 21449 115091 21515 115094
rect 23013 115091 23079 115094
rect 24025 115154 24091 115157
rect 29361 115154 29427 115157
rect 24025 115152 29427 115154
rect 24025 115096 24030 115152
rect 24086 115096 29366 115152
rect 29422 115096 29427 115152
rect 24025 115094 29427 115096
rect 24025 115091 24091 115094
rect 29361 115091 29427 115094
rect 35341 115152 35450 115157
rect 35341 115096 35346 115152
rect 35402 115096 35450 115152
rect 35341 115094 35450 115096
rect 37365 115154 37431 115157
rect 39200 115154 40800 115184
rect 37365 115152 40800 115154
rect 37365 115096 37370 115152
rect 37426 115096 40800 115152
rect 37365 115094 40800 115096
rect 35341 115091 35407 115094
rect 37365 115091 37431 115094
rect 39200 115064 40800 115094
rect 26417 115018 26483 115021
rect 28809 115018 28875 115021
rect 26417 115016 28875 115018
rect 26417 114960 26422 115016
rect 26478 114960 28814 115016
rect 28870 114960 28875 115016
rect 26417 114958 28875 114960
rect 26417 114955 26483 114958
rect 28809 114955 28875 114958
rect 19568 114816 19888 114817
rect 19568 114752 19576 114816
rect 19640 114752 19656 114816
rect 19720 114752 19736 114816
rect 19800 114752 19816 114816
rect 19880 114752 19888 114816
rect 19568 114751 19888 114752
rect 36537 114746 36603 114749
rect 39200 114746 40800 114776
rect 36537 114744 40800 114746
rect 36537 114688 36542 114744
rect 36598 114688 40800 114744
rect 36537 114686 40800 114688
rect 36537 114683 36603 114686
rect 39200 114656 40800 114686
rect -800 114610 800 114640
rect 2037 114610 2103 114613
rect -800 114608 2103 114610
rect -800 114552 2042 114608
rect 2098 114552 2103 114608
rect -800 114550 2103 114552
rect -800 114520 800 114550
rect 2037 114547 2103 114550
rect 37917 114338 37983 114341
rect 39200 114338 40800 114368
rect 37917 114336 40800 114338
rect 37917 114280 37922 114336
rect 37978 114280 40800 114336
rect 37917 114278 40800 114280
rect 37917 114275 37983 114278
rect 4208 114272 4528 114273
rect 4208 114208 4216 114272
rect 4280 114208 4296 114272
rect 4360 114208 4376 114272
rect 4440 114208 4456 114272
rect 4520 114208 4528 114272
rect 4208 114207 4528 114208
rect 34928 114272 35248 114273
rect 34928 114208 34936 114272
rect 35000 114208 35016 114272
rect 35080 114208 35096 114272
rect 35160 114208 35176 114272
rect 35240 114208 35248 114272
rect 39200 114248 40800 114278
rect 34928 114207 35248 114208
rect -800 113794 800 113824
rect 1853 113794 1919 113797
rect -800 113792 1919 113794
rect -800 113736 1858 113792
rect 1914 113736 1919 113792
rect -800 113734 1919 113736
rect -800 113704 800 113734
rect 1853 113731 1919 113734
rect 37917 113794 37983 113797
rect 39200 113794 40800 113824
rect 37917 113792 40800 113794
rect 37917 113736 37922 113792
rect 37978 113736 40800 113792
rect 37917 113734 40800 113736
rect 37917 113731 37983 113734
rect 19568 113728 19888 113729
rect 19568 113664 19576 113728
rect 19640 113664 19656 113728
rect 19720 113664 19736 113728
rect 19800 113664 19816 113728
rect 19880 113664 19888 113728
rect 39200 113704 40800 113734
rect 19568 113663 19888 113664
rect 37181 113386 37247 113389
rect 39200 113386 40800 113416
rect 37181 113384 40800 113386
rect 37181 113328 37186 113384
rect 37242 113328 40800 113384
rect 37181 113326 40800 113328
rect 37181 113323 37247 113326
rect 39200 113296 40800 113326
rect 4208 113184 4528 113185
rect -800 113114 800 113144
rect 4208 113120 4216 113184
rect 4280 113120 4296 113184
rect 4360 113120 4376 113184
rect 4440 113120 4456 113184
rect 4520 113120 4528 113184
rect 4208 113119 4528 113120
rect 34928 113184 35248 113185
rect 34928 113120 34936 113184
rect 35000 113120 35016 113184
rect 35080 113120 35096 113184
rect 35160 113120 35176 113184
rect 35240 113120 35248 113184
rect 34928 113119 35248 113120
rect 1945 113114 2011 113117
rect -800 113112 2011 113114
rect -800 113056 1950 113112
rect 2006 113056 2011 113112
rect -800 113054 2011 113056
rect -800 113024 800 113054
rect 1945 113051 2011 113054
rect 37917 112978 37983 112981
rect 39200 112978 40800 113008
rect 37917 112976 40800 112978
rect 37917 112920 37922 112976
rect 37978 112920 40800 112976
rect 37917 112918 40800 112920
rect 37917 112915 37983 112918
rect 39200 112888 40800 112918
rect 19568 112640 19888 112641
rect 19568 112576 19576 112640
rect 19640 112576 19656 112640
rect 19720 112576 19736 112640
rect 19800 112576 19816 112640
rect 19880 112576 19888 112640
rect 19568 112575 19888 112576
rect 37089 112570 37155 112573
rect 39200 112570 40800 112600
rect 37089 112568 40800 112570
rect 37089 112512 37094 112568
rect 37150 112512 40800 112568
rect 37089 112510 40800 112512
rect 37089 112507 37155 112510
rect 39200 112480 40800 112510
rect -800 112298 800 112328
rect 2037 112298 2103 112301
rect -800 112296 2103 112298
rect -800 112240 2042 112296
rect 2098 112240 2103 112296
rect -800 112238 2103 112240
rect -800 112208 800 112238
rect 2037 112235 2103 112238
rect 4208 112096 4528 112097
rect 4208 112032 4216 112096
rect 4280 112032 4296 112096
rect 4360 112032 4376 112096
rect 4440 112032 4456 112096
rect 4520 112032 4528 112096
rect 4208 112031 4528 112032
rect 34928 112096 35248 112097
rect 34928 112032 34936 112096
rect 35000 112032 35016 112096
rect 35080 112032 35096 112096
rect 35160 112032 35176 112096
rect 35240 112032 35248 112096
rect 34928 112031 35248 112032
rect 37089 112026 37155 112029
rect 39200 112026 40800 112056
rect 37089 112024 40800 112026
rect 37089 111968 37094 112024
rect 37150 111968 40800 112024
rect 37089 111966 40800 111968
rect 37089 111963 37155 111966
rect 39200 111936 40800 111966
rect 37825 111618 37891 111621
rect 39200 111618 40800 111648
rect 37825 111616 40800 111618
rect 37825 111560 37830 111616
rect 37886 111560 40800 111616
rect 37825 111558 40800 111560
rect 37825 111555 37891 111558
rect 19568 111552 19888 111553
rect -800 111482 800 111512
rect 19568 111488 19576 111552
rect 19640 111488 19656 111552
rect 19720 111488 19736 111552
rect 19800 111488 19816 111552
rect 19880 111488 19888 111552
rect 39200 111528 40800 111558
rect 19568 111487 19888 111488
rect 1945 111482 2011 111485
rect -800 111480 2011 111482
rect -800 111424 1950 111480
rect 2006 111424 2011 111480
rect -800 111422 2011 111424
rect -800 111392 800 111422
rect 1945 111419 2011 111422
rect 37089 111210 37155 111213
rect 39200 111210 40800 111240
rect 37089 111208 40800 111210
rect 37089 111152 37094 111208
rect 37150 111152 40800 111208
rect 37089 111150 40800 111152
rect 37089 111147 37155 111150
rect 39200 111120 40800 111150
rect 4208 111008 4528 111009
rect 4208 110944 4216 111008
rect 4280 110944 4296 111008
rect 4360 110944 4376 111008
rect 4440 110944 4456 111008
rect 4520 110944 4528 111008
rect 4208 110943 4528 110944
rect 34928 111008 35248 111009
rect 34928 110944 34936 111008
rect 35000 110944 35016 111008
rect 35080 110944 35096 111008
rect 35160 110944 35176 111008
rect 35240 110944 35248 111008
rect 34928 110943 35248 110944
rect -800 110666 800 110696
rect 2037 110666 2103 110669
rect -800 110664 2103 110666
rect -800 110608 2042 110664
rect 2098 110608 2103 110664
rect -800 110606 2103 110608
rect -800 110576 800 110606
rect 2037 110603 2103 110606
rect 37825 110666 37891 110669
rect 39200 110666 40800 110696
rect 37825 110664 40800 110666
rect 37825 110608 37830 110664
rect 37886 110608 40800 110664
rect 37825 110606 40800 110608
rect 37825 110603 37891 110606
rect 39200 110576 40800 110606
rect 19568 110464 19888 110465
rect 19568 110400 19576 110464
rect 19640 110400 19656 110464
rect 19720 110400 19736 110464
rect 19800 110400 19816 110464
rect 19880 110400 19888 110464
rect 19568 110399 19888 110400
rect 37089 110258 37155 110261
rect 39200 110258 40800 110288
rect 37089 110256 40800 110258
rect 37089 110200 37094 110256
rect 37150 110200 40800 110256
rect 37089 110198 40800 110200
rect 37089 110195 37155 110198
rect 39200 110168 40800 110198
rect 35801 110122 35867 110125
rect 35574 110120 35867 110122
rect 35574 110064 35806 110120
rect 35862 110064 35867 110120
rect 35574 110062 35867 110064
rect 4208 109920 4528 109921
rect -800 109850 800 109880
rect 4208 109856 4216 109920
rect 4280 109856 4296 109920
rect 4360 109856 4376 109920
rect 4440 109856 4456 109920
rect 4520 109856 4528 109920
rect 4208 109855 4528 109856
rect 34928 109920 35248 109921
rect 34928 109856 34936 109920
rect 35000 109856 35016 109920
rect 35080 109856 35096 109920
rect 35160 109856 35176 109920
rect 35240 109856 35248 109920
rect 34928 109855 35248 109856
rect 1945 109850 2011 109853
rect -800 109848 2011 109850
rect -800 109792 1950 109848
rect 2006 109792 2011 109848
rect -800 109790 2011 109792
rect -800 109760 800 109790
rect 1945 109787 2011 109790
rect 35433 109714 35499 109717
rect 35574 109714 35634 110062
rect 35801 110059 35867 110062
rect 37089 109850 37155 109853
rect 39200 109850 40800 109880
rect 37089 109848 40800 109850
rect 37089 109792 37094 109848
rect 37150 109792 40800 109848
rect 37089 109790 40800 109792
rect 37089 109787 37155 109790
rect 39200 109760 40800 109790
rect 35433 109712 35634 109714
rect 35433 109656 35438 109712
rect 35494 109656 35634 109712
rect 35433 109654 35634 109656
rect 35433 109651 35499 109654
rect 37825 109442 37891 109445
rect 39200 109442 40800 109472
rect 37825 109440 40800 109442
rect 37825 109384 37830 109440
rect 37886 109384 40800 109440
rect 37825 109382 40800 109384
rect 37825 109379 37891 109382
rect 19568 109376 19888 109377
rect 19568 109312 19576 109376
rect 19640 109312 19656 109376
rect 19720 109312 19736 109376
rect 19800 109312 19816 109376
rect 19880 109312 19888 109376
rect 39200 109352 40800 109382
rect 19568 109311 19888 109312
rect -800 109034 800 109064
rect 1853 109034 1919 109037
rect -800 109032 1919 109034
rect -800 108976 1858 109032
rect 1914 108976 1919 109032
rect -800 108974 1919 108976
rect -800 108944 800 108974
rect 1853 108971 1919 108974
rect 37089 108898 37155 108901
rect 39200 108898 40800 108928
rect 37089 108896 40800 108898
rect 37089 108840 37094 108896
rect 37150 108840 40800 108896
rect 37089 108838 40800 108840
rect 37089 108835 37155 108838
rect 4208 108832 4528 108833
rect 4208 108768 4216 108832
rect 4280 108768 4296 108832
rect 4360 108768 4376 108832
rect 4440 108768 4456 108832
rect 4520 108768 4528 108832
rect 4208 108767 4528 108768
rect 34928 108832 35248 108833
rect 34928 108768 34936 108832
rect 35000 108768 35016 108832
rect 35080 108768 35096 108832
rect 35160 108768 35176 108832
rect 35240 108768 35248 108832
rect 39200 108808 40800 108838
rect 34928 108767 35248 108768
rect 37825 108490 37891 108493
rect 39200 108490 40800 108520
rect 37825 108488 40800 108490
rect 37825 108432 37830 108488
rect 37886 108432 40800 108488
rect 37825 108430 40800 108432
rect 37825 108427 37891 108430
rect 39200 108400 40800 108430
rect 19568 108288 19888 108289
rect -800 108218 800 108248
rect 19568 108224 19576 108288
rect 19640 108224 19656 108288
rect 19720 108224 19736 108288
rect 19800 108224 19816 108288
rect 19880 108224 19888 108288
rect 19568 108223 19888 108224
rect 1945 108218 2011 108221
rect -800 108216 2011 108218
rect -800 108160 1950 108216
rect 2006 108160 2011 108216
rect -800 108158 2011 108160
rect -800 108128 800 108158
rect 1945 108155 2011 108158
rect 37181 108082 37247 108085
rect 39200 108082 40800 108112
rect 37181 108080 40800 108082
rect 37181 108024 37186 108080
rect 37242 108024 40800 108080
rect 37181 108022 40800 108024
rect 37181 108019 37247 108022
rect 39200 107992 40800 108022
rect 4208 107744 4528 107745
rect 4208 107680 4216 107744
rect 4280 107680 4296 107744
rect 4360 107680 4376 107744
rect 4440 107680 4456 107744
rect 4520 107680 4528 107744
rect 4208 107679 4528 107680
rect 34928 107744 35248 107745
rect 34928 107680 34936 107744
rect 35000 107680 35016 107744
rect 35080 107680 35096 107744
rect 35160 107680 35176 107744
rect 35240 107680 35248 107744
rect 34928 107679 35248 107680
rect 37181 107538 37247 107541
rect 39200 107538 40800 107568
rect 37181 107536 40800 107538
rect 37181 107480 37186 107536
rect 37242 107480 40800 107536
rect 37181 107478 40800 107480
rect 37181 107475 37247 107478
rect 39200 107448 40800 107478
rect -800 107402 800 107432
rect 2037 107402 2103 107405
rect -800 107400 2103 107402
rect -800 107344 2042 107400
rect 2098 107344 2103 107400
rect -800 107342 2103 107344
rect -800 107312 800 107342
rect 2037 107339 2103 107342
rect 19568 107200 19888 107201
rect 19568 107136 19576 107200
rect 19640 107136 19656 107200
rect 19720 107136 19736 107200
rect 19800 107136 19816 107200
rect 19880 107136 19888 107200
rect 19568 107135 19888 107136
rect 37917 107130 37983 107133
rect 39200 107130 40800 107160
rect 37917 107128 40800 107130
rect 37917 107072 37922 107128
rect 37978 107072 40800 107128
rect 37917 107070 40800 107072
rect 37917 107067 37983 107070
rect 39200 107040 40800 107070
rect -800 106722 800 106752
rect 1945 106722 2011 106725
rect -800 106720 2011 106722
rect -800 106664 1950 106720
rect 2006 106664 2011 106720
rect -800 106662 2011 106664
rect -800 106632 800 106662
rect 1945 106659 2011 106662
rect 37181 106722 37247 106725
rect 39200 106722 40800 106752
rect 37181 106720 40800 106722
rect 37181 106664 37186 106720
rect 37242 106664 40800 106720
rect 37181 106662 40800 106664
rect 37181 106659 37247 106662
rect 4208 106656 4528 106657
rect 4208 106592 4216 106656
rect 4280 106592 4296 106656
rect 4360 106592 4376 106656
rect 4440 106592 4456 106656
rect 4520 106592 4528 106656
rect 4208 106591 4528 106592
rect 34928 106656 35248 106657
rect 34928 106592 34936 106656
rect 35000 106592 35016 106656
rect 35080 106592 35096 106656
rect 35160 106592 35176 106656
rect 35240 106592 35248 106656
rect 39200 106632 40800 106662
rect 34928 106591 35248 106592
rect 37917 106178 37983 106181
rect 39200 106178 40800 106208
rect 37917 106176 40800 106178
rect 37917 106120 37922 106176
rect 37978 106120 40800 106176
rect 37917 106118 40800 106120
rect 37917 106115 37983 106118
rect 19568 106112 19888 106113
rect 19568 106048 19576 106112
rect 19640 106048 19656 106112
rect 19720 106048 19736 106112
rect 19800 106048 19816 106112
rect 19880 106048 19888 106112
rect 39200 106088 40800 106118
rect 19568 106047 19888 106048
rect -800 105906 800 105936
rect 1393 105906 1459 105909
rect -800 105904 1459 105906
rect -800 105848 1398 105904
rect 1454 105848 1459 105904
rect -800 105846 1459 105848
rect -800 105816 800 105846
rect 1393 105843 1459 105846
rect 37181 105770 37247 105773
rect 39200 105770 40800 105800
rect 37181 105768 40800 105770
rect 37181 105712 37186 105768
rect 37242 105712 40800 105768
rect 37181 105710 40800 105712
rect 37181 105707 37247 105710
rect 39200 105680 40800 105710
rect 4208 105568 4528 105569
rect 4208 105504 4216 105568
rect 4280 105504 4296 105568
rect 4360 105504 4376 105568
rect 4440 105504 4456 105568
rect 4520 105504 4528 105568
rect 4208 105503 4528 105504
rect 34928 105568 35248 105569
rect 34928 105504 34936 105568
rect 35000 105504 35016 105568
rect 35080 105504 35096 105568
rect 35160 105504 35176 105568
rect 35240 105504 35248 105568
rect 34928 105503 35248 105504
rect 37917 105362 37983 105365
rect 39200 105362 40800 105392
rect 37917 105360 40800 105362
rect 37917 105304 37922 105360
rect 37978 105304 40800 105360
rect 37917 105302 40800 105304
rect 37917 105299 37983 105302
rect 39200 105272 40800 105302
rect -800 105090 800 105120
rect 1945 105090 2011 105093
rect -800 105088 2011 105090
rect -800 105032 1950 105088
rect 2006 105032 2011 105088
rect -800 105030 2011 105032
rect -800 105000 800 105030
rect 1945 105027 2011 105030
rect 19568 105024 19888 105025
rect 19568 104960 19576 105024
rect 19640 104960 19656 105024
rect 19720 104960 19736 105024
rect 19800 104960 19816 105024
rect 19880 104960 19888 105024
rect 19568 104959 19888 104960
rect 37181 104954 37247 104957
rect 39200 104954 40800 104984
rect 37181 104952 40800 104954
rect 37181 104896 37186 104952
rect 37242 104896 40800 104952
rect 37181 104894 40800 104896
rect 37181 104891 37247 104894
rect 39200 104864 40800 104894
rect 4208 104480 4528 104481
rect 4208 104416 4216 104480
rect 4280 104416 4296 104480
rect 4360 104416 4376 104480
rect 4440 104416 4456 104480
rect 4520 104416 4528 104480
rect 4208 104415 4528 104416
rect 34928 104480 35248 104481
rect 34928 104416 34936 104480
rect 35000 104416 35016 104480
rect 35080 104416 35096 104480
rect 35160 104416 35176 104480
rect 35240 104416 35248 104480
rect 34928 104415 35248 104416
rect 37181 104410 37247 104413
rect 39200 104410 40800 104440
rect 37181 104408 40800 104410
rect 37181 104352 37186 104408
rect 37242 104352 40800 104408
rect 37181 104350 40800 104352
rect 37181 104347 37247 104350
rect 39200 104320 40800 104350
rect -800 104274 800 104304
rect 1485 104274 1551 104277
rect -800 104272 1551 104274
rect -800 104216 1490 104272
rect 1546 104216 1551 104272
rect -800 104214 1551 104216
rect -800 104184 800 104214
rect 1485 104211 1551 104214
rect 37917 104002 37983 104005
rect 39200 104002 40800 104032
rect 37917 104000 40800 104002
rect 37917 103944 37922 104000
rect 37978 103944 40800 104000
rect 37917 103942 40800 103944
rect 37917 103939 37983 103942
rect 19568 103936 19888 103937
rect 19568 103872 19576 103936
rect 19640 103872 19656 103936
rect 19720 103872 19736 103936
rect 19800 103872 19816 103936
rect 19880 103872 19888 103936
rect 39200 103912 40800 103942
rect 19568 103871 19888 103872
rect 37181 103594 37247 103597
rect 39200 103594 40800 103624
rect 37181 103592 40800 103594
rect 37181 103536 37186 103592
rect 37242 103536 40800 103592
rect 37181 103534 40800 103536
rect 37181 103531 37247 103534
rect 39200 103504 40800 103534
rect -800 103458 800 103488
rect 2037 103458 2103 103461
rect -800 103456 2103 103458
rect -800 103400 2042 103456
rect 2098 103400 2103 103456
rect -800 103398 2103 103400
rect -800 103368 800 103398
rect 2037 103395 2103 103398
rect 4208 103392 4528 103393
rect 4208 103328 4216 103392
rect 4280 103328 4296 103392
rect 4360 103328 4376 103392
rect 4440 103328 4456 103392
rect 4520 103328 4528 103392
rect 4208 103327 4528 103328
rect 34928 103392 35248 103393
rect 34928 103328 34936 103392
rect 35000 103328 35016 103392
rect 35080 103328 35096 103392
rect 35160 103328 35176 103392
rect 35240 103328 35248 103392
rect 34928 103327 35248 103328
rect 37917 103050 37983 103053
rect 39200 103050 40800 103080
rect 37917 103048 40800 103050
rect 37917 102992 37922 103048
rect 37978 102992 40800 103048
rect 37917 102990 40800 102992
rect 37917 102987 37983 102990
rect 39200 102960 40800 102990
rect 19568 102848 19888 102849
rect 19568 102784 19576 102848
rect 19640 102784 19656 102848
rect 19720 102784 19736 102848
rect 19800 102784 19816 102848
rect 19880 102784 19888 102848
rect 19568 102783 19888 102784
rect -800 102642 800 102672
rect 2037 102642 2103 102645
rect -800 102640 2103 102642
rect -800 102584 2042 102640
rect 2098 102584 2103 102640
rect -800 102582 2103 102584
rect -800 102552 800 102582
rect 2037 102579 2103 102582
rect 37181 102642 37247 102645
rect 39200 102642 40800 102672
rect 37181 102640 40800 102642
rect 37181 102584 37186 102640
rect 37242 102584 40800 102640
rect 37181 102582 40800 102584
rect 37181 102579 37247 102582
rect 39200 102552 40800 102582
rect 4208 102304 4528 102305
rect 4208 102240 4216 102304
rect 4280 102240 4296 102304
rect 4360 102240 4376 102304
rect 4440 102240 4456 102304
rect 4520 102240 4528 102304
rect 4208 102239 4528 102240
rect 34928 102304 35248 102305
rect 34928 102240 34936 102304
rect 35000 102240 35016 102304
rect 35080 102240 35096 102304
rect 35160 102240 35176 102304
rect 35240 102240 35248 102304
rect 34928 102239 35248 102240
rect 37181 102234 37247 102237
rect 39200 102234 40800 102264
rect 37181 102232 40800 102234
rect 37181 102176 37186 102232
rect 37242 102176 40800 102232
rect 37181 102174 40800 102176
rect 37181 102171 37247 102174
rect 39200 102144 40800 102174
rect -800 101826 800 101856
rect 1393 101826 1459 101829
rect -800 101824 1459 101826
rect -800 101768 1398 101824
rect 1454 101768 1459 101824
rect -800 101766 1459 101768
rect -800 101736 800 101766
rect 1393 101763 1459 101766
rect 37917 101826 37983 101829
rect 39200 101826 40800 101856
rect 37917 101824 40800 101826
rect 37917 101768 37922 101824
rect 37978 101768 40800 101824
rect 37917 101766 40800 101768
rect 37917 101763 37983 101766
rect 19568 101760 19888 101761
rect 19568 101696 19576 101760
rect 19640 101696 19656 101760
rect 19720 101696 19736 101760
rect 19800 101696 19816 101760
rect 19880 101696 19888 101760
rect 39200 101736 40800 101766
rect 19568 101695 19888 101696
rect 37181 101282 37247 101285
rect 39200 101282 40800 101312
rect 37181 101280 40800 101282
rect 37181 101224 37186 101280
rect 37242 101224 40800 101280
rect 37181 101222 40800 101224
rect 37181 101219 37247 101222
rect 4208 101216 4528 101217
rect 4208 101152 4216 101216
rect 4280 101152 4296 101216
rect 4360 101152 4376 101216
rect 4440 101152 4456 101216
rect 4520 101152 4528 101216
rect 4208 101151 4528 101152
rect 34928 101216 35248 101217
rect 34928 101152 34936 101216
rect 35000 101152 35016 101216
rect 35080 101152 35096 101216
rect 35160 101152 35176 101216
rect 35240 101152 35248 101216
rect 39200 101192 40800 101222
rect 34928 101151 35248 101152
rect -800 101010 800 101040
rect 1393 101010 1459 101013
rect -800 101008 1459 101010
rect -800 100952 1398 101008
rect 1454 100952 1459 101008
rect -800 100950 1459 100952
rect -800 100920 800 100950
rect 1393 100947 1459 100950
rect 37917 100874 37983 100877
rect 39200 100874 40800 100904
rect 37917 100872 40800 100874
rect 37917 100816 37922 100872
rect 37978 100816 40800 100872
rect 37917 100814 40800 100816
rect 37917 100811 37983 100814
rect 39200 100784 40800 100814
rect 19568 100672 19888 100673
rect 19568 100608 19576 100672
rect 19640 100608 19656 100672
rect 19720 100608 19736 100672
rect 19800 100608 19816 100672
rect 19880 100608 19888 100672
rect 19568 100607 19888 100608
rect 37181 100466 37247 100469
rect 39200 100466 40800 100496
rect 37181 100464 40800 100466
rect 37181 100408 37186 100464
rect 37242 100408 40800 100464
rect 37181 100406 40800 100408
rect 37181 100403 37247 100406
rect 39200 100376 40800 100406
rect -800 100330 800 100360
rect 1393 100330 1459 100333
rect -800 100328 1459 100330
rect -800 100272 1398 100328
rect 1454 100272 1459 100328
rect -800 100270 1459 100272
rect -800 100240 800 100270
rect 1393 100267 1459 100270
rect 4208 100128 4528 100129
rect 4208 100064 4216 100128
rect 4280 100064 4296 100128
rect 4360 100064 4376 100128
rect 4440 100064 4456 100128
rect 4520 100064 4528 100128
rect 4208 100063 4528 100064
rect 34928 100128 35248 100129
rect 34928 100064 34936 100128
rect 35000 100064 35016 100128
rect 35080 100064 35096 100128
rect 35160 100064 35176 100128
rect 35240 100064 35248 100128
rect 34928 100063 35248 100064
rect 37273 99922 37339 99925
rect 39200 99922 40800 99952
rect 37273 99920 40800 99922
rect 37273 99864 37278 99920
rect 37334 99864 40800 99920
rect 37273 99862 40800 99864
rect 37273 99859 37339 99862
rect 39200 99832 40800 99862
rect 19568 99584 19888 99585
rect -800 99514 800 99544
rect 19568 99520 19576 99584
rect 19640 99520 19656 99584
rect 19720 99520 19736 99584
rect 19800 99520 19816 99584
rect 19880 99520 19888 99584
rect 19568 99519 19888 99520
rect 1393 99514 1459 99517
rect -800 99512 1459 99514
rect -800 99456 1398 99512
rect 1454 99456 1459 99512
rect -800 99454 1459 99456
rect -800 99424 800 99454
rect 1393 99451 1459 99454
rect 37181 99514 37247 99517
rect 39200 99514 40800 99544
rect 37181 99512 40800 99514
rect 37181 99456 37186 99512
rect 37242 99456 40800 99512
rect 37181 99454 40800 99456
rect 37181 99451 37247 99454
rect 39200 99424 40800 99454
rect 37917 99106 37983 99109
rect 39200 99106 40800 99136
rect 37917 99104 40800 99106
rect 37917 99048 37922 99104
rect 37978 99048 40800 99104
rect 37917 99046 40800 99048
rect 37917 99043 37983 99046
rect 4208 99040 4528 99041
rect 4208 98976 4216 99040
rect 4280 98976 4296 99040
rect 4360 98976 4376 99040
rect 4440 98976 4456 99040
rect 4520 98976 4528 99040
rect 4208 98975 4528 98976
rect 34928 99040 35248 99041
rect 34928 98976 34936 99040
rect 35000 98976 35016 99040
rect 35080 98976 35096 99040
rect 35160 98976 35176 99040
rect 35240 98976 35248 99040
rect 39200 99016 40800 99046
rect 34928 98975 35248 98976
rect -800 98698 800 98728
rect 1393 98698 1459 98701
rect -800 98696 1459 98698
rect -800 98640 1398 98696
rect 1454 98640 1459 98696
rect -800 98638 1459 98640
rect -800 98608 800 98638
rect 1393 98635 1459 98638
rect 37917 98698 37983 98701
rect 39200 98698 40800 98728
rect 37917 98696 40800 98698
rect 37917 98640 37922 98696
rect 37978 98640 40800 98696
rect 37917 98638 40800 98640
rect 37917 98635 37983 98638
rect 39200 98608 40800 98638
rect 19568 98496 19888 98497
rect 19568 98432 19576 98496
rect 19640 98432 19656 98496
rect 19720 98432 19736 98496
rect 19800 98432 19816 98496
rect 19880 98432 19888 98496
rect 19568 98431 19888 98432
rect 37089 98154 37155 98157
rect 39200 98154 40800 98184
rect 37089 98152 40800 98154
rect 37089 98096 37094 98152
rect 37150 98096 40800 98152
rect 37089 98094 40800 98096
rect 37089 98091 37155 98094
rect 39200 98064 40800 98094
rect 4208 97952 4528 97953
rect -800 97882 800 97912
rect 4208 97888 4216 97952
rect 4280 97888 4296 97952
rect 4360 97888 4376 97952
rect 4440 97888 4456 97952
rect 4520 97888 4528 97952
rect 4208 97887 4528 97888
rect 34928 97952 35248 97953
rect 34928 97888 34936 97952
rect 35000 97888 35016 97952
rect 35080 97888 35096 97952
rect 35160 97888 35176 97952
rect 35240 97888 35248 97952
rect 34928 97887 35248 97888
rect 1393 97882 1459 97885
rect -800 97880 1459 97882
rect -800 97824 1398 97880
rect 1454 97824 1459 97880
rect -800 97822 1459 97824
rect -800 97792 800 97822
rect 1393 97819 1459 97822
rect 37825 97746 37891 97749
rect 39200 97746 40800 97776
rect 37825 97744 40800 97746
rect 37825 97688 37830 97744
rect 37886 97688 40800 97744
rect 37825 97686 40800 97688
rect 37825 97683 37891 97686
rect 39200 97656 40800 97686
rect 19568 97408 19888 97409
rect 19568 97344 19576 97408
rect 19640 97344 19656 97408
rect 19720 97344 19736 97408
rect 19800 97344 19816 97408
rect 19880 97344 19888 97408
rect 19568 97343 19888 97344
rect 37089 97338 37155 97341
rect 39200 97338 40800 97368
rect 37089 97336 40800 97338
rect 37089 97280 37094 97336
rect 37150 97280 40800 97336
rect 37089 97278 40800 97280
rect 37089 97275 37155 97278
rect 39200 97248 40800 97278
rect -800 97066 800 97096
rect 1393 97066 1459 97069
rect -800 97064 1459 97066
rect -800 97008 1398 97064
rect 1454 97008 1459 97064
rect -800 97006 1459 97008
rect -800 96976 800 97006
rect 1393 97003 1459 97006
rect 4208 96864 4528 96865
rect 4208 96800 4216 96864
rect 4280 96800 4296 96864
rect 4360 96800 4376 96864
rect 4440 96800 4456 96864
rect 4520 96800 4528 96864
rect 4208 96799 4528 96800
rect 34928 96864 35248 96865
rect 34928 96800 34936 96864
rect 35000 96800 35016 96864
rect 35080 96800 35096 96864
rect 35160 96800 35176 96864
rect 35240 96800 35248 96864
rect 34928 96799 35248 96800
rect 37089 96794 37155 96797
rect 39200 96794 40800 96824
rect 37089 96792 40800 96794
rect 37089 96736 37094 96792
rect 37150 96736 40800 96792
rect 37089 96734 40800 96736
rect 37089 96731 37155 96734
rect 39200 96704 40800 96734
rect 37917 96386 37983 96389
rect 39200 96386 40800 96416
rect 37917 96384 40800 96386
rect 37917 96328 37922 96384
rect 37978 96328 40800 96384
rect 37917 96326 40800 96328
rect 37917 96323 37983 96326
rect 19568 96320 19888 96321
rect -800 96250 800 96280
rect 19568 96256 19576 96320
rect 19640 96256 19656 96320
rect 19720 96256 19736 96320
rect 19800 96256 19816 96320
rect 19880 96256 19888 96320
rect 39200 96296 40800 96326
rect 19568 96255 19888 96256
rect 1393 96250 1459 96253
rect -800 96248 1459 96250
rect -800 96192 1398 96248
rect 1454 96192 1459 96248
rect -800 96190 1459 96192
rect -800 96160 800 96190
rect 1393 96187 1459 96190
rect 37181 95978 37247 95981
rect 39200 95978 40800 96008
rect 37181 95976 40800 95978
rect 37181 95920 37186 95976
rect 37242 95920 40800 95976
rect 37181 95918 40800 95920
rect 37181 95915 37247 95918
rect 39200 95888 40800 95918
rect 4208 95776 4528 95777
rect 4208 95712 4216 95776
rect 4280 95712 4296 95776
rect 4360 95712 4376 95776
rect 4440 95712 4456 95776
rect 4520 95712 4528 95776
rect 4208 95711 4528 95712
rect 34928 95776 35248 95777
rect 34928 95712 34936 95776
rect 35000 95712 35016 95776
rect 35080 95712 35096 95776
rect 35160 95712 35176 95776
rect 35240 95712 35248 95776
rect 34928 95711 35248 95712
rect -800 95434 800 95464
rect 1393 95434 1459 95437
rect -800 95432 1459 95434
rect -800 95376 1398 95432
rect 1454 95376 1459 95432
rect -800 95374 1459 95376
rect -800 95344 800 95374
rect 1393 95371 1459 95374
rect 37917 95434 37983 95437
rect 39200 95434 40800 95464
rect 37917 95432 40800 95434
rect 37917 95376 37922 95432
rect 37978 95376 40800 95432
rect 37917 95374 40800 95376
rect 37917 95371 37983 95374
rect 39200 95344 40800 95374
rect 19568 95232 19888 95233
rect 19568 95168 19576 95232
rect 19640 95168 19656 95232
rect 19720 95168 19736 95232
rect 19800 95168 19816 95232
rect 19880 95168 19888 95232
rect 19568 95167 19888 95168
rect 37181 95026 37247 95029
rect 39200 95026 40800 95056
rect 37181 95024 40800 95026
rect 37181 94968 37186 95024
rect 37242 94968 40800 95024
rect 37181 94966 40800 94968
rect 37181 94963 37247 94966
rect 39200 94936 40800 94966
rect 4208 94688 4528 94689
rect -800 94618 800 94648
rect 4208 94624 4216 94688
rect 4280 94624 4296 94688
rect 4360 94624 4376 94688
rect 4440 94624 4456 94688
rect 4520 94624 4528 94688
rect 4208 94623 4528 94624
rect 34928 94688 35248 94689
rect 34928 94624 34936 94688
rect 35000 94624 35016 94688
rect 35080 94624 35096 94688
rect 35160 94624 35176 94688
rect 35240 94624 35248 94688
rect 34928 94623 35248 94624
rect 1393 94618 1459 94621
rect -800 94616 1459 94618
rect -800 94560 1398 94616
rect 1454 94560 1459 94616
rect -800 94558 1459 94560
rect -800 94528 800 94558
rect 1393 94555 1459 94558
rect 37181 94618 37247 94621
rect 39200 94618 40800 94648
rect 37181 94616 40800 94618
rect 37181 94560 37186 94616
rect 37242 94560 40800 94616
rect 37181 94558 40800 94560
rect 37181 94555 37247 94558
rect 39200 94528 40800 94558
rect 37917 94210 37983 94213
rect 39200 94210 40800 94240
rect 37917 94208 40800 94210
rect 37917 94152 37922 94208
rect 37978 94152 40800 94208
rect 37917 94150 40800 94152
rect 37917 94147 37983 94150
rect 19568 94144 19888 94145
rect 19568 94080 19576 94144
rect 19640 94080 19656 94144
rect 19720 94080 19736 94144
rect 19800 94080 19816 94144
rect 19880 94080 19888 94144
rect 39200 94120 40800 94150
rect 19568 94079 19888 94080
rect -800 93802 800 93832
rect 1393 93802 1459 93805
rect -800 93800 1459 93802
rect -800 93744 1398 93800
rect 1454 93744 1459 93800
rect -800 93742 1459 93744
rect -800 93712 800 93742
rect 1393 93739 1459 93742
rect 37181 93666 37247 93669
rect 39200 93666 40800 93696
rect 37181 93664 40800 93666
rect 37181 93608 37186 93664
rect 37242 93608 40800 93664
rect 37181 93606 40800 93608
rect 37181 93603 37247 93606
rect 4208 93600 4528 93601
rect 4208 93536 4216 93600
rect 4280 93536 4296 93600
rect 4360 93536 4376 93600
rect 4440 93536 4456 93600
rect 4520 93536 4528 93600
rect 4208 93535 4528 93536
rect 34928 93600 35248 93601
rect 34928 93536 34936 93600
rect 35000 93536 35016 93600
rect 35080 93536 35096 93600
rect 35160 93536 35176 93600
rect 35240 93536 35248 93600
rect 39200 93576 40800 93606
rect 34928 93535 35248 93536
rect 37273 93258 37339 93261
rect 39200 93258 40800 93288
rect 37273 93256 40800 93258
rect 37273 93200 37278 93256
rect 37334 93200 40800 93256
rect 37273 93198 40800 93200
rect 37273 93195 37339 93198
rect 39200 93168 40800 93198
rect -800 93122 800 93152
rect 1393 93122 1459 93125
rect -800 93120 1459 93122
rect -800 93064 1398 93120
rect 1454 93064 1459 93120
rect -800 93062 1459 93064
rect -800 93032 800 93062
rect 1393 93059 1459 93062
rect 19568 93056 19888 93057
rect 19568 92992 19576 93056
rect 19640 92992 19656 93056
rect 19720 92992 19736 93056
rect 19800 92992 19816 93056
rect 19880 92992 19888 93056
rect 19568 92991 19888 92992
rect 37917 92850 37983 92853
rect 39200 92850 40800 92880
rect 37917 92848 40800 92850
rect 37917 92792 37922 92848
rect 37978 92792 40800 92848
rect 37917 92790 40800 92792
rect 37917 92787 37983 92790
rect 39200 92760 40800 92790
rect 4208 92512 4528 92513
rect 4208 92448 4216 92512
rect 4280 92448 4296 92512
rect 4360 92448 4376 92512
rect 4440 92448 4456 92512
rect 4520 92448 4528 92512
rect 4208 92447 4528 92448
rect 34928 92512 35248 92513
rect 34928 92448 34936 92512
rect 35000 92448 35016 92512
rect 35080 92448 35096 92512
rect 35160 92448 35176 92512
rect 35240 92448 35248 92512
rect 34928 92447 35248 92448
rect -800 92306 800 92336
rect 1393 92306 1459 92309
rect -800 92304 1459 92306
rect -800 92248 1398 92304
rect 1454 92248 1459 92304
rect -800 92246 1459 92248
rect -800 92216 800 92246
rect 1393 92243 1459 92246
rect 37273 92306 37339 92309
rect 39200 92306 40800 92336
rect 37273 92304 40800 92306
rect 37273 92248 37278 92304
rect 37334 92248 40800 92304
rect 37273 92246 40800 92248
rect 37273 92243 37339 92246
rect 39200 92216 40800 92246
rect 19568 91968 19888 91969
rect 19568 91904 19576 91968
rect 19640 91904 19656 91968
rect 19720 91904 19736 91968
rect 19800 91904 19816 91968
rect 19880 91904 19888 91968
rect 19568 91903 19888 91904
rect 37181 91898 37247 91901
rect 39200 91898 40800 91928
rect 37181 91896 40800 91898
rect 37181 91840 37186 91896
rect 37242 91840 40800 91896
rect 37181 91838 40800 91840
rect 37181 91835 37247 91838
rect 39200 91808 40800 91838
rect -800 91490 800 91520
rect 1393 91490 1459 91493
rect -800 91488 1459 91490
rect -800 91432 1398 91488
rect 1454 91432 1459 91488
rect -800 91430 1459 91432
rect -800 91400 800 91430
rect 1393 91427 1459 91430
rect 37917 91490 37983 91493
rect 39200 91490 40800 91520
rect 37917 91488 40800 91490
rect 37917 91432 37922 91488
rect 37978 91432 40800 91488
rect 37917 91430 40800 91432
rect 37917 91427 37983 91430
rect 4208 91424 4528 91425
rect 4208 91360 4216 91424
rect 4280 91360 4296 91424
rect 4360 91360 4376 91424
rect 4440 91360 4456 91424
rect 4520 91360 4528 91424
rect 4208 91359 4528 91360
rect 34928 91424 35248 91425
rect 34928 91360 34936 91424
rect 35000 91360 35016 91424
rect 35080 91360 35096 91424
rect 35160 91360 35176 91424
rect 35240 91360 35248 91424
rect 39200 91400 40800 91430
rect 34928 91359 35248 91360
rect 37181 91082 37247 91085
rect 39200 91082 40800 91112
rect 37181 91080 40800 91082
rect 37181 91024 37186 91080
rect 37242 91024 40800 91080
rect 37181 91022 40800 91024
rect 37181 91019 37247 91022
rect 39200 90992 40800 91022
rect 19568 90880 19888 90881
rect 19568 90816 19576 90880
rect 19640 90816 19656 90880
rect 19720 90816 19736 90880
rect 19800 90816 19816 90880
rect 19880 90816 19888 90880
rect 19568 90815 19888 90816
rect -800 90674 800 90704
rect 2037 90674 2103 90677
rect -800 90672 2103 90674
rect -800 90616 2042 90672
rect 2098 90616 2103 90672
rect -800 90614 2103 90616
rect -800 90584 800 90614
rect 2037 90611 2103 90614
rect 37917 90538 37983 90541
rect 39200 90538 40800 90568
rect 37917 90536 40800 90538
rect 37917 90480 37922 90536
rect 37978 90480 40800 90536
rect 37917 90478 40800 90480
rect 37917 90475 37983 90478
rect 39200 90448 40800 90478
rect 4208 90336 4528 90337
rect 4208 90272 4216 90336
rect 4280 90272 4296 90336
rect 4360 90272 4376 90336
rect 4440 90272 4456 90336
rect 4520 90272 4528 90336
rect 4208 90271 4528 90272
rect 34928 90336 35248 90337
rect 34928 90272 34936 90336
rect 35000 90272 35016 90336
rect 35080 90272 35096 90336
rect 35160 90272 35176 90336
rect 35240 90272 35248 90336
rect 34928 90271 35248 90272
rect 37273 90130 37339 90133
rect 39200 90130 40800 90160
rect 37273 90128 40800 90130
rect 37273 90072 37278 90128
rect 37334 90072 40800 90128
rect 37273 90070 40800 90072
rect 37273 90067 37339 90070
rect 39200 90040 40800 90070
rect -800 89858 800 89888
rect 1393 89858 1459 89861
rect -800 89856 1459 89858
rect -800 89800 1398 89856
rect 1454 89800 1459 89856
rect -800 89798 1459 89800
rect -800 89768 800 89798
rect 1393 89795 1459 89798
rect 19568 89792 19888 89793
rect 19568 89728 19576 89792
rect 19640 89728 19656 89792
rect 19720 89728 19736 89792
rect 19800 89728 19816 89792
rect 19880 89728 19888 89792
rect 19568 89727 19888 89728
rect 37181 89722 37247 89725
rect 39200 89722 40800 89752
rect 37181 89720 40800 89722
rect 37181 89664 37186 89720
rect 37242 89664 40800 89720
rect 37181 89662 40800 89664
rect 37181 89659 37247 89662
rect 39200 89632 40800 89662
rect 4208 89248 4528 89249
rect 4208 89184 4216 89248
rect 4280 89184 4296 89248
rect 4360 89184 4376 89248
rect 4440 89184 4456 89248
rect 4520 89184 4528 89248
rect 4208 89183 4528 89184
rect 34928 89248 35248 89249
rect 34928 89184 34936 89248
rect 35000 89184 35016 89248
rect 35080 89184 35096 89248
rect 35160 89184 35176 89248
rect 35240 89184 35248 89248
rect 34928 89183 35248 89184
rect 37917 89178 37983 89181
rect 39200 89178 40800 89208
rect 37917 89176 40800 89178
rect 37917 89120 37922 89176
rect 37978 89120 40800 89176
rect 37917 89118 40800 89120
rect 37917 89115 37983 89118
rect 39200 89088 40800 89118
rect -800 89042 800 89072
rect 1393 89042 1459 89045
rect -800 89040 1459 89042
rect -800 88984 1398 89040
rect 1454 88984 1459 89040
rect -800 88982 1459 88984
rect -800 88952 800 88982
rect 1393 88979 1459 88982
rect 37273 88770 37339 88773
rect 39200 88770 40800 88800
rect 37273 88768 40800 88770
rect 37273 88712 37278 88768
rect 37334 88712 40800 88768
rect 37273 88710 40800 88712
rect 37273 88707 37339 88710
rect 19568 88704 19888 88705
rect 19568 88640 19576 88704
rect 19640 88640 19656 88704
rect 19720 88640 19736 88704
rect 19800 88640 19816 88704
rect 19880 88640 19888 88704
rect 39200 88680 40800 88710
rect 19568 88639 19888 88640
rect 37917 88362 37983 88365
rect 39200 88362 40800 88392
rect 37917 88360 40800 88362
rect 37917 88304 37922 88360
rect 37978 88304 40800 88360
rect 37917 88302 40800 88304
rect 37917 88299 37983 88302
rect 39200 88272 40800 88302
rect -800 88226 800 88256
rect 1393 88226 1459 88229
rect -800 88224 1459 88226
rect -800 88168 1398 88224
rect 1454 88168 1459 88224
rect -800 88166 1459 88168
rect -800 88136 800 88166
rect 1393 88163 1459 88166
rect 4208 88160 4528 88161
rect 4208 88096 4216 88160
rect 4280 88096 4296 88160
rect 4360 88096 4376 88160
rect 4440 88096 4456 88160
rect 4520 88096 4528 88160
rect 4208 88095 4528 88096
rect 34928 88160 35248 88161
rect 34928 88096 34936 88160
rect 35000 88096 35016 88160
rect 35080 88096 35096 88160
rect 35160 88096 35176 88160
rect 35240 88096 35248 88160
rect 34928 88095 35248 88096
rect 37273 87954 37339 87957
rect 39200 87954 40800 87984
rect 37273 87952 40800 87954
rect 37273 87896 37278 87952
rect 37334 87896 40800 87952
rect 37273 87894 40800 87896
rect 37273 87891 37339 87894
rect 39200 87864 40800 87894
rect 19568 87616 19888 87617
rect 19568 87552 19576 87616
rect 19640 87552 19656 87616
rect 19720 87552 19736 87616
rect 19800 87552 19816 87616
rect 19880 87552 19888 87616
rect 19568 87551 19888 87552
rect -800 87410 800 87440
rect 1393 87410 1459 87413
rect -800 87408 1459 87410
rect -800 87352 1398 87408
rect 1454 87352 1459 87408
rect -800 87350 1459 87352
rect -800 87320 800 87350
rect 1393 87347 1459 87350
rect 37181 87410 37247 87413
rect 39200 87410 40800 87440
rect 37181 87408 40800 87410
rect 37181 87352 37186 87408
rect 37242 87352 40800 87408
rect 37181 87350 40800 87352
rect 37181 87347 37247 87350
rect 39200 87320 40800 87350
rect 34789 87274 34855 87277
rect 34654 87272 34855 87274
rect 34654 87216 34794 87272
rect 34850 87216 34855 87272
rect 34654 87214 34855 87216
rect 4208 87072 4528 87073
rect 4208 87008 4216 87072
rect 4280 87008 4296 87072
rect 4360 87008 4376 87072
rect 4440 87008 4456 87072
rect 4520 87008 4528 87072
rect 4208 87007 4528 87008
rect 34654 87002 34714 87214
rect 34789 87211 34855 87214
rect 36813 87274 36879 87277
rect 36813 87272 37106 87274
rect 36813 87216 36818 87272
rect 36874 87216 37106 87272
rect 36813 87214 37106 87216
rect 36813 87211 36879 87214
rect 36721 87138 36787 87141
rect 36905 87138 36971 87141
rect 36721 87136 36971 87138
rect 36721 87080 36726 87136
rect 36782 87080 36910 87136
rect 36966 87080 36971 87136
rect 36721 87078 36971 87080
rect 36721 87075 36787 87078
rect 36905 87075 36971 87078
rect 34928 87072 35248 87073
rect 34928 87008 34936 87072
rect 35000 87008 35016 87072
rect 35080 87008 35096 87072
rect 35160 87008 35176 87072
rect 35240 87008 35248 87072
rect 34928 87007 35248 87008
rect 34789 87002 34855 87005
rect 34654 87000 34855 87002
rect 34654 86944 34794 87000
rect 34850 86944 34855 87000
rect 34654 86942 34855 86944
rect 34789 86939 34855 86942
rect 36813 87002 36879 87005
rect 37046 87002 37106 87214
rect 36813 87000 37106 87002
rect 36813 86944 36818 87000
rect 36874 86944 37106 87000
rect 36813 86942 37106 86944
rect 37917 87002 37983 87005
rect 39200 87002 40800 87032
rect 37917 87000 40800 87002
rect 37917 86944 37922 87000
rect 37978 86944 40800 87000
rect 37917 86942 40800 86944
rect 36813 86939 36879 86942
rect 37917 86939 37983 86942
rect 39200 86912 40800 86942
rect -800 86730 800 86760
rect 1393 86730 1459 86733
rect -800 86728 1459 86730
rect -800 86672 1398 86728
rect 1454 86672 1459 86728
rect -800 86670 1459 86672
rect -800 86640 800 86670
rect 1393 86667 1459 86670
rect 37273 86594 37339 86597
rect 39200 86594 40800 86624
rect 37273 86592 40800 86594
rect 37273 86536 37278 86592
rect 37334 86536 40800 86592
rect 37273 86534 40800 86536
rect 37273 86531 37339 86534
rect 19568 86528 19888 86529
rect 19568 86464 19576 86528
rect 19640 86464 19656 86528
rect 19720 86464 19736 86528
rect 19800 86464 19816 86528
rect 19880 86464 19888 86528
rect 39200 86504 40800 86534
rect 19568 86463 19888 86464
rect 29637 86322 29703 86325
rect 34329 86322 34395 86325
rect 29637 86320 34395 86322
rect 29637 86264 29642 86320
rect 29698 86264 34334 86320
rect 34390 86264 34395 86320
rect 29637 86262 34395 86264
rect 29637 86259 29703 86262
rect 34329 86259 34395 86262
rect 37917 86050 37983 86053
rect 39200 86050 40800 86080
rect 37917 86048 40800 86050
rect 37917 85992 37922 86048
rect 37978 85992 40800 86048
rect 37917 85990 40800 85992
rect 37917 85987 37983 85990
rect 4208 85984 4528 85985
rect -800 85914 800 85944
rect 4208 85920 4216 85984
rect 4280 85920 4296 85984
rect 4360 85920 4376 85984
rect 4440 85920 4456 85984
rect 4520 85920 4528 85984
rect 4208 85919 4528 85920
rect 34928 85984 35248 85985
rect 34928 85920 34936 85984
rect 35000 85920 35016 85984
rect 35080 85920 35096 85984
rect 35160 85920 35176 85984
rect 35240 85920 35248 85984
rect 39200 85960 40800 85990
rect 34928 85919 35248 85920
rect 1393 85914 1459 85917
rect -800 85912 1459 85914
rect -800 85856 1398 85912
rect 1454 85856 1459 85912
rect -800 85854 1459 85856
rect -800 85824 800 85854
rect 1393 85851 1459 85854
rect 37273 85642 37339 85645
rect 39200 85642 40800 85672
rect 37273 85640 40800 85642
rect 37273 85584 37278 85640
rect 37334 85584 40800 85640
rect 37273 85582 40800 85584
rect 37273 85579 37339 85582
rect 39200 85552 40800 85582
rect 19568 85440 19888 85441
rect 19568 85376 19576 85440
rect 19640 85376 19656 85440
rect 19720 85376 19736 85440
rect 19800 85376 19816 85440
rect 19880 85376 19888 85440
rect 19568 85375 19888 85376
rect 37917 85234 37983 85237
rect 39200 85234 40800 85264
rect 37917 85232 40800 85234
rect 37917 85176 37922 85232
rect 37978 85176 40800 85232
rect 37917 85174 40800 85176
rect 37917 85171 37983 85174
rect 39200 85144 40800 85174
rect -800 85098 800 85128
rect 1393 85098 1459 85101
rect -800 85096 1459 85098
rect -800 85040 1398 85096
rect 1454 85040 1459 85096
rect -800 85038 1459 85040
rect -800 85008 800 85038
rect 1393 85035 1459 85038
rect 4208 84896 4528 84897
rect 4208 84832 4216 84896
rect 4280 84832 4296 84896
rect 4360 84832 4376 84896
rect 4440 84832 4456 84896
rect 4520 84832 4528 84896
rect 4208 84831 4528 84832
rect 34928 84896 35248 84897
rect 34928 84832 34936 84896
rect 35000 84832 35016 84896
rect 35080 84832 35096 84896
rect 35160 84832 35176 84896
rect 35240 84832 35248 84896
rect 34928 84831 35248 84832
rect 37273 84826 37339 84829
rect 39200 84826 40800 84856
rect 37273 84824 40800 84826
rect 37273 84768 37278 84824
rect 37334 84768 40800 84824
rect 37273 84766 40800 84768
rect 37273 84763 37339 84766
rect 39200 84736 40800 84766
rect 19568 84352 19888 84353
rect -800 84282 800 84312
rect 19568 84288 19576 84352
rect 19640 84288 19656 84352
rect 19720 84288 19736 84352
rect 19800 84288 19816 84352
rect 19880 84288 19888 84352
rect 19568 84287 19888 84288
rect 1393 84282 1459 84285
rect -800 84280 1459 84282
rect -800 84224 1398 84280
rect 1454 84224 1459 84280
rect -800 84222 1459 84224
rect -800 84192 800 84222
rect 1393 84219 1459 84222
rect 37181 84282 37247 84285
rect 39200 84282 40800 84312
rect 37181 84280 40800 84282
rect 37181 84224 37186 84280
rect 37242 84224 40800 84280
rect 37181 84222 40800 84224
rect 37181 84219 37247 84222
rect 39200 84192 40800 84222
rect 37917 83874 37983 83877
rect 39200 83874 40800 83904
rect 37917 83872 40800 83874
rect 37917 83816 37922 83872
rect 37978 83816 40800 83872
rect 37917 83814 40800 83816
rect 37917 83811 37983 83814
rect 4208 83808 4528 83809
rect 4208 83744 4216 83808
rect 4280 83744 4296 83808
rect 4360 83744 4376 83808
rect 4440 83744 4456 83808
rect 4520 83744 4528 83808
rect 4208 83743 4528 83744
rect 34928 83808 35248 83809
rect 34928 83744 34936 83808
rect 35000 83744 35016 83808
rect 35080 83744 35096 83808
rect 35160 83744 35176 83808
rect 35240 83744 35248 83808
rect 39200 83784 40800 83814
rect 34928 83743 35248 83744
rect -800 83466 800 83496
rect 1393 83466 1459 83469
rect -800 83464 1459 83466
rect -800 83408 1398 83464
rect 1454 83408 1459 83464
rect -800 83406 1459 83408
rect -800 83376 800 83406
rect 1393 83403 1459 83406
rect 37273 83466 37339 83469
rect 39200 83466 40800 83496
rect 37273 83464 40800 83466
rect 37273 83408 37278 83464
rect 37334 83408 40800 83464
rect 37273 83406 40800 83408
rect 37273 83403 37339 83406
rect 39200 83376 40800 83406
rect 19568 83264 19888 83265
rect 19568 83200 19576 83264
rect 19640 83200 19656 83264
rect 19720 83200 19736 83264
rect 19800 83200 19816 83264
rect 19880 83200 19888 83264
rect 19568 83199 19888 83200
rect 37917 82922 37983 82925
rect 39200 82922 40800 82952
rect 37917 82920 40800 82922
rect 37917 82864 37922 82920
rect 37978 82864 40800 82920
rect 37917 82862 40800 82864
rect 37917 82859 37983 82862
rect 39200 82832 40800 82862
rect 4208 82720 4528 82721
rect -800 82650 800 82680
rect 4208 82656 4216 82720
rect 4280 82656 4296 82720
rect 4360 82656 4376 82720
rect 4440 82656 4456 82720
rect 4520 82656 4528 82720
rect 4208 82655 4528 82656
rect 34928 82720 35248 82721
rect 34928 82656 34936 82720
rect 35000 82656 35016 82720
rect 35080 82656 35096 82720
rect 35160 82656 35176 82720
rect 35240 82656 35248 82720
rect 34928 82655 35248 82656
rect 1393 82650 1459 82653
rect -800 82648 1459 82650
rect -800 82592 1398 82648
rect 1454 82592 1459 82648
rect -800 82590 1459 82592
rect -800 82560 800 82590
rect 1393 82587 1459 82590
rect 37273 82514 37339 82517
rect 39200 82514 40800 82544
rect 37273 82512 40800 82514
rect 37273 82456 37278 82512
rect 37334 82456 40800 82512
rect 37273 82454 40800 82456
rect 37273 82451 37339 82454
rect 39200 82424 40800 82454
rect 19568 82176 19888 82177
rect 19568 82112 19576 82176
rect 19640 82112 19656 82176
rect 19720 82112 19736 82176
rect 19800 82112 19816 82176
rect 19880 82112 19888 82176
rect 19568 82111 19888 82112
rect 37181 82106 37247 82109
rect 39200 82106 40800 82136
rect 37181 82104 40800 82106
rect 37181 82048 37186 82104
rect 37242 82048 40800 82104
rect 37181 82046 40800 82048
rect 37181 82043 37247 82046
rect 39200 82016 40800 82046
rect 33041 81970 33107 81973
rect 32998 81968 33107 81970
rect 32998 81912 33046 81968
rect 33102 81912 33107 81968
rect 32998 81907 33107 81912
rect -800 81834 800 81864
rect 1393 81834 1459 81837
rect -800 81832 1459 81834
rect -800 81776 1398 81832
rect 1454 81776 1459 81832
rect -800 81774 1459 81776
rect -800 81744 800 81774
rect 1393 81771 1459 81774
rect 4208 81632 4528 81633
rect 4208 81568 4216 81632
rect 4280 81568 4296 81632
rect 4360 81568 4376 81632
rect 4440 81568 4456 81632
rect 4520 81568 4528 81632
rect 4208 81567 4528 81568
rect 32765 81562 32831 81565
rect 32998 81562 33058 81907
rect 34928 81632 35248 81633
rect 34928 81568 34936 81632
rect 35000 81568 35016 81632
rect 35080 81568 35096 81632
rect 35160 81568 35176 81632
rect 35240 81568 35248 81632
rect 34928 81567 35248 81568
rect 32765 81560 33058 81562
rect 32765 81504 32770 81560
rect 32826 81504 33058 81560
rect 32765 81502 33058 81504
rect 37917 81562 37983 81565
rect 39200 81562 40800 81592
rect 37917 81560 40800 81562
rect 37917 81504 37922 81560
rect 37978 81504 40800 81560
rect 37917 81502 40800 81504
rect 32765 81499 32831 81502
rect 37917 81499 37983 81502
rect 39200 81472 40800 81502
rect 37273 81154 37339 81157
rect 39200 81154 40800 81184
rect 37273 81152 40800 81154
rect 37273 81096 37278 81152
rect 37334 81096 40800 81152
rect 37273 81094 40800 81096
rect 37273 81091 37339 81094
rect 19568 81088 19888 81089
rect -800 81018 800 81048
rect 19568 81024 19576 81088
rect 19640 81024 19656 81088
rect 19720 81024 19736 81088
rect 19800 81024 19816 81088
rect 19880 81024 19888 81088
rect 39200 81064 40800 81094
rect 19568 81023 19888 81024
rect 1393 81018 1459 81021
rect -800 81016 1459 81018
rect -800 80960 1398 81016
rect 1454 80960 1459 81016
rect -800 80958 1459 80960
rect -800 80928 800 80958
rect 1393 80955 1459 80958
rect 37917 80746 37983 80749
rect 39200 80746 40800 80776
rect 37917 80744 40800 80746
rect 37917 80688 37922 80744
rect 37978 80688 40800 80744
rect 37917 80686 40800 80688
rect 37917 80683 37983 80686
rect 39200 80656 40800 80686
rect 4208 80544 4528 80545
rect 4208 80480 4216 80544
rect 4280 80480 4296 80544
rect 4360 80480 4376 80544
rect 4440 80480 4456 80544
rect 4520 80480 4528 80544
rect 4208 80479 4528 80480
rect 34928 80544 35248 80545
rect 34928 80480 34936 80544
rect 35000 80480 35016 80544
rect 35080 80480 35096 80544
rect 35160 80480 35176 80544
rect 35240 80480 35248 80544
rect 34928 80479 35248 80480
rect -800 80338 800 80368
rect 1393 80338 1459 80341
rect -800 80336 1459 80338
rect -800 80280 1398 80336
rect 1454 80280 1459 80336
rect -800 80278 1459 80280
rect -800 80248 800 80278
rect 1393 80275 1459 80278
rect 37273 80338 37339 80341
rect 39200 80338 40800 80368
rect 37273 80336 40800 80338
rect 37273 80280 37278 80336
rect 37334 80280 40800 80336
rect 37273 80278 40800 80280
rect 37273 80275 37339 80278
rect 39200 80248 40800 80278
rect 19568 80000 19888 80001
rect 19568 79936 19576 80000
rect 19640 79936 19656 80000
rect 19720 79936 19736 80000
rect 19800 79936 19816 80000
rect 19880 79936 19888 80000
rect 19568 79935 19888 79936
rect 37181 79794 37247 79797
rect 39200 79794 40800 79824
rect 37181 79792 40800 79794
rect 37181 79736 37186 79792
rect 37242 79736 40800 79792
rect 37181 79734 40800 79736
rect 37181 79731 37247 79734
rect 39200 79704 40800 79734
rect -800 79522 800 79552
rect 1393 79522 1459 79525
rect -800 79520 1459 79522
rect -800 79464 1398 79520
rect 1454 79464 1459 79520
rect -800 79462 1459 79464
rect -800 79432 800 79462
rect 1393 79459 1459 79462
rect 4208 79456 4528 79457
rect 4208 79392 4216 79456
rect 4280 79392 4296 79456
rect 4360 79392 4376 79456
rect 4440 79392 4456 79456
rect 4520 79392 4528 79456
rect 4208 79391 4528 79392
rect 34928 79456 35248 79457
rect 34928 79392 34936 79456
rect 35000 79392 35016 79456
rect 35080 79392 35096 79456
rect 35160 79392 35176 79456
rect 35240 79392 35248 79456
rect 34928 79391 35248 79392
rect 37917 79386 37983 79389
rect 39200 79386 40800 79416
rect 37917 79384 40800 79386
rect 37917 79328 37922 79384
rect 37978 79328 40800 79384
rect 37917 79326 40800 79328
rect 37917 79323 37983 79326
rect 39200 79296 40800 79326
rect 37273 78978 37339 78981
rect 39200 78978 40800 79008
rect 37273 78976 40800 78978
rect 37273 78920 37278 78976
rect 37334 78920 40800 78976
rect 37273 78918 40800 78920
rect 37273 78915 37339 78918
rect 19568 78912 19888 78913
rect 19568 78848 19576 78912
rect 19640 78848 19656 78912
rect 19720 78848 19736 78912
rect 19800 78848 19816 78912
rect 19880 78848 19888 78912
rect 39200 78888 40800 78918
rect 19568 78847 19888 78848
rect -800 78706 800 78736
rect 1393 78706 1459 78709
rect -800 78704 1459 78706
rect -800 78648 1398 78704
rect 1454 78648 1459 78704
rect -800 78646 1459 78648
rect -800 78616 800 78646
rect 1393 78643 1459 78646
rect 37917 78434 37983 78437
rect 39200 78434 40800 78464
rect 37917 78432 40800 78434
rect 37917 78376 37922 78432
rect 37978 78376 40800 78432
rect 37917 78374 40800 78376
rect 37917 78371 37983 78374
rect 4208 78368 4528 78369
rect 4208 78304 4216 78368
rect 4280 78304 4296 78368
rect 4360 78304 4376 78368
rect 4440 78304 4456 78368
rect 4520 78304 4528 78368
rect 4208 78303 4528 78304
rect 34928 78368 35248 78369
rect 34928 78304 34936 78368
rect 35000 78304 35016 78368
rect 35080 78304 35096 78368
rect 35160 78304 35176 78368
rect 35240 78304 35248 78368
rect 39200 78344 40800 78374
rect 34928 78303 35248 78304
rect 37273 78026 37339 78029
rect 39200 78026 40800 78056
rect 37273 78024 40800 78026
rect 37273 77968 37278 78024
rect 37334 77968 40800 78024
rect 37273 77966 40800 77968
rect 37273 77963 37339 77966
rect 39200 77936 40800 77966
rect -800 77890 800 77920
rect 1393 77890 1459 77893
rect -800 77888 1459 77890
rect -800 77832 1398 77888
rect 1454 77832 1459 77888
rect -800 77830 1459 77832
rect -800 77800 800 77830
rect 1393 77827 1459 77830
rect 19568 77824 19888 77825
rect 19568 77760 19576 77824
rect 19640 77760 19656 77824
rect 19720 77760 19736 77824
rect 19800 77760 19816 77824
rect 19880 77760 19888 77824
rect 19568 77759 19888 77760
rect 37917 77618 37983 77621
rect 39200 77618 40800 77648
rect 37917 77616 40800 77618
rect 37917 77560 37922 77616
rect 37978 77560 40800 77616
rect 37917 77558 40800 77560
rect 37917 77555 37983 77558
rect 39200 77528 40800 77558
rect 4208 77280 4528 77281
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 77215 4528 77216
rect 34928 77280 35248 77281
rect 34928 77216 34936 77280
rect 35000 77216 35016 77280
rect 35080 77216 35096 77280
rect 35160 77216 35176 77280
rect 35240 77216 35248 77280
rect 34928 77215 35248 77216
rect 37273 77210 37339 77213
rect 39200 77210 40800 77240
rect 37273 77208 40800 77210
rect 37273 77152 37278 77208
rect 37334 77152 40800 77208
rect 37273 77150 40800 77152
rect 37273 77147 37339 77150
rect 39200 77120 40800 77150
rect -800 77074 800 77104
rect 1393 77074 1459 77077
rect -800 77072 1459 77074
rect -800 77016 1398 77072
rect 1454 77016 1459 77072
rect -800 77014 1459 77016
rect -800 76984 800 77014
rect 1393 77011 1459 77014
rect 19568 76736 19888 76737
rect 19568 76672 19576 76736
rect 19640 76672 19656 76736
rect 19720 76672 19736 76736
rect 19800 76672 19816 76736
rect 19880 76672 19888 76736
rect 19568 76671 19888 76672
rect 37917 76666 37983 76669
rect 39200 76666 40800 76696
rect 37917 76664 40800 76666
rect 37917 76608 37922 76664
rect 37978 76608 40800 76664
rect 37917 76606 40800 76608
rect 37917 76603 37983 76606
rect 39200 76576 40800 76606
rect -800 76258 800 76288
rect 1393 76258 1459 76261
rect -800 76256 1459 76258
rect -800 76200 1398 76256
rect 1454 76200 1459 76256
rect -800 76198 1459 76200
rect -800 76168 800 76198
rect 1393 76195 1459 76198
rect 38009 76258 38075 76261
rect 39200 76258 40800 76288
rect 38009 76256 40800 76258
rect 38009 76200 38014 76256
rect 38070 76200 40800 76256
rect 38009 76198 40800 76200
rect 38009 76195 38075 76198
rect 4208 76192 4528 76193
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 76127 4528 76128
rect 34928 76192 35248 76193
rect 34928 76128 34936 76192
rect 35000 76128 35016 76192
rect 35080 76128 35096 76192
rect 35160 76128 35176 76192
rect 35240 76128 35248 76192
rect 39200 76168 40800 76198
rect 34928 76127 35248 76128
rect 37273 75850 37339 75853
rect 39200 75850 40800 75880
rect 37273 75848 40800 75850
rect 37273 75792 37278 75848
rect 37334 75792 40800 75848
rect 37273 75790 40800 75792
rect 37273 75787 37339 75790
rect 39200 75760 40800 75790
rect 19568 75648 19888 75649
rect 19568 75584 19576 75648
rect 19640 75584 19656 75648
rect 19720 75584 19736 75648
rect 19800 75584 19816 75648
rect 19880 75584 19888 75648
rect 19568 75583 19888 75584
rect -800 75442 800 75472
rect 1393 75442 1459 75445
rect -800 75440 1459 75442
rect -800 75384 1398 75440
rect 1454 75384 1459 75440
rect -800 75382 1459 75384
rect -800 75352 800 75382
rect 1393 75379 1459 75382
rect 37181 75306 37247 75309
rect 39200 75306 40800 75336
rect 37181 75304 40800 75306
rect 37181 75248 37186 75304
rect 37242 75248 40800 75304
rect 37181 75246 40800 75248
rect 37181 75243 37247 75246
rect 39200 75216 40800 75246
rect 4208 75104 4528 75105
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 4208 75039 4528 75040
rect 34928 75104 35248 75105
rect 34928 75040 34936 75104
rect 35000 75040 35016 75104
rect 35080 75040 35096 75104
rect 35160 75040 35176 75104
rect 35240 75040 35248 75104
rect 34928 75039 35248 75040
rect 37273 74898 37339 74901
rect 39200 74898 40800 74928
rect 37273 74896 40800 74898
rect 37273 74840 37278 74896
rect 37334 74840 40800 74896
rect 37273 74838 40800 74840
rect 37273 74835 37339 74838
rect 39200 74808 40800 74838
rect -800 74626 800 74656
rect 1393 74626 1459 74629
rect -800 74624 1459 74626
rect -800 74568 1398 74624
rect 1454 74568 1459 74624
rect -800 74566 1459 74568
rect -800 74536 800 74566
rect 1393 74563 1459 74566
rect 19568 74560 19888 74561
rect 19568 74496 19576 74560
rect 19640 74496 19656 74560
rect 19720 74496 19736 74560
rect 19800 74496 19816 74560
rect 19880 74496 19888 74560
rect 19568 74495 19888 74496
rect 37181 74490 37247 74493
rect 39200 74490 40800 74520
rect 37181 74488 40800 74490
rect 37181 74432 37186 74488
rect 37242 74432 40800 74488
rect 37181 74430 40800 74432
rect 37181 74427 37247 74430
rect 39200 74400 40800 74430
rect 37917 74082 37983 74085
rect 39200 74082 40800 74112
rect 37917 74080 40800 74082
rect 37917 74024 37922 74080
rect 37978 74024 40800 74080
rect 37917 74022 40800 74024
rect 37917 74019 37983 74022
rect 4208 74016 4528 74017
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 73951 4528 73952
rect 34928 74016 35248 74017
rect 34928 73952 34936 74016
rect 35000 73952 35016 74016
rect 35080 73952 35096 74016
rect 35160 73952 35176 74016
rect 35240 73952 35248 74016
rect 39200 73992 40800 74022
rect 34928 73951 35248 73952
rect -800 73810 800 73840
rect 1393 73810 1459 73813
rect -800 73808 1459 73810
rect -800 73752 1398 73808
rect 1454 73752 1459 73808
rect -800 73750 1459 73752
rect -800 73720 800 73750
rect 1393 73747 1459 73750
rect 37273 73538 37339 73541
rect 39200 73538 40800 73568
rect 37273 73536 40800 73538
rect 37273 73480 37278 73536
rect 37334 73480 40800 73536
rect 37273 73478 40800 73480
rect 37273 73475 37339 73478
rect 19568 73472 19888 73473
rect 19568 73408 19576 73472
rect 19640 73408 19656 73472
rect 19720 73408 19736 73472
rect 19800 73408 19816 73472
rect 19880 73408 19888 73472
rect 39200 73448 40800 73478
rect 19568 73407 19888 73408
rect -800 73130 800 73160
rect 1393 73130 1459 73133
rect -800 73128 1459 73130
rect -800 73072 1398 73128
rect 1454 73072 1459 73128
rect -800 73070 1459 73072
rect -800 73040 800 73070
rect 1393 73067 1459 73070
rect 37917 73130 37983 73133
rect 39200 73130 40800 73160
rect 37917 73128 40800 73130
rect 37917 73072 37922 73128
rect 37978 73072 40800 73128
rect 37917 73070 40800 73072
rect 37917 73067 37983 73070
rect 39200 73040 40800 73070
rect 4208 72928 4528 72929
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 72863 4528 72864
rect 34928 72928 35248 72929
rect 34928 72864 34936 72928
rect 35000 72864 35016 72928
rect 35080 72864 35096 72928
rect 35160 72864 35176 72928
rect 35240 72864 35248 72928
rect 34928 72863 35248 72864
rect 37273 72722 37339 72725
rect 39200 72722 40800 72752
rect 37273 72720 40800 72722
rect 37273 72664 37278 72720
rect 37334 72664 40800 72720
rect 37273 72662 40800 72664
rect 37273 72659 37339 72662
rect 39200 72632 40800 72662
rect 19568 72384 19888 72385
rect -800 72314 800 72344
rect 19568 72320 19576 72384
rect 19640 72320 19656 72384
rect 19720 72320 19736 72384
rect 19800 72320 19816 72384
rect 19880 72320 19888 72384
rect 19568 72319 19888 72320
rect 1393 72314 1459 72317
rect -800 72312 1459 72314
rect -800 72256 1398 72312
rect 1454 72256 1459 72312
rect -800 72254 1459 72256
rect -800 72224 800 72254
rect 1393 72251 1459 72254
rect 37181 72178 37247 72181
rect 39200 72178 40800 72208
rect 37181 72176 40800 72178
rect 37181 72120 37186 72176
rect 37242 72120 40800 72176
rect 37181 72118 40800 72120
rect 37181 72115 37247 72118
rect 39200 72088 40800 72118
rect 4208 71840 4528 71841
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 71775 4528 71776
rect 34928 71840 35248 71841
rect 34928 71776 34936 71840
rect 35000 71776 35016 71840
rect 35080 71776 35096 71840
rect 35160 71776 35176 71840
rect 35240 71776 35248 71840
rect 34928 71775 35248 71776
rect 38929 71770 38995 71773
rect 39200 71770 40800 71800
rect 38929 71768 40800 71770
rect 38929 71712 38934 71768
rect 38990 71712 40800 71768
rect 38929 71710 40800 71712
rect 38929 71707 38995 71710
rect 39200 71680 40800 71710
rect -800 71498 800 71528
rect 1393 71498 1459 71501
rect -800 71496 1459 71498
rect -800 71440 1398 71496
rect 1454 71440 1459 71496
rect -800 71438 1459 71440
rect -800 71408 800 71438
rect 1393 71435 1459 71438
rect 37457 71362 37523 71365
rect 39200 71362 40800 71392
rect 37457 71360 40800 71362
rect 37457 71304 37462 71360
rect 37518 71304 40800 71360
rect 37457 71302 40800 71304
rect 37457 71299 37523 71302
rect 19568 71296 19888 71297
rect 19568 71232 19576 71296
rect 19640 71232 19656 71296
rect 19720 71232 19736 71296
rect 19800 71232 19816 71296
rect 19880 71232 19888 71296
rect 39200 71272 40800 71302
rect 19568 71231 19888 71232
rect 37365 70818 37431 70821
rect 39200 70818 40800 70848
rect 37365 70816 40800 70818
rect 37365 70760 37370 70816
rect 37426 70760 40800 70816
rect 37365 70758 40800 70760
rect 37365 70755 37431 70758
rect 4208 70752 4528 70753
rect -800 70682 800 70712
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 70687 4528 70688
rect 34928 70752 35248 70753
rect 34928 70688 34936 70752
rect 35000 70688 35016 70752
rect 35080 70688 35096 70752
rect 35160 70688 35176 70752
rect 35240 70688 35248 70752
rect 39200 70728 40800 70758
rect 34928 70687 35248 70688
rect 1393 70682 1459 70685
rect -800 70680 1459 70682
rect -800 70624 1398 70680
rect 1454 70624 1459 70680
rect -800 70622 1459 70624
rect -800 70592 800 70622
rect 1393 70619 1459 70622
rect 37917 70410 37983 70413
rect 38101 70410 38167 70413
rect 37917 70408 38026 70410
rect 37917 70352 37922 70408
rect 37978 70352 38026 70408
rect 37917 70347 38026 70352
rect 38101 70408 39130 70410
rect 38101 70352 38106 70408
rect 38162 70380 39130 70408
rect 39200 70380 40800 70440
rect 38162 70352 40800 70380
rect 38101 70350 40800 70352
rect 38101 70347 38167 70350
rect 19568 70208 19888 70209
rect 19568 70144 19576 70208
rect 19640 70144 19656 70208
rect 19720 70144 19736 70208
rect 19800 70144 19816 70208
rect 19880 70144 19888 70208
rect 19568 70143 19888 70144
rect 37966 70138 38026 70347
rect 39070 70320 40800 70350
rect 38561 70138 38627 70141
rect 37966 70136 38627 70138
rect 37966 70080 38566 70136
rect 38622 70080 38627 70136
rect 37966 70078 38627 70080
rect 38561 70075 38627 70078
rect 36721 70002 36787 70005
rect 39200 70002 40800 70032
rect 36721 70000 40800 70002
rect 36721 69944 36726 70000
rect 36782 69944 40800 70000
rect 36721 69942 40800 69944
rect 36721 69939 36787 69942
rect 39200 69912 40800 69942
rect -800 69866 800 69896
rect 1393 69866 1459 69869
rect -800 69864 1459 69866
rect -800 69808 1398 69864
rect 1454 69808 1459 69864
rect -800 69806 1459 69808
rect -800 69776 800 69806
rect 1393 69803 1459 69806
rect 36905 69866 36971 69869
rect 36905 69864 37290 69866
rect 36905 69808 36910 69864
rect 36966 69808 37290 69864
rect 36905 69806 37290 69808
rect 36905 69803 36971 69806
rect 4208 69664 4528 69665
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 69599 4528 69600
rect 34928 69664 35248 69665
rect 34928 69600 34936 69664
rect 35000 69600 35016 69664
rect 35080 69600 35096 69664
rect 35160 69600 35176 69664
rect 35240 69600 35248 69664
rect 34928 69599 35248 69600
rect 37230 69458 37290 69806
rect 37457 69594 37523 69597
rect 39200 69594 40800 69624
rect 37457 69592 40800 69594
rect 37457 69536 37462 69592
rect 37518 69536 40800 69592
rect 37457 69534 40800 69536
rect 37457 69531 37523 69534
rect 39200 69504 40800 69534
rect 37457 69458 37523 69461
rect 37230 69456 37523 69458
rect 37230 69400 37462 69456
rect 37518 69400 37523 69456
rect 37230 69398 37523 69400
rect 37457 69395 37523 69398
rect 19568 69120 19888 69121
rect -800 69050 800 69080
rect 19568 69056 19576 69120
rect 19640 69056 19656 69120
rect 19720 69056 19736 69120
rect 19800 69056 19816 69120
rect 19880 69056 19888 69120
rect 19568 69055 19888 69056
rect 1393 69050 1459 69053
rect -800 69048 1459 69050
rect -800 68992 1398 69048
rect 1454 68992 1459 69048
rect -800 68990 1459 68992
rect -800 68960 800 68990
rect 1393 68987 1459 68990
rect 37365 69050 37431 69053
rect 39200 69050 40800 69080
rect 37365 69048 40800 69050
rect 37365 68992 37370 69048
rect 37426 68992 40800 69048
rect 37365 68990 40800 68992
rect 37365 68987 37431 68990
rect 39200 68960 40800 68990
rect 37181 68914 37247 68917
rect 37046 68912 37247 68914
rect 37046 68856 37186 68912
rect 37242 68856 37247 68912
rect 37046 68854 37247 68856
rect 37046 68645 37106 68854
rect 37181 68851 37247 68854
rect 36997 68640 37106 68645
rect 36997 68584 37002 68640
rect 37058 68584 37106 68640
rect 36997 68582 37106 68584
rect 38285 68642 38351 68645
rect 39200 68642 40800 68672
rect 38285 68640 40800 68642
rect 38285 68584 38290 68640
rect 38346 68584 40800 68640
rect 38285 68582 40800 68584
rect 36997 68579 37063 68582
rect 38285 68579 38351 68582
rect 4208 68576 4528 68577
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 68511 4528 68512
rect 34928 68576 35248 68577
rect 34928 68512 34936 68576
rect 35000 68512 35016 68576
rect 35080 68512 35096 68576
rect 35160 68512 35176 68576
rect 35240 68512 35248 68576
rect 39200 68552 40800 68582
rect 34928 68511 35248 68512
rect 35341 68506 35407 68509
rect 37365 68506 37431 68509
rect 35341 68504 37431 68506
rect 35341 68448 35346 68504
rect 35402 68448 37370 68504
rect 37426 68448 37431 68504
rect 35341 68446 37431 68448
rect 35341 68443 35407 68446
rect 37365 68443 37431 68446
rect -800 68234 800 68264
rect 1393 68234 1459 68237
rect -800 68232 1459 68234
rect -800 68176 1398 68232
rect 1454 68176 1459 68232
rect -800 68174 1459 68176
rect -800 68144 800 68174
rect 1393 68171 1459 68174
rect 35801 68234 35867 68237
rect 39200 68234 40800 68264
rect 35801 68232 40800 68234
rect 35801 68176 35806 68232
rect 35862 68176 40800 68232
rect 35801 68174 40800 68176
rect 35801 68171 35867 68174
rect 39200 68144 40800 68174
rect 19568 68032 19888 68033
rect 19568 67968 19576 68032
rect 19640 67968 19656 68032
rect 19720 67968 19736 68032
rect 19800 67968 19816 68032
rect 19880 67968 19888 68032
rect 19568 67967 19888 67968
rect 36261 67690 36327 67693
rect 39200 67690 40800 67720
rect 36261 67688 40800 67690
rect 36261 67632 36266 67688
rect 36322 67632 40800 67688
rect 36261 67630 40800 67632
rect 36261 67627 36327 67630
rect 39200 67600 40800 67630
rect 4208 67488 4528 67489
rect -800 67418 800 67448
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 67423 4528 67424
rect 34928 67488 35248 67489
rect 34928 67424 34936 67488
rect 35000 67424 35016 67488
rect 35080 67424 35096 67488
rect 35160 67424 35176 67488
rect 35240 67424 35248 67488
rect 34928 67423 35248 67424
rect 1393 67418 1459 67421
rect -800 67416 1459 67418
rect -800 67360 1398 67416
rect 1454 67360 1459 67416
rect -800 67358 1459 67360
rect -800 67328 800 67358
rect 1393 67355 1459 67358
rect 38377 67282 38443 67285
rect 39200 67282 40800 67312
rect 38377 67280 40800 67282
rect 38377 67224 38382 67280
rect 38438 67224 40800 67280
rect 38377 67222 40800 67224
rect 38377 67219 38443 67222
rect 39200 67192 40800 67222
rect 19568 66944 19888 66945
rect 19568 66880 19576 66944
rect 19640 66880 19656 66944
rect 19720 66880 19736 66944
rect 19800 66880 19816 66944
rect 19880 66880 19888 66944
rect 19568 66879 19888 66880
rect 34789 66874 34855 66877
rect 39200 66874 40800 66904
rect 34789 66872 40800 66874
rect 34789 66816 34794 66872
rect 34850 66816 40800 66872
rect 34789 66814 40800 66816
rect 34789 66811 34855 66814
rect 39200 66784 40800 66814
rect -800 66738 800 66768
rect 1393 66738 1459 66741
rect -800 66736 1459 66738
rect -800 66680 1398 66736
rect 1454 66680 1459 66736
rect -800 66678 1459 66680
rect -800 66648 800 66678
rect 1393 66675 1459 66678
rect 35341 66466 35407 66469
rect 39200 66466 40800 66496
rect 35341 66464 40800 66466
rect 35341 66408 35346 66464
rect 35402 66408 40800 66464
rect 35341 66406 40800 66408
rect 35341 66403 35407 66406
rect 4208 66400 4528 66401
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 66335 4528 66336
rect 34928 66400 35248 66401
rect 34928 66336 34936 66400
rect 35000 66336 35016 66400
rect 35080 66336 35096 66400
rect 35160 66336 35176 66400
rect 35240 66336 35248 66400
rect 39200 66376 40800 66406
rect 34928 66335 35248 66336
rect -800 65922 800 65952
rect 1393 65922 1459 65925
rect -800 65920 1459 65922
rect -800 65864 1398 65920
rect 1454 65864 1459 65920
rect -800 65862 1459 65864
rect -800 65832 800 65862
rect 1393 65859 1459 65862
rect 38193 65922 38259 65925
rect 39200 65922 40800 65952
rect 38193 65920 40800 65922
rect 38193 65864 38198 65920
rect 38254 65864 40800 65920
rect 38193 65862 40800 65864
rect 38193 65859 38259 65862
rect 19568 65856 19888 65857
rect 19568 65792 19576 65856
rect 19640 65792 19656 65856
rect 19720 65792 19736 65856
rect 19800 65792 19816 65856
rect 19880 65792 19888 65856
rect 39200 65832 40800 65862
rect 19568 65791 19888 65792
rect 35065 65514 35131 65517
rect 39200 65514 40800 65544
rect 35065 65512 40800 65514
rect 35065 65456 35070 65512
rect 35126 65456 40800 65512
rect 35065 65454 40800 65456
rect 35065 65451 35131 65454
rect 39200 65424 40800 65454
rect 4208 65312 4528 65313
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 65247 4528 65248
rect 34928 65312 35248 65313
rect 34928 65248 34936 65312
rect 35000 65248 35016 65312
rect 35080 65248 35096 65312
rect 35160 65248 35176 65312
rect 35240 65248 35248 65312
rect 34928 65247 35248 65248
rect -800 65106 800 65136
rect 1393 65106 1459 65109
rect -800 65104 1459 65106
rect -800 65048 1398 65104
rect 1454 65048 1459 65104
rect -800 65046 1459 65048
rect -800 65016 800 65046
rect 1393 65043 1459 65046
rect 34789 65106 34855 65109
rect 39200 65106 40800 65136
rect 34789 65104 40800 65106
rect 34789 65048 34794 65104
rect 34850 65048 40800 65104
rect 34789 65046 40800 65048
rect 34789 65043 34855 65046
rect 39200 65016 40800 65046
rect 35065 64970 35131 64973
rect 37641 64970 37707 64973
rect 35065 64968 37707 64970
rect 35065 64912 35070 64968
rect 35126 64912 37646 64968
rect 37702 64912 37707 64968
rect 35065 64910 37707 64912
rect 35065 64907 35131 64910
rect 37641 64907 37707 64910
rect 35249 64834 35315 64837
rect 35206 64832 35315 64834
rect 35206 64776 35254 64832
rect 35310 64776 35315 64832
rect 35206 64771 35315 64776
rect 36905 64834 36971 64837
rect 38653 64834 38719 64837
rect 36905 64832 38719 64834
rect 36905 64776 36910 64832
rect 36966 64776 38658 64832
rect 38714 64776 38719 64832
rect 36905 64774 38719 64776
rect 36905 64771 36971 64774
rect 38653 64771 38719 64774
rect 19568 64768 19888 64769
rect 19568 64704 19576 64768
rect 19640 64704 19656 64768
rect 19720 64704 19736 64768
rect 19800 64704 19816 64768
rect 19880 64704 19888 64768
rect 19568 64703 19888 64704
rect 35206 64565 35266 64771
rect 35433 64698 35499 64701
rect 37549 64698 37615 64701
rect 35433 64696 37615 64698
rect 35433 64640 35438 64696
rect 35494 64640 37554 64696
rect 37610 64640 37615 64696
rect 35433 64638 37615 64640
rect 35433 64635 35499 64638
rect 37549 64635 37615 64638
rect 35206 64560 35315 64565
rect 35206 64504 35254 64560
rect 35310 64504 35315 64560
rect 35206 64502 35315 64504
rect 35249 64499 35315 64502
rect 35709 64562 35775 64565
rect 39200 64562 40800 64592
rect 35709 64560 40800 64562
rect 35709 64504 35714 64560
rect 35770 64504 40800 64560
rect 35709 64502 40800 64504
rect 35709 64499 35775 64502
rect 39200 64472 40800 64502
rect 34881 64426 34947 64429
rect 34470 64424 34947 64426
rect 34470 64368 34886 64424
rect 34942 64368 34947 64424
rect 34470 64366 34947 64368
rect -800 64290 800 64320
rect 1393 64290 1459 64293
rect -800 64288 1459 64290
rect -800 64232 1398 64288
rect 1454 64232 1459 64288
rect -800 64230 1459 64232
rect -800 64200 800 64230
rect 1393 64227 1459 64230
rect 4208 64224 4528 64225
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 64159 4528 64160
rect 34470 63882 34530 64366
rect 34881 64363 34947 64366
rect 36077 64426 36143 64429
rect 36353 64426 36419 64429
rect 36077 64424 36419 64426
rect 36077 64368 36082 64424
rect 36138 64368 36358 64424
rect 36414 64368 36419 64424
rect 36077 64366 36419 64368
rect 36077 64363 36143 64366
rect 36353 64363 36419 64366
rect 34928 64224 35248 64225
rect 34928 64160 34936 64224
rect 35000 64160 35016 64224
rect 35080 64160 35096 64224
rect 35160 64160 35176 64224
rect 35240 64160 35248 64224
rect 34928 64159 35248 64160
rect 35341 64154 35407 64157
rect 39200 64154 40800 64184
rect 35341 64152 40800 64154
rect 35341 64096 35346 64152
rect 35402 64096 40800 64152
rect 35341 64094 40800 64096
rect 35341 64091 35407 64094
rect 39200 64064 40800 64094
rect 34605 64018 34671 64021
rect 36905 64018 36971 64021
rect 34605 64016 36971 64018
rect 34605 63960 34610 64016
rect 34666 63960 36910 64016
rect 36966 63960 36971 64016
rect 34605 63958 36971 63960
rect 34605 63955 34671 63958
rect 36905 63955 36971 63958
rect 35157 63882 35223 63885
rect 34470 63880 35223 63882
rect 34470 63824 35162 63880
rect 35218 63824 35223 63880
rect 34470 63822 35223 63824
rect 35157 63819 35223 63822
rect 35525 63882 35591 63885
rect 37273 63882 37339 63885
rect 35525 63880 37339 63882
rect 35525 63824 35530 63880
rect 35586 63824 37278 63880
rect 37334 63824 37339 63880
rect 35525 63822 37339 63824
rect 35525 63819 35591 63822
rect 37273 63819 37339 63822
rect 36445 63746 36511 63749
rect 39200 63746 40800 63776
rect 36445 63744 40800 63746
rect 36445 63688 36450 63744
rect 36506 63688 40800 63744
rect 36445 63686 40800 63688
rect 36445 63683 36511 63686
rect 19568 63680 19888 63681
rect 19568 63616 19576 63680
rect 19640 63616 19656 63680
rect 19720 63616 19736 63680
rect 19800 63616 19816 63680
rect 19880 63616 19888 63680
rect 39200 63656 40800 63686
rect 19568 63615 19888 63616
rect 35801 63610 35867 63613
rect 36721 63610 36787 63613
rect 37641 63610 37707 63613
rect 35801 63608 37707 63610
rect 35801 63552 35806 63608
rect 35862 63552 36726 63608
rect 36782 63552 37646 63608
rect 37702 63552 37707 63608
rect 35801 63550 37707 63552
rect 35801 63547 35867 63550
rect 36721 63547 36787 63550
rect 37641 63547 37707 63550
rect -800 63474 800 63504
rect 1393 63474 1459 63477
rect -800 63472 1459 63474
rect -800 63416 1398 63472
rect 1454 63416 1459 63472
rect -800 63414 1459 63416
rect -800 63384 800 63414
rect 1393 63411 1459 63414
rect 35801 63474 35867 63477
rect 37549 63474 37615 63477
rect 35801 63472 37615 63474
rect 35801 63416 35806 63472
rect 35862 63416 37554 63472
rect 37610 63416 37615 63472
rect 35801 63414 37615 63416
rect 35801 63411 35867 63414
rect 37549 63411 37615 63414
rect 34789 63338 34855 63341
rect 39200 63338 40800 63368
rect 34789 63336 40800 63338
rect 34789 63280 34794 63336
rect 34850 63280 40800 63336
rect 34789 63278 40800 63280
rect 34789 63275 34855 63278
rect 39200 63248 40800 63278
rect 4208 63136 4528 63137
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 63071 4528 63072
rect 34928 63136 35248 63137
rect 34928 63072 34936 63136
rect 35000 63072 35016 63136
rect 35080 63072 35096 63136
rect 35160 63072 35176 63136
rect 35240 63072 35248 63136
rect 34928 63071 35248 63072
rect 36077 63066 36143 63069
rect 39757 63066 39823 63069
rect 36077 63064 39823 63066
rect 36077 63008 36082 63064
rect 36138 63008 39762 63064
rect 39818 63008 39823 63064
rect 36077 63006 39823 63008
rect 36077 63003 36143 63006
rect 39757 63003 39823 63006
rect 33593 62930 33659 62933
rect 37273 62930 37339 62933
rect 33593 62928 37339 62930
rect 33593 62872 33598 62928
rect 33654 62872 37278 62928
rect 37334 62872 37339 62928
rect 33593 62870 37339 62872
rect 33593 62867 33659 62870
rect 37273 62867 37339 62870
rect 35709 62794 35775 62797
rect 39200 62794 40800 62824
rect 35709 62792 40800 62794
rect 35709 62736 35714 62792
rect 35770 62736 40800 62792
rect 35709 62734 40800 62736
rect 35709 62731 35775 62734
rect 39200 62704 40800 62734
rect -800 62658 800 62688
rect 1393 62658 1459 62661
rect -800 62656 1459 62658
rect -800 62600 1398 62656
rect 1454 62600 1459 62656
rect -800 62598 1459 62600
rect -800 62568 800 62598
rect 1393 62595 1459 62598
rect 19568 62592 19888 62593
rect 19568 62528 19576 62592
rect 19640 62528 19656 62592
rect 19720 62528 19736 62592
rect 19800 62528 19816 62592
rect 19880 62528 19888 62592
rect 19568 62527 19888 62528
rect 36261 62386 36327 62389
rect 39200 62386 40800 62416
rect 36261 62384 40800 62386
rect 36261 62328 36266 62384
rect 36322 62328 40800 62384
rect 36261 62326 40800 62328
rect 36261 62323 36327 62326
rect 39200 62296 40800 62326
rect 36721 62250 36787 62253
rect 37457 62250 37523 62253
rect 36721 62248 37523 62250
rect 36721 62192 36726 62248
rect 36782 62192 37462 62248
rect 37518 62192 37523 62248
rect 36721 62190 37523 62192
rect 36721 62187 36787 62190
rect 37457 62187 37523 62190
rect 4208 62048 4528 62049
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 61983 4528 61984
rect 34928 62048 35248 62049
rect 34928 61984 34936 62048
rect 35000 61984 35016 62048
rect 35080 61984 35096 62048
rect 35160 61984 35176 62048
rect 35240 61984 35248 62048
rect 34928 61983 35248 61984
rect 36721 61978 36787 61981
rect 39200 61978 40800 62008
rect 36721 61976 40800 61978
rect 36721 61920 36726 61976
rect 36782 61920 40800 61976
rect 36721 61918 40800 61920
rect 36721 61915 36787 61918
rect 39200 61888 40800 61918
rect -800 61842 800 61872
rect 1393 61842 1459 61845
rect -800 61840 1459 61842
rect -800 61784 1398 61840
rect 1454 61784 1459 61840
rect -800 61782 1459 61784
rect -800 61752 800 61782
rect 1393 61779 1459 61782
rect 19568 61504 19888 61505
rect 19568 61440 19576 61504
rect 19640 61440 19656 61504
rect 19720 61440 19736 61504
rect 19800 61440 19816 61504
rect 19880 61440 19888 61504
rect 19568 61439 19888 61440
rect 34881 61434 34947 61437
rect 39200 61434 40800 61464
rect 34881 61432 40800 61434
rect 34881 61376 34886 61432
rect 34942 61376 40800 61432
rect 34881 61374 40800 61376
rect 34881 61371 34947 61374
rect 39200 61344 40800 61374
rect -800 61026 800 61056
rect 1393 61026 1459 61029
rect -800 61024 1459 61026
rect -800 60968 1398 61024
rect 1454 60968 1459 61024
rect -800 60966 1459 60968
rect -800 60936 800 60966
rect 1393 60963 1459 60966
rect 35801 61026 35867 61029
rect 39200 61026 40800 61056
rect 35801 61024 40800 61026
rect 35801 60968 35806 61024
rect 35862 60968 40800 61024
rect 35801 60966 40800 60968
rect 35801 60963 35867 60966
rect 4208 60960 4528 60961
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 60895 4528 60896
rect 34928 60960 35248 60961
rect 34928 60896 34936 60960
rect 35000 60896 35016 60960
rect 35080 60896 35096 60960
rect 35160 60896 35176 60960
rect 35240 60896 35248 60960
rect 39200 60936 40800 60966
rect 34928 60895 35248 60896
rect 35157 60618 35223 60621
rect 39200 60618 40800 60648
rect 35157 60616 40800 60618
rect 35157 60560 35162 60616
rect 35218 60560 40800 60616
rect 35157 60558 40800 60560
rect 35157 60555 35223 60558
rect 39200 60528 40800 60558
rect 19568 60416 19888 60417
rect -800 60346 800 60376
rect 19568 60352 19576 60416
rect 19640 60352 19656 60416
rect 19720 60352 19736 60416
rect 19800 60352 19816 60416
rect 19880 60352 19888 60416
rect 19568 60351 19888 60352
rect 1393 60346 1459 60349
rect -800 60344 1459 60346
rect -800 60288 1398 60344
rect 1454 60288 1459 60344
rect -800 60286 1459 60288
rect -800 60256 800 60286
rect 1393 60283 1459 60286
rect 35157 60210 35223 60213
rect 39200 60210 40800 60240
rect 35157 60208 40800 60210
rect 35157 60152 35162 60208
rect 35218 60152 40800 60208
rect 35157 60150 40800 60152
rect 35157 60147 35223 60150
rect 39200 60120 40800 60150
rect 4208 59872 4528 59873
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 59807 4528 59808
rect 34928 59872 35248 59873
rect 34928 59808 34936 59872
rect 35000 59808 35016 59872
rect 35080 59808 35096 59872
rect 35160 59808 35176 59872
rect 35240 59808 35248 59872
rect 34928 59807 35248 59808
rect 34789 59666 34855 59669
rect 39200 59666 40800 59696
rect 34789 59664 40800 59666
rect 34789 59608 34794 59664
rect 34850 59608 40800 59664
rect 34789 59606 40800 59608
rect 34789 59603 34855 59606
rect 39200 59576 40800 59606
rect -800 59530 800 59560
rect 1393 59530 1459 59533
rect -800 59528 1459 59530
rect -800 59472 1398 59528
rect 1454 59472 1459 59528
rect -800 59470 1459 59472
rect -800 59440 800 59470
rect 1393 59467 1459 59470
rect 35249 59530 35315 59533
rect 37825 59530 37891 59533
rect 35249 59528 37891 59530
rect 35249 59472 35254 59528
rect 35310 59472 37830 59528
rect 37886 59472 37891 59528
rect 35249 59470 37891 59472
rect 35249 59467 35315 59470
rect 37825 59467 37891 59470
rect 19568 59328 19888 59329
rect 19568 59264 19576 59328
rect 19640 59264 19656 59328
rect 19720 59264 19736 59328
rect 19800 59264 19816 59328
rect 19880 59264 19888 59328
rect 19568 59263 19888 59264
rect 35801 59258 35867 59261
rect 39200 59258 40800 59288
rect 35801 59256 40800 59258
rect 35801 59200 35806 59256
rect 35862 59200 40800 59256
rect 35801 59198 40800 59200
rect 35801 59195 35867 59198
rect 39200 59168 40800 59198
rect 36813 58850 36879 58853
rect 39200 58850 40800 58880
rect 36813 58848 40800 58850
rect 36813 58792 36818 58848
rect 36874 58792 40800 58848
rect 36813 58790 40800 58792
rect 36813 58787 36879 58790
rect 4208 58784 4528 58785
rect -800 58714 800 58744
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 58719 4528 58720
rect 34928 58784 35248 58785
rect 34928 58720 34936 58784
rect 35000 58720 35016 58784
rect 35080 58720 35096 58784
rect 35160 58720 35176 58784
rect 35240 58720 35248 58784
rect 39200 58760 40800 58790
rect 34928 58719 35248 58720
rect 1393 58714 1459 58717
rect -800 58712 1459 58714
rect -800 58656 1398 58712
rect 1454 58656 1459 58712
rect -800 58654 1459 58656
rect -800 58624 800 58654
rect 1393 58651 1459 58654
rect 36261 58578 36327 58581
rect 36445 58578 36511 58581
rect 36261 58576 36511 58578
rect 36261 58520 36266 58576
rect 36322 58520 36450 58576
rect 36506 58520 36511 58576
rect 36261 58518 36511 58520
rect 36261 58515 36327 58518
rect 36445 58515 36511 58518
rect 36721 58306 36787 58309
rect 39200 58306 40800 58336
rect 36721 58304 40800 58306
rect 36721 58248 36726 58304
rect 36782 58248 40800 58304
rect 36721 58246 40800 58248
rect 36721 58243 36787 58246
rect 19568 58240 19888 58241
rect 19568 58176 19576 58240
rect 19640 58176 19656 58240
rect 19720 58176 19736 58240
rect 19800 58176 19816 58240
rect 19880 58176 19888 58240
rect 39200 58216 40800 58246
rect 19568 58175 19888 58176
rect -800 57898 800 57928
rect 1393 57898 1459 57901
rect -800 57896 1459 57898
rect -800 57840 1398 57896
rect 1454 57840 1459 57896
rect -800 57838 1459 57840
rect -800 57808 800 57838
rect 1393 57835 1459 57838
rect 37181 57898 37247 57901
rect 39200 57898 40800 57928
rect 37181 57896 40800 57898
rect 37181 57840 37186 57896
rect 37242 57840 40800 57896
rect 37181 57838 40800 57840
rect 37181 57835 37247 57838
rect 39200 57808 40800 57838
rect 4208 57696 4528 57697
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 57631 4528 57632
rect 34928 57696 35248 57697
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 57631 35248 57632
rect 37457 57490 37523 57493
rect 39200 57490 40800 57520
rect 37457 57488 40800 57490
rect 37457 57432 37462 57488
rect 37518 57432 40800 57488
rect 37457 57430 40800 57432
rect 37457 57427 37523 57430
rect 39200 57400 40800 57430
rect 19568 57152 19888 57153
rect -800 57082 800 57112
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 19568 57087 19888 57088
rect 1393 57082 1459 57085
rect -800 57080 1459 57082
rect -800 57024 1398 57080
rect 1454 57024 1459 57080
rect -800 57022 1459 57024
rect -800 56992 800 57022
rect 1393 57019 1459 57022
rect 37917 56946 37983 56949
rect 39200 56946 40800 56976
rect 37917 56944 40800 56946
rect 37917 56888 37922 56944
rect 37978 56888 40800 56944
rect 37917 56886 40800 56888
rect 37917 56883 37983 56886
rect 39200 56856 40800 56886
rect 4208 56608 4528 56609
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 56543 4528 56544
rect 34928 56608 35248 56609
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 34928 56543 35248 56544
rect 37917 56538 37983 56541
rect 39200 56538 40800 56568
rect 37917 56536 40800 56538
rect 37917 56480 37922 56536
rect 37978 56480 40800 56536
rect 37917 56478 40800 56480
rect 37917 56475 37983 56478
rect 39200 56448 40800 56478
rect -800 56266 800 56296
rect 1393 56266 1459 56269
rect -800 56264 1459 56266
rect -800 56208 1398 56264
rect 1454 56208 1459 56264
rect -800 56206 1459 56208
rect -800 56176 800 56206
rect 1393 56203 1459 56206
rect 37457 56130 37523 56133
rect 39200 56130 40800 56160
rect 37457 56128 40800 56130
rect 37457 56072 37462 56128
rect 37518 56072 40800 56128
rect 37457 56070 40800 56072
rect 37457 56067 37523 56070
rect 19568 56064 19888 56065
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 39200 56040 40800 56070
rect 19568 55999 19888 56000
rect 37181 55722 37247 55725
rect 39200 55722 40800 55752
rect 37181 55720 40800 55722
rect 37181 55664 37186 55720
rect 37242 55664 40800 55720
rect 37181 55662 40800 55664
rect 37181 55659 37247 55662
rect 39200 55632 40800 55662
rect 4208 55520 4528 55521
rect -800 55450 800 55480
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 55455 4528 55456
rect 34928 55520 35248 55521
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 55455 35248 55456
rect 1393 55450 1459 55453
rect -800 55448 1459 55450
rect -800 55392 1398 55448
rect 1454 55392 1459 55448
rect -800 55390 1459 55392
rect -800 55360 800 55390
rect 1393 55387 1459 55390
rect 37917 55178 37983 55181
rect 39200 55178 40800 55208
rect 37917 55176 40800 55178
rect 37917 55120 37922 55176
rect 37978 55120 40800 55176
rect 37917 55118 40800 55120
rect 37917 55115 37983 55118
rect 39200 55088 40800 55118
rect 19568 54976 19888 54977
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 19568 54911 19888 54912
rect 37457 54770 37523 54773
rect 39200 54770 40800 54800
rect 37457 54768 40800 54770
rect 37457 54712 37462 54768
rect 37518 54712 40800 54768
rect 37457 54710 40800 54712
rect 37457 54707 37523 54710
rect 39200 54680 40800 54710
rect -800 54634 800 54664
rect 1393 54634 1459 54637
rect -800 54632 1459 54634
rect -800 54576 1398 54632
rect 1454 54576 1459 54632
rect -800 54574 1459 54576
rect -800 54544 800 54574
rect 1393 54571 1459 54574
rect 4208 54432 4528 54433
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 54367 4528 54368
rect 34928 54432 35248 54433
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 34928 54367 35248 54368
rect 37181 54362 37247 54365
rect 39200 54362 40800 54392
rect 37181 54360 40800 54362
rect 37181 54304 37186 54360
rect 37242 54304 40800 54360
rect 37181 54302 40800 54304
rect 37181 54299 37247 54302
rect 39200 54272 40800 54302
rect 19568 53888 19888 53889
rect -800 53818 800 53848
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 53823 19888 53824
rect 1393 53818 1459 53821
rect -800 53816 1459 53818
rect -800 53760 1398 53816
rect 1454 53760 1459 53816
rect -800 53758 1459 53760
rect -800 53728 800 53758
rect 1393 53755 1459 53758
rect 37181 53818 37247 53821
rect 39200 53818 40800 53848
rect 37181 53816 40800 53818
rect 37181 53760 37186 53816
rect 37242 53760 40800 53816
rect 37181 53758 40800 53760
rect 37181 53755 37247 53758
rect 39200 53728 40800 53758
rect 36721 53410 36787 53413
rect 39200 53410 40800 53440
rect 36721 53408 40800 53410
rect 36721 53352 36726 53408
rect 36782 53352 40800 53408
rect 36721 53350 40800 53352
rect 36721 53347 36787 53350
rect 4208 53344 4528 53345
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 53279 4528 53280
rect 34928 53344 35248 53345
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 39200 53320 40800 53350
rect 34928 53279 35248 53280
rect -800 53138 800 53168
rect 1393 53138 1459 53141
rect -800 53136 1459 53138
rect -800 53080 1398 53136
rect 1454 53080 1459 53136
rect -800 53078 1459 53080
rect -800 53048 800 53078
rect 1393 53075 1459 53078
rect 37273 53002 37339 53005
rect 39200 53002 40800 53032
rect 37273 53000 40800 53002
rect 37273 52944 37278 53000
rect 37334 52944 40800 53000
rect 37273 52942 40800 52944
rect 37273 52939 37339 52942
rect 39200 52912 40800 52942
rect 19568 52800 19888 52801
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 19568 52735 19888 52736
rect 37917 52594 37983 52597
rect 39200 52594 40800 52624
rect 37917 52592 40800 52594
rect 37917 52536 37922 52592
rect 37978 52536 40800 52592
rect 37917 52534 40800 52536
rect 37917 52531 37983 52534
rect 39200 52504 40800 52534
rect -800 52322 800 52352
rect 1393 52322 1459 52325
rect -800 52320 1459 52322
rect -800 52264 1398 52320
rect 1454 52264 1459 52320
rect -800 52262 1459 52264
rect -800 52232 800 52262
rect 1393 52259 1459 52262
rect 4208 52256 4528 52257
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 52191 4528 52192
rect 34928 52256 35248 52257
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 34928 52191 35248 52192
rect 37457 52050 37523 52053
rect 39200 52050 40800 52080
rect 37457 52048 40800 52050
rect 37457 51992 37462 52048
rect 37518 51992 40800 52048
rect 37457 51990 40800 51992
rect 37457 51987 37523 51990
rect 39200 51960 40800 51990
rect 19568 51712 19888 51713
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 51647 19888 51648
rect 37181 51642 37247 51645
rect 39200 51642 40800 51672
rect 37181 51640 40800 51642
rect 37181 51584 37186 51640
rect 37242 51584 40800 51640
rect 37181 51582 40800 51584
rect 37181 51579 37247 51582
rect 39200 51552 40800 51582
rect -800 51506 800 51536
rect 1393 51506 1459 51509
rect -800 51504 1459 51506
rect -800 51448 1398 51504
rect 1454 51448 1459 51504
rect -800 51446 1459 51448
rect -800 51416 800 51446
rect 1393 51443 1459 51446
rect 37917 51234 37983 51237
rect 39200 51234 40800 51264
rect 37917 51232 40800 51234
rect 37917 51176 37922 51232
rect 37978 51176 40800 51232
rect 37917 51174 40800 51176
rect 37917 51171 37983 51174
rect 4208 51168 4528 51169
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 51103 4528 51104
rect 34928 51168 35248 51169
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 39200 51144 40800 51174
rect 34928 51103 35248 51104
rect -800 50690 800 50720
rect 1853 50690 1919 50693
rect -800 50688 1919 50690
rect -800 50632 1858 50688
rect 1914 50632 1919 50688
rect -800 50630 1919 50632
rect -800 50600 800 50630
rect 1853 50627 1919 50630
rect 37457 50690 37523 50693
rect 39200 50690 40800 50720
rect 37457 50688 40800 50690
rect 37457 50632 37462 50688
rect 37518 50632 40800 50688
rect 37457 50630 40800 50632
rect 37457 50627 37523 50630
rect 19568 50624 19888 50625
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 39200 50600 40800 50630
rect 19568 50559 19888 50560
rect 37917 50282 37983 50285
rect 39200 50282 40800 50312
rect 37917 50280 40800 50282
rect 37917 50224 37922 50280
rect 37978 50224 40800 50280
rect 37917 50222 40800 50224
rect 37917 50219 37983 50222
rect 39200 50192 40800 50222
rect 4208 50080 4528 50081
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 50015 4528 50016
rect 34928 50080 35248 50081
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 50015 35248 50016
rect -800 49874 800 49904
rect 1853 49874 1919 49877
rect -800 49872 1919 49874
rect -800 49816 1858 49872
rect 1914 49816 1919 49872
rect -800 49814 1919 49816
rect -800 49784 800 49814
rect 1853 49811 1919 49814
rect 37917 49874 37983 49877
rect 39200 49874 40800 49904
rect 37917 49872 40800 49874
rect 37917 49816 37922 49872
rect 37978 49816 40800 49872
rect 37917 49814 40800 49816
rect 37917 49811 37983 49814
rect 39200 49784 40800 49814
rect 19568 49536 19888 49537
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 49471 19888 49472
rect 37365 49466 37431 49469
rect 39200 49466 40800 49496
rect 37365 49464 40800 49466
rect 37365 49408 37370 49464
rect 37426 49408 40800 49464
rect 37365 49406 40800 49408
rect 37365 49403 37431 49406
rect 39200 49376 40800 49406
rect -800 49058 800 49088
rect 1853 49058 1919 49061
rect -800 49056 1919 49058
rect -800 49000 1858 49056
rect 1914 49000 1919 49056
rect -800 48998 1919 49000
rect -800 48968 800 48998
rect 1853 48995 1919 48998
rect 4208 48992 4528 48993
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 48927 4528 48928
rect 34928 48992 35248 48993
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 34928 48927 35248 48928
rect 37273 48922 37339 48925
rect 39200 48922 40800 48952
rect 37273 48920 40800 48922
rect 37273 48864 37278 48920
rect 37334 48864 40800 48920
rect 37273 48862 40800 48864
rect 37273 48859 37339 48862
rect 39200 48832 40800 48862
rect 37917 48514 37983 48517
rect 39200 48514 40800 48544
rect 37917 48512 40800 48514
rect 37917 48456 37922 48512
rect 37978 48456 40800 48512
rect 37917 48454 40800 48456
rect 37917 48451 37983 48454
rect 19568 48448 19888 48449
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 39200 48424 40800 48454
rect 19568 48383 19888 48384
rect -800 48242 800 48272
rect 1853 48242 1919 48245
rect -800 48240 1919 48242
rect -800 48184 1858 48240
rect 1914 48184 1919 48240
rect -800 48182 1919 48184
rect -800 48152 800 48182
rect 1853 48179 1919 48182
rect 37365 48106 37431 48109
rect 39200 48106 40800 48136
rect 37365 48104 40800 48106
rect 37365 48048 37370 48104
rect 37426 48048 40800 48104
rect 37365 48046 40800 48048
rect 37365 48043 37431 48046
rect 39200 48016 40800 48046
rect 4208 47904 4528 47905
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 47839 4528 47840
rect 34928 47904 35248 47905
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 47839 35248 47840
rect 37273 47562 37339 47565
rect 39200 47562 40800 47592
rect 37273 47560 40800 47562
rect 37273 47504 37278 47560
rect 37334 47504 40800 47560
rect 37273 47502 40800 47504
rect 37273 47499 37339 47502
rect 39200 47472 40800 47502
rect -800 47426 800 47456
rect 1853 47426 1919 47429
rect -800 47424 1919 47426
rect -800 47368 1858 47424
rect 1914 47368 1919 47424
rect -800 47366 1919 47368
rect -800 47336 800 47366
rect 1853 47363 1919 47366
rect 19568 47360 19888 47361
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 47295 19888 47296
rect 37917 47154 37983 47157
rect 39200 47154 40800 47184
rect 37917 47152 40800 47154
rect 37917 47096 37922 47152
rect 37978 47096 40800 47152
rect 37917 47094 40800 47096
rect 37917 47091 37983 47094
rect 39200 47064 40800 47094
rect 4208 46816 4528 46817
rect -800 46746 800 46776
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 34928 46816 35248 46817
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 46751 35248 46752
rect 1853 46746 1919 46749
rect -800 46744 1919 46746
rect -800 46688 1858 46744
rect 1914 46688 1919 46744
rect -800 46686 1919 46688
rect -800 46656 800 46686
rect 1853 46683 1919 46686
rect 35341 46746 35407 46749
rect 35801 46746 35867 46749
rect 35341 46744 35867 46746
rect 35341 46688 35346 46744
rect 35402 46688 35806 46744
rect 35862 46688 35867 46744
rect 35341 46686 35867 46688
rect 35341 46683 35407 46686
rect 35801 46683 35867 46686
rect 37457 46746 37523 46749
rect 39200 46746 40800 46776
rect 37457 46744 40800 46746
rect 37457 46688 37462 46744
rect 37518 46688 40800 46744
rect 37457 46686 40800 46688
rect 37457 46683 37523 46686
rect 39200 46656 40800 46686
rect 19568 46272 19888 46273
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 46207 19888 46208
rect 37181 46202 37247 46205
rect 39200 46202 40800 46232
rect 37181 46200 40800 46202
rect 37181 46144 37186 46200
rect 37242 46144 40800 46200
rect 37181 46142 40800 46144
rect 37181 46139 37247 46142
rect 39200 46112 40800 46142
rect -800 45930 800 45960
rect 1853 45930 1919 45933
rect -800 45928 1919 45930
rect -800 45872 1858 45928
rect 1914 45872 1919 45928
rect -800 45870 1919 45872
rect -800 45840 800 45870
rect 1853 45867 1919 45870
rect 37917 45794 37983 45797
rect 39200 45794 40800 45824
rect 37917 45792 40800 45794
rect 37917 45736 37922 45792
rect 37978 45736 40800 45792
rect 37917 45734 40800 45736
rect 37917 45731 37983 45734
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 34928 45728 35248 45729
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 39200 45704 40800 45734
rect 34928 45663 35248 45664
rect 37457 45386 37523 45389
rect 39200 45386 40800 45416
rect 37457 45384 40800 45386
rect 37457 45328 37462 45384
rect 37518 45328 40800 45384
rect 37457 45326 40800 45328
rect 37457 45323 37523 45326
rect 39200 45296 40800 45326
rect 19568 45184 19888 45185
rect -800 45114 800 45144
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 45119 19888 45120
rect 1853 45114 1919 45117
rect -800 45112 1919 45114
rect -800 45056 1858 45112
rect 1914 45056 1919 45112
rect -800 45054 1919 45056
rect -800 45024 800 45054
rect 1853 45051 1919 45054
rect 37917 44978 37983 44981
rect 39200 44978 40800 45008
rect 37917 44976 40800 44978
rect 37917 44920 37922 44976
rect 37978 44920 40800 44976
rect 37917 44918 40800 44920
rect 37917 44915 37983 44918
rect 39200 44888 40800 44918
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 34928 44640 35248 44641
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 44575 35248 44576
rect 37917 44434 37983 44437
rect 39200 44434 40800 44464
rect 37917 44432 40800 44434
rect 37917 44376 37922 44432
rect 37978 44376 40800 44432
rect 37917 44374 40800 44376
rect 37917 44371 37983 44374
rect 39200 44344 40800 44374
rect -800 44298 800 44328
rect 1853 44298 1919 44301
rect -800 44296 1919 44298
rect -800 44240 1858 44296
rect 1914 44240 1919 44296
rect -800 44238 1919 44240
rect -800 44208 800 44238
rect 1853 44235 1919 44238
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 44031 19888 44032
rect 37181 44026 37247 44029
rect 39200 44026 40800 44056
rect 37181 44024 40800 44026
rect 37181 43968 37186 44024
rect 37242 43968 40800 44024
rect 37181 43966 40800 43968
rect 37181 43963 37247 43966
rect 39200 43936 40800 43966
rect 37181 43618 37247 43621
rect 39200 43618 40800 43648
rect 37181 43616 40800 43618
rect 37181 43560 37186 43616
rect 37242 43560 40800 43616
rect 37181 43558 40800 43560
rect 37181 43555 37247 43558
rect 4208 43552 4528 43553
rect -800 43482 800 43512
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 39200 43528 40800 43558
rect 34928 43487 35248 43488
rect 1853 43482 1919 43485
rect -800 43480 1919 43482
rect -800 43424 1858 43480
rect 1914 43424 1919 43480
rect -800 43422 1919 43424
rect -800 43392 800 43422
rect 1853 43419 1919 43422
rect 37917 43074 37983 43077
rect 39200 43074 40800 43104
rect 37917 43072 40800 43074
rect 37917 43016 37922 43072
rect 37978 43016 40800 43072
rect 37917 43014 40800 43016
rect 37917 43011 37983 43014
rect 19568 43008 19888 43009
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 39200 42984 40800 43014
rect 19568 42943 19888 42944
rect -800 42666 800 42696
rect 1853 42666 1919 42669
rect -800 42664 1919 42666
rect -800 42608 1858 42664
rect 1914 42608 1919 42664
rect -800 42606 1919 42608
rect -800 42576 800 42606
rect 1853 42603 1919 42606
rect 37365 42666 37431 42669
rect 39200 42666 40800 42696
rect 37365 42664 40800 42666
rect 37365 42608 37370 42664
rect 37426 42608 40800 42664
rect 37365 42606 40800 42608
rect 37365 42603 37431 42606
rect 39200 42576 40800 42606
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 42399 35248 42400
rect 37273 42258 37339 42261
rect 39200 42258 40800 42288
rect 37273 42256 40800 42258
rect 37273 42200 37278 42256
rect 37334 42200 40800 42256
rect 37273 42198 40800 42200
rect 37273 42195 37339 42198
rect 39200 42168 40800 42198
rect 19568 41920 19888 41921
rect -800 41850 800 41880
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 41855 19888 41856
rect 1853 41850 1919 41853
rect -800 41848 1919 41850
rect -800 41792 1858 41848
rect 1914 41792 1919 41848
rect -800 41790 1919 41792
rect -800 41760 800 41790
rect 1853 41787 1919 41790
rect 37917 41850 37983 41853
rect 39200 41850 40800 41880
rect 37917 41848 40800 41850
rect 37917 41792 37922 41848
rect 37978 41792 40800 41848
rect 37917 41790 40800 41792
rect 37917 41787 37983 41790
rect 39200 41760 40800 41790
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 41311 35248 41312
rect 37181 41306 37247 41309
rect 39200 41306 40800 41336
rect 37181 41304 40800 41306
rect 37181 41248 37186 41304
rect 37242 41248 40800 41304
rect 37181 41246 40800 41248
rect 37181 41243 37247 41246
rect 39200 41216 40800 41246
rect -800 41034 800 41064
rect 1853 41034 1919 41037
rect -800 41032 1919 41034
rect -800 40976 1858 41032
rect 1914 40976 1919 41032
rect -800 40974 1919 40976
rect -800 40944 800 40974
rect 1853 40971 1919 40974
rect 37273 40898 37339 40901
rect 39200 40898 40800 40928
rect 37273 40896 40800 40898
rect 37273 40840 37278 40896
rect 37334 40840 40800 40896
rect 37273 40838 40800 40840
rect 37273 40835 37339 40838
rect 19568 40832 19888 40833
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 39200 40808 40800 40838
rect 19568 40767 19888 40768
rect 37917 40490 37983 40493
rect 39200 40490 40800 40520
rect 37917 40488 40800 40490
rect 37917 40432 37922 40488
rect 37978 40432 40800 40488
rect 37917 40430 40800 40432
rect 37917 40427 37983 40430
rect 39200 40400 40800 40430
rect -800 40354 800 40384
rect 1853 40354 1919 40357
rect -800 40352 1919 40354
rect -800 40296 1858 40352
rect 1914 40296 1919 40352
rect -800 40294 1919 40296
rect -800 40264 800 40294
rect 1853 40291 1919 40294
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 40223 35248 40224
rect 37457 39946 37523 39949
rect 39200 39946 40800 39976
rect 37457 39944 40800 39946
rect 37457 39888 37462 39944
rect 37518 39888 40800 39944
rect 37457 39886 40800 39888
rect 37457 39883 37523 39886
rect 39200 39856 40800 39886
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 39679 19888 39680
rect -800 39538 800 39568
rect 1853 39538 1919 39541
rect -800 39536 1919 39538
rect -800 39480 1858 39536
rect 1914 39480 1919 39536
rect -800 39478 1919 39480
rect -800 39448 800 39478
rect 1853 39475 1919 39478
rect 37917 39538 37983 39541
rect 39200 39538 40800 39568
rect 37917 39536 40800 39538
rect 37917 39480 37922 39536
rect 37978 39480 40800 39536
rect 37917 39478 40800 39480
rect 37917 39475 37983 39478
rect 39200 39448 40800 39478
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 37917 39130 37983 39133
rect 39200 39130 40800 39160
rect 37917 39128 40800 39130
rect 37917 39072 37922 39128
rect 37978 39072 40800 39128
rect 37917 39070 40800 39072
rect 37917 39067 37983 39070
rect 39200 39040 40800 39070
rect -800 38722 800 38752
rect 1853 38722 1919 38725
rect -800 38720 1919 38722
rect -800 38664 1858 38720
rect 1914 38664 1919 38720
rect -800 38662 1919 38664
rect -800 38632 800 38662
rect 1853 38659 1919 38662
rect 37457 38722 37523 38725
rect 39200 38722 40800 38752
rect 37457 38720 40800 38722
rect 37457 38664 37462 38720
rect 37518 38664 40800 38720
rect 37457 38662 40800 38664
rect 37457 38659 37523 38662
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 39200 38632 40800 38662
rect 19568 38591 19888 38592
rect 37181 38178 37247 38181
rect 39200 38178 40800 38208
rect 37181 38176 40800 38178
rect 37181 38120 37186 38176
rect 37242 38120 40800 38176
rect 37181 38118 40800 38120
rect 37181 38115 37247 38118
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 39200 38088 40800 38118
rect 34928 38047 35248 38048
rect -800 37906 800 37936
rect 1853 37906 1919 37909
rect -800 37904 1919 37906
rect -800 37848 1858 37904
rect 1914 37848 1919 37904
rect -800 37846 1919 37848
rect -800 37816 800 37846
rect 1853 37843 1919 37846
rect 37917 37770 37983 37773
rect 39200 37770 40800 37800
rect 37917 37768 40800 37770
rect 37917 37712 37922 37768
rect 37978 37712 40800 37768
rect 37917 37710 40800 37712
rect 37917 37707 37983 37710
rect 39200 37680 40800 37710
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 37365 37362 37431 37365
rect 39200 37362 40800 37392
rect 37365 37360 40800 37362
rect 37365 37304 37370 37360
rect 37426 37304 40800 37360
rect 37365 37302 40800 37304
rect 37365 37299 37431 37302
rect 39200 37272 40800 37302
rect -800 37090 800 37120
rect 1853 37090 1919 37093
rect -800 37088 1919 37090
rect -800 37032 1858 37088
rect 1914 37032 1919 37088
rect -800 37030 1919 37032
rect -800 37000 800 37030
rect 1853 37027 1919 37030
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 35709 36816 35775 36821
rect 35709 36760 35714 36816
rect 35770 36760 35775 36816
rect 35709 36755 35775 36760
rect 37273 36818 37339 36821
rect 39200 36818 40800 36848
rect 37273 36816 40800 36818
rect 37273 36760 37278 36816
rect 37334 36760 40800 36816
rect 37273 36758 40800 36760
rect 37273 36755 37339 36758
rect 35712 36549 35772 36755
rect 39200 36728 40800 36758
rect 35709 36544 35775 36549
rect 35709 36488 35714 36544
rect 35770 36488 35775 36544
rect 35709 36483 35775 36488
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 34697 36410 34763 36413
rect 35525 36410 35591 36413
rect 34697 36408 35591 36410
rect 34697 36352 34702 36408
rect 34758 36352 35530 36408
rect 35586 36352 35591 36408
rect 34697 36350 35591 36352
rect 34697 36347 34763 36350
rect 35525 36347 35591 36350
rect 37917 36410 37983 36413
rect 39200 36410 40800 36440
rect 37917 36408 40800 36410
rect 37917 36352 37922 36408
rect 37978 36352 40800 36408
rect 37917 36350 40800 36352
rect 37917 36347 37983 36350
rect 39200 36320 40800 36350
rect -800 36274 800 36304
rect 1853 36274 1919 36277
rect -800 36272 1919 36274
rect -800 36216 1858 36272
rect 1914 36216 1919 36272
rect -800 36214 1919 36216
rect -800 36184 800 36214
rect 1853 36211 1919 36214
rect 32397 36138 32463 36141
rect 33777 36138 33843 36141
rect 34881 36138 34947 36141
rect 32397 36136 34947 36138
rect 32397 36080 32402 36136
rect 32458 36080 33782 36136
rect 33838 36080 34886 36136
rect 34942 36080 34947 36136
rect 32397 36078 34947 36080
rect 32397 36075 32463 36078
rect 33777 36075 33843 36078
rect 34881 36075 34947 36078
rect 37365 36002 37431 36005
rect 39200 36002 40800 36032
rect 37365 36000 40800 36002
rect 37365 35944 37370 36000
rect 37426 35944 40800 36000
rect 37365 35942 40800 35944
rect 37365 35939 37431 35942
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 39200 35912 40800 35942
rect 34928 35871 35248 35872
rect -800 35458 800 35488
rect 1853 35458 1919 35461
rect -800 35456 1919 35458
rect -800 35400 1858 35456
rect 1914 35400 1919 35456
rect -800 35398 1919 35400
rect -800 35368 800 35398
rect 1853 35395 1919 35398
rect 37273 35458 37339 35461
rect 39200 35458 40800 35488
rect 37273 35456 40800 35458
rect 37273 35400 37278 35456
rect 37334 35400 40800 35456
rect 37273 35398 40800 35400
rect 37273 35395 37339 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 39200 35368 40800 35398
rect 19568 35327 19888 35328
rect 37917 35050 37983 35053
rect 39200 35050 40800 35080
rect 37917 35048 40800 35050
rect 37917 34992 37922 35048
rect 37978 34992 40800 35048
rect 37917 34990 40800 34992
rect 37917 34987 37983 34990
rect 39200 34960 40800 34990
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect -800 34642 800 34672
rect 1853 34642 1919 34645
rect -800 34640 1919 34642
rect -800 34584 1858 34640
rect 1914 34584 1919 34640
rect -800 34582 1919 34584
rect -800 34552 800 34582
rect 1853 34579 1919 34582
rect 37457 34642 37523 34645
rect 39200 34642 40800 34672
rect 37457 34640 40800 34642
rect 37457 34584 37462 34640
rect 37518 34584 40800 34640
rect 37457 34582 40800 34584
rect 37457 34579 37523 34582
rect 39200 34552 40800 34582
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 37917 34234 37983 34237
rect 39200 34234 40800 34264
rect 37917 34232 40800 34234
rect 37917 34176 37922 34232
rect 37978 34176 40800 34232
rect 37917 34174 40800 34176
rect 37917 34171 37983 34174
rect 39200 34144 40800 34174
rect -800 33826 800 33856
rect 1853 33826 1919 33829
rect -800 33824 1919 33826
rect -800 33768 1858 33824
rect 1914 33768 1919 33824
rect -800 33766 1919 33768
rect -800 33736 800 33766
rect 1853 33763 1919 33766
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 37917 33690 37983 33693
rect 39200 33690 40800 33720
rect 37917 33688 40800 33690
rect 37917 33632 37922 33688
rect 37978 33632 40800 33688
rect 37917 33630 40800 33632
rect 37917 33627 37983 33630
rect 39200 33600 40800 33630
rect 37457 33282 37523 33285
rect 39200 33282 40800 33312
rect 37457 33280 40800 33282
rect 37457 33224 37462 33280
rect 37518 33224 40800 33280
rect 37457 33222 40800 33224
rect 37457 33219 37523 33222
rect 19568 33216 19888 33217
rect -800 33146 800 33176
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 39200 33192 40800 33222
rect 19568 33151 19888 33152
rect 1853 33146 1919 33149
rect -800 33144 1919 33146
rect -800 33088 1858 33144
rect 1914 33088 1919 33144
rect -800 33086 1919 33088
rect -800 33056 800 33086
rect 1853 33083 1919 33086
rect 37181 32874 37247 32877
rect 39200 32874 40800 32904
rect 37181 32872 40800 32874
rect 37181 32816 37186 32872
rect 37242 32816 40800 32872
rect 37181 32814 40800 32816
rect 37181 32811 37247 32814
rect 39200 32784 40800 32814
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect -800 32330 800 32360
rect 1853 32330 1919 32333
rect -800 32328 1919 32330
rect -800 32272 1858 32328
rect 1914 32272 1919 32328
rect -800 32270 1919 32272
rect -800 32240 800 32270
rect 1853 32267 1919 32270
rect 37917 32330 37983 32333
rect 39200 32330 40800 32360
rect 37917 32328 40800 32330
rect 37917 32272 37922 32328
rect 37978 32272 40800 32328
rect 37917 32270 40800 32272
rect 37917 32267 37983 32270
rect 39200 32240 40800 32270
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 37365 31922 37431 31925
rect 39200 31922 40800 31952
rect 37365 31920 40800 31922
rect 37365 31864 37370 31920
rect 37426 31864 40800 31920
rect 37365 31862 40800 31864
rect 37365 31859 37431 31862
rect 39200 31832 40800 31862
rect 4208 31584 4528 31585
rect -800 31514 800 31544
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 1853 31514 1919 31517
rect -800 31512 1919 31514
rect -800 31456 1858 31512
rect 1914 31456 1919 31512
rect -800 31454 1919 31456
rect -800 31424 800 31454
rect 1853 31451 1919 31454
rect 37273 31514 37339 31517
rect 39200 31514 40800 31544
rect 37273 31512 40800 31514
rect 37273 31456 37278 31512
rect 37334 31456 40800 31512
rect 37273 31454 40800 31456
rect 37273 31451 37339 31454
rect 39200 31424 40800 31454
rect 37917 31106 37983 31109
rect 39200 31106 40800 31136
rect 37917 31104 40800 31106
rect 37917 31048 37922 31104
rect 37978 31048 40800 31104
rect 37917 31046 40800 31048
rect 37917 31043 37983 31046
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 39200 31016 40800 31046
rect 19568 30975 19888 30976
rect -800 30698 800 30728
rect 1853 30698 1919 30701
rect -800 30696 1919 30698
rect -800 30640 1858 30696
rect 1914 30640 1919 30696
rect -800 30638 1919 30640
rect -800 30608 800 30638
rect 1853 30635 1919 30638
rect 37365 30562 37431 30565
rect 39200 30562 40800 30592
rect 37365 30560 40800 30562
rect 37365 30504 37370 30560
rect 37426 30504 40800 30560
rect 37365 30502 40800 30504
rect 37365 30499 37431 30502
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 39200 30472 40800 30502
rect 34928 30431 35248 30432
rect 37273 30154 37339 30157
rect 39200 30154 40800 30184
rect 37273 30152 40800 30154
rect 37273 30096 37278 30152
rect 37334 30096 40800 30152
rect 37273 30094 40800 30096
rect 37273 30091 37339 30094
rect 39200 30064 40800 30094
rect 19568 29952 19888 29953
rect -800 29882 800 29912
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 1853 29882 1919 29885
rect -800 29880 1919 29882
rect -800 29824 1858 29880
rect 1914 29824 1919 29880
rect -800 29822 1919 29824
rect -800 29792 800 29822
rect 1853 29819 1919 29822
rect 37917 29746 37983 29749
rect 39200 29746 40800 29776
rect 37917 29744 40800 29746
rect 37917 29688 37922 29744
rect 37978 29688 40800 29744
rect 37917 29686 40800 29688
rect 37917 29683 37983 29686
rect 39200 29656 40800 29686
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 37457 29202 37523 29205
rect 39200 29202 40800 29232
rect 37457 29200 40800 29202
rect 37457 29144 37462 29200
rect 37518 29144 40800 29200
rect 37457 29142 40800 29144
rect 37457 29139 37523 29142
rect 39200 29112 40800 29142
rect -800 29066 800 29096
rect 1853 29066 1919 29069
rect -800 29064 1919 29066
rect -800 29008 1858 29064
rect 1914 29008 1919 29064
rect -800 29006 1919 29008
rect -800 28976 800 29006
rect 1853 29003 1919 29006
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 38009 28794 38075 28797
rect 39200 28794 40800 28824
rect 38009 28792 40800 28794
rect 38009 28736 38014 28792
rect 38070 28736 40800 28792
rect 38009 28734 40800 28736
rect 38009 28731 38075 28734
rect 39200 28704 40800 28734
rect 37917 28386 37983 28389
rect 39200 28386 40800 28416
rect 37917 28384 40800 28386
rect 37917 28328 37922 28384
rect 37978 28328 40800 28384
rect 37917 28326 40800 28328
rect 37917 28323 37983 28326
rect 4208 28320 4528 28321
rect -800 28250 800 28280
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 39200 28296 40800 28326
rect 34928 28255 35248 28256
rect 1853 28250 1919 28253
rect -800 28248 1919 28250
rect -800 28192 1858 28248
rect 1914 28192 1919 28248
rect -800 28190 1919 28192
rect -800 28160 800 28190
rect 1853 28187 1919 28190
rect 37457 27978 37523 27981
rect 39200 27978 40800 28008
rect 37457 27976 40800 27978
rect 37457 27920 37462 27976
rect 37518 27920 40800 27976
rect 37457 27918 40800 27920
rect 37457 27915 37523 27918
rect 39200 27888 40800 27918
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect -800 27434 800 27464
rect 1853 27434 1919 27437
rect -800 27432 1919 27434
rect -800 27376 1858 27432
rect 1914 27376 1919 27432
rect -800 27374 1919 27376
rect -800 27344 800 27374
rect 1853 27371 1919 27374
rect 37181 27434 37247 27437
rect 39200 27434 40800 27464
rect 37181 27432 40800 27434
rect 37181 27376 37186 27432
rect 37242 27376 40800 27432
rect 37181 27374 40800 27376
rect 37181 27371 37247 27374
rect 39200 27344 40800 27374
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 37917 27026 37983 27029
rect 39200 27026 40800 27056
rect 37917 27024 40800 27026
rect 37917 26968 37922 27024
rect 37978 26968 40800 27024
rect 37917 26966 40800 26968
rect 37917 26963 37983 26966
rect 39200 26936 40800 26966
rect -800 26754 800 26784
rect 1853 26754 1919 26757
rect -800 26752 1919 26754
rect -800 26696 1858 26752
rect 1914 26696 1919 26752
rect -800 26694 1919 26696
rect -800 26664 800 26694
rect 1853 26691 1919 26694
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 37365 26618 37431 26621
rect 39200 26618 40800 26648
rect 37365 26616 40800 26618
rect 37365 26560 37370 26616
rect 37426 26560 40800 26616
rect 37365 26558 40800 26560
rect 37365 26555 37431 26558
rect 39200 26528 40800 26558
rect 34605 26482 34671 26485
rect 34605 26480 34714 26482
rect 34605 26424 34610 26480
rect 34666 26424 34714 26480
rect 34605 26419 34714 26424
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect -800 25938 800 25968
rect 1853 25938 1919 25941
rect -800 25936 1919 25938
rect -800 25880 1858 25936
rect 1914 25880 1919 25936
rect -800 25878 1919 25880
rect 34654 25938 34714 26419
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 37273 26074 37339 26077
rect 39200 26074 40800 26104
rect 37273 26072 40800 26074
rect 37273 26016 37278 26072
rect 37334 26016 40800 26072
rect 37273 26014 40800 26016
rect 37273 26011 37339 26014
rect 39200 25984 40800 26014
rect 34881 25938 34947 25941
rect 34654 25936 34947 25938
rect 34654 25880 34886 25936
rect 34942 25880 34947 25936
rect 34654 25878 34947 25880
rect -800 25848 800 25878
rect 1853 25875 1919 25878
rect 34881 25875 34947 25878
rect 37917 25666 37983 25669
rect 39200 25666 40800 25696
rect 37917 25664 40800 25666
rect 37917 25608 37922 25664
rect 37978 25608 40800 25664
rect 37917 25606 40800 25608
rect 37917 25603 37983 25606
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 39200 25576 40800 25606
rect 19568 25535 19888 25536
rect 34237 25530 34303 25533
rect 38101 25530 38167 25533
rect 34237 25528 38167 25530
rect 34237 25472 34242 25528
rect 34298 25472 38106 25528
rect 38162 25472 38167 25528
rect 34237 25470 38167 25472
rect 34237 25467 34303 25470
rect 38101 25467 38167 25470
rect 34973 25394 35039 25397
rect 37733 25394 37799 25397
rect 34973 25392 37799 25394
rect 34973 25336 34978 25392
rect 35034 25336 37738 25392
rect 37794 25336 37799 25392
rect 34973 25334 37799 25336
rect 34973 25331 35039 25334
rect 37733 25331 37799 25334
rect 34513 25258 34579 25261
rect 34697 25258 34763 25261
rect 34513 25256 34763 25258
rect 34513 25200 34518 25256
rect 34574 25200 34702 25256
rect 34758 25200 34763 25256
rect 34513 25198 34763 25200
rect 34513 25195 34579 25198
rect 34697 25195 34763 25198
rect 34881 25258 34947 25261
rect 37181 25258 37247 25261
rect 39200 25258 40800 25288
rect 34881 25256 35450 25258
rect 34881 25200 34886 25256
rect 34942 25200 35450 25256
rect 34881 25198 35450 25200
rect 34881 25195 34947 25198
rect -800 25122 800 25152
rect 1853 25122 1919 25125
rect -800 25120 1919 25122
rect -800 25064 1858 25120
rect 1914 25064 1919 25120
rect -800 25062 1919 25064
rect -800 25032 800 25062
rect 1853 25059 1919 25062
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 35157 24884 35223 24887
rect 35390 24884 35450 25198
rect 37181 25256 40800 25258
rect 37181 25200 37186 25256
rect 37242 25200 40800 25256
rect 37181 25198 40800 25200
rect 37181 25195 37247 25198
rect 39200 25168 40800 25198
rect 35157 24882 35450 24884
rect 35157 24826 35162 24882
rect 35218 24826 35450 24882
rect 35157 24824 35450 24826
rect 37273 24850 37339 24853
rect 39200 24850 40800 24880
rect 37273 24848 40800 24850
rect 35157 24821 35223 24824
rect 37273 24792 37278 24848
rect 37334 24792 40800 24848
rect 37273 24790 40800 24792
rect 37273 24787 37339 24790
rect 39200 24760 40800 24790
rect 32949 24578 33015 24581
rect 34329 24578 34395 24581
rect 32949 24576 34395 24578
rect 32949 24520 32954 24576
rect 33010 24520 34334 24576
rect 34390 24520 34395 24576
rect 32949 24518 34395 24520
rect 32949 24515 33015 24518
rect 34329 24515 34395 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect -800 24306 800 24336
rect 1853 24306 1919 24309
rect -800 24304 1919 24306
rect -800 24248 1858 24304
rect 1914 24248 1919 24304
rect -800 24246 1919 24248
rect -800 24216 800 24246
rect 1853 24243 1919 24246
rect 37917 24306 37983 24309
rect 39200 24306 40800 24336
rect 37917 24304 40800 24306
rect 37917 24248 37922 24304
rect 37978 24248 40800 24304
rect 37917 24246 40800 24248
rect 37917 24243 37983 24246
rect 39200 24216 40800 24246
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 37365 23898 37431 23901
rect 39200 23898 40800 23928
rect 37365 23896 40800 23898
rect 37365 23840 37370 23896
rect 37426 23840 40800 23896
rect 37365 23838 40800 23840
rect 37365 23835 37431 23838
rect 39200 23808 40800 23838
rect -800 23490 800 23520
rect 1853 23490 1919 23493
rect -800 23488 1919 23490
rect -800 23432 1858 23488
rect 1914 23432 1919 23488
rect -800 23430 1919 23432
rect -800 23400 800 23430
rect 1853 23427 1919 23430
rect 34605 23490 34671 23493
rect 35617 23490 35683 23493
rect 34605 23488 35683 23490
rect 34605 23432 34610 23488
rect 34666 23432 35622 23488
rect 35678 23432 35683 23488
rect 34605 23430 35683 23432
rect 34605 23427 34671 23430
rect 35617 23427 35683 23430
rect 37273 23490 37339 23493
rect 39200 23490 40800 23520
rect 37273 23488 40800 23490
rect 37273 23432 37278 23488
rect 37334 23432 40800 23488
rect 37273 23430 40800 23432
rect 37273 23427 37339 23430
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 39200 23400 40800 23430
rect 19568 23359 19888 23360
rect 31477 23082 31543 23085
rect 33685 23082 33751 23085
rect 31477 23080 33751 23082
rect 31477 23024 31482 23080
rect 31538 23024 33690 23080
rect 33746 23024 33751 23080
rect 31477 23022 33751 23024
rect 31477 23019 31543 23022
rect 33685 23019 33751 23022
rect 33869 23082 33935 23085
rect 33869 23080 33978 23082
rect 33869 23024 33874 23080
rect 33930 23024 33978 23080
rect 33869 23019 33978 23024
rect 34605 23080 34671 23085
rect 34605 23024 34610 23080
rect 34666 23024 34671 23080
rect 34605 23019 34671 23024
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect -800 22674 800 22704
rect 1853 22674 1919 22677
rect -800 22672 1919 22674
rect -800 22616 1858 22672
rect 1914 22616 1919 22672
rect -800 22614 1919 22616
rect -800 22584 800 22614
rect 1853 22611 1919 22614
rect 32857 22536 32923 22541
rect 32857 22480 32862 22536
rect 32918 22480 32923 22536
rect 32857 22475 32923 22480
rect 32860 22402 32920 22475
rect 33317 22402 33383 22405
rect 32860 22400 33383 22402
rect 32860 22344 33322 22400
rect 33378 22344 33383 22400
rect 32860 22342 33383 22344
rect 33317 22339 33383 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 32305 22264 32371 22269
rect 32305 22208 32310 22264
rect 32366 22208 32371 22264
rect 32305 22203 32371 22208
rect 32308 21994 32368 22203
rect 33041 22130 33107 22133
rect 33918 22130 33978 23019
rect 34421 22946 34487 22949
rect 34608 22946 34668 23019
rect 34421 22944 34668 22946
rect 34421 22888 34426 22944
rect 34482 22888 34668 22944
rect 34421 22886 34668 22888
rect 37917 22946 37983 22949
rect 39200 22946 40800 22976
rect 37917 22944 40800 22946
rect 37917 22888 37922 22944
rect 37978 22888 40800 22944
rect 37917 22886 40800 22888
rect 34421 22883 34487 22886
rect 37917 22883 37983 22886
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 39200 22856 40800 22886
rect 34928 22815 35248 22816
rect 35065 22536 35131 22541
rect 35065 22480 35070 22536
rect 35126 22480 35131 22536
rect 35065 22475 35131 22480
rect 37273 22538 37339 22541
rect 39200 22538 40800 22568
rect 37273 22536 40800 22538
rect 37273 22480 37278 22536
rect 37334 22480 40800 22536
rect 37273 22478 40800 22480
rect 37273 22475 37339 22478
rect 34145 22266 34211 22269
rect 35068 22266 35128 22475
rect 39200 22448 40800 22478
rect 34145 22264 35128 22266
rect 34145 22208 34150 22264
rect 34206 22208 35128 22264
rect 34145 22206 35128 22208
rect 34145 22203 34211 22206
rect 34329 22130 34395 22133
rect 33041 22128 33426 22130
rect 33041 22072 33046 22128
rect 33102 22072 33426 22128
rect 33041 22070 33426 22072
rect 33918 22128 34395 22130
rect 33918 22072 34334 22128
rect 34390 22072 34395 22128
rect 33918 22070 34395 22072
rect 33041 22067 33107 22070
rect 33225 21994 33291 21997
rect 32308 21992 33291 21994
rect 32308 21936 33230 21992
rect 33286 21936 33291 21992
rect 32308 21934 33291 21936
rect 33225 21931 33291 21934
rect -800 21858 800 21888
rect 1853 21858 1919 21861
rect -800 21856 1919 21858
rect -800 21800 1858 21856
rect 1914 21800 1919 21856
rect -800 21798 1919 21800
rect -800 21768 800 21798
rect 1853 21795 1919 21798
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 32029 21722 32095 21725
rect 32029 21720 32828 21722
rect 32029 21664 32034 21720
rect 32090 21664 32828 21720
rect 32029 21662 32828 21664
rect 32029 21659 32095 21662
rect 32213 21586 32279 21589
rect 32489 21586 32555 21589
rect 32213 21584 32322 21586
rect 32213 21528 32218 21584
rect 32274 21528 32322 21584
rect 32213 21523 32322 21528
rect 32489 21584 32690 21586
rect 32489 21528 32494 21584
rect 32550 21528 32690 21584
rect 32489 21526 32690 21528
rect 32489 21523 32555 21526
rect 32262 21450 32322 21523
rect 32262 21390 32506 21450
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect -800 21042 800 21072
rect 1853 21042 1919 21045
rect -800 21040 1919 21042
rect -800 20984 1858 21040
rect 1914 20984 1919 21040
rect -800 20982 1919 20984
rect -800 20952 800 20982
rect 1853 20979 1919 20982
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 32446 20634 32506 21390
rect 32630 20770 32690 21526
rect 32768 20909 32828 21662
rect 33366 21181 33426 22070
rect 34329 22067 34395 22070
rect 35065 22130 35131 22133
rect 37457 22130 37523 22133
rect 35065 22128 37523 22130
rect 35065 22072 35070 22128
rect 35126 22072 37462 22128
rect 37518 22072 37523 22128
rect 35065 22070 37523 22072
rect 35065 22067 35131 22070
rect 37457 22067 37523 22070
rect 37917 22130 37983 22133
rect 39200 22130 40800 22160
rect 37917 22128 40800 22130
rect 37917 22072 37922 22128
rect 37978 22072 40800 22128
rect 37917 22070 40800 22072
rect 37917 22067 37983 22070
rect 39200 22040 40800 22070
rect 33685 21994 33751 21997
rect 34421 21994 34487 21997
rect 34881 21994 34947 21997
rect 33685 21992 34487 21994
rect 33685 21936 33690 21992
rect 33746 21936 34426 21992
rect 34482 21936 34487 21992
rect 33685 21934 34487 21936
rect 33685 21931 33751 21934
rect 34421 21931 34487 21934
rect 34608 21992 34947 21994
rect 34608 21936 34886 21992
rect 34942 21936 34947 21992
rect 34608 21934 34947 21936
rect 34053 21858 34119 21861
rect 34608 21858 34668 21934
rect 34881 21931 34947 21934
rect 35617 21994 35683 21997
rect 35893 21994 35959 21997
rect 35617 21992 35959 21994
rect 35617 21936 35622 21992
rect 35678 21936 35898 21992
rect 35954 21936 35959 21992
rect 35617 21934 35959 21936
rect 35617 21931 35683 21934
rect 35893 21931 35959 21934
rect 34053 21856 34668 21858
rect 34053 21800 34058 21856
rect 34114 21800 34668 21856
rect 34053 21798 34668 21800
rect 34053 21795 34119 21798
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 37917 21586 37983 21589
rect 39200 21586 40800 21616
rect 37917 21584 40800 21586
rect 37917 21528 37922 21584
rect 37978 21528 40800 21584
rect 37917 21526 40800 21528
rect 37917 21523 37983 21526
rect 39200 21496 40800 21526
rect 34329 21450 34395 21453
rect 34286 21448 34395 21450
rect 34286 21392 34334 21448
rect 34390 21392 34395 21448
rect 34286 21387 34395 21392
rect 33317 21176 33426 21181
rect 33317 21120 33322 21176
rect 33378 21120 33426 21176
rect 33317 21118 33426 21120
rect 34145 21178 34211 21181
rect 34286 21178 34346 21387
rect 35341 21178 35407 21181
rect 34145 21176 34346 21178
rect 34145 21120 34150 21176
rect 34206 21120 34346 21176
rect 34145 21118 34346 21120
rect 34516 21176 35407 21178
rect 34516 21120 35346 21176
rect 35402 21120 35407 21176
rect 34516 21118 35407 21120
rect 33317 21115 33383 21118
rect 34145 21115 34211 21118
rect 32765 20904 32831 20909
rect 32765 20848 32770 20904
rect 32826 20848 32831 20904
rect 32765 20843 32831 20848
rect 33133 20770 33199 20773
rect 32630 20768 33199 20770
rect 32630 20712 33138 20768
rect 33194 20712 33199 20768
rect 32630 20710 33199 20712
rect 33133 20707 33199 20710
rect 32446 20574 32690 20634
rect -800 20362 800 20392
rect 1853 20362 1919 20365
rect -800 20360 1919 20362
rect -800 20304 1858 20360
rect 1914 20304 1919 20360
rect -800 20302 1919 20304
rect 32630 20362 32690 20574
rect 34516 20501 34576 21118
rect 35341 21115 35407 21118
rect 37273 21178 37339 21181
rect 39200 21178 40800 21208
rect 37273 21176 40800 21178
rect 37273 21120 37278 21176
rect 37334 21120 40800 21176
rect 37273 21118 40800 21120
rect 37273 21115 37339 21118
rect 39200 21088 40800 21118
rect 35157 20906 35223 20909
rect 35433 20906 35499 20909
rect 35157 20904 35499 20906
rect 35157 20848 35162 20904
rect 35218 20848 35438 20904
rect 35494 20848 35499 20904
rect 35157 20846 35499 20848
rect 35157 20843 35223 20846
rect 35433 20843 35499 20846
rect 37181 20770 37247 20773
rect 39200 20770 40800 20800
rect 37181 20768 40800 20770
rect 37181 20712 37186 20768
rect 37242 20712 40800 20768
rect 37181 20710 40800 20712
rect 37181 20707 37247 20710
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 39200 20680 40800 20710
rect 34928 20639 35248 20640
rect 34513 20496 34579 20501
rect 34513 20440 34518 20496
rect 34574 20440 34579 20496
rect 34513 20435 34579 20440
rect 32857 20362 32923 20365
rect 32630 20360 32923 20362
rect 32630 20304 32862 20360
rect 32918 20304 32923 20360
rect 32630 20302 32923 20304
rect -800 20272 800 20302
rect 1853 20299 1919 20302
rect 32857 20299 32923 20302
rect 33317 20362 33383 20365
rect 34881 20362 34947 20365
rect 33317 20360 34947 20362
rect 33317 20304 33322 20360
rect 33378 20304 34886 20360
rect 34942 20304 34947 20360
rect 33317 20302 34947 20304
rect 33317 20299 33383 20302
rect 34881 20299 34947 20302
rect 37917 20362 37983 20365
rect 39200 20362 40800 20392
rect 37917 20360 40800 20362
rect 37917 20304 37922 20360
rect 37978 20304 40800 20360
rect 37917 20302 40800 20304
rect 37917 20299 37983 20302
rect 39200 20272 40800 20302
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 30925 20090 30991 20093
rect 35893 20090 35959 20093
rect 30925 20088 35959 20090
rect 30925 20032 30930 20088
rect 30986 20032 35898 20088
rect 35954 20032 35959 20088
rect 30925 20030 35959 20032
rect 30925 20027 30991 20030
rect 35893 20027 35959 20030
rect 33317 19954 33383 19957
rect 33317 19952 33610 19954
rect 33317 19896 33322 19952
rect 33378 19896 33610 19952
rect 33317 19894 33610 19896
rect 33317 19891 33383 19894
rect 30557 19818 30623 19821
rect 30741 19818 30807 19821
rect 30557 19816 30807 19818
rect 30557 19760 30562 19816
rect 30618 19760 30746 19816
rect 30802 19760 30807 19816
rect 30557 19758 30807 19760
rect 33550 19818 33610 19894
rect 34513 19952 34579 19957
rect 34513 19896 34518 19952
rect 34574 19896 34579 19952
rect 34513 19891 34579 19896
rect 33869 19818 33935 19821
rect 33550 19816 33935 19818
rect 33550 19760 33874 19816
rect 33930 19760 33935 19816
rect 33550 19758 33935 19760
rect 30557 19755 30623 19758
rect 30741 19755 30807 19758
rect 33869 19755 33935 19758
rect 4208 19616 4528 19617
rect -800 19546 800 19576
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 1853 19546 1919 19549
rect -800 19544 1919 19546
rect -800 19488 1858 19544
rect 1914 19488 1919 19544
rect -800 19486 1919 19488
rect -800 19456 800 19486
rect 1853 19483 1919 19486
rect 32765 19544 32831 19549
rect 32765 19488 32770 19544
rect 32826 19488 32831 19544
rect 32765 19483 32831 19488
rect 34053 19546 34119 19549
rect 34516 19546 34576 19891
rect 34881 19818 34947 19821
rect 34053 19544 34576 19546
rect 34053 19488 34058 19544
rect 34114 19488 34576 19544
rect 34053 19486 34576 19488
rect 34700 19816 34947 19818
rect 34700 19760 34886 19816
rect 34942 19760 34947 19816
rect 34700 19758 34947 19760
rect 34053 19483 34119 19486
rect 32305 19410 32371 19413
rect 32768 19410 32828 19483
rect 32305 19408 32828 19410
rect 32305 19352 32310 19408
rect 32366 19352 32828 19408
rect 32305 19350 32828 19352
rect 34700 19410 34760 19758
rect 34881 19755 34947 19758
rect 37181 19818 37247 19821
rect 39200 19818 40800 19848
rect 37181 19816 40800 19818
rect 37181 19760 37186 19816
rect 37242 19760 40800 19816
rect 37181 19758 40800 19760
rect 37181 19755 37247 19758
rect 39200 19728 40800 19758
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 34881 19410 34947 19413
rect 34700 19408 34947 19410
rect 34700 19352 34886 19408
rect 34942 19352 34947 19408
rect 34700 19350 34947 19352
rect 32305 19347 32371 19350
rect 34881 19347 34947 19350
rect 37273 19410 37339 19413
rect 39200 19410 40800 19440
rect 37273 19408 40800 19410
rect 37273 19352 37278 19408
rect 37334 19352 40800 19408
rect 37273 19350 40800 19352
rect 37273 19347 37339 19350
rect 39200 19320 40800 19350
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 37917 19002 37983 19005
rect 39200 19002 40800 19032
rect 37917 19000 40800 19002
rect 37917 18944 37922 19000
rect 37978 18944 40800 19000
rect 37917 18942 40800 18944
rect 37917 18939 37983 18942
rect 39200 18912 40800 18942
rect -800 18730 800 18760
rect 1853 18730 1919 18733
rect -800 18728 1919 18730
rect -800 18672 1858 18728
rect 1914 18672 1919 18728
rect -800 18670 1919 18672
rect -800 18640 800 18670
rect 1853 18667 1919 18670
rect 25129 18730 25195 18733
rect 26601 18730 26667 18733
rect 28257 18730 28323 18733
rect 35065 18730 35131 18733
rect 25129 18728 28323 18730
rect 25129 18672 25134 18728
rect 25190 18672 26606 18728
rect 26662 18672 28262 18728
rect 28318 18672 28323 18728
rect 25129 18670 28323 18672
rect 25129 18667 25195 18670
rect 26601 18667 26667 18670
rect 28257 18667 28323 18670
rect 34700 18728 35131 18730
rect 34700 18672 35070 18728
rect 35126 18672 35131 18728
rect 34700 18670 35131 18672
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 29545 18456 29611 18461
rect 29545 18400 29550 18456
rect 29606 18400 29611 18456
rect 29545 18395 29611 18400
rect 29548 18186 29608 18395
rect 34700 18322 34760 18670
rect 35065 18667 35131 18670
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 37181 18458 37247 18461
rect 39200 18458 40800 18488
rect 37181 18456 40800 18458
rect 37181 18400 37186 18456
rect 37242 18400 40800 18456
rect 37181 18398 40800 18400
rect 37181 18395 37247 18398
rect 39200 18368 40800 18398
rect 34881 18322 34947 18325
rect 34700 18320 34947 18322
rect 34700 18264 34886 18320
rect 34942 18264 34947 18320
rect 34700 18262 34947 18264
rect 34881 18259 34947 18262
rect 29134 18126 29608 18186
rect 19568 17984 19888 17985
rect -800 17914 800 17944
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 1853 17914 1919 17917
rect -800 17912 1919 17914
rect -800 17856 1858 17912
rect 1914 17856 1919 17912
rect -800 17854 1919 17856
rect -800 17824 800 17854
rect 1853 17851 1919 17854
rect 28993 17642 29059 17645
rect 29134 17642 29194 18126
rect 37273 18050 37339 18053
rect 39200 18050 40800 18080
rect 37273 18048 40800 18050
rect 37273 17992 37278 18048
rect 37334 17992 40800 18048
rect 37273 17990 40800 17992
rect 37273 17987 37339 17990
rect 39200 17960 40800 17990
rect 30189 17642 30255 17645
rect 28993 17640 30255 17642
rect 28993 17584 28998 17640
rect 29054 17584 30194 17640
rect 30250 17584 30255 17640
rect 28993 17582 30255 17584
rect 28993 17579 29059 17582
rect 30189 17579 30255 17582
rect 37917 17642 37983 17645
rect 39200 17642 40800 17672
rect 37917 17640 40800 17642
rect 37917 17584 37922 17640
rect 37978 17584 40800 17640
rect 37917 17582 40800 17584
rect 37917 17579 37983 17582
rect 39200 17552 40800 17582
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 37273 17234 37339 17237
rect 39200 17234 40800 17264
rect 37273 17232 40800 17234
rect 37273 17176 37278 17232
rect 37334 17176 40800 17232
rect 37273 17174 40800 17176
rect 37273 17171 37339 17174
rect 39200 17144 40800 17174
rect -800 17098 800 17128
rect 1853 17098 1919 17101
rect -800 17096 1919 17098
rect -800 17040 1858 17096
rect 1914 17040 1919 17096
rect -800 17038 1919 17040
rect -800 17008 800 17038
rect 1853 17035 1919 17038
rect 33961 17098 34027 17101
rect 33961 17096 34162 17098
rect 33961 17040 33966 17096
rect 34022 17040 34162 17096
rect 33961 17038 34162 17040
rect 33961 17035 34027 17038
rect 33317 16962 33383 16965
rect 33961 16962 34027 16965
rect 33317 16960 34027 16962
rect 33317 16904 33322 16960
rect 33378 16904 33966 16960
rect 34022 16904 34027 16960
rect 33317 16902 34027 16904
rect 34102 16962 34162 17038
rect 34329 16962 34395 16965
rect 34102 16960 34395 16962
rect 34102 16904 34334 16960
rect 34390 16904 34395 16960
rect 34102 16902 34395 16904
rect 33317 16899 33383 16902
rect 33961 16899 34027 16902
rect 34329 16899 34395 16902
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 37917 16690 37983 16693
rect 39200 16690 40800 16720
rect 37917 16688 40800 16690
rect 37917 16632 37922 16688
rect 37978 16632 40800 16688
rect 37917 16630 40800 16632
rect 37917 16627 37983 16630
rect 39200 16600 40800 16630
rect 30281 16554 30347 16557
rect 31753 16554 31819 16557
rect 30281 16552 31819 16554
rect 30281 16496 30286 16552
rect 30342 16496 31758 16552
rect 31814 16496 31819 16552
rect 30281 16494 31819 16496
rect 30281 16491 30347 16494
rect 31753 16491 31819 16494
rect 34145 16554 34211 16557
rect 36169 16554 36235 16557
rect 34145 16552 36235 16554
rect 34145 16496 34150 16552
rect 34206 16496 36174 16552
rect 36230 16496 36235 16552
rect 34145 16494 36235 16496
rect 34145 16491 34211 16494
rect 36169 16491 36235 16494
rect 4208 16352 4528 16353
rect -800 16282 800 16312
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 1853 16282 1919 16285
rect -800 16280 1919 16282
rect -800 16224 1858 16280
rect 1914 16224 1919 16280
rect -800 16222 1919 16224
rect -800 16192 800 16222
rect 1853 16219 1919 16222
rect 37917 16282 37983 16285
rect 39200 16282 40800 16312
rect 37917 16280 40800 16282
rect 37917 16224 37922 16280
rect 37978 16224 40800 16280
rect 37917 16222 40800 16224
rect 37917 16219 37983 16222
rect 39200 16192 40800 16222
rect 32305 16010 32371 16013
rect 34329 16010 34395 16013
rect 32305 16008 34395 16010
rect 32305 15952 32310 16008
rect 32366 15952 34334 16008
rect 34390 15952 34395 16008
rect 32305 15950 34395 15952
rect 32305 15947 32371 15950
rect 34329 15947 34395 15950
rect 37273 15874 37339 15877
rect 39200 15874 40800 15904
rect 37273 15872 40800 15874
rect 37273 15816 37278 15872
rect 37334 15816 40800 15872
rect 37273 15814 40800 15816
rect 37273 15811 37339 15814
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 39200 15784 40800 15814
rect 19568 15743 19888 15744
rect 33961 15602 34027 15605
rect 35433 15602 35499 15605
rect 33961 15600 34162 15602
rect 33961 15544 33966 15600
rect 34022 15544 34162 15600
rect 33961 15542 34162 15544
rect 33961 15539 34027 15542
rect -800 15466 800 15496
rect 1853 15466 1919 15469
rect -800 15464 1919 15466
rect -800 15408 1858 15464
rect 1914 15408 1919 15464
rect -800 15406 1919 15408
rect -800 15376 800 15406
rect 1853 15403 1919 15406
rect 27889 15466 27955 15469
rect 31385 15466 31451 15469
rect 27889 15464 31451 15466
rect 27889 15408 27894 15464
rect 27950 15408 31390 15464
rect 31446 15408 31451 15464
rect 27889 15406 31451 15408
rect 27889 15403 27955 15406
rect 31385 15403 31451 15406
rect 31661 15330 31727 15333
rect 33961 15330 34027 15333
rect 31661 15328 34027 15330
rect 31661 15272 31666 15328
rect 31722 15272 33966 15328
rect 34022 15272 34027 15328
rect 31661 15270 34027 15272
rect 31661 15267 31727 15270
rect 33961 15267 34027 15270
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34102 15194 34162 15542
rect 35433 15600 35680 15602
rect 35433 15544 35438 15600
rect 35494 15544 35680 15600
rect 35433 15542 35680 15544
rect 35433 15539 35499 15542
rect 35620 15469 35680 15542
rect 35617 15464 35683 15469
rect 35617 15408 35622 15464
rect 35678 15408 35683 15464
rect 35617 15403 35683 15408
rect 37181 15330 37247 15333
rect 39200 15330 40800 15360
rect 37181 15328 40800 15330
rect 37181 15272 37186 15328
rect 37242 15272 40800 15328
rect 37181 15270 40800 15272
rect 37181 15267 37247 15270
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 39200 15240 40800 15270
rect 34928 15199 35248 15200
rect 34329 15194 34395 15197
rect 34102 15192 34395 15194
rect 34102 15136 34334 15192
rect 34390 15136 34395 15192
rect 34102 15134 34395 15136
rect 34329 15131 34395 15134
rect 28901 14922 28967 14925
rect 30373 14922 30439 14925
rect 28901 14920 30439 14922
rect 28901 14864 28906 14920
rect 28962 14864 30378 14920
rect 30434 14864 30439 14920
rect 28901 14862 30439 14864
rect 28901 14859 28967 14862
rect 30373 14859 30439 14862
rect 37917 14922 37983 14925
rect 39200 14922 40800 14952
rect 37917 14920 40800 14922
rect 37917 14864 37922 14920
rect 37978 14864 40800 14920
rect 37917 14862 40800 14864
rect 37917 14859 37983 14862
rect 39200 14832 40800 14862
rect 23565 14786 23631 14789
rect 25129 14786 25195 14789
rect 27429 14786 27495 14789
rect 23565 14784 27495 14786
rect 23565 14728 23570 14784
rect 23626 14728 25134 14784
rect 25190 14728 27434 14784
rect 27490 14728 27495 14784
rect 23565 14726 27495 14728
rect 23565 14723 23631 14726
rect 25129 14723 25195 14726
rect 27429 14723 27495 14726
rect 28901 14786 28967 14789
rect 29729 14786 29795 14789
rect 28901 14784 29795 14786
rect 28901 14728 28906 14784
rect 28962 14728 29734 14784
rect 29790 14728 29795 14784
rect 28901 14726 29795 14728
rect 28901 14723 28967 14726
rect 29729 14723 29795 14726
rect 19568 14720 19888 14721
rect -800 14650 800 14680
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 1853 14650 1919 14653
rect -800 14648 1919 14650
rect -800 14592 1858 14648
rect 1914 14592 1919 14648
rect -800 14590 1919 14592
rect -800 14560 800 14590
rect 1853 14587 1919 14590
rect 23473 14514 23539 14517
rect 26049 14514 26115 14517
rect 27797 14514 27863 14517
rect 23473 14512 27863 14514
rect 23473 14456 23478 14512
rect 23534 14456 26054 14512
rect 26110 14456 27802 14512
rect 27858 14456 27863 14512
rect 23473 14454 27863 14456
rect 23473 14451 23539 14454
rect 26049 14451 26115 14454
rect 27797 14451 27863 14454
rect 33317 14514 33383 14517
rect 34329 14514 34395 14517
rect 33317 14512 34395 14514
rect 33317 14456 33322 14512
rect 33378 14456 34334 14512
rect 34390 14456 34395 14512
rect 33317 14454 34395 14456
rect 33317 14451 33383 14454
rect 34329 14451 34395 14454
rect 37181 14514 37247 14517
rect 39200 14514 40800 14544
rect 37181 14512 40800 14514
rect 37181 14456 37186 14512
rect 37242 14456 40800 14512
rect 37181 14454 40800 14456
rect 37181 14451 37247 14454
rect 39200 14424 40800 14454
rect 23657 14378 23723 14381
rect 29177 14378 29243 14381
rect 23657 14376 29243 14378
rect 23657 14320 23662 14376
rect 23718 14320 29182 14376
rect 29238 14320 29243 14376
rect 23657 14318 29243 14320
rect 23657 14315 23723 14318
rect 29177 14315 29243 14318
rect 32949 14378 33015 14381
rect 35525 14378 35591 14381
rect 32949 14376 35591 14378
rect 32949 14320 32954 14376
rect 33010 14320 35530 14376
rect 35586 14320 35591 14376
rect 32949 14318 35591 14320
rect 32949 14315 33015 14318
rect 35525 14315 35591 14318
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 37273 14106 37339 14109
rect 39200 14106 40800 14136
rect 37273 14104 40800 14106
rect 37273 14048 37278 14104
rect 37334 14048 40800 14104
rect 37273 14046 40800 14048
rect 37273 14043 37339 14046
rect 39200 14016 40800 14046
rect -800 13834 800 13864
rect 1853 13834 1919 13837
rect -800 13832 1919 13834
rect -800 13776 1858 13832
rect 1914 13776 1919 13832
rect -800 13774 1919 13776
rect -800 13744 800 13774
rect 1853 13771 1919 13774
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 24209 13562 24275 13565
rect 27613 13562 27679 13565
rect 24209 13560 27679 13562
rect 24209 13504 24214 13560
rect 24270 13504 27618 13560
rect 27674 13504 27679 13560
rect 24209 13502 27679 13504
rect 24209 13499 24275 13502
rect 27613 13499 27679 13502
rect 37181 13562 37247 13565
rect 39200 13562 40800 13592
rect 37181 13560 40800 13562
rect 37181 13504 37186 13560
rect 37242 13504 40800 13560
rect 37181 13502 40800 13504
rect 37181 13499 37247 13502
rect 39200 13472 40800 13502
rect -800 13154 800 13184
rect 1853 13154 1919 13157
rect -800 13152 1919 13154
rect -800 13096 1858 13152
rect 1914 13096 1919 13152
rect -800 13094 1919 13096
rect -800 13064 800 13094
rect 1853 13091 1919 13094
rect 37917 13154 37983 13157
rect 39200 13154 40800 13184
rect 37917 13152 40800 13154
rect 37917 13096 37922 13152
rect 37978 13096 40800 13152
rect 37917 13094 40800 13096
rect 37917 13091 37983 13094
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 39200 13064 40800 13094
rect 34928 13023 35248 13024
rect 37273 12746 37339 12749
rect 39200 12746 40800 12776
rect 37273 12744 40800 12746
rect 37273 12688 37278 12744
rect 37334 12688 40800 12744
rect 37273 12686 40800 12688
rect 37273 12683 37339 12686
rect 39200 12656 40800 12686
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect -800 12338 800 12368
rect 1853 12338 1919 12341
rect -800 12336 1919 12338
rect -800 12280 1858 12336
rect 1914 12280 1919 12336
rect -800 12278 1919 12280
rect -800 12248 800 12278
rect 1853 12275 1919 12278
rect 37917 12202 37983 12205
rect 39200 12202 40800 12232
rect 37917 12200 40800 12202
rect 37917 12144 37922 12200
rect 37978 12144 40800 12200
rect 37917 12142 40800 12144
rect 37917 12139 37983 12142
rect 39200 12112 40800 12142
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 37273 11794 37339 11797
rect 39200 11794 40800 11824
rect 37273 11792 40800 11794
rect 37273 11736 37278 11792
rect 37334 11736 40800 11792
rect 37273 11734 40800 11736
rect 37273 11731 37339 11734
rect 39200 11704 40800 11734
rect -800 11522 800 11552
rect 1853 11522 1919 11525
rect -800 11520 1919 11522
rect -800 11464 1858 11520
rect 1914 11464 1919 11520
rect -800 11462 1919 11464
rect -800 11432 800 11462
rect 1853 11459 1919 11462
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 37181 11386 37247 11389
rect 39200 11386 40800 11416
rect 37181 11384 40800 11386
rect 37181 11328 37186 11384
rect 37242 11328 40800 11384
rect 37181 11326 40800 11328
rect 37181 11323 37247 11326
rect 39200 11296 40800 11326
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 38929 10842 38995 10845
rect 39200 10842 40800 10872
rect 38929 10840 40800 10842
rect 38929 10784 38934 10840
rect 38990 10784 40800 10840
rect 38929 10782 40800 10784
rect 38929 10779 38995 10782
rect 39200 10752 40800 10782
rect -800 10706 800 10736
rect 1853 10706 1919 10709
rect -800 10704 1919 10706
rect -800 10648 1858 10704
rect 1914 10648 1919 10704
rect -800 10646 1919 10648
rect -800 10616 800 10646
rect 1853 10643 1919 10646
rect 37273 10434 37339 10437
rect 39200 10434 40800 10464
rect 37273 10432 40800 10434
rect 37273 10376 37278 10432
rect 37334 10376 40800 10432
rect 37273 10374 40800 10376
rect 37273 10371 37339 10374
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 39200 10344 40800 10374
rect 19568 10303 19888 10304
rect 37917 10026 37983 10029
rect 39200 10026 40800 10056
rect 37917 10024 40800 10026
rect 37917 9968 37922 10024
rect 37978 9968 40800 10024
rect 37917 9966 40800 9968
rect 37917 9963 37983 9966
rect 39200 9936 40800 9966
rect -800 9890 800 9920
rect 1853 9890 1919 9893
rect -800 9888 1919 9890
rect -800 9832 1858 9888
rect 1914 9832 1919 9888
rect -800 9830 1919 9832
rect -800 9800 800 9830
rect 1853 9827 1919 9830
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 37273 9618 37339 9621
rect 39200 9618 40800 9648
rect 37273 9616 40800 9618
rect 37273 9560 37278 9616
rect 37334 9560 40800 9616
rect 37273 9558 40800 9560
rect 37273 9555 37339 9558
rect 39200 9528 40800 9558
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect -800 9074 800 9104
rect 1853 9074 1919 9077
rect -800 9072 1919 9074
rect -800 9016 1858 9072
rect 1914 9016 1919 9072
rect -800 9014 1919 9016
rect -800 8984 800 9014
rect 1853 9011 1919 9014
rect 37181 9074 37247 9077
rect 39200 9074 40800 9104
rect 37181 9072 40800 9074
rect 37181 9016 37186 9072
rect 37242 9016 40800 9072
rect 37181 9014 40800 9016
rect 37181 9011 37247 9014
rect 39200 8984 40800 9014
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 37917 8666 37983 8669
rect 39200 8666 40800 8696
rect 37917 8664 40800 8666
rect 37917 8608 37922 8664
rect 37978 8608 40800 8664
rect 37917 8606 40800 8608
rect 37917 8603 37983 8606
rect 39200 8576 40800 8606
rect -800 8258 800 8288
rect 1853 8258 1919 8261
rect -800 8256 1919 8258
rect -800 8200 1858 8256
rect 1914 8200 1919 8256
rect -800 8198 1919 8200
rect -800 8168 800 8198
rect 1853 8195 1919 8198
rect 37181 8258 37247 8261
rect 39200 8258 40800 8288
rect 37181 8256 40800 8258
rect 37181 8200 37186 8256
rect 37242 8200 40800 8256
rect 37181 8198 40800 8200
rect 37181 8195 37247 8198
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 39200 8168 40800 8198
rect 19568 8127 19888 8128
rect 37917 7714 37983 7717
rect 39200 7714 40800 7744
rect 37917 7712 40800 7714
rect 37917 7656 37922 7712
rect 37978 7656 40800 7712
rect 37917 7654 40800 7656
rect 37917 7651 37983 7654
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 39200 7624 40800 7654
rect 34928 7583 35248 7584
rect -800 7442 800 7472
rect 1853 7442 1919 7445
rect -800 7440 1919 7442
rect -800 7384 1858 7440
rect 1914 7384 1919 7440
rect -800 7382 1919 7384
rect -800 7352 800 7382
rect 1853 7379 1919 7382
rect 37273 7306 37339 7309
rect 39200 7306 40800 7336
rect 37273 7304 40800 7306
rect 37273 7248 37278 7304
rect 37334 7248 40800 7304
rect 37273 7246 40800 7248
rect 37273 7243 37339 7246
rect 39200 7216 40800 7246
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 37181 6898 37247 6901
rect 39200 6898 40800 6928
rect 37181 6896 40800 6898
rect 37181 6840 37186 6896
rect 37242 6840 40800 6896
rect 37181 6838 40800 6840
rect 37181 6835 37247 6838
rect 39200 6808 40800 6838
rect -800 6762 800 6792
rect 1853 6762 1919 6765
rect -800 6760 1919 6762
rect -800 6704 1858 6760
rect 1914 6704 1919 6760
rect -800 6702 1919 6704
rect -800 6672 800 6702
rect 1853 6699 1919 6702
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 37917 6490 37983 6493
rect 39200 6490 40800 6520
rect 37917 6488 40800 6490
rect 37917 6432 37922 6488
rect 37978 6432 40800 6488
rect 37917 6430 40800 6432
rect 37917 6427 37983 6430
rect 39200 6400 40800 6430
rect 19568 6016 19888 6017
rect -800 5946 800 5976
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 1853 5946 1919 5949
rect -800 5944 1919 5946
rect -800 5888 1858 5944
rect 1914 5888 1919 5944
rect -800 5886 1919 5888
rect -800 5856 800 5886
rect 1853 5883 1919 5886
rect 37273 5946 37339 5949
rect 39200 5946 40800 5976
rect 37273 5944 40800 5946
rect 37273 5888 37278 5944
rect 37334 5888 40800 5944
rect 37273 5886 40800 5888
rect 37273 5883 37339 5886
rect 39200 5856 40800 5886
rect 37181 5538 37247 5541
rect 39200 5538 40800 5568
rect 37181 5536 40800 5538
rect 37181 5480 37186 5536
rect 37242 5480 40800 5536
rect 37181 5478 40800 5480
rect 37181 5475 37247 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 39200 5448 40800 5478
rect 34928 5407 35248 5408
rect -800 5130 800 5160
rect 1853 5130 1919 5133
rect -800 5128 1919 5130
rect -800 5072 1858 5128
rect 1914 5072 1919 5128
rect -800 5070 1919 5072
rect -800 5040 800 5070
rect 1853 5067 1919 5070
rect 38929 5130 38995 5133
rect 39200 5130 40800 5160
rect 38929 5128 40800 5130
rect 38929 5072 38934 5128
rect 38990 5072 40800 5128
rect 38929 5070 40800 5072
rect 38929 5067 38995 5070
rect 39200 5040 40800 5070
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 36445 4586 36511 4589
rect 39200 4586 40800 4616
rect 36445 4584 40800 4586
rect 36445 4528 36450 4584
rect 36506 4528 40800 4584
rect 36445 4526 40800 4528
rect 36445 4523 36511 4526
rect 39200 4496 40800 4526
rect 4208 4384 4528 4385
rect -800 4314 800 4344
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 1853 4314 1919 4317
rect -800 4312 1919 4314
rect -800 4256 1858 4312
rect 1914 4256 1919 4312
rect -800 4254 1919 4256
rect -800 4224 800 4254
rect 1853 4251 1919 4254
rect 34605 4178 34671 4181
rect 39200 4178 40800 4208
rect 34605 4176 40800 4178
rect 34605 4120 34610 4176
rect 34666 4120 40800 4176
rect 34605 4118 40800 4120
rect 34605 4115 34671 4118
rect 39200 4088 40800 4118
rect 31845 4042 31911 4045
rect 31710 4040 31911 4042
rect 31710 3984 31850 4040
rect 31906 3984 31911 4040
rect 31710 3982 31911 3984
rect 31710 3909 31770 3982
rect 31845 3979 31911 3982
rect 29361 3906 29427 3909
rect 31017 3906 31083 3909
rect 29361 3904 31083 3906
rect 29361 3848 29366 3904
rect 29422 3848 31022 3904
rect 31078 3848 31083 3904
rect 29361 3846 31083 3848
rect 29361 3843 29427 3846
rect 31017 3843 31083 3846
rect 31661 3904 31770 3909
rect 31661 3848 31666 3904
rect 31722 3848 31770 3904
rect 31661 3846 31770 3848
rect 31661 3843 31727 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 26325 3770 26391 3773
rect 31385 3770 31451 3773
rect 26325 3768 31451 3770
rect 26325 3712 26330 3768
rect 26386 3712 31390 3768
rect 31446 3712 31451 3768
rect 26325 3710 31451 3712
rect 26325 3707 26391 3710
rect 31385 3707 31451 3710
rect 35525 3770 35591 3773
rect 39200 3770 40800 3800
rect 35525 3768 40800 3770
rect 35525 3712 35530 3768
rect 35586 3712 40800 3768
rect 35525 3710 40800 3712
rect 35525 3707 35591 3710
rect 39200 3680 40800 3710
rect 30005 3634 30071 3637
rect 31109 3634 31175 3637
rect 30005 3632 31175 3634
rect 30005 3576 30010 3632
rect 30066 3576 31114 3632
rect 31170 3576 31175 3632
rect 30005 3574 31175 3576
rect 30005 3571 30071 3574
rect 31109 3571 31175 3574
rect -800 3498 800 3528
rect 1853 3498 1919 3501
rect -800 3496 1919 3498
rect -800 3440 1858 3496
rect 1914 3440 1919 3496
rect -800 3438 1919 3440
rect -800 3408 800 3438
rect 1853 3435 1919 3438
rect 25037 3498 25103 3501
rect 31569 3498 31635 3501
rect 25037 3496 31635 3498
rect 25037 3440 25042 3496
rect 25098 3440 31574 3496
rect 31630 3440 31635 3496
rect 25037 3438 31635 3440
rect 25037 3435 25103 3438
rect 31569 3435 31635 3438
rect 35893 3362 35959 3365
rect 39200 3362 40800 3392
rect 35893 3360 40800 3362
rect 35893 3304 35898 3360
rect 35954 3304 40800 3360
rect 35893 3302 40800 3304
rect 35893 3299 35959 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 39200 3272 40800 3302
rect 34928 3231 35248 3232
rect 26601 3226 26667 3229
rect 28625 3226 28691 3229
rect 26601 3224 28691 3226
rect 26601 3168 26606 3224
rect 26662 3168 28630 3224
rect 28686 3168 28691 3224
rect 26601 3166 28691 3168
rect 26601 3163 26667 3166
rect 28625 3163 28691 3166
rect 28993 3090 29059 3093
rect 30465 3090 30531 3093
rect 28993 3088 30531 3090
rect 28993 3032 28998 3088
rect 29054 3032 30470 3088
rect 30526 3032 30531 3088
rect 28993 3030 30531 3032
rect 28993 3027 29059 3030
rect 30465 3027 30531 3030
rect 30649 3090 30715 3093
rect 37917 3090 37983 3093
rect 30649 3088 37983 3090
rect 30649 3032 30654 3088
rect 30710 3032 37922 3088
rect 37978 3032 37983 3088
rect 30649 3030 37983 3032
rect 30649 3027 30715 3030
rect 37917 3027 37983 3030
rect 26325 2954 26391 2957
rect 29177 2954 29243 2957
rect 26325 2952 29243 2954
rect 26325 2896 26330 2952
rect 26386 2896 29182 2952
rect 29238 2896 29243 2952
rect 26325 2894 29243 2896
rect 26325 2891 26391 2894
rect 29177 2891 29243 2894
rect 36905 2818 36971 2821
rect 39200 2818 40800 2848
rect 36905 2816 40800 2818
rect 36905 2760 36910 2816
rect 36966 2760 40800 2816
rect 36905 2758 40800 2760
rect 36905 2755 36971 2758
rect 19568 2752 19888 2753
rect -800 2682 800 2712
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 39200 2728 40800 2758
rect 19568 2687 19888 2688
rect 1393 2682 1459 2685
rect -800 2680 1459 2682
rect -800 2624 1398 2680
rect 1454 2624 1459 2680
rect -800 2622 1459 2624
rect -800 2592 800 2622
rect 1393 2619 1459 2622
rect 34605 2410 34671 2413
rect 39200 2410 40800 2440
rect 34605 2408 40800 2410
rect 34605 2352 34610 2408
rect 34666 2352 40800 2408
rect 34605 2350 40800 2352
rect 34605 2347 34671 2350
rect 39200 2320 40800 2350
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 35617 2002 35683 2005
rect 39200 2002 40800 2032
rect 35617 2000 40800 2002
rect 35617 1944 35622 2000
rect 35678 1944 40800 2000
rect 35617 1942 40800 1944
rect 35617 1939 35683 1942
rect 39200 1912 40800 1942
rect -800 1866 800 1896
rect 2773 1866 2839 1869
rect -800 1864 2839 1866
rect -800 1808 2778 1864
rect 2834 1808 2839 1864
rect -800 1806 2839 1808
rect -800 1776 800 1806
rect 2773 1803 2839 1806
rect 36077 1458 36143 1461
rect 39200 1458 40800 1488
rect 36077 1456 40800 1458
rect 36077 1400 36082 1456
rect 36138 1400 40800 1456
rect 36077 1398 40800 1400
rect 36077 1395 36143 1398
rect 39200 1368 40800 1398
rect -800 1050 800 1080
rect 1853 1050 1919 1053
rect -800 1048 1919 1050
rect -800 992 1858 1048
rect 1914 992 1919 1048
rect -800 990 1919 992
rect -800 960 800 990
rect 1853 987 1919 990
rect 35801 1050 35867 1053
rect 39200 1050 40800 1080
rect 35801 1048 40800 1050
rect 35801 992 35806 1048
rect 35862 992 40800 1048
rect 35801 990 40800 992
rect 35801 987 35867 990
rect 39200 960 40800 990
rect 36721 642 36787 645
rect 39200 642 40800 672
rect 36721 640 40800 642
rect 36721 584 36726 640
rect 36782 584 40800 640
rect 36721 582 40800 584
rect 36721 579 36787 582
rect 39200 552 40800 582
rect -800 370 800 400
rect 2865 370 2931 373
rect -800 368 2931 370
rect -800 312 2870 368
rect 2926 312 2931 368
rect -800 310 2931 312
rect -800 280 800 310
rect 2865 307 2931 310
rect 37089 234 37155 237
rect 39200 234 40800 264
rect 37089 232 40800 234
rect 37089 176 37094 232
rect 37150 176 40800 232
rect 37089 174 40800 176
rect 37089 171 37155 174
rect 39200 144 40800 174
<< via3 >>
rect 4216 117532 4280 117536
rect 4216 117476 4220 117532
rect 4220 117476 4276 117532
rect 4276 117476 4280 117532
rect 4216 117472 4280 117476
rect 4296 117532 4360 117536
rect 4296 117476 4300 117532
rect 4300 117476 4356 117532
rect 4356 117476 4360 117532
rect 4296 117472 4360 117476
rect 4376 117532 4440 117536
rect 4376 117476 4380 117532
rect 4380 117476 4436 117532
rect 4436 117476 4440 117532
rect 4376 117472 4440 117476
rect 4456 117532 4520 117536
rect 4456 117476 4460 117532
rect 4460 117476 4516 117532
rect 4516 117476 4520 117532
rect 4456 117472 4520 117476
rect 34936 117532 35000 117536
rect 34936 117476 34940 117532
rect 34940 117476 34996 117532
rect 34996 117476 35000 117532
rect 34936 117472 35000 117476
rect 35016 117532 35080 117536
rect 35016 117476 35020 117532
rect 35020 117476 35076 117532
rect 35076 117476 35080 117532
rect 35016 117472 35080 117476
rect 35096 117532 35160 117536
rect 35096 117476 35100 117532
rect 35100 117476 35156 117532
rect 35156 117476 35160 117532
rect 35096 117472 35160 117476
rect 35176 117532 35240 117536
rect 35176 117476 35180 117532
rect 35180 117476 35236 117532
rect 35236 117476 35240 117532
rect 35176 117472 35240 117476
rect 19576 116988 19640 116992
rect 19576 116932 19580 116988
rect 19580 116932 19636 116988
rect 19636 116932 19640 116988
rect 19576 116928 19640 116932
rect 19656 116988 19720 116992
rect 19656 116932 19660 116988
rect 19660 116932 19716 116988
rect 19716 116932 19720 116988
rect 19656 116928 19720 116932
rect 19736 116988 19800 116992
rect 19736 116932 19740 116988
rect 19740 116932 19796 116988
rect 19796 116932 19800 116988
rect 19736 116928 19800 116932
rect 19816 116988 19880 116992
rect 19816 116932 19820 116988
rect 19820 116932 19876 116988
rect 19876 116932 19880 116988
rect 19816 116928 19880 116932
rect 4216 116444 4280 116448
rect 4216 116388 4220 116444
rect 4220 116388 4276 116444
rect 4276 116388 4280 116444
rect 4216 116384 4280 116388
rect 4296 116444 4360 116448
rect 4296 116388 4300 116444
rect 4300 116388 4356 116444
rect 4356 116388 4360 116444
rect 4296 116384 4360 116388
rect 4376 116444 4440 116448
rect 4376 116388 4380 116444
rect 4380 116388 4436 116444
rect 4436 116388 4440 116444
rect 4376 116384 4440 116388
rect 4456 116444 4520 116448
rect 4456 116388 4460 116444
rect 4460 116388 4516 116444
rect 4516 116388 4520 116444
rect 4456 116384 4520 116388
rect 34936 116444 35000 116448
rect 34936 116388 34940 116444
rect 34940 116388 34996 116444
rect 34996 116388 35000 116444
rect 34936 116384 35000 116388
rect 35016 116444 35080 116448
rect 35016 116388 35020 116444
rect 35020 116388 35076 116444
rect 35076 116388 35080 116444
rect 35016 116384 35080 116388
rect 35096 116444 35160 116448
rect 35096 116388 35100 116444
rect 35100 116388 35156 116444
rect 35156 116388 35160 116444
rect 35096 116384 35160 116388
rect 35176 116444 35240 116448
rect 35176 116388 35180 116444
rect 35180 116388 35236 116444
rect 35236 116388 35240 116444
rect 35176 116384 35240 116388
rect 19576 115900 19640 115904
rect 19576 115844 19580 115900
rect 19580 115844 19636 115900
rect 19636 115844 19640 115900
rect 19576 115840 19640 115844
rect 19656 115900 19720 115904
rect 19656 115844 19660 115900
rect 19660 115844 19716 115900
rect 19716 115844 19720 115900
rect 19656 115840 19720 115844
rect 19736 115900 19800 115904
rect 19736 115844 19740 115900
rect 19740 115844 19796 115900
rect 19796 115844 19800 115900
rect 19736 115840 19800 115844
rect 19816 115900 19880 115904
rect 19816 115844 19820 115900
rect 19820 115844 19876 115900
rect 19876 115844 19880 115900
rect 19816 115840 19880 115844
rect 4216 115356 4280 115360
rect 4216 115300 4220 115356
rect 4220 115300 4276 115356
rect 4276 115300 4280 115356
rect 4216 115296 4280 115300
rect 4296 115356 4360 115360
rect 4296 115300 4300 115356
rect 4300 115300 4356 115356
rect 4356 115300 4360 115356
rect 4296 115296 4360 115300
rect 4376 115356 4440 115360
rect 4376 115300 4380 115356
rect 4380 115300 4436 115356
rect 4436 115300 4440 115356
rect 4376 115296 4440 115300
rect 4456 115356 4520 115360
rect 4456 115300 4460 115356
rect 4460 115300 4516 115356
rect 4516 115300 4520 115356
rect 4456 115296 4520 115300
rect 34936 115356 35000 115360
rect 34936 115300 34940 115356
rect 34940 115300 34996 115356
rect 34996 115300 35000 115356
rect 34936 115296 35000 115300
rect 35016 115356 35080 115360
rect 35016 115300 35020 115356
rect 35020 115300 35076 115356
rect 35076 115300 35080 115356
rect 35016 115296 35080 115300
rect 35096 115356 35160 115360
rect 35096 115300 35100 115356
rect 35100 115300 35156 115356
rect 35156 115300 35160 115356
rect 35096 115296 35160 115300
rect 35176 115356 35240 115360
rect 35176 115300 35180 115356
rect 35180 115300 35236 115356
rect 35236 115300 35240 115356
rect 35176 115296 35240 115300
rect 19576 114812 19640 114816
rect 19576 114756 19580 114812
rect 19580 114756 19636 114812
rect 19636 114756 19640 114812
rect 19576 114752 19640 114756
rect 19656 114812 19720 114816
rect 19656 114756 19660 114812
rect 19660 114756 19716 114812
rect 19716 114756 19720 114812
rect 19656 114752 19720 114756
rect 19736 114812 19800 114816
rect 19736 114756 19740 114812
rect 19740 114756 19796 114812
rect 19796 114756 19800 114812
rect 19736 114752 19800 114756
rect 19816 114812 19880 114816
rect 19816 114756 19820 114812
rect 19820 114756 19876 114812
rect 19876 114756 19880 114812
rect 19816 114752 19880 114756
rect 4216 114268 4280 114272
rect 4216 114212 4220 114268
rect 4220 114212 4276 114268
rect 4276 114212 4280 114268
rect 4216 114208 4280 114212
rect 4296 114268 4360 114272
rect 4296 114212 4300 114268
rect 4300 114212 4356 114268
rect 4356 114212 4360 114268
rect 4296 114208 4360 114212
rect 4376 114268 4440 114272
rect 4376 114212 4380 114268
rect 4380 114212 4436 114268
rect 4436 114212 4440 114268
rect 4376 114208 4440 114212
rect 4456 114268 4520 114272
rect 4456 114212 4460 114268
rect 4460 114212 4516 114268
rect 4516 114212 4520 114268
rect 4456 114208 4520 114212
rect 34936 114268 35000 114272
rect 34936 114212 34940 114268
rect 34940 114212 34996 114268
rect 34996 114212 35000 114268
rect 34936 114208 35000 114212
rect 35016 114268 35080 114272
rect 35016 114212 35020 114268
rect 35020 114212 35076 114268
rect 35076 114212 35080 114268
rect 35016 114208 35080 114212
rect 35096 114268 35160 114272
rect 35096 114212 35100 114268
rect 35100 114212 35156 114268
rect 35156 114212 35160 114268
rect 35096 114208 35160 114212
rect 35176 114268 35240 114272
rect 35176 114212 35180 114268
rect 35180 114212 35236 114268
rect 35236 114212 35240 114268
rect 35176 114208 35240 114212
rect 19576 113724 19640 113728
rect 19576 113668 19580 113724
rect 19580 113668 19636 113724
rect 19636 113668 19640 113724
rect 19576 113664 19640 113668
rect 19656 113724 19720 113728
rect 19656 113668 19660 113724
rect 19660 113668 19716 113724
rect 19716 113668 19720 113724
rect 19656 113664 19720 113668
rect 19736 113724 19800 113728
rect 19736 113668 19740 113724
rect 19740 113668 19796 113724
rect 19796 113668 19800 113724
rect 19736 113664 19800 113668
rect 19816 113724 19880 113728
rect 19816 113668 19820 113724
rect 19820 113668 19876 113724
rect 19876 113668 19880 113724
rect 19816 113664 19880 113668
rect 4216 113180 4280 113184
rect 4216 113124 4220 113180
rect 4220 113124 4276 113180
rect 4276 113124 4280 113180
rect 4216 113120 4280 113124
rect 4296 113180 4360 113184
rect 4296 113124 4300 113180
rect 4300 113124 4356 113180
rect 4356 113124 4360 113180
rect 4296 113120 4360 113124
rect 4376 113180 4440 113184
rect 4376 113124 4380 113180
rect 4380 113124 4436 113180
rect 4436 113124 4440 113180
rect 4376 113120 4440 113124
rect 4456 113180 4520 113184
rect 4456 113124 4460 113180
rect 4460 113124 4516 113180
rect 4516 113124 4520 113180
rect 4456 113120 4520 113124
rect 34936 113180 35000 113184
rect 34936 113124 34940 113180
rect 34940 113124 34996 113180
rect 34996 113124 35000 113180
rect 34936 113120 35000 113124
rect 35016 113180 35080 113184
rect 35016 113124 35020 113180
rect 35020 113124 35076 113180
rect 35076 113124 35080 113180
rect 35016 113120 35080 113124
rect 35096 113180 35160 113184
rect 35096 113124 35100 113180
rect 35100 113124 35156 113180
rect 35156 113124 35160 113180
rect 35096 113120 35160 113124
rect 35176 113180 35240 113184
rect 35176 113124 35180 113180
rect 35180 113124 35236 113180
rect 35236 113124 35240 113180
rect 35176 113120 35240 113124
rect 19576 112636 19640 112640
rect 19576 112580 19580 112636
rect 19580 112580 19636 112636
rect 19636 112580 19640 112636
rect 19576 112576 19640 112580
rect 19656 112636 19720 112640
rect 19656 112580 19660 112636
rect 19660 112580 19716 112636
rect 19716 112580 19720 112636
rect 19656 112576 19720 112580
rect 19736 112636 19800 112640
rect 19736 112580 19740 112636
rect 19740 112580 19796 112636
rect 19796 112580 19800 112636
rect 19736 112576 19800 112580
rect 19816 112636 19880 112640
rect 19816 112580 19820 112636
rect 19820 112580 19876 112636
rect 19876 112580 19880 112636
rect 19816 112576 19880 112580
rect 4216 112092 4280 112096
rect 4216 112036 4220 112092
rect 4220 112036 4276 112092
rect 4276 112036 4280 112092
rect 4216 112032 4280 112036
rect 4296 112092 4360 112096
rect 4296 112036 4300 112092
rect 4300 112036 4356 112092
rect 4356 112036 4360 112092
rect 4296 112032 4360 112036
rect 4376 112092 4440 112096
rect 4376 112036 4380 112092
rect 4380 112036 4436 112092
rect 4436 112036 4440 112092
rect 4376 112032 4440 112036
rect 4456 112092 4520 112096
rect 4456 112036 4460 112092
rect 4460 112036 4516 112092
rect 4516 112036 4520 112092
rect 4456 112032 4520 112036
rect 34936 112092 35000 112096
rect 34936 112036 34940 112092
rect 34940 112036 34996 112092
rect 34996 112036 35000 112092
rect 34936 112032 35000 112036
rect 35016 112092 35080 112096
rect 35016 112036 35020 112092
rect 35020 112036 35076 112092
rect 35076 112036 35080 112092
rect 35016 112032 35080 112036
rect 35096 112092 35160 112096
rect 35096 112036 35100 112092
rect 35100 112036 35156 112092
rect 35156 112036 35160 112092
rect 35096 112032 35160 112036
rect 35176 112092 35240 112096
rect 35176 112036 35180 112092
rect 35180 112036 35236 112092
rect 35236 112036 35240 112092
rect 35176 112032 35240 112036
rect 19576 111548 19640 111552
rect 19576 111492 19580 111548
rect 19580 111492 19636 111548
rect 19636 111492 19640 111548
rect 19576 111488 19640 111492
rect 19656 111548 19720 111552
rect 19656 111492 19660 111548
rect 19660 111492 19716 111548
rect 19716 111492 19720 111548
rect 19656 111488 19720 111492
rect 19736 111548 19800 111552
rect 19736 111492 19740 111548
rect 19740 111492 19796 111548
rect 19796 111492 19800 111548
rect 19736 111488 19800 111492
rect 19816 111548 19880 111552
rect 19816 111492 19820 111548
rect 19820 111492 19876 111548
rect 19876 111492 19880 111548
rect 19816 111488 19880 111492
rect 4216 111004 4280 111008
rect 4216 110948 4220 111004
rect 4220 110948 4276 111004
rect 4276 110948 4280 111004
rect 4216 110944 4280 110948
rect 4296 111004 4360 111008
rect 4296 110948 4300 111004
rect 4300 110948 4356 111004
rect 4356 110948 4360 111004
rect 4296 110944 4360 110948
rect 4376 111004 4440 111008
rect 4376 110948 4380 111004
rect 4380 110948 4436 111004
rect 4436 110948 4440 111004
rect 4376 110944 4440 110948
rect 4456 111004 4520 111008
rect 4456 110948 4460 111004
rect 4460 110948 4516 111004
rect 4516 110948 4520 111004
rect 4456 110944 4520 110948
rect 34936 111004 35000 111008
rect 34936 110948 34940 111004
rect 34940 110948 34996 111004
rect 34996 110948 35000 111004
rect 34936 110944 35000 110948
rect 35016 111004 35080 111008
rect 35016 110948 35020 111004
rect 35020 110948 35076 111004
rect 35076 110948 35080 111004
rect 35016 110944 35080 110948
rect 35096 111004 35160 111008
rect 35096 110948 35100 111004
rect 35100 110948 35156 111004
rect 35156 110948 35160 111004
rect 35096 110944 35160 110948
rect 35176 111004 35240 111008
rect 35176 110948 35180 111004
rect 35180 110948 35236 111004
rect 35236 110948 35240 111004
rect 35176 110944 35240 110948
rect 19576 110460 19640 110464
rect 19576 110404 19580 110460
rect 19580 110404 19636 110460
rect 19636 110404 19640 110460
rect 19576 110400 19640 110404
rect 19656 110460 19720 110464
rect 19656 110404 19660 110460
rect 19660 110404 19716 110460
rect 19716 110404 19720 110460
rect 19656 110400 19720 110404
rect 19736 110460 19800 110464
rect 19736 110404 19740 110460
rect 19740 110404 19796 110460
rect 19796 110404 19800 110460
rect 19736 110400 19800 110404
rect 19816 110460 19880 110464
rect 19816 110404 19820 110460
rect 19820 110404 19876 110460
rect 19876 110404 19880 110460
rect 19816 110400 19880 110404
rect 4216 109916 4280 109920
rect 4216 109860 4220 109916
rect 4220 109860 4276 109916
rect 4276 109860 4280 109916
rect 4216 109856 4280 109860
rect 4296 109916 4360 109920
rect 4296 109860 4300 109916
rect 4300 109860 4356 109916
rect 4356 109860 4360 109916
rect 4296 109856 4360 109860
rect 4376 109916 4440 109920
rect 4376 109860 4380 109916
rect 4380 109860 4436 109916
rect 4436 109860 4440 109916
rect 4376 109856 4440 109860
rect 4456 109916 4520 109920
rect 4456 109860 4460 109916
rect 4460 109860 4516 109916
rect 4516 109860 4520 109916
rect 4456 109856 4520 109860
rect 34936 109916 35000 109920
rect 34936 109860 34940 109916
rect 34940 109860 34996 109916
rect 34996 109860 35000 109916
rect 34936 109856 35000 109860
rect 35016 109916 35080 109920
rect 35016 109860 35020 109916
rect 35020 109860 35076 109916
rect 35076 109860 35080 109916
rect 35016 109856 35080 109860
rect 35096 109916 35160 109920
rect 35096 109860 35100 109916
rect 35100 109860 35156 109916
rect 35156 109860 35160 109916
rect 35096 109856 35160 109860
rect 35176 109916 35240 109920
rect 35176 109860 35180 109916
rect 35180 109860 35236 109916
rect 35236 109860 35240 109916
rect 35176 109856 35240 109860
rect 19576 109372 19640 109376
rect 19576 109316 19580 109372
rect 19580 109316 19636 109372
rect 19636 109316 19640 109372
rect 19576 109312 19640 109316
rect 19656 109372 19720 109376
rect 19656 109316 19660 109372
rect 19660 109316 19716 109372
rect 19716 109316 19720 109372
rect 19656 109312 19720 109316
rect 19736 109372 19800 109376
rect 19736 109316 19740 109372
rect 19740 109316 19796 109372
rect 19796 109316 19800 109372
rect 19736 109312 19800 109316
rect 19816 109372 19880 109376
rect 19816 109316 19820 109372
rect 19820 109316 19876 109372
rect 19876 109316 19880 109372
rect 19816 109312 19880 109316
rect 4216 108828 4280 108832
rect 4216 108772 4220 108828
rect 4220 108772 4276 108828
rect 4276 108772 4280 108828
rect 4216 108768 4280 108772
rect 4296 108828 4360 108832
rect 4296 108772 4300 108828
rect 4300 108772 4356 108828
rect 4356 108772 4360 108828
rect 4296 108768 4360 108772
rect 4376 108828 4440 108832
rect 4376 108772 4380 108828
rect 4380 108772 4436 108828
rect 4436 108772 4440 108828
rect 4376 108768 4440 108772
rect 4456 108828 4520 108832
rect 4456 108772 4460 108828
rect 4460 108772 4516 108828
rect 4516 108772 4520 108828
rect 4456 108768 4520 108772
rect 34936 108828 35000 108832
rect 34936 108772 34940 108828
rect 34940 108772 34996 108828
rect 34996 108772 35000 108828
rect 34936 108768 35000 108772
rect 35016 108828 35080 108832
rect 35016 108772 35020 108828
rect 35020 108772 35076 108828
rect 35076 108772 35080 108828
rect 35016 108768 35080 108772
rect 35096 108828 35160 108832
rect 35096 108772 35100 108828
rect 35100 108772 35156 108828
rect 35156 108772 35160 108828
rect 35096 108768 35160 108772
rect 35176 108828 35240 108832
rect 35176 108772 35180 108828
rect 35180 108772 35236 108828
rect 35236 108772 35240 108828
rect 35176 108768 35240 108772
rect 19576 108284 19640 108288
rect 19576 108228 19580 108284
rect 19580 108228 19636 108284
rect 19636 108228 19640 108284
rect 19576 108224 19640 108228
rect 19656 108284 19720 108288
rect 19656 108228 19660 108284
rect 19660 108228 19716 108284
rect 19716 108228 19720 108284
rect 19656 108224 19720 108228
rect 19736 108284 19800 108288
rect 19736 108228 19740 108284
rect 19740 108228 19796 108284
rect 19796 108228 19800 108284
rect 19736 108224 19800 108228
rect 19816 108284 19880 108288
rect 19816 108228 19820 108284
rect 19820 108228 19876 108284
rect 19876 108228 19880 108284
rect 19816 108224 19880 108228
rect 4216 107740 4280 107744
rect 4216 107684 4220 107740
rect 4220 107684 4276 107740
rect 4276 107684 4280 107740
rect 4216 107680 4280 107684
rect 4296 107740 4360 107744
rect 4296 107684 4300 107740
rect 4300 107684 4356 107740
rect 4356 107684 4360 107740
rect 4296 107680 4360 107684
rect 4376 107740 4440 107744
rect 4376 107684 4380 107740
rect 4380 107684 4436 107740
rect 4436 107684 4440 107740
rect 4376 107680 4440 107684
rect 4456 107740 4520 107744
rect 4456 107684 4460 107740
rect 4460 107684 4516 107740
rect 4516 107684 4520 107740
rect 4456 107680 4520 107684
rect 34936 107740 35000 107744
rect 34936 107684 34940 107740
rect 34940 107684 34996 107740
rect 34996 107684 35000 107740
rect 34936 107680 35000 107684
rect 35016 107740 35080 107744
rect 35016 107684 35020 107740
rect 35020 107684 35076 107740
rect 35076 107684 35080 107740
rect 35016 107680 35080 107684
rect 35096 107740 35160 107744
rect 35096 107684 35100 107740
rect 35100 107684 35156 107740
rect 35156 107684 35160 107740
rect 35096 107680 35160 107684
rect 35176 107740 35240 107744
rect 35176 107684 35180 107740
rect 35180 107684 35236 107740
rect 35236 107684 35240 107740
rect 35176 107680 35240 107684
rect 19576 107196 19640 107200
rect 19576 107140 19580 107196
rect 19580 107140 19636 107196
rect 19636 107140 19640 107196
rect 19576 107136 19640 107140
rect 19656 107196 19720 107200
rect 19656 107140 19660 107196
rect 19660 107140 19716 107196
rect 19716 107140 19720 107196
rect 19656 107136 19720 107140
rect 19736 107196 19800 107200
rect 19736 107140 19740 107196
rect 19740 107140 19796 107196
rect 19796 107140 19800 107196
rect 19736 107136 19800 107140
rect 19816 107196 19880 107200
rect 19816 107140 19820 107196
rect 19820 107140 19876 107196
rect 19876 107140 19880 107196
rect 19816 107136 19880 107140
rect 4216 106652 4280 106656
rect 4216 106596 4220 106652
rect 4220 106596 4276 106652
rect 4276 106596 4280 106652
rect 4216 106592 4280 106596
rect 4296 106652 4360 106656
rect 4296 106596 4300 106652
rect 4300 106596 4356 106652
rect 4356 106596 4360 106652
rect 4296 106592 4360 106596
rect 4376 106652 4440 106656
rect 4376 106596 4380 106652
rect 4380 106596 4436 106652
rect 4436 106596 4440 106652
rect 4376 106592 4440 106596
rect 4456 106652 4520 106656
rect 4456 106596 4460 106652
rect 4460 106596 4516 106652
rect 4516 106596 4520 106652
rect 4456 106592 4520 106596
rect 34936 106652 35000 106656
rect 34936 106596 34940 106652
rect 34940 106596 34996 106652
rect 34996 106596 35000 106652
rect 34936 106592 35000 106596
rect 35016 106652 35080 106656
rect 35016 106596 35020 106652
rect 35020 106596 35076 106652
rect 35076 106596 35080 106652
rect 35016 106592 35080 106596
rect 35096 106652 35160 106656
rect 35096 106596 35100 106652
rect 35100 106596 35156 106652
rect 35156 106596 35160 106652
rect 35096 106592 35160 106596
rect 35176 106652 35240 106656
rect 35176 106596 35180 106652
rect 35180 106596 35236 106652
rect 35236 106596 35240 106652
rect 35176 106592 35240 106596
rect 19576 106108 19640 106112
rect 19576 106052 19580 106108
rect 19580 106052 19636 106108
rect 19636 106052 19640 106108
rect 19576 106048 19640 106052
rect 19656 106108 19720 106112
rect 19656 106052 19660 106108
rect 19660 106052 19716 106108
rect 19716 106052 19720 106108
rect 19656 106048 19720 106052
rect 19736 106108 19800 106112
rect 19736 106052 19740 106108
rect 19740 106052 19796 106108
rect 19796 106052 19800 106108
rect 19736 106048 19800 106052
rect 19816 106108 19880 106112
rect 19816 106052 19820 106108
rect 19820 106052 19876 106108
rect 19876 106052 19880 106108
rect 19816 106048 19880 106052
rect 4216 105564 4280 105568
rect 4216 105508 4220 105564
rect 4220 105508 4276 105564
rect 4276 105508 4280 105564
rect 4216 105504 4280 105508
rect 4296 105564 4360 105568
rect 4296 105508 4300 105564
rect 4300 105508 4356 105564
rect 4356 105508 4360 105564
rect 4296 105504 4360 105508
rect 4376 105564 4440 105568
rect 4376 105508 4380 105564
rect 4380 105508 4436 105564
rect 4436 105508 4440 105564
rect 4376 105504 4440 105508
rect 4456 105564 4520 105568
rect 4456 105508 4460 105564
rect 4460 105508 4516 105564
rect 4516 105508 4520 105564
rect 4456 105504 4520 105508
rect 34936 105564 35000 105568
rect 34936 105508 34940 105564
rect 34940 105508 34996 105564
rect 34996 105508 35000 105564
rect 34936 105504 35000 105508
rect 35016 105564 35080 105568
rect 35016 105508 35020 105564
rect 35020 105508 35076 105564
rect 35076 105508 35080 105564
rect 35016 105504 35080 105508
rect 35096 105564 35160 105568
rect 35096 105508 35100 105564
rect 35100 105508 35156 105564
rect 35156 105508 35160 105564
rect 35096 105504 35160 105508
rect 35176 105564 35240 105568
rect 35176 105508 35180 105564
rect 35180 105508 35236 105564
rect 35236 105508 35240 105564
rect 35176 105504 35240 105508
rect 19576 105020 19640 105024
rect 19576 104964 19580 105020
rect 19580 104964 19636 105020
rect 19636 104964 19640 105020
rect 19576 104960 19640 104964
rect 19656 105020 19720 105024
rect 19656 104964 19660 105020
rect 19660 104964 19716 105020
rect 19716 104964 19720 105020
rect 19656 104960 19720 104964
rect 19736 105020 19800 105024
rect 19736 104964 19740 105020
rect 19740 104964 19796 105020
rect 19796 104964 19800 105020
rect 19736 104960 19800 104964
rect 19816 105020 19880 105024
rect 19816 104964 19820 105020
rect 19820 104964 19876 105020
rect 19876 104964 19880 105020
rect 19816 104960 19880 104964
rect 4216 104476 4280 104480
rect 4216 104420 4220 104476
rect 4220 104420 4276 104476
rect 4276 104420 4280 104476
rect 4216 104416 4280 104420
rect 4296 104476 4360 104480
rect 4296 104420 4300 104476
rect 4300 104420 4356 104476
rect 4356 104420 4360 104476
rect 4296 104416 4360 104420
rect 4376 104476 4440 104480
rect 4376 104420 4380 104476
rect 4380 104420 4436 104476
rect 4436 104420 4440 104476
rect 4376 104416 4440 104420
rect 4456 104476 4520 104480
rect 4456 104420 4460 104476
rect 4460 104420 4516 104476
rect 4516 104420 4520 104476
rect 4456 104416 4520 104420
rect 34936 104476 35000 104480
rect 34936 104420 34940 104476
rect 34940 104420 34996 104476
rect 34996 104420 35000 104476
rect 34936 104416 35000 104420
rect 35016 104476 35080 104480
rect 35016 104420 35020 104476
rect 35020 104420 35076 104476
rect 35076 104420 35080 104476
rect 35016 104416 35080 104420
rect 35096 104476 35160 104480
rect 35096 104420 35100 104476
rect 35100 104420 35156 104476
rect 35156 104420 35160 104476
rect 35096 104416 35160 104420
rect 35176 104476 35240 104480
rect 35176 104420 35180 104476
rect 35180 104420 35236 104476
rect 35236 104420 35240 104476
rect 35176 104416 35240 104420
rect 19576 103932 19640 103936
rect 19576 103876 19580 103932
rect 19580 103876 19636 103932
rect 19636 103876 19640 103932
rect 19576 103872 19640 103876
rect 19656 103932 19720 103936
rect 19656 103876 19660 103932
rect 19660 103876 19716 103932
rect 19716 103876 19720 103932
rect 19656 103872 19720 103876
rect 19736 103932 19800 103936
rect 19736 103876 19740 103932
rect 19740 103876 19796 103932
rect 19796 103876 19800 103932
rect 19736 103872 19800 103876
rect 19816 103932 19880 103936
rect 19816 103876 19820 103932
rect 19820 103876 19876 103932
rect 19876 103876 19880 103932
rect 19816 103872 19880 103876
rect 4216 103388 4280 103392
rect 4216 103332 4220 103388
rect 4220 103332 4276 103388
rect 4276 103332 4280 103388
rect 4216 103328 4280 103332
rect 4296 103388 4360 103392
rect 4296 103332 4300 103388
rect 4300 103332 4356 103388
rect 4356 103332 4360 103388
rect 4296 103328 4360 103332
rect 4376 103388 4440 103392
rect 4376 103332 4380 103388
rect 4380 103332 4436 103388
rect 4436 103332 4440 103388
rect 4376 103328 4440 103332
rect 4456 103388 4520 103392
rect 4456 103332 4460 103388
rect 4460 103332 4516 103388
rect 4516 103332 4520 103388
rect 4456 103328 4520 103332
rect 34936 103388 35000 103392
rect 34936 103332 34940 103388
rect 34940 103332 34996 103388
rect 34996 103332 35000 103388
rect 34936 103328 35000 103332
rect 35016 103388 35080 103392
rect 35016 103332 35020 103388
rect 35020 103332 35076 103388
rect 35076 103332 35080 103388
rect 35016 103328 35080 103332
rect 35096 103388 35160 103392
rect 35096 103332 35100 103388
rect 35100 103332 35156 103388
rect 35156 103332 35160 103388
rect 35096 103328 35160 103332
rect 35176 103388 35240 103392
rect 35176 103332 35180 103388
rect 35180 103332 35236 103388
rect 35236 103332 35240 103388
rect 35176 103328 35240 103332
rect 19576 102844 19640 102848
rect 19576 102788 19580 102844
rect 19580 102788 19636 102844
rect 19636 102788 19640 102844
rect 19576 102784 19640 102788
rect 19656 102844 19720 102848
rect 19656 102788 19660 102844
rect 19660 102788 19716 102844
rect 19716 102788 19720 102844
rect 19656 102784 19720 102788
rect 19736 102844 19800 102848
rect 19736 102788 19740 102844
rect 19740 102788 19796 102844
rect 19796 102788 19800 102844
rect 19736 102784 19800 102788
rect 19816 102844 19880 102848
rect 19816 102788 19820 102844
rect 19820 102788 19876 102844
rect 19876 102788 19880 102844
rect 19816 102784 19880 102788
rect 4216 102300 4280 102304
rect 4216 102244 4220 102300
rect 4220 102244 4276 102300
rect 4276 102244 4280 102300
rect 4216 102240 4280 102244
rect 4296 102300 4360 102304
rect 4296 102244 4300 102300
rect 4300 102244 4356 102300
rect 4356 102244 4360 102300
rect 4296 102240 4360 102244
rect 4376 102300 4440 102304
rect 4376 102244 4380 102300
rect 4380 102244 4436 102300
rect 4436 102244 4440 102300
rect 4376 102240 4440 102244
rect 4456 102300 4520 102304
rect 4456 102244 4460 102300
rect 4460 102244 4516 102300
rect 4516 102244 4520 102300
rect 4456 102240 4520 102244
rect 34936 102300 35000 102304
rect 34936 102244 34940 102300
rect 34940 102244 34996 102300
rect 34996 102244 35000 102300
rect 34936 102240 35000 102244
rect 35016 102300 35080 102304
rect 35016 102244 35020 102300
rect 35020 102244 35076 102300
rect 35076 102244 35080 102300
rect 35016 102240 35080 102244
rect 35096 102300 35160 102304
rect 35096 102244 35100 102300
rect 35100 102244 35156 102300
rect 35156 102244 35160 102300
rect 35096 102240 35160 102244
rect 35176 102300 35240 102304
rect 35176 102244 35180 102300
rect 35180 102244 35236 102300
rect 35236 102244 35240 102300
rect 35176 102240 35240 102244
rect 19576 101756 19640 101760
rect 19576 101700 19580 101756
rect 19580 101700 19636 101756
rect 19636 101700 19640 101756
rect 19576 101696 19640 101700
rect 19656 101756 19720 101760
rect 19656 101700 19660 101756
rect 19660 101700 19716 101756
rect 19716 101700 19720 101756
rect 19656 101696 19720 101700
rect 19736 101756 19800 101760
rect 19736 101700 19740 101756
rect 19740 101700 19796 101756
rect 19796 101700 19800 101756
rect 19736 101696 19800 101700
rect 19816 101756 19880 101760
rect 19816 101700 19820 101756
rect 19820 101700 19876 101756
rect 19876 101700 19880 101756
rect 19816 101696 19880 101700
rect 4216 101212 4280 101216
rect 4216 101156 4220 101212
rect 4220 101156 4276 101212
rect 4276 101156 4280 101212
rect 4216 101152 4280 101156
rect 4296 101212 4360 101216
rect 4296 101156 4300 101212
rect 4300 101156 4356 101212
rect 4356 101156 4360 101212
rect 4296 101152 4360 101156
rect 4376 101212 4440 101216
rect 4376 101156 4380 101212
rect 4380 101156 4436 101212
rect 4436 101156 4440 101212
rect 4376 101152 4440 101156
rect 4456 101212 4520 101216
rect 4456 101156 4460 101212
rect 4460 101156 4516 101212
rect 4516 101156 4520 101212
rect 4456 101152 4520 101156
rect 34936 101212 35000 101216
rect 34936 101156 34940 101212
rect 34940 101156 34996 101212
rect 34996 101156 35000 101212
rect 34936 101152 35000 101156
rect 35016 101212 35080 101216
rect 35016 101156 35020 101212
rect 35020 101156 35076 101212
rect 35076 101156 35080 101212
rect 35016 101152 35080 101156
rect 35096 101212 35160 101216
rect 35096 101156 35100 101212
rect 35100 101156 35156 101212
rect 35156 101156 35160 101212
rect 35096 101152 35160 101156
rect 35176 101212 35240 101216
rect 35176 101156 35180 101212
rect 35180 101156 35236 101212
rect 35236 101156 35240 101212
rect 35176 101152 35240 101156
rect 19576 100668 19640 100672
rect 19576 100612 19580 100668
rect 19580 100612 19636 100668
rect 19636 100612 19640 100668
rect 19576 100608 19640 100612
rect 19656 100668 19720 100672
rect 19656 100612 19660 100668
rect 19660 100612 19716 100668
rect 19716 100612 19720 100668
rect 19656 100608 19720 100612
rect 19736 100668 19800 100672
rect 19736 100612 19740 100668
rect 19740 100612 19796 100668
rect 19796 100612 19800 100668
rect 19736 100608 19800 100612
rect 19816 100668 19880 100672
rect 19816 100612 19820 100668
rect 19820 100612 19876 100668
rect 19876 100612 19880 100668
rect 19816 100608 19880 100612
rect 4216 100124 4280 100128
rect 4216 100068 4220 100124
rect 4220 100068 4276 100124
rect 4276 100068 4280 100124
rect 4216 100064 4280 100068
rect 4296 100124 4360 100128
rect 4296 100068 4300 100124
rect 4300 100068 4356 100124
rect 4356 100068 4360 100124
rect 4296 100064 4360 100068
rect 4376 100124 4440 100128
rect 4376 100068 4380 100124
rect 4380 100068 4436 100124
rect 4436 100068 4440 100124
rect 4376 100064 4440 100068
rect 4456 100124 4520 100128
rect 4456 100068 4460 100124
rect 4460 100068 4516 100124
rect 4516 100068 4520 100124
rect 4456 100064 4520 100068
rect 34936 100124 35000 100128
rect 34936 100068 34940 100124
rect 34940 100068 34996 100124
rect 34996 100068 35000 100124
rect 34936 100064 35000 100068
rect 35016 100124 35080 100128
rect 35016 100068 35020 100124
rect 35020 100068 35076 100124
rect 35076 100068 35080 100124
rect 35016 100064 35080 100068
rect 35096 100124 35160 100128
rect 35096 100068 35100 100124
rect 35100 100068 35156 100124
rect 35156 100068 35160 100124
rect 35096 100064 35160 100068
rect 35176 100124 35240 100128
rect 35176 100068 35180 100124
rect 35180 100068 35236 100124
rect 35236 100068 35240 100124
rect 35176 100064 35240 100068
rect 19576 99580 19640 99584
rect 19576 99524 19580 99580
rect 19580 99524 19636 99580
rect 19636 99524 19640 99580
rect 19576 99520 19640 99524
rect 19656 99580 19720 99584
rect 19656 99524 19660 99580
rect 19660 99524 19716 99580
rect 19716 99524 19720 99580
rect 19656 99520 19720 99524
rect 19736 99580 19800 99584
rect 19736 99524 19740 99580
rect 19740 99524 19796 99580
rect 19796 99524 19800 99580
rect 19736 99520 19800 99524
rect 19816 99580 19880 99584
rect 19816 99524 19820 99580
rect 19820 99524 19876 99580
rect 19876 99524 19880 99580
rect 19816 99520 19880 99524
rect 4216 99036 4280 99040
rect 4216 98980 4220 99036
rect 4220 98980 4276 99036
rect 4276 98980 4280 99036
rect 4216 98976 4280 98980
rect 4296 99036 4360 99040
rect 4296 98980 4300 99036
rect 4300 98980 4356 99036
rect 4356 98980 4360 99036
rect 4296 98976 4360 98980
rect 4376 99036 4440 99040
rect 4376 98980 4380 99036
rect 4380 98980 4436 99036
rect 4436 98980 4440 99036
rect 4376 98976 4440 98980
rect 4456 99036 4520 99040
rect 4456 98980 4460 99036
rect 4460 98980 4516 99036
rect 4516 98980 4520 99036
rect 4456 98976 4520 98980
rect 34936 99036 35000 99040
rect 34936 98980 34940 99036
rect 34940 98980 34996 99036
rect 34996 98980 35000 99036
rect 34936 98976 35000 98980
rect 35016 99036 35080 99040
rect 35016 98980 35020 99036
rect 35020 98980 35076 99036
rect 35076 98980 35080 99036
rect 35016 98976 35080 98980
rect 35096 99036 35160 99040
rect 35096 98980 35100 99036
rect 35100 98980 35156 99036
rect 35156 98980 35160 99036
rect 35096 98976 35160 98980
rect 35176 99036 35240 99040
rect 35176 98980 35180 99036
rect 35180 98980 35236 99036
rect 35236 98980 35240 99036
rect 35176 98976 35240 98980
rect 19576 98492 19640 98496
rect 19576 98436 19580 98492
rect 19580 98436 19636 98492
rect 19636 98436 19640 98492
rect 19576 98432 19640 98436
rect 19656 98492 19720 98496
rect 19656 98436 19660 98492
rect 19660 98436 19716 98492
rect 19716 98436 19720 98492
rect 19656 98432 19720 98436
rect 19736 98492 19800 98496
rect 19736 98436 19740 98492
rect 19740 98436 19796 98492
rect 19796 98436 19800 98492
rect 19736 98432 19800 98436
rect 19816 98492 19880 98496
rect 19816 98436 19820 98492
rect 19820 98436 19876 98492
rect 19876 98436 19880 98492
rect 19816 98432 19880 98436
rect 4216 97948 4280 97952
rect 4216 97892 4220 97948
rect 4220 97892 4276 97948
rect 4276 97892 4280 97948
rect 4216 97888 4280 97892
rect 4296 97948 4360 97952
rect 4296 97892 4300 97948
rect 4300 97892 4356 97948
rect 4356 97892 4360 97948
rect 4296 97888 4360 97892
rect 4376 97948 4440 97952
rect 4376 97892 4380 97948
rect 4380 97892 4436 97948
rect 4436 97892 4440 97948
rect 4376 97888 4440 97892
rect 4456 97948 4520 97952
rect 4456 97892 4460 97948
rect 4460 97892 4516 97948
rect 4516 97892 4520 97948
rect 4456 97888 4520 97892
rect 34936 97948 35000 97952
rect 34936 97892 34940 97948
rect 34940 97892 34996 97948
rect 34996 97892 35000 97948
rect 34936 97888 35000 97892
rect 35016 97948 35080 97952
rect 35016 97892 35020 97948
rect 35020 97892 35076 97948
rect 35076 97892 35080 97948
rect 35016 97888 35080 97892
rect 35096 97948 35160 97952
rect 35096 97892 35100 97948
rect 35100 97892 35156 97948
rect 35156 97892 35160 97948
rect 35096 97888 35160 97892
rect 35176 97948 35240 97952
rect 35176 97892 35180 97948
rect 35180 97892 35236 97948
rect 35236 97892 35240 97948
rect 35176 97888 35240 97892
rect 19576 97404 19640 97408
rect 19576 97348 19580 97404
rect 19580 97348 19636 97404
rect 19636 97348 19640 97404
rect 19576 97344 19640 97348
rect 19656 97404 19720 97408
rect 19656 97348 19660 97404
rect 19660 97348 19716 97404
rect 19716 97348 19720 97404
rect 19656 97344 19720 97348
rect 19736 97404 19800 97408
rect 19736 97348 19740 97404
rect 19740 97348 19796 97404
rect 19796 97348 19800 97404
rect 19736 97344 19800 97348
rect 19816 97404 19880 97408
rect 19816 97348 19820 97404
rect 19820 97348 19876 97404
rect 19876 97348 19880 97404
rect 19816 97344 19880 97348
rect 4216 96860 4280 96864
rect 4216 96804 4220 96860
rect 4220 96804 4276 96860
rect 4276 96804 4280 96860
rect 4216 96800 4280 96804
rect 4296 96860 4360 96864
rect 4296 96804 4300 96860
rect 4300 96804 4356 96860
rect 4356 96804 4360 96860
rect 4296 96800 4360 96804
rect 4376 96860 4440 96864
rect 4376 96804 4380 96860
rect 4380 96804 4436 96860
rect 4436 96804 4440 96860
rect 4376 96800 4440 96804
rect 4456 96860 4520 96864
rect 4456 96804 4460 96860
rect 4460 96804 4516 96860
rect 4516 96804 4520 96860
rect 4456 96800 4520 96804
rect 34936 96860 35000 96864
rect 34936 96804 34940 96860
rect 34940 96804 34996 96860
rect 34996 96804 35000 96860
rect 34936 96800 35000 96804
rect 35016 96860 35080 96864
rect 35016 96804 35020 96860
rect 35020 96804 35076 96860
rect 35076 96804 35080 96860
rect 35016 96800 35080 96804
rect 35096 96860 35160 96864
rect 35096 96804 35100 96860
rect 35100 96804 35156 96860
rect 35156 96804 35160 96860
rect 35096 96800 35160 96804
rect 35176 96860 35240 96864
rect 35176 96804 35180 96860
rect 35180 96804 35236 96860
rect 35236 96804 35240 96860
rect 35176 96800 35240 96804
rect 19576 96316 19640 96320
rect 19576 96260 19580 96316
rect 19580 96260 19636 96316
rect 19636 96260 19640 96316
rect 19576 96256 19640 96260
rect 19656 96316 19720 96320
rect 19656 96260 19660 96316
rect 19660 96260 19716 96316
rect 19716 96260 19720 96316
rect 19656 96256 19720 96260
rect 19736 96316 19800 96320
rect 19736 96260 19740 96316
rect 19740 96260 19796 96316
rect 19796 96260 19800 96316
rect 19736 96256 19800 96260
rect 19816 96316 19880 96320
rect 19816 96260 19820 96316
rect 19820 96260 19876 96316
rect 19876 96260 19880 96316
rect 19816 96256 19880 96260
rect 4216 95772 4280 95776
rect 4216 95716 4220 95772
rect 4220 95716 4276 95772
rect 4276 95716 4280 95772
rect 4216 95712 4280 95716
rect 4296 95772 4360 95776
rect 4296 95716 4300 95772
rect 4300 95716 4356 95772
rect 4356 95716 4360 95772
rect 4296 95712 4360 95716
rect 4376 95772 4440 95776
rect 4376 95716 4380 95772
rect 4380 95716 4436 95772
rect 4436 95716 4440 95772
rect 4376 95712 4440 95716
rect 4456 95772 4520 95776
rect 4456 95716 4460 95772
rect 4460 95716 4516 95772
rect 4516 95716 4520 95772
rect 4456 95712 4520 95716
rect 34936 95772 35000 95776
rect 34936 95716 34940 95772
rect 34940 95716 34996 95772
rect 34996 95716 35000 95772
rect 34936 95712 35000 95716
rect 35016 95772 35080 95776
rect 35016 95716 35020 95772
rect 35020 95716 35076 95772
rect 35076 95716 35080 95772
rect 35016 95712 35080 95716
rect 35096 95772 35160 95776
rect 35096 95716 35100 95772
rect 35100 95716 35156 95772
rect 35156 95716 35160 95772
rect 35096 95712 35160 95716
rect 35176 95772 35240 95776
rect 35176 95716 35180 95772
rect 35180 95716 35236 95772
rect 35236 95716 35240 95772
rect 35176 95712 35240 95716
rect 19576 95228 19640 95232
rect 19576 95172 19580 95228
rect 19580 95172 19636 95228
rect 19636 95172 19640 95228
rect 19576 95168 19640 95172
rect 19656 95228 19720 95232
rect 19656 95172 19660 95228
rect 19660 95172 19716 95228
rect 19716 95172 19720 95228
rect 19656 95168 19720 95172
rect 19736 95228 19800 95232
rect 19736 95172 19740 95228
rect 19740 95172 19796 95228
rect 19796 95172 19800 95228
rect 19736 95168 19800 95172
rect 19816 95228 19880 95232
rect 19816 95172 19820 95228
rect 19820 95172 19876 95228
rect 19876 95172 19880 95228
rect 19816 95168 19880 95172
rect 4216 94684 4280 94688
rect 4216 94628 4220 94684
rect 4220 94628 4276 94684
rect 4276 94628 4280 94684
rect 4216 94624 4280 94628
rect 4296 94684 4360 94688
rect 4296 94628 4300 94684
rect 4300 94628 4356 94684
rect 4356 94628 4360 94684
rect 4296 94624 4360 94628
rect 4376 94684 4440 94688
rect 4376 94628 4380 94684
rect 4380 94628 4436 94684
rect 4436 94628 4440 94684
rect 4376 94624 4440 94628
rect 4456 94684 4520 94688
rect 4456 94628 4460 94684
rect 4460 94628 4516 94684
rect 4516 94628 4520 94684
rect 4456 94624 4520 94628
rect 34936 94684 35000 94688
rect 34936 94628 34940 94684
rect 34940 94628 34996 94684
rect 34996 94628 35000 94684
rect 34936 94624 35000 94628
rect 35016 94684 35080 94688
rect 35016 94628 35020 94684
rect 35020 94628 35076 94684
rect 35076 94628 35080 94684
rect 35016 94624 35080 94628
rect 35096 94684 35160 94688
rect 35096 94628 35100 94684
rect 35100 94628 35156 94684
rect 35156 94628 35160 94684
rect 35096 94624 35160 94628
rect 35176 94684 35240 94688
rect 35176 94628 35180 94684
rect 35180 94628 35236 94684
rect 35236 94628 35240 94684
rect 35176 94624 35240 94628
rect 19576 94140 19640 94144
rect 19576 94084 19580 94140
rect 19580 94084 19636 94140
rect 19636 94084 19640 94140
rect 19576 94080 19640 94084
rect 19656 94140 19720 94144
rect 19656 94084 19660 94140
rect 19660 94084 19716 94140
rect 19716 94084 19720 94140
rect 19656 94080 19720 94084
rect 19736 94140 19800 94144
rect 19736 94084 19740 94140
rect 19740 94084 19796 94140
rect 19796 94084 19800 94140
rect 19736 94080 19800 94084
rect 19816 94140 19880 94144
rect 19816 94084 19820 94140
rect 19820 94084 19876 94140
rect 19876 94084 19880 94140
rect 19816 94080 19880 94084
rect 4216 93596 4280 93600
rect 4216 93540 4220 93596
rect 4220 93540 4276 93596
rect 4276 93540 4280 93596
rect 4216 93536 4280 93540
rect 4296 93596 4360 93600
rect 4296 93540 4300 93596
rect 4300 93540 4356 93596
rect 4356 93540 4360 93596
rect 4296 93536 4360 93540
rect 4376 93596 4440 93600
rect 4376 93540 4380 93596
rect 4380 93540 4436 93596
rect 4436 93540 4440 93596
rect 4376 93536 4440 93540
rect 4456 93596 4520 93600
rect 4456 93540 4460 93596
rect 4460 93540 4516 93596
rect 4516 93540 4520 93596
rect 4456 93536 4520 93540
rect 34936 93596 35000 93600
rect 34936 93540 34940 93596
rect 34940 93540 34996 93596
rect 34996 93540 35000 93596
rect 34936 93536 35000 93540
rect 35016 93596 35080 93600
rect 35016 93540 35020 93596
rect 35020 93540 35076 93596
rect 35076 93540 35080 93596
rect 35016 93536 35080 93540
rect 35096 93596 35160 93600
rect 35096 93540 35100 93596
rect 35100 93540 35156 93596
rect 35156 93540 35160 93596
rect 35096 93536 35160 93540
rect 35176 93596 35240 93600
rect 35176 93540 35180 93596
rect 35180 93540 35236 93596
rect 35236 93540 35240 93596
rect 35176 93536 35240 93540
rect 19576 93052 19640 93056
rect 19576 92996 19580 93052
rect 19580 92996 19636 93052
rect 19636 92996 19640 93052
rect 19576 92992 19640 92996
rect 19656 93052 19720 93056
rect 19656 92996 19660 93052
rect 19660 92996 19716 93052
rect 19716 92996 19720 93052
rect 19656 92992 19720 92996
rect 19736 93052 19800 93056
rect 19736 92996 19740 93052
rect 19740 92996 19796 93052
rect 19796 92996 19800 93052
rect 19736 92992 19800 92996
rect 19816 93052 19880 93056
rect 19816 92996 19820 93052
rect 19820 92996 19876 93052
rect 19876 92996 19880 93052
rect 19816 92992 19880 92996
rect 4216 92508 4280 92512
rect 4216 92452 4220 92508
rect 4220 92452 4276 92508
rect 4276 92452 4280 92508
rect 4216 92448 4280 92452
rect 4296 92508 4360 92512
rect 4296 92452 4300 92508
rect 4300 92452 4356 92508
rect 4356 92452 4360 92508
rect 4296 92448 4360 92452
rect 4376 92508 4440 92512
rect 4376 92452 4380 92508
rect 4380 92452 4436 92508
rect 4436 92452 4440 92508
rect 4376 92448 4440 92452
rect 4456 92508 4520 92512
rect 4456 92452 4460 92508
rect 4460 92452 4516 92508
rect 4516 92452 4520 92508
rect 4456 92448 4520 92452
rect 34936 92508 35000 92512
rect 34936 92452 34940 92508
rect 34940 92452 34996 92508
rect 34996 92452 35000 92508
rect 34936 92448 35000 92452
rect 35016 92508 35080 92512
rect 35016 92452 35020 92508
rect 35020 92452 35076 92508
rect 35076 92452 35080 92508
rect 35016 92448 35080 92452
rect 35096 92508 35160 92512
rect 35096 92452 35100 92508
rect 35100 92452 35156 92508
rect 35156 92452 35160 92508
rect 35096 92448 35160 92452
rect 35176 92508 35240 92512
rect 35176 92452 35180 92508
rect 35180 92452 35236 92508
rect 35236 92452 35240 92508
rect 35176 92448 35240 92452
rect 19576 91964 19640 91968
rect 19576 91908 19580 91964
rect 19580 91908 19636 91964
rect 19636 91908 19640 91964
rect 19576 91904 19640 91908
rect 19656 91964 19720 91968
rect 19656 91908 19660 91964
rect 19660 91908 19716 91964
rect 19716 91908 19720 91964
rect 19656 91904 19720 91908
rect 19736 91964 19800 91968
rect 19736 91908 19740 91964
rect 19740 91908 19796 91964
rect 19796 91908 19800 91964
rect 19736 91904 19800 91908
rect 19816 91964 19880 91968
rect 19816 91908 19820 91964
rect 19820 91908 19876 91964
rect 19876 91908 19880 91964
rect 19816 91904 19880 91908
rect 4216 91420 4280 91424
rect 4216 91364 4220 91420
rect 4220 91364 4276 91420
rect 4276 91364 4280 91420
rect 4216 91360 4280 91364
rect 4296 91420 4360 91424
rect 4296 91364 4300 91420
rect 4300 91364 4356 91420
rect 4356 91364 4360 91420
rect 4296 91360 4360 91364
rect 4376 91420 4440 91424
rect 4376 91364 4380 91420
rect 4380 91364 4436 91420
rect 4436 91364 4440 91420
rect 4376 91360 4440 91364
rect 4456 91420 4520 91424
rect 4456 91364 4460 91420
rect 4460 91364 4516 91420
rect 4516 91364 4520 91420
rect 4456 91360 4520 91364
rect 34936 91420 35000 91424
rect 34936 91364 34940 91420
rect 34940 91364 34996 91420
rect 34996 91364 35000 91420
rect 34936 91360 35000 91364
rect 35016 91420 35080 91424
rect 35016 91364 35020 91420
rect 35020 91364 35076 91420
rect 35076 91364 35080 91420
rect 35016 91360 35080 91364
rect 35096 91420 35160 91424
rect 35096 91364 35100 91420
rect 35100 91364 35156 91420
rect 35156 91364 35160 91420
rect 35096 91360 35160 91364
rect 35176 91420 35240 91424
rect 35176 91364 35180 91420
rect 35180 91364 35236 91420
rect 35236 91364 35240 91420
rect 35176 91360 35240 91364
rect 19576 90876 19640 90880
rect 19576 90820 19580 90876
rect 19580 90820 19636 90876
rect 19636 90820 19640 90876
rect 19576 90816 19640 90820
rect 19656 90876 19720 90880
rect 19656 90820 19660 90876
rect 19660 90820 19716 90876
rect 19716 90820 19720 90876
rect 19656 90816 19720 90820
rect 19736 90876 19800 90880
rect 19736 90820 19740 90876
rect 19740 90820 19796 90876
rect 19796 90820 19800 90876
rect 19736 90816 19800 90820
rect 19816 90876 19880 90880
rect 19816 90820 19820 90876
rect 19820 90820 19876 90876
rect 19876 90820 19880 90876
rect 19816 90816 19880 90820
rect 4216 90332 4280 90336
rect 4216 90276 4220 90332
rect 4220 90276 4276 90332
rect 4276 90276 4280 90332
rect 4216 90272 4280 90276
rect 4296 90332 4360 90336
rect 4296 90276 4300 90332
rect 4300 90276 4356 90332
rect 4356 90276 4360 90332
rect 4296 90272 4360 90276
rect 4376 90332 4440 90336
rect 4376 90276 4380 90332
rect 4380 90276 4436 90332
rect 4436 90276 4440 90332
rect 4376 90272 4440 90276
rect 4456 90332 4520 90336
rect 4456 90276 4460 90332
rect 4460 90276 4516 90332
rect 4516 90276 4520 90332
rect 4456 90272 4520 90276
rect 34936 90332 35000 90336
rect 34936 90276 34940 90332
rect 34940 90276 34996 90332
rect 34996 90276 35000 90332
rect 34936 90272 35000 90276
rect 35016 90332 35080 90336
rect 35016 90276 35020 90332
rect 35020 90276 35076 90332
rect 35076 90276 35080 90332
rect 35016 90272 35080 90276
rect 35096 90332 35160 90336
rect 35096 90276 35100 90332
rect 35100 90276 35156 90332
rect 35156 90276 35160 90332
rect 35096 90272 35160 90276
rect 35176 90332 35240 90336
rect 35176 90276 35180 90332
rect 35180 90276 35236 90332
rect 35236 90276 35240 90332
rect 35176 90272 35240 90276
rect 19576 89788 19640 89792
rect 19576 89732 19580 89788
rect 19580 89732 19636 89788
rect 19636 89732 19640 89788
rect 19576 89728 19640 89732
rect 19656 89788 19720 89792
rect 19656 89732 19660 89788
rect 19660 89732 19716 89788
rect 19716 89732 19720 89788
rect 19656 89728 19720 89732
rect 19736 89788 19800 89792
rect 19736 89732 19740 89788
rect 19740 89732 19796 89788
rect 19796 89732 19800 89788
rect 19736 89728 19800 89732
rect 19816 89788 19880 89792
rect 19816 89732 19820 89788
rect 19820 89732 19876 89788
rect 19876 89732 19880 89788
rect 19816 89728 19880 89732
rect 4216 89244 4280 89248
rect 4216 89188 4220 89244
rect 4220 89188 4276 89244
rect 4276 89188 4280 89244
rect 4216 89184 4280 89188
rect 4296 89244 4360 89248
rect 4296 89188 4300 89244
rect 4300 89188 4356 89244
rect 4356 89188 4360 89244
rect 4296 89184 4360 89188
rect 4376 89244 4440 89248
rect 4376 89188 4380 89244
rect 4380 89188 4436 89244
rect 4436 89188 4440 89244
rect 4376 89184 4440 89188
rect 4456 89244 4520 89248
rect 4456 89188 4460 89244
rect 4460 89188 4516 89244
rect 4516 89188 4520 89244
rect 4456 89184 4520 89188
rect 34936 89244 35000 89248
rect 34936 89188 34940 89244
rect 34940 89188 34996 89244
rect 34996 89188 35000 89244
rect 34936 89184 35000 89188
rect 35016 89244 35080 89248
rect 35016 89188 35020 89244
rect 35020 89188 35076 89244
rect 35076 89188 35080 89244
rect 35016 89184 35080 89188
rect 35096 89244 35160 89248
rect 35096 89188 35100 89244
rect 35100 89188 35156 89244
rect 35156 89188 35160 89244
rect 35096 89184 35160 89188
rect 35176 89244 35240 89248
rect 35176 89188 35180 89244
rect 35180 89188 35236 89244
rect 35236 89188 35240 89244
rect 35176 89184 35240 89188
rect 19576 88700 19640 88704
rect 19576 88644 19580 88700
rect 19580 88644 19636 88700
rect 19636 88644 19640 88700
rect 19576 88640 19640 88644
rect 19656 88700 19720 88704
rect 19656 88644 19660 88700
rect 19660 88644 19716 88700
rect 19716 88644 19720 88700
rect 19656 88640 19720 88644
rect 19736 88700 19800 88704
rect 19736 88644 19740 88700
rect 19740 88644 19796 88700
rect 19796 88644 19800 88700
rect 19736 88640 19800 88644
rect 19816 88700 19880 88704
rect 19816 88644 19820 88700
rect 19820 88644 19876 88700
rect 19876 88644 19880 88700
rect 19816 88640 19880 88644
rect 4216 88156 4280 88160
rect 4216 88100 4220 88156
rect 4220 88100 4276 88156
rect 4276 88100 4280 88156
rect 4216 88096 4280 88100
rect 4296 88156 4360 88160
rect 4296 88100 4300 88156
rect 4300 88100 4356 88156
rect 4356 88100 4360 88156
rect 4296 88096 4360 88100
rect 4376 88156 4440 88160
rect 4376 88100 4380 88156
rect 4380 88100 4436 88156
rect 4436 88100 4440 88156
rect 4376 88096 4440 88100
rect 4456 88156 4520 88160
rect 4456 88100 4460 88156
rect 4460 88100 4516 88156
rect 4516 88100 4520 88156
rect 4456 88096 4520 88100
rect 34936 88156 35000 88160
rect 34936 88100 34940 88156
rect 34940 88100 34996 88156
rect 34996 88100 35000 88156
rect 34936 88096 35000 88100
rect 35016 88156 35080 88160
rect 35016 88100 35020 88156
rect 35020 88100 35076 88156
rect 35076 88100 35080 88156
rect 35016 88096 35080 88100
rect 35096 88156 35160 88160
rect 35096 88100 35100 88156
rect 35100 88100 35156 88156
rect 35156 88100 35160 88156
rect 35096 88096 35160 88100
rect 35176 88156 35240 88160
rect 35176 88100 35180 88156
rect 35180 88100 35236 88156
rect 35236 88100 35240 88156
rect 35176 88096 35240 88100
rect 19576 87612 19640 87616
rect 19576 87556 19580 87612
rect 19580 87556 19636 87612
rect 19636 87556 19640 87612
rect 19576 87552 19640 87556
rect 19656 87612 19720 87616
rect 19656 87556 19660 87612
rect 19660 87556 19716 87612
rect 19716 87556 19720 87612
rect 19656 87552 19720 87556
rect 19736 87612 19800 87616
rect 19736 87556 19740 87612
rect 19740 87556 19796 87612
rect 19796 87556 19800 87612
rect 19736 87552 19800 87556
rect 19816 87612 19880 87616
rect 19816 87556 19820 87612
rect 19820 87556 19876 87612
rect 19876 87556 19880 87612
rect 19816 87552 19880 87556
rect 4216 87068 4280 87072
rect 4216 87012 4220 87068
rect 4220 87012 4276 87068
rect 4276 87012 4280 87068
rect 4216 87008 4280 87012
rect 4296 87068 4360 87072
rect 4296 87012 4300 87068
rect 4300 87012 4356 87068
rect 4356 87012 4360 87068
rect 4296 87008 4360 87012
rect 4376 87068 4440 87072
rect 4376 87012 4380 87068
rect 4380 87012 4436 87068
rect 4436 87012 4440 87068
rect 4376 87008 4440 87012
rect 4456 87068 4520 87072
rect 4456 87012 4460 87068
rect 4460 87012 4516 87068
rect 4516 87012 4520 87068
rect 4456 87008 4520 87012
rect 34936 87068 35000 87072
rect 34936 87012 34940 87068
rect 34940 87012 34996 87068
rect 34996 87012 35000 87068
rect 34936 87008 35000 87012
rect 35016 87068 35080 87072
rect 35016 87012 35020 87068
rect 35020 87012 35076 87068
rect 35076 87012 35080 87068
rect 35016 87008 35080 87012
rect 35096 87068 35160 87072
rect 35096 87012 35100 87068
rect 35100 87012 35156 87068
rect 35156 87012 35160 87068
rect 35096 87008 35160 87012
rect 35176 87068 35240 87072
rect 35176 87012 35180 87068
rect 35180 87012 35236 87068
rect 35236 87012 35240 87068
rect 35176 87008 35240 87012
rect 19576 86524 19640 86528
rect 19576 86468 19580 86524
rect 19580 86468 19636 86524
rect 19636 86468 19640 86524
rect 19576 86464 19640 86468
rect 19656 86524 19720 86528
rect 19656 86468 19660 86524
rect 19660 86468 19716 86524
rect 19716 86468 19720 86524
rect 19656 86464 19720 86468
rect 19736 86524 19800 86528
rect 19736 86468 19740 86524
rect 19740 86468 19796 86524
rect 19796 86468 19800 86524
rect 19736 86464 19800 86468
rect 19816 86524 19880 86528
rect 19816 86468 19820 86524
rect 19820 86468 19876 86524
rect 19876 86468 19880 86524
rect 19816 86464 19880 86468
rect 4216 85980 4280 85984
rect 4216 85924 4220 85980
rect 4220 85924 4276 85980
rect 4276 85924 4280 85980
rect 4216 85920 4280 85924
rect 4296 85980 4360 85984
rect 4296 85924 4300 85980
rect 4300 85924 4356 85980
rect 4356 85924 4360 85980
rect 4296 85920 4360 85924
rect 4376 85980 4440 85984
rect 4376 85924 4380 85980
rect 4380 85924 4436 85980
rect 4436 85924 4440 85980
rect 4376 85920 4440 85924
rect 4456 85980 4520 85984
rect 4456 85924 4460 85980
rect 4460 85924 4516 85980
rect 4516 85924 4520 85980
rect 4456 85920 4520 85924
rect 34936 85980 35000 85984
rect 34936 85924 34940 85980
rect 34940 85924 34996 85980
rect 34996 85924 35000 85980
rect 34936 85920 35000 85924
rect 35016 85980 35080 85984
rect 35016 85924 35020 85980
rect 35020 85924 35076 85980
rect 35076 85924 35080 85980
rect 35016 85920 35080 85924
rect 35096 85980 35160 85984
rect 35096 85924 35100 85980
rect 35100 85924 35156 85980
rect 35156 85924 35160 85980
rect 35096 85920 35160 85924
rect 35176 85980 35240 85984
rect 35176 85924 35180 85980
rect 35180 85924 35236 85980
rect 35236 85924 35240 85980
rect 35176 85920 35240 85924
rect 19576 85436 19640 85440
rect 19576 85380 19580 85436
rect 19580 85380 19636 85436
rect 19636 85380 19640 85436
rect 19576 85376 19640 85380
rect 19656 85436 19720 85440
rect 19656 85380 19660 85436
rect 19660 85380 19716 85436
rect 19716 85380 19720 85436
rect 19656 85376 19720 85380
rect 19736 85436 19800 85440
rect 19736 85380 19740 85436
rect 19740 85380 19796 85436
rect 19796 85380 19800 85436
rect 19736 85376 19800 85380
rect 19816 85436 19880 85440
rect 19816 85380 19820 85436
rect 19820 85380 19876 85436
rect 19876 85380 19880 85436
rect 19816 85376 19880 85380
rect 4216 84892 4280 84896
rect 4216 84836 4220 84892
rect 4220 84836 4276 84892
rect 4276 84836 4280 84892
rect 4216 84832 4280 84836
rect 4296 84892 4360 84896
rect 4296 84836 4300 84892
rect 4300 84836 4356 84892
rect 4356 84836 4360 84892
rect 4296 84832 4360 84836
rect 4376 84892 4440 84896
rect 4376 84836 4380 84892
rect 4380 84836 4436 84892
rect 4436 84836 4440 84892
rect 4376 84832 4440 84836
rect 4456 84892 4520 84896
rect 4456 84836 4460 84892
rect 4460 84836 4516 84892
rect 4516 84836 4520 84892
rect 4456 84832 4520 84836
rect 34936 84892 35000 84896
rect 34936 84836 34940 84892
rect 34940 84836 34996 84892
rect 34996 84836 35000 84892
rect 34936 84832 35000 84836
rect 35016 84892 35080 84896
rect 35016 84836 35020 84892
rect 35020 84836 35076 84892
rect 35076 84836 35080 84892
rect 35016 84832 35080 84836
rect 35096 84892 35160 84896
rect 35096 84836 35100 84892
rect 35100 84836 35156 84892
rect 35156 84836 35160 84892
rect 35096 84832 35160 84836
rect 35176 84892 35240 84896
rect 35176 84836 35180 84892
rect 35180 84836 35236 84892
rect 35236 84836 35240 84892
rect 35176 84832 35240 84836
rect 19576 84348 19640 84352
rect 19576 84292 19580 84348
rect 19580 84292 19636 84348
rect 19636 84292 19640 84348
rect 19576 84288 19640 84292
rect 19656 84348 19720 84352
rect 19656 84292 19660 84348
rect 19660 84292 19716 84348
rect 19716 84292 19720 84348
rect 19656 84288 19720 84292
rect 19736 84348 19800 84352
rect 19736 84292 19740 84348
rect 19740 84292 19796 84348
rect 19796 84292 19800 84348
rect 19736 84288 19800 84292
rect 19816 84348 19880 84352
rect 19816 84292 19820 84348
rect 19820 84292 19876 84348
rect 19876 84292 19880 84348
rect 19816 84288 19880 84292
rect 4216 83804 4280 83808
rect 4216 83748 4220 83804
rect 4220 83748 4276 83804
rect 4276 83748 4280 83804
rect 4216 83744 4280 83748
rect 4296 83804 4360 83808
rect 4296 83748 4300 83804
rect 4300 83748 4356 83804
rect 4356 83748 4360 83804
rect 4296 83744 4360 83748
rect 4376 83804 4440 83808
rect 4376 83748 4380 83804
rect 4380 83748 4436 83804
rect 4436 83748 4440 83804
rect 4376 83744 4440 83748
rect 4456 83804 4520 83808
rect 4456 83748 4460 83804
rect 4460 83748 4516 83804
rect 4516 83748 4520 83804
rect 4456 83744 4520 83748
rect 34936 83804 35000 83808
rect 34936 83748 34940 83804
rect 34940 83748 34996 83804
rect 34996 83748 35000 83804
rect 34936 83744 35000 83748
rect 35016 83804 35080 83808
rect 35016 83748 35020 83804
rect 35020 83748 35076 83804
rect 35076 83748 35080 83804
rect 35016 83744 35080 83748
rect 35096 83804 35160 83808
rect 35096 83748 35100 83804
rect 35100 83748 35156 83804
rect 35156 83748 35160 83804
rect 35096 83744 35160 83748
rect 35176 83804 35240 83808
rect 35176 83748 35180 83804
rect 35180 83748 35236 83804
rect 35236 83748 35240 83804
rect 35176 83744 35240 83748
rect 19576 83260 19640 83264
rect 19576 83204 19580 83260
rect 19580 83204 19636 83260
rect 19636 83204 19640 83260
rect 19576 83200 19640 83204
rect 19656 83260 19720 83264
rect 19656 83204 19660 83260
rect 19660 83204 19716 83260
rect 19716 83204 19720 83260
rect 19656 83200 19720 83204
rect 19736 83260 19800 83264
rect 19736 83204 19740 83260
rect 19740 83204 19796 83260
rect 19796 83204 19800 83260
rect 19736 83200 19800 83204
rect 19816 83260 19880 83264
rect 19816 83204 19820 83260
rect 19820 83204 19876 83260
rect 19876 83204 19880 83260
rect 19816 83200 19880 83204
rect 4216 82716 4280 82720
rect 4216 82660 4220 82716
rect 4220 82660 4276 82716
rect 4276 82660 4280 82716
rect 4216 82656 4280 82660
rect 4296 82716 4360 82720
rect 4296 82660 4300 82716
rect 4300 82660 4356 82716
rect 4356 82660 4360 82716
rect 4296 82656 4360 82660
rect 4376 82716 4440 82720
rect 4376 82660 4380 82716
rect 4380 82660 4436 82716
rect 4436 82660 4440 82716
rect 4376 82656 4440 82660
rect 4456 82716 4520 82720
rect 4456 82660 4460 82716
rect 4460 82660 4516 82716
rect 4516 82660 4520 82716
rect 4456 82656 4520 82660
rect 34936 82716 35000 82720
rect 34936 82660 34940 82716
rect 34940 82660 34996 82716
rect 34996 82660 35000 82716
rect 34936 82656 35000 82660
rect 35016 82716 35080 82720
rect 35016 82660 35020 82716
rect 35020 82660 35076 82716
rect 35076 82660 35080 82716
rect 35016 82656 35080 82660
rect 35096 82716 35160 82720
rect 35096 82660 35100 82716
rect 35100 82660 35156 82716
rect 35156 82660 35160 82716
rect 35096 82656 35160 82660
rect 35176 82716 35240 82720
rect 35176 82660 35180 82716
rect 35180 82660 35236 82716
rect 35236 82660 35240 82716
rect 35176 82656 35240 82660
rect 19576 82172 19640 82176
rect 19576 82116 19580 82172
rect 19580 82116 19636 82172
rect 19636 82116 19640 82172
rect 19576 82112 19640 82116
rect 19656 82172 19720 82176
rect 19656 82116 19660 82172
rect 19660 82116 19716 82172
rect 19716 82116 19720 82172
rect 19656 82112 19720 82116
rect 19736 82172 19800 82176
rect 19736 82116 19740 82172
rect 19740 82116 19796 82172
rect 19796 82116 19800 82172
rect 19736 82112 19800 82116
rect 19816 82172 19880 82176
rect 19816 82116 19820 82172
rect 19820 82116 19876 82172
rect 19876 82116 19880 82172
rect 19816 82112 19880 82116
rect 4216 81628 4280 81632
rect 4216 81572 4220 81628
rect 4220 81572 4276 81628
rect 4276 81572 4280 81628
rect 4216 81568 4280 81572
rect 4296 81628 4360 81632
rect 4296 81572 4300 81628
rect 4300 81572 4356 81628
rect 4356 81572 4360 81628
rect 4296 81568 4360 81572
rect 4376 81628 4440 81632
rect 4376 81572 4380 81628
rect 4380 81572 4436 81628
rect 4436 81572 4440 81628
rect 4376 81568 4440 81572
rect 4456 81628 4520 81632
rect 4456 81572 4460 81628
rect 4460 81572 4516 81628
rect 4516 81572 4520 81628
rect 4456 81568 4520 81572
rect 34936 81628 35000 81632
rect 34936 81572 34940 81628
rect 34940 81572 34996 81628
rect 34996 81572 35000 81628
rect 34936 81568 35000 81572
rect 35016 81628 35080 81632
rect 35016 81572 35020 81628
rect 35020 81572 35076 81628
rect 35076 81572 35080 81628
rect 35016 81568 35080 81572
rect 35096 81628 35160 81632
rect 35096 81572 35100 81628
rect 35100 81572 35156 81628
rect 35156 81572 35160 81628
rect 35096 81568 35160 81572
rect 35176 81628 35240 81632
rect 35176 81572 35180 81628
rect 35180 81572 35236 81628
rect 35236 81572 35240 81628
rect 35176 81568 35240 81572
rect 19576 81084 19640 81088
rect 19576 81028 19580 81084
rect 19580 81028 19636 81084
rect 19636 81028 19640 81084
rect 19576 81024 19640 81028
rect 19656 81084 19720 81088
rect 19656 81028 19660 81084
rect 19660 81028 19716 81084
rect 19716 81028 19720 81084
rect 19656 81024 19720 81028
rect 19736 81084 19800 81088
rect 19736 81028 19740 81084
rect 19740 81028 19796 81084
rect 19796 81028 19800 81084
rect 19736 81024 19800 81028
rect 19816 81084 19880 81088
rect 19816 81028 19820 81084
rect 19820 81028 19876 81084
rect 19876 81028 19880 81084
rect 19816 81024 19880 81028
rect 4216 80540 4280 80544
rect 4216 80484 4220 80540
rect 4220 80484 4276 80540
rect 4276 80484 4280 80540
rect 4216 80480 4280 80484
rect 4296 80540 4360 80544
rect 4296 80484 4300 80540
rect 4300 80484 4356 80540
rect 4356 80484 4360 80540
rect 4296 80480 4360 80484
rect 4376 80540 4440 80544
rect 4376 80484 4380 80540
rect 4380 80484 4436 80540
rect 4436 80484 4440 80540
rect 4376 80480 4440 80484
rect 4456 80540 4520 80544
rect 4456 80484 4460 80540
rect 4460 80484 4516 80540
rect 4516 80484 4520 80540
rect 4456 80480 4520 80484
rect 34936 80540 35000 80544
rect 34936 80484 34940 80540
rect 34940 80484 34996 80540
rect 34996 80484 35000 80540
rect 34936 80480 35000 80484
rect 35016 80540 35080 80544
rect 35016 80484 35020 80540
rect 35020 80484 35076 80540
rect 35076 80484 35080 80540
rect 35016 80480 35080 80484
rect 35096 80540 35160 80544
rect 35096 80484 35100 80540
rect 35100 80484 35156 80540
rect 35156 80484 35160 80540
rect 35096 80480 35160 80484
rect 35176 80540 35240 80544
rect 35176 80484 35180 80540
rect 35180 80484 35236 80540
rect 35236 80484 35240 80540
rect 35176 80480 35240 80484
rect 19576 79996 19640 80000
rect 19576 79940 19580 79996
rect 19580 79940 19636 79996
rect 19636 79940 19640 79996
rect 19576 79936 19640 79940
rect 19656 79996 19720 80000
rect 19656 79940 19660 79996
rect 19660 79940 19716 79996
rect 19716 79940 19720 79996
rect 19656 79936 19720 79940
rect 19736 79996 19800 80000
rect 19736 79940 19740 79996
rect 19740 79940 19796 79996
rect 19796 79940 19800 79996
rect 19736 79936 19800 79940
rect 19816 79996 19880 80000
rect 19816 79940 19820 79996
rect 19820 79940 19876 79996
rect 19876 79940 19880 79996
rect 19816 79936 19880 79940
rect 4216 79452 4280 79456
rect 4216 79396 4220 79452
rect 4220 79396 4276 79452
rect 4276 79396 4280 79452
rect 4216 79392 4280 79396
rect 4296 79452 4360 79456
rect 4296 79396 4300 79452
rect 4300 79396 4356 79452
rect 4356 79396 4360 79452
rect 4296 79392 4360 79396
rect 4376 79452 4440 79456
rect 4376 79396 4380 79452
rect 4380 79396 4436 79452
rect 4436 79396 4440 79452
rect 4376 79392 4440 79396
rect 4456 79452 4520 79456
rect 4456 79396 4460 79452
rect 4460 79396 4516 79452
rect 4516 79396 4520 79452
rect 4456 79392 4520 79396
rect 34936 79452 35000 79456
rect 34936 79396 34940 79452
rect 34940 79396 34996 79452
rect 34996 79396 35000 79452
rect 34936 79392 35000 79396
rect 35016 79452 35080 79456
rect 35016 79396 35020 79452
rect 35020 79396 35076 79452
rect 35076 79396 35080 79452
rect 35016 79392 35080 79396
rect 35096 79452 35160 79456
rect 35096 79396 35100 79452
rect 35100 79396 35156 79452
rect 35156 79396 35160 79452
rect 35096 79392 35160 79396
rect 35176 79452 35240 79456
rect 35176 79396 35180 79452
rect 35180 79396 35236 79452
rect 35236 79396 35240 79452
rect 35176 79392 35240 79396
rect 19576 78908 19640 78912
rect 19576 78852 19580 78908
rect 19580 78852 19636 78908
rect 19636 78852 19640 78908
rect 19576 78848 19640 78852
rect 19656 78908 19720 78912
rect 19656 78852 19660 78908
rect 19660 78852 19716 78908
rect 19716 78852 19720 78908
rect 19656 78848 19720 78852
rect 19736 78908 19800 78912
rect 19736 78852 19740 78908
rect 19740 78852 19796 78908
rect 19796 78852 19800 78908
rect 19736 78848 19800 78852
rect 19816 78908 19880 78912
rect 19816 78852 19820 78908
rect 19820 78852 19876 78908
rect 19876 78852 19880 78908
rect 19816 78848 19880 78852
rect 4216 78364 4280 78368
rect 4216 78308 4220 78364
rect 4220 78308 4276 78364
rect 4276 78308 4280 78364
rect 4216 78304 4280 78308
rect 4296 78364 4360 78368
rect 4296 78308 4300 78364
rect 4300 78308 4356 78364
rect 4356 78308 4360 78364
rect 4296 78304 4360 78308
rect 4376 78364 4440 78368
rect 4376 78308 4380 78364
rect 4380 78308 4436 78364
rect 4436 78308 4440 78364
rect 4376 78304 4440 78308
rect 4456 78364 4520 78368
rect 4456 78308 4460 78364
rect 4460 78308 4516 78364
rect 4516 78308 4520 78364
rect 4456 78304 4520 78308
rect 34936 78364 35000 78368
rect 34936 78308 34940 78364
rect 34940 78308 34996 78364
rect 34996 78308 35000 78364
rect 34936 78304 35000 78308
rect 35016 78364 35080 78368
rect 35016 78308 35020 78364
rect 35020 78308 35076 78364
rect 35076 78308 35080 78364
rect 35016 78304 35080 78308
rect 35096 78364 35160 78368
rect 35096 78308 35100 78364
rect 35100 78308 35156 78364
rect 35156 78308 35160 78364
rect 35096 78304 35160 78308
rect 35176 78364 35240 78368
rect 35176 78308 35180 78364
rect 35180 78308 35236 78364
rect 35236 78308 35240 78364
rect 35176 78304 35240 78308
rect 19576 77820 19640 77824
rect 19576 77764 19580 77820
rect 19580 77764 19636 77820
rect 19636 77764 19640 77820
rect 19576 77760 19640 77764
rect 19656 77820 19720 77824
rect 19656 77764 19660 77820
rect 19660 77764 19716 77820
rect 19716 77764 19720 77820
rect 19656 77760 19720 77764
rect 19736 77820 19800 77824
rect 19736 77764 19740 77820
rect 19740 77764 19796 77820
rect 19796 77764 19800 77820
rect 19736 77760 19800 77764
rect 19816 77820 19880 77824
rect 19816 77764 19820 77820
rect 19820 77764 19876 77820
rect 19876 77764 19880 77820
rect 19816 77760 19880 77764
rect 4216 77276 4280 77280
rect 4216 77220 4220 77276
rect 4220 77220 4276 77276
rect 4276 77220 4280 77276
rect 4216 77216 4280 77220
rect 4296 77276 4360 77280
rect 4296 77220 4300 77276
rect 4300 77220 4356 77276
rect 4356 77220 4360 77276
rect 4296 77216 4360 77220
rect 4376 77276 4440 77280
rect 4376 77220 4380 77276
rect 4380 77220 4436 77276
rect 4436 77220 4440 77276
rect 4376 77216 4440 77220
rect 4456 77276 4520 77280
rect 4456 77220 4460 77276
rect 4460 77220 4516 77276
rect 4516 77220 4520 77276
rect 4456 77216 4520 77220
rect 34936 77276 35000 77280
rect 34936 77220 34940 77276
rect 34940 77220 34996 77276
rect 34996 77220 35000 77276
rect 34936 77216 35000 77220
rect 35016 77276 35080 77280
rect 35016 77220 35020 77276
rect 35020 77220 35076 77276
rect 35076 77220 35080 77276
rect 35016 77216 35080 77220
rect 35096 77276 35160 77280
rect 35096 77220 35100 77276
rect 35100 77220 35156 77276
rect 35156 77220 35160 77276
rect 35096 77216 35160 77220
rect 35176 77276 35240 77280
rect 35176 77220 35180 77276
rect 35180 77220 35236 77276
rect 35236 77220 35240 77276
rect 35176 77216 35240 77220
rect 19576 76732 19640 76736
rect 19576 76676 19580 76732
rect 19580 76676 19636 76732
rect 19636 76676 19640 76732
rect 19576 76672 19640 76676
rect 19656 76732 19720 76736
rect 19656 76676 19660 76732
rect 19660 76676 19716 76732
rect 19716 76676 19720 76732
rect 19656 76672 19720 76676
rect 19736 76732 19800 76736
rect 19736 76676 19740 76732
rect 19740 76676 19796 76732
rect 19796 76676 19800 76732
rect 19736 76672 19800 76676
rect 19816 76732 19880 76736
rect 19816 76676 19820 76732
rect 19820 76676 19876 76732
rect 19876 76676 19880 76732
rect 19816 76672 19880 76676
rect 4216 76188 4280 76192
rect 4216 76132 4220 76188
rect 4220 76132 4276 76188
rect 4276 76132 4280 76188
rect 4216 76128 4280 76132
rect 4296 76188 4360 76192
rect 4296 76132 4300 76188
rect 4300 76132 4356 76188
rect 4356 76132 4360 76188
rect 4296 76128 4360 76132
rect 4376 76188 4440 76192
rect 4376 76132 4380 76188
rect 4380 76132 4436 76188
rect 4436 76132 4440 76188
rect 4376 76128 4440 76132
rect 4456 76188 4520 76192
rect 4456 76132 4460 76188
rect 4460 76132 4516 76188
rect 4516 76132 4520 76188
rect 4456 76128 4520 76132
rect 34936 76188 35000 76192
rect 34936 76132 34940 76188
rect 34940 76132 34996 76188
rect 34996 76132 35000 76188
rect 34936 76128 35000 76132
rect 35016 76188 35080 76192
rect 35016 76132 35020 76188
rect 35020 76132 35076 76188
rect 35076 76132 35080 76188
rect 35016 76128 35080 76132
rect 35096 76188 35160 76192
rect 35096 76132 35100 76188
rect 35100 76132 35156 76188
rect 35156 76132 35160 76188
rect 35096 76128 35160 76132
rect 35176 76188 35240 76192
rect 35176 76132 35180 76188
rect 35180 76132 35236 76188
rect 35236 76132 35240 76188
rect 35176 76128 35240 76132
rect 19576 75644 19640 75648
rect 19576 75588 19580 75644
rect 19580 75588 19636 75644
rect 19636 75588 19640 75644
rect 19576 75584 19640 75588
rect 19656 75644 19720 75648
rect 19656 75588 19660 75644
rect 19660 75588 19716 75644
rect 19716 75588 19720 75644
rect 19656 75584 19720 75588
rect 19736 75644 19800 75648
rect 19736 75588 19740 75644
rect 19740 75588 19796 75644
rect 19796 75588 19800 75644
rect 19736 75584 19800 75588
rect 19816 75644 19880 75648
rect 19816 75588 19820 75644
rect 19820 75588 19876 75644
rect 19876 75588 19880 75644
rect 19816 75584 19880 75588
rect 4216 75100 4280 75104
rect 4216 75044 4220 75100
rect 4220 75044 4276 75100
rect 4276 75044 4280 75100
rect 4216 75040 4280 75044
rect 4296 75100 4360 75104
rect 4296 75044 4300 75100
rect 4300 75044 4356 75100
rect 4356 75044 4360 75100
rect 4296 75040 4360 75044
rect 4376 75100 4440 75104
rect 4376 75044 4380 75100
rect 4380 75044 4436 75100
rect 4436 75044 4440 75100
rect 4376 75040 4440 75044
rect 4456 75100 4520 75104
rect 4456 75044 4460 75100
rect 4460 75044 4516 75100
rect 4516 75044 4520 75100
rect 4456 75040 4520 75044
rect 34936 75100 35000 75104
rect 34936 75044 34940 75100
rect 34940 75044 34996 75100
rect 34996 75044 35000 75100
rect 34936 75040 35000 75044
rect 35016 75100 35080 75104
rect 35016 75044 35020 75100
rect 35020 75044 35076 75100
rect 35076 75044 35080 75100
rect 35016 75040 35080 75044
rect 35096 75100 35160 75104
rect 35096 75044 35100 75100
rect 35100 75044 35156 75100
rect 35156 75044 35160 75100
rect 35096 75040 35160 75044
rect 35176 75100 35240 75104
rect 35176 75044 35180 75100
rect 35180 75044 35236 75100
rect 35236 75044 35240 75100
rect 35176 75040 35240 75044
rect 19576 74556 19640 74560
rect 19576 74500 19580 74556
rect 19580 74500 19636 74556
rect 19636 74500 19640 74556
rect 19576 74496 19640 74500
rect 19656 74556 19720 74560
rect 19656 74500 19660 74556
rect 19660 74500 19716 74556
rect 19716 74500 19720 74556
rect 19656 74496 19720 74500
rect 19736 74556 19800 74560
rect 19736 74500 19740 74556
rect 19740 74500 19796 74556
rect 19796 74500 19800 74556
rect 19736 74496 19800 74500
rect 19816 74556 19880 74560
rect 19816 74500 19820 74556
rect 19820 74500 19876 74556
rect 19876 74500 19880 74556
rect 19816 74496 19880 74500
rect 4216 74012 4280 74016
rect 4216 73956 4220 74012
rect 4220 73956 4276 74012
rect 4276 73956 4280 74012
rect 4216 73952 4280 73956
rect 4296 74012 4360 74016
rect 4296 73956 4300 74012
rect 4300 73956 4356 74012
rect 4356 73956 4360 74012
rect 4296 73952 4360 73956
rect 4376 74012 4440 74016
rect 4376 73956 4380 74012
rect 4380 73956 4436 74012
rect 4436 73956 4440 74012
rect 4376 73952 4440 73956
rect 4456 74012 4520 74016
rect 4456 73956 4460 74012
rect 4460 73956 4516 74012
rect 4516 73956 4520 74012
rect 4456 73952 4520 73956
rect 34936 74012 35000 74016
rect 34936 73956 34940 74012
rect 34940 73956 34996 74012
rect 34996 73956 35000 74012
rect 34936 73952 35000 73956
rect 35016 74012 35080 74016
rect 35016 73956 35020 74012
rect 35020 73956 35076 74012
rect 35076 73956 35080 74012
rect 35016 73952 35080 73956
rect 35096 74012 35160 74016
rect 35096 73956 35100 74012
rect 35100 73956 35156 74012
rect 35156 73956 35160 74012
rect 35096 73952 35160 73956
rect 35176 74012 35240 74016
rect 35176 73956 35180 74012
rect 35180 73956 35236 74012
rect 35236 73956 35240 74012
rect 35176 73952 35240 73956
rect 19576 73468 19640 73472
rect 19576 73412 19580 73468
rect 19580 73412 19636 73468
rect 19636 73412 19640 73468
rect 19576 73408 19640 73412
rect 19656 73468 19720 73472
rect 19656 73412 19660 73468
rect 19660 73412 19716 73468
rect 19716 73412 19720 73468
rect 19656 73408 19720 73412
rect 19736 73468 19800 73472
rect 19736 73412 19740 73468
rect 19740 73412 19796 73468
rect 19796 73412 19800 73468
rect 19736 73408 19800 73412
rect 19816 73468 19880 73472
rect 19816 73412 19820 73468
rect 19820 73412 19876 73468
rect 19876 73412 19880 73468
rect 19816 73408 19880 73412
rect 4216 72924 4280 72928
rect 4216 72868 4220 72924
rect 4220 72868 4276 72924
rect 4276 72868 4280 72924
rect 4216 72864 4280 72868
rect 4296 72924 4360 72928
rect 4296 72868 4300 72924
rect 4300 72868 4356 72924
rect 4356 72868 4360 72924
rect 4296 72864 4360 72868
rect 4376 72924 4440 72928
rect 4376 72868 4380 72924
rect 4380 72868 4436 72924
rect 4436 72868 4440 72924
rect 4376 72864 4440 72868
rect 4456 72924 4520 72928
rect 4456 72868 4460 72924
rect 4460 72868 4516 72924
rect 4516 72868 4520 72924
rect 4456 72864 4520 72868
rect 34936 72924 35000 72928
rect 34936 72868 34940 72924
rect 34940 72868 34996 72924
rect 34996 72868 35000 72924
rect 34936 72864 35000 72868
rect 35016 72924 35080 72928
rect 35016 72868 35020 72924
rect 35020 72868 35076 72924
rect 35076 72868 35080 72924
rect 35016 72864 35080 72868
rect 35096 72924 35160 72928
rect 35096 72868 35100 72924
rect 35100 72868 35156 72924
rect 35156 72868 35160 72924
rect 35096 72864 35160 72868
rect 35176 72924 35240 72928
rect 35176 72868 35180 72924
rect 35180 72868 35236 72924
rect 35236 72868 35240 72924
rect 35176 72864 35240 72868
rect 19576 72380 19640 72384
rect 19576 72324 19580 72380
rect 19580 72324 19636 72380
rect 19636 72324 19640 72380
rect 19576 72320 19640 72324
rect 19656 72380 19720 72384
rect 19656 72324 19660 72380
rect 19660 72324 19716 72380
rect 19716 72324 19720 72380
rect 19656 72320 19720 72324
rect 19736 72380 19800 72384
rect 19736 72324 19740 72380
rect 19740 72324 19796 72380
rect 19796 72324 19800 72380
rect 19736 72320 19800 72324
rect 19816 72380 19880 72384
rect 19816 72324 19820 72380
rect 19820 72324 19876 72380
rect 19876 72324 19880 72380
rect 19816 72320 19880 72324
rect 4216 71836 4280 71840
rect 4216 71780 4220 71836
rect 4220 71780 4276 71836
rect 4276 71780 4280 71836
rect 4216 71776 4280 71780
rect 4296 71836 4360 71840
rect 4296 71780 4300 71836
rect 4300 71780 4356 71836
rect 4356 71780 4360 71836
rect 4296 71776 4360 71780
rect 4376 71836 4440 71840
rect 4376 71780 4380 71836
rect 4380 71780 4436 71836
rect 4436 71780 4440 71836
rect 4376 71776 4440 71780
rect 4456 71836 4520 71840
rect 4456 71780 4460 71836
rect 4460 71780 4516 71836
rect 4516 71780 4520 71836
rect 4456 71776 4520 71780
rect 34936 71836 35000 71840
rect 34936 71780 34940 71836
rect 34940 71780 34996 71836
rect 34996 71780 35000 71836
rect 34936 71776 35000 71780
rect 35016 71836 35080 71840
rect 35016 71780 35020 71836
rect 35020 71780 35076 71836
rect 35076 71780 35080 71836
rect 35016 71776 35080 71780
rect 35096 71836 35160 71840
rect 35096 71780 35100 71836
rect 35100 71780 35156 71836
rect 35156 71780 35160 71836
rect 35096 71776 35160 71780
rect 35176 71836 35240 71840
rect 35176 71780 35180 71836
rect 35180 71780 35236 71836
rect 35236 71780 35240 71836
rect 35176 71776 35240 71780
rect 19576 71292 19640 71296
rect 19576 71236 19580 71292
rect 19580 71236 19636 71292
rect 19636 71236 19640 71292
rect 19576 71232 19640 71236
rect 19656 71292 19720 71296
rect 19656 71236 19660 71292
rect 19660 71236 19716 71292
rect 19716 71236 19720 71292
rect 19656 71232 19720 71236
rect 19736 71292 19800 71296
rect 19736 71236 19740 71292
rect 19740 71236 19796 71292
rect 19796 71236 19800 71292
rect 19736 71232 19800 71236
rect 19816 71292 19880 71296
rect 19816 71236 19820 71292
rect 19820 71236 19876 71292
rect 19876 71236 19880 71292
rect 19816 71232 19880 71236
rect 4216 70748 4280 70752
rect 4216 70692 4220 70748
rect 4220 70692 4276 70748
rect 4276 70692 4280 70748
rect 4216 70688 4280 70692
rect 4296 70748 4360 70752
rect 4296 70692 4300 70748
rect 4300 70692 4356 70748
rect 4356 70692 4360 70748
rect 4296 70688 4360 70692
rect 4376 70748 4440 70752
rect 4376 70692 4380 70748
rect 4380 70692 4436 70748
rect 4436 70692 4440 70748
rect 4376 70688 4440 70692
rect 4456 70748 4520 70752
rect 4456 70692 4460 70748
rect 4460 70692 4516 70748
rect 4516 70692 4520 70748
rect 4456 70688 4520 70692
rect 34936 70748 35000 70752
rect 34936 70692 34940 70748
rect 34940 70692 34996 70748
rect 34996 70692 35000 70748
rect 34936 70688 35000 70692
rect 35016 70748 35080 70752
rect 35016 70692 35020 70748
rect 35020 70692 35076 70748
rect 35076 70692 35080 70748
rect 35016 70688 35080 70692
rect 35096 70748 35160 70752
rect 35096 70692 35100 70748
rect 35100 70692 35156 70748
rect 35156 70692 35160 70748
rect 35096 70688 35160 70692
rect 35176 70748 35240 70752
rect 35176 70692 35180 70748
rect 35180 70692 35236 70748
rect 35236 70692 35240 70748
rect 35176 70688 35240 70692
rect 19576 70204 19640 70208
rect 19576 70148 19580 70204
rect 19580 70148 19636 70204
rect 19636 70148 19640 70204
rect 19576 70144 19640 70148
rect 19656 70204 19720 70208
rect 19656 70148 19660 70204
rect 19660 70148 19716 70204
rect 19716 70148 19720 70204
rect 19656 70144 19720 70148
rect 19736 70204 19800 70208
rect 19736 70148 19740 70204
rect 19740 70148 19796 70204
rect 19796 70148 19800 70204
rect 19736 70144 19800 70148
rect 19816 70204 19880 70208
rect 19816 70148 19820 70204
rect 19820 70148 19876 70204
rect 19876 70148 19880 70204
rect 19816 70144 19880 70148
rect 4216 69660 4280 69664
rect 4216 69604 4220 69660
rect 4220 69604 4276 69660
rect 4276 69604 4280 69660
rect 4216 69600 4280 69604
rect 4296 69660 4360 69664
rect 4296 69604 4300 69660
rect 4300 69604 4356 69660
rect 4356 69604 4360 69660
rect 4296 69600 4360 69604
rect 4376 69660 4440 69664
rect 4376 69604 4380 69660
rect 4380 69604 4436 69660
rect 4436 69604 4440 69660
rect 4376 69600 4440 69604
rect 4456 69660 4520 69664
rect 4456 69604 4460 69660
rect 4460 69604 4516 69660
rect 4516 69604 4520 69660
rect 4456 69600 4520 69604
rect 34936 69660 35000 69664
rect 34936 69604 34940 69660
rect 34940 69604 34996 69660
rect 34996 69604 35000 69660
rect 34936 69600 35000 69604
rect 35016 69660 35080 69664
rect 35016 69604 35020 69660
rect 35020 69604 35076 69660
rect 35076 69604 35080 69660
rect 35016 69600 35080 69604
rect 35096 69660 35160 69664
rect 35096 69604 35100 69660
rect 35100 69604 35156 69660
rect 35156 69604 35160 69660
rect 35096 69600 35160 69604
rect 35176 69660 35240 69664
rect 35176 69604 35180 69660
rect 35180 69604 35236 69660
rect 35236 69604 35240 69660
rect 35176 69600 35240 69604
rect 19576 69116 19640 69120
rect 19576 69060 19580 69116
rect 19580 69060 19636 69116
rect 19636 69060 19640 69116
rect 19576 69056 19640 69060
rect 19656 69116 19720 69120
rect 19656 69060 19660 69116
rect 19660 69060 19716 69116
rect 19716 69060 19720 69116
rect 19656 69056 19720 69060
rect 19736 69116 19800 69120
rect 19736 69060 19740 69116
rect 19740 69060 19796 69116
rect 19796 69060 19800 69116
rect 19736 69056 19800 69060
rect 19816 69116 19880 69120
rect 19816 69060 19820 69116
rect 19820 69060 19876 69116
rect 19876 69060 19880 69116
rect 19816 69056 19880 69060
rect 4216 68572 4280 68576
rect 4216 68516 4220 68572
rect 4220 68516 4276 68572
rect 4276 68516 4280 68572
rect 4216 68512 4280 68516
rect 4296 68572 4360 68576
rect 4296 68516 4300 68572
rect 4300 68516 4356 68572
rect 4356 68516 4360 68572
rect 4296 68512 4360 68516
rect 4376 68572 4440 68576
rect 4376 68516 4380 68572
rect 4380 68516 4436 68572
rect 4436 68516 4440 68572
rect 4376 68512 4440 68516
rect 4456 68572 4520 68576
rect 4456 68516 4460 68572
rect 4460 68516 4516 68572
rect 4516 68516 4520 68572
rect 4456 68512 4520 68516
rect 34936 68572 35000 68576
rect 34936 68516 34940 68572
rect 34940 68516 34996 68572
rect 34996 68516 35000 68572
rect 34936 68512 35000 68516
rect 35016 68572 35080 68576
rect 35016 68516 35020 68572
rect 35020 68516 35076 68572
rect 35076 68516 35080 68572
rect 35016 68512 35080 68516
rect 35096 68572 35160 68576
rect 35096 68516 35100 68572
rect 35100 68516 35156 68572
rect 35156 68516 35160 68572
rect 35096 68512 35160 68516
rect 35176 68572 35240 68576
rect 35176 68516 35180 68572
rect 35180 68516 35236 68572
rect 35236 68516 35240 68572
rect 35176 68512 35240 68516
rect 19576 68028 19640 68032
rect 19576 67972 19580 68028
rect 19580 67972 19636 68028
rect 19636 67972 19640 68028
rect 19576 67968 19640 67972
rect 19656 68028 19720 68032
rect 19656 67972 19660 68028
rect 19660 67972 19716 68028
rect 19716 67972 19720 68028
rect 19656 67968 19720 67972
rect 19736 68028 19800 68032
rect 19736 67972 19740 68028
rect 19740 67972 19796 68028
rect 19796 67972 19800 68028
rect 19736 67968 19800 67972
rect 19816 68028 19880 68032
rect 19816 67972 19820 68028
rect 19820 67972 19876 68028
rect 19876 67972 19880 68028
rect 19816 67968 19880 67972
rect 4216 67484 4280 67488
rect 4216 67428 4220 67484
rect 4220 67428 4276 67484
rect 4276 67428 4280 67484
rect 4216 67424 4280 67428
rect 4296 67484 4360 67488
rect 4296 67428 4300 67484
rect 4300 67428 4356 67484
rect 4356 67428 4360 67484
rect 4296 67424 4360 67428
rect 4376 67484 4440 67488
rect 4376 67428 4380 67484
rect 4380 67428 4436 67484
rect 4436 67428 4440 67484
rect 4376 67424 4440 67428
rect 4456 67484 4520 67488
rect 4456 67428 4460 67484
rect 4460 67428 4516 67484
rect 4516 67428 4520 67484
rect 4456 67424 4520 67428
rect 34936 67484 35000 67488
rect 34936 67428 34940 67484
rect 34940 67428 34996 67484
rect 34996 67428 35000 67484
rect 34936 67424 35000 67428
rect 35016 67484 35080 67488
rect 35016 67428 35020 67484
rect 35020 67428 35076 67484
rect 35076 67428 35080 67484
rect 35016 67424 35080 67428
rect 35096 67484 35160 67488
rect 35096 67428 35100 67484
rect 35100 67428 35156 67484
rect 35156 67428 35160 67484
rect 35096 67424 35160 67428
rect 35176 67484 35240 67488
rect 35176 67428 35180 67484
rect 35180 67428 35236 67484
rect 35236 67428 35240 67484
rect 35176 67424 35240 67428
rect 19576 66940 19640 66944
rect 19576 66884 19580 66940
rect 19580 66884 19636 66940
rect 19636 66884 19640 66940
rect 19576 66880 19640 66884
rect 19656 66940 19720 66944
rect 19656 66884 19660 66940
rect 19660 66884 19716 66940
rect 19716 66884 19720 66940
rect 19656 66880 19720 66884
rect 19736 66940 19800 66944
rect 19736 66884 19740 66940
rect 19740 66884 19796 66940
rect 19796 66884 19800 66940
rect 19736 66880 19800 66884
rect 19816 66940 19880 66944
rect 19816 66884 19820 66940
rect 19820 66884 19876 66940
rect 19876 66884 19880 66940
rect 19816 66880 19880 66884
rect 4216 66396 4280 66400
rect 4216 66340 4220 66396
rect 4220 66340 4276 66396
rect 4276 66340 4280 66396
rect 4216 66336 4280 66340
rect 4296 66396 4360 66400
rect 4296 66340 4300 66396
rect 4300 66340 4356 66396
rect 4356 66340 4360 66396
rect 4296 66336 4360 66340
rect 4376 66396 4440 66400
rect 4376 66340 4380 66396
rect 4380 66340 4436 66396
rect 4436 66340 4440 66396
rect 4376 66336 4440 66340
rect 4456 66396 4520 66400
rect 4456 66340 4460 66396
rect 4460 66340 4516 66396
rect 4516 66340 4520 66396
rect 4456 66336 4520 66340
rect 34936 66396 35000 66400
rect 34936 66340 34940 66396
rect 34940 66340 34996 66396
rect 34996 66340 35000 66396
rect 34936 66336 35000 66340
rect 35016 66396 35080 66400
rect 35016 66340 35020 66396
rect 35020 66340 35076 66396
rect 35076 66340 35080 66396
rect 35016 66336 35080 66340
rect 35096 66396 35160 66400
rect 35096 66340 35100 66396
rect 35100 66340 35156 66396
rect 35156 66340 35160 66396
rect 35096 66336 35160 66340
rect 35176 66396 35240 66400
rect 35176 66340 35180 66396
rect 35180 66340 35236 66396
rect 35236 66340 35240 66396
rect 35176 66336 35240 66340
rect 19576 65852 19640 65856
rect 19576 65796 19580 65852
rect 19580 65796 19636 65852
rect 19636 65796 19640 65852
rect 19576 65792 19640 65796
rect 19656 65852 19720 65856
rect 19656 65796 19660 65852
rect 19660 65796 19716 65852
rect 19716 65796 19720 65852
rect 19656 65792 19720 65796
rect 19736 65852 19800 65856
rect 19736 65796 19740 65852
rect 19740 65796 19796 65852
rect 19796 65796 19800 65852
rect 19736 65792 19800 65796
rect 19816 65852 19880 65856
rect 19816 65796 19820 65852
rect 19820 65796 19876 65852
rect 19876 65796 19880 65852
rect 19816 65792 19880 65796
rect 4216 65308 4280 65312
rect 4216 65252 4220 65308
rect 4220 65252 4276 65308
rect 4276 65252 4280 65308
rect 4216 65248 4280 65252
rect 4296 65308 4360 65312
rect 4296 65252 4300 65308
rect 4300 65252 4356 65308
rect 4356 65252 4360 65308
rect 4296 65248 4360 65252
rect 4376 65308 4440 65312
rect 4376 65252 4380 65308
rect 4380 65252 4436 65308
rect 4436 65252 4440 65308
rect 4376 65248 4440 65252
rect 4456 65308 4520 65312
rect 4456 65252 4460 65308
rect 4460 65252 4516 65308
rect 4516 65252 4520 65308
rect 4456 65248 4520 65252
rect 34936 65308 35000 65312
rect 34936 65252 34940 65308
rect 34940 65252 34996 65308
rect 34996 65252 35000 65308
rect 34936 65248 35000 65252
rect 35016 65308 35080 65312
rect 35016 65252 35020 65308
rect 35020 65252 35076 65308
rect 35076 65252 35080 65308
rect 35016 65248 35080 65252
rect 35096 65308 35160 65312
rect 35096 65252 35100 65308
rect 35100 65252 35156 65308
rect 35156 65252 35160 65308
rect 35096 65248 35160 65252
rect 35176 65308 35240 65312
rect 35176 65252 35180 65308
rect 35180 65252 35236 65308
rect 35236 65252 35240 65308
rect 35176 65248 35240 65252
rect 19576 64764 19640 64768
rect 19576 64708 19580 64764
rect 19580 64708 19636 64764
rect 19636 64708 19640 64764
rect 19576 64704 19640 64708
rect 19656 64764 19720 64768
rect 19656 64708 19660 64764
rect 19660 64708 19716 64764
rect 19716 64708 19720 64764
rect 19656 64704 19720 64708
rect 19736 64764 19800 64768
rect 19736 64708 19740 64764
rect 19740 64708 19796 64764
rect 19796 64708 19800 64764
rect 19736 64704 19800 64708
rect 19816 64764 19880 64768
rect 19816 64708 19820 64764
rect 19820 64708 19876 64764
rect 19876 64708 19880 64764
rect 19816 64704 19880 64708
rect 4216 64220 4280 64224
rect 4216 64164 4220 64220
rect 4220 64164 4276 64220
rect 4276 64164 4280 64220
rect 4216 64160 4280 64164
rect 4296 64220 4360 64224
rect 4296 64164 4300 64220
rect 4300 64164 4356 64220
rect 4356 64164 4360 64220
rect 4296 64160 4360 64164
rect 4376 64220 4440 64224
rect 4376 64164 4380 64220
rect 4380 64164 4436 64220
rect 4436 64164 4440 64220
rect 4376 64160 4440 64164
rect 4456 64220 4520 64224
rect 4456 64164 4460 64220
rect 4460 64164 4516 64220
rect 4516 64164 4520 64220
rect 4456 64160 4520 64164
rect 34936 64220 35000 64224
rect 34936 64164 34940 64220
rect 34940 64164 34996 64220
rect 34996 64164 35000 64220
rect 34936 64160 35000 64164
rect 35016 64220 35080 64224
rect 35016 64164 35020 64220
rect 35020 64164 35076 64220
rect 35076 64164 35080 64220
rect 35016 64160 35080 64164
rect 35096 64220 35160 64224
rect 35096 64164 35100 64220
rect 35100 64164 35156 64220
rect 35156 64164 35160 64220
rect 35096 64160 35160 64164
rect 35176 64220 35240 64224
rect 35176 64164 35180 64220
rect 35180 64164 35236 64220
rect 35236 64164 35240 64220
rect 35176 64160 35240 64164
rect 19576 63676 19640 63680
rect 19576 63620 19580 63676
rect 19580 63620 19636 63676
rect 19636 63620 19640 63676
rect 19576 63616 19640 63620
rect 19656 63676 19720 63680
rect 19656 63620 19660 63676
rect 19660 63620 19716 63676
rect 19716 63620 19720 63676
rect 19656 63616 19720 63620
rect 19736 63676 19800 63680
rect 19736 63620 19740 63676
rect 19740 63620 19796 63676
rect 19796 63620 19800 63676
rect 19736 63616 19800 63620
rect 19816 63676 19880 63680
rect 19816 63620 19820 63676
rect 19820 63620 19876 63676
rect 19876 63620 19880 63676
rect 19816 63616 19880 63620
rect 4216 63132 4280 63136
rect 4216 63076 4220 63132
rect 4220 63076 4276 63132
rect 4276 63076 4280 63132
rect 4216 63072 4280 63076
rect 4296 63132 4360 63136
rect 4296 63076 4300 63132
rect 4300 63076 4356 63132
rect 4356 63076 4360 63132
rect 4296 63072 4360 63076
rect 4376 63132 4440 63136
rect 4376 63076 4380 63132
rect 4380 63076 4436 63132
rect 4436 63076 4440 63132
rect 4376 63072 4440 63076
rect 4456 63132 4520 63136
rect 4456 63076 4460 63132
rect 4460 63076 4516 63132
rect 4516 63076 4520 63132
rect 4456 63072 4520 63076
rect 34936 63132 35000 63136
rect 34936 63076 34940 63132
rect 34940 63076 34996 63132
rect 34996 63076 35000 63132
rect 34936 63072 35000 63076
rect 35016 63132 35080 63136
rect 35016 63076 35020 63132
rect 35020 63076 35076 63132
rect 35076 63076 35080 63132
rect 35016 63072 35080 63076
rect 35096 63132 35160 63136
rect 35096 63076 35100 63132
rect 35100 63076 35156 63132
rect 35156 63076 35160 63132
rect 35096 63072 35160 63076
rect 35176 63132 35240 63136
rect 35176 63076 35180 63132
rect 35180 63076 35236 63132
rect 35236 63076 35240 63132
rect 35176 63072 35240 63076
rect 19576 62588 19640 62592
rect 19576 62532 19580 62588
rect 19580 62532 19636 62588
rect 19636 62532 19640 62588
rect 19576 62528 19640 62532
rect 19656 62588 19720 62592
rect 19656 62532 19660 62588
rect 19660 62532 19716 62588
rect 19716 62532 19720 62588
rect 19656 62528 19720 62532
rect 19736 62588 19800 62592
rect 19736 62532 19740 62588
rect 19740 62532 19796 62588
rect 19796 62532 19800 62588
rect 19736 62528 19800 62532
rect 19816 62588 19880 62592
rect 19816 62532 19820 62588
rect 19820 62532 19876 62588
rect 19876 62532 19880 62588
rect 19816 62528 19880 62532
rect 4216 62044 4280 62048
rect 4216 61988 4220 62044
rect 4220 61988 4276 62044
rect 4276 61988 4280 62044
rect 4216 61984 4280 61988
rect 4296 62044 4360 62048
rect 4296 61988 4300 62044
rect 4300 61988 4356 62044
rect 4356 61988 4360 62044
rect 4296 61984 4360 61988
rect 4376 62044 4440 62048
rect 4376 61988 4380 62044
rect 4380 61988 4436 62044
rect 4436 61988 4440 62044
rect 4376 61984 4440 61988
rect 4456 62044 4520 62048
rect 4456 61988 4460 62044
rect 4460 61988 4516 62044
rect 4516 61988 4520 62044
rect 4456 61984 4520 61988
rect 34936 62044 35000 62048
rect 34936 61988 34940 62044
rect 34940 61988 34996 62044
rect 34996 61988 35000 62044
rect 34936 61984 35000 61988
rect 35016 62044 35080 62048
rect 35016 61988 35020 62044
rect 35020 61988 35076 62044
rect 35076 61988 35080 62044
rect 35016 61984 35080 61988
rect 35096 62044 35160 62048
rect 35096 61988 35100 62044
rect 35100 61988 35156 62044
rect 35156 61988 35160 62044
rect 35096 61984 35160 61988
rect 35176 62044 35240 62048
rect 35176 61988 35180 62044
rect 35180 61988 35236 62044
rect 35236 61988 35240 62044
rect 35176 61984 35240 61988
rect 19576 61500 19640 61504
rect 19576 61444 19580 61500
rect 19580 61444 19636 61500
rect 19636 61444 19640 61500
rect 19576 61440 19640 61444
rect 19656 61500 19720 61504
rect 19656 61444 19660 61500
rect 19660 61444 19716 61500
rect 19716 61444 19720 61500
rect 19656 61440 19720 61444
rect 19736 61500 19800 61504
rect 19736 61444 19740 61500
rect 19740 61444 19796 61500
rect 19796 61444 19800 61500
rect 19736 61440 19800 61444
rect 19816 61500 19880 61504
rect 19816 61444 19820 61500
rect 19820 61444 19876 61500
rect 19876 61444 19880 61500
rect 19816 61440 19880 61444
rect 4216 60956 4280 60960
rect 4216 60900 4220 60956
rect 4220 60900 4276 60956
rect 4276 60900 4280 60956
rect 4216 60896 4280 60900
rect 4296 60956 4360 60960
rect 4296 60900 4300 60956
rect 4300 60900 4356 60956
rect 4356 60900 4360 60956
rect 4296 60896 4360 60900
rect 4376 60956 4440 60960
rect 4376 60900 4380 60956
rect 4380 60900 4436 60956
rect 4436 60900 4440 60956
rect 4376 60896 4440 60900
rect 4456 60956 4520 60960
rect 4456 60900 4460 60956
rect 4460 60900 4516 60956
rect 4516 60900 4520 60956
rect 4456 60896 4520 60900
rect 34936 60956 35000 60960
rect 34936 60900 34940 60956
rect 34940 60900 34996 60956
rect 34996 60900 35000 60956
rect 34936 60896 35000 60900
rect 35016 60956 35080 60960
rect 35016 60900 35020 60956
rect 35020 60900 35076 60956
rect 35076 60900 35080 60956
rect 35016 60896 35080 60900
rect 35096 60956 35160 60960
rect 35096 60900 35100 60956
rect 35100 60900 35156 60956
rect 35156 60900 35160 60956
rect 35096 60896 35160 60900
rect 35176 60956 35240 60960
rect 35176 60900 35180 60956
rect 35180 60900 35236 60956
rect 35236 60900 35240 60956
rect 35176 60896 35240 60900
rect 19576 60412 19640 60416
rect 19576 60356 19580 60412
rect 19580 60356 19636 60412
rect 19636 60356 19640 60412
rect 19576 60352 19640 60356
rect 19656 60412 19720 60416
rect 19656 60356 19660 60412
rect 19660 60356 19716 60412
rect 19716 60356 19720 60412
rect 19656 60352 19720 60356
rect 19736 60412 19800 60416
rect 19736 60356 19740 60412
rect 19740 60356 19796 60412
rect 19796 60356 19800 60412
rect 19736 60352 19800 60356
rect 19816 60412 19880 60416
rect 19816 60356 19820 60412
rect 19820 60356 19876 60412
rect 19876 60356 19880 60412
rect 19816 60352 19880 60356
rect 4216 59868 4280 59872
rect 4216 59812 4220 59868
rect 4220 59812 4276 59868
rect 4276 59812 4280 59868
rect 4216 59808 4280 59812
rect 4296 59868 4360 59872
rect 4296 59812 4300 59868
rect 4300 59812 4356 59868
rect 4356 59812 4360 59868
rect 4296 59808 4360 59812
rect 4376 59868 4440 59872
rect 4376 59812 4380 59868
rect 4380 59812 4436 59868
rect 4436 59812 4440 59868
rect 4376 59808 4440 59812
rect 4456 59868 4520 59872
rect 4456 59812 4460 59868
rect 4460 59812 4516 59868
rect 4516 59812 4520 59868
rect 4456 59808 4520 59812
rect 34936 59868 35000 59872
rect 34936 59812 34940 59868
rect 34940 59812 34996 59868
rect 34996 59812 35000 59868
rect 34936 59808 35000 59812
rect 35016 59868 35080 59872
rect 35016 59812 35020 59868
rect 35020 59812 35076 59868
rect 35076 59812 35080 59868
rect 35016 59808 35080 59812
rect 35096 59868 35160 59872
rect 35096 59812 35100 59868
rect 35100 59812 35156 59868
rect 35156 59812 35160 59868
rect 35096 59808 35160 59812
rect 35176 59868 35240 59872
rect 35176 59812 35180 59868
rect 35180 59812 35236 59868
rect 35236 59812 35240 59868
rect 35176 59808 35240 59812
rect 19576 59324 19640 59328
rect 19576 59268 19580 59324
rect 19580 59268 19636 59324
rect 19636 59268 19640 59324
rect 19576 59264 19640 59268
rect 19656 59324 19720 59328
rect 19656 59268 19660 59324
rect 19660 59268 19716 59324
rect 19716 59268 19720 59324
rect 19656 59264 19720 59268
rect 19736 59324 19800 59328
rect 19736 59268 19740 59324
rect 19740 59268 19796 59324
rect 19796 59268 19800 59324
rect 19736 59264 19800 59268
rect 19816 59324 19880 59328
rect 19816 59268 19820 59324
rect 19820 59268 19876 59324
rect 19876 59268 19880 59324
rect 19816 59264 19880 59268
rect 4216 58780 4280 58784
rect 4216 58724 4220 58780
rect 4220 58724 4276 58780
rect 4276 58724 4280 58780
rect 4216 58720 4280 58724
rect 4296 58780 4360 58784
rect 4296 58724 4300 58780
rect 4300 58724 4356 58780
rect 4356 58724 4360 58780
rect 4296 58720 4360 58724
rect 4376 58780 4440 58784
rect 4376 58724 4380 58780
rect 4380 58724 4436 58780
rect 4436 58724 4440 58780
rect 4376 58720 4440 58724
rect 4456 58780 4520 58784
rect 4456 58724 4460 58780
rect 4460 58724 4516 58780
rect 4516 58724 4520 58780
rect 4456 58720 4520 58724
rect 34936 58780 35000 58784
rect 34936 58724 34940 58780
rect 34940 58724 34996 58780
rect 34996 58724 35000 58780
rect 34936 58720 35000 58724
rect 35016 58780 35080 58784
rect 35016 58724 35020 58780
rect 35020 58724 35076 58780
rect 35076 58724 35080 58780
rect 35016 58720 35080 58724
rect 35096 58780 35160 58784
rect 35096 58724 35100 58780
rect 35100 58724 35156 58780
rect 35156 58724 35160 58780
rect 35096 58720 35160 58724
rect 35176 58780 35240 58784
rect 35176 58724 35180 58780
rect 35180 58724 35236 58780
rect 35236 58724 35240 58780
rect 35176 58720 35240 58724
rect 19576 58236 19640 58240
rect 19576 58180 19580 58236
rect 19580 58180 19636 58236
rect 19636 58180 19640 58236
rect 19576 58176 19640 58180
rect 19656 58236 19720 58240
rect 19656 58180 19660 58236
rect 19660 58180 19716 58236
rect 19716 58180 19720 58236
rect 19656 58176 19720 58180
rect 19736 58236 19800 58240
rect 19736 58180 19740 58236
rect 19740 58180 19796 58236
rect 19796 58180 19800 58236
rect 19736 58176 19800 58180
rect 19816 58236 19880 58240
rect 19816 58180 19820 58236
rect 19820 58180 19876 58236
rect 19876 58180 19880 58236
rect 19816 58176 19880 58180
rect 4216 57692 4280 57696
rect 4216 57636 4220 57692
rect 4220 57636 4276 57692
rect 4276 57636 4280 57692
rect 4216 57632 4280 57636
rect 4296 57692 4360 57696
rect 4296 57636 4300 57692
rect 4300 57636 4356 57692
rect 4356 57636 4360 57692
rect 4296 57632 4360 57636
rect 4376 57692 4440 57696
rect 4376 57636 4380 57692
rect 4380 57636 4436 57692
rect 4436 57636 4440 57692
rect 4376 57632 4440 57636
rect 4456 57692 4520 57696
rect 4456 57636 4460 57692
rect 4460 57636 4516 57692
rect 4516 57636 4520 57692
rect 4456 57632 4520 57636
rect 34936 57692 35000 57696
rect 34936 57636 34940 57692
rect 34940 57636 34996 57692
rect 34996 57636 35000 57692
rect 34936 57632 35000 57636
rect 35016 57692 35080 57696
rect 35016 57636 35020 57692
rect 35020 57636 35076 57692
rect 35076 57636 35080 57692
rect 35016 57632 35080 57636
rect 35096 57692 35160 57696
rect 35096 57636 35100 57692
rect 35100 57636 35156 57692
rect 35156 57636 35160 57692
rect 35096 57632 35160 57636
rect 35176 57692 35240 57696
rect 35176 57636 35180 57692
rect 35180 57636 35236 57692
rect 35236 57636 35240 57692
rect 35176 57632 35240 57636
rect 19576 57148 19640 57152
rect 19576 57092 19580 57148
rect 19580 57092 19636 57148
rect 19636 57092 19640 57148
rect 19576 57088 19640 57092
rect 19656 57148 19720 57152
rect 19656 57092 19660 57148
rect 19660 57092 19716 57148
rect 19716 57092 19720 57148
rect 19656 57088 19720 57092
rect 19736 57148 19800 57152
rect 19736 57092 19740 57148
rect 19740 57092 19796 57148
rect 19796 57092 19800 57148
rect 19736 57088 19800 57092
rect 19816 57148 19880 57152
rect 19816 57092 19820 57148
rect 19820 57092 19876 57148
rect 19876 57092 19880 57148
rect 19816 57088 19880 57092
rect 4216 56604 4280 56608
rect 4216 56548 4220 56604
rect 4220 56548 4276 56604
rect 4276 56548 4280 56604
rect 4216 56544 4280 56548
rect 4296 56604 4360 56608
rect 4296 56548 4300 56604
rect 4300 56548 4356 56604
rect 4356 56548 4360 56604
rect 4296 56544 4360 56548
rect 4376 56604 4440 56608
rect 4376 56548 4380 56604
rect 4380 56548 4436 56604
rect 4436 56548 4440 56604
rect 4376 56544 4440 56548
rect 4456 56604 4520 56608
rect 4456 56548 4460 56604
rect 4460 56548 4516 56604
rect 4516 56548 4520 56604
rect 4456 56544 4520 56548
rect 34936 56604 35000 56608
rect 34936 56548 34940 56604
rect 34940 56548 34996 56604
rect 34996 56548 35000 56604
rect 34936 56544 35000 56548
rect 35016 56604 35080 56608
rect 35016 56548 35020 56604
rect 35020 56548 35076 56604
rect 35076 56548 35080 56604
rect 35016 56544 35080 56548
rect 35096 56604 35160 56608
rect 35096 56548 35100 56604
rect 35100 56548 35156 56604
rect 35156 56548 35160 56604
rect 35096 56544 35160 56548
rect 35176 56604 35240 56608
rect 35176 56548 35180 56604
rect 35180 56548 35236 56604
rect 35236 56548 35240 56604
rect 35176 56544 35240 56548
rect 19576 56060 19640 56064
rect 19576 56004 19580 56060
rect 19580 56004 19636 56060
rect 19636 56004 19640 56060
rect 19576 56000 19640 56004
rect 19656 56060 19720 56064
rect 19656 56004 19660 56060
rect 19660 56004 19716 56060
rect 19716 56004 19720 56060
rect 19656 56000 19720 56004
rect 19736 56060 19800 56064
rect 19736 56004 19740 56060
rect 19740 56004 19796 56060
rect 19796 56004 19800 56060
rect 19736 56000 19800 56004
rect 19816 56060 19880 56064
rect 19816 56004 19820 56060
rect 19820 56004 19876 56060
rect 19876 56004 19880 56060
rect 19816 56000 19880 56004
rect 4216 55516 4280 55520
rect 4216 55460 4220 55516
rect 4220 55460 4276 55516
rect 4276 55460 4280 55516
rect 4216 55456 4280 55460
rect 4296 55516 4360 55520
rect 4296 55460 4300 55516
rect 4300 55460 4356 55516
rect 4356 55460 4360 55516
rect 4296 55456 4360 55460
rect 4376 55516 4440 55520
rect 4376 55460 4380 55516
rect 4380 55460 4436 55516
rect 4436 55460 4440 55516
rect 4376 55456 4440 55460
rect 4456 55516 4520 55520
rect 4456 55460 4460 55516
rect 4460 55460 4516 55516
rect 4516 55460 4520 55516
rect 4456 55456 4520 55460
rect 34936 55516 35000 55520
rect 34936 55460 34940 55516
rect 34940 55460 34996 55516
rect 34996 55460 35000 55516
rect 34936 55456 35000 55460
rect 35016 55516 35080 55520
rect 35016 55460 35020 55516
rect 35020 55460 35076 55516
rect 35076 55460 35080 55516
rect 35016 55456 35080 55460
rect 35096 55516 35160 55520
rect 35096 55460 35100 55516
rect 35100 55460 35156 55516
rect 35156 55460 35160 55516
rect 35096 55456 35160 55460
rect 35176 55516 35240 55520
rect 35176 55460 35180 55516
rect 35180 55460 35236 55516
rect 35236 55460 35240 55516
rect 35176 55456 35240 55460
rect 19576 54972 19640 54976
rect 19576 54916 19580 54972
rect 19580 54916 19636 54972
rect 19636 54916 19640 54972
rect 19576 54912 19640 54916
rect 19656 54972 19720 54976
rect 19656 54916 19660 54972
rect 19660 54916 19716 54972
rect 19716 54916 19720 54972
rect 19656 54912 19720 54916
rect 19736 54972 19800 54976
rect 19736 54916 19740 54972
rect 19740 54916 19796 54972
rect 19796 54916 19800 54972
rect 19736 54912 19800 54916
rect 19816 54972 19880 54976
rect 19816 54916 19820 54972
rect 19820 54916 19876 54972
rect 19876 54916 19880 54972
rect 19816 54912 19880 54916
rect 4216 54428 4280 54432
rect 4216 54372 4220 54428
rect 4220 54372 4276 54428
rect 4276 54372 4280 54428
rect 4216 54368 4280 54372
rect 4296 54428 4360 54432
rect 4296 54372 4300 54428
rect 4300 54372 4356 54428
rect 4356 54372 4360 54428
rect 4296 54368 4360 54372
rect 4376 54428 4440 54432
rect 4376 54372 4380 54428
rect 4380 54372 4436 54428
rect 4436 54372 4440 54428
rect 4376 54368 4440 54372
rect 4456 54428 4520 54432
rect 4456 54372 4460 54428
rect 4460 54372 4516 54428
rect 4516 54372 4520 54428
rect 4456 54368 4520 54372
rect 34936 54428 35000 54432
rect 34936 54372 34940 54428
rect 34940 54372 34996 54428
rect 34996 54372 35000 54428
rect 34936 54368 35000 54372
rect 35016 54428 35080 54432
rect 35016 54372 35020 54428
rect 35020 54372 35076 54428
rect 35076 54372 35080 54428
rect 35016 54368 35080 54372
rect 35096 54428 35160 54432
rect 35096 54372 35100 54428
rect 35100 54372 35156 54428
rect 35156 54372 35160 54428
rect 35096 54368 35160 54372
rect 35176 54428 35240 54432
rect 35176 54372 35180 54428
rect 35180 54372 35236 54428
rect 35236 54372 35240 54428
rect 35176 54368 35240 54372
rect 19576 53884 19640 53888
rect 19576 53828 19580 53884
rect 19580 53828 19636 53884
rect 19636 53828 19640 53884
rect 19576 53824 19640 53828
rect 19656 53884 19720 53888
rect 19656 53828 19660 53884
rect 19660 53828 19716 53884
rect 19716 53828 19720 53884
rect 19656 53824 19720 53828
rect 19736 53884 19800 53888
rect 19736 53828 19740 53884
rect 19740 53828 19796 53884
rect 19796 53828 19800 53884
rect 19736 53824 19800 53828
rect 19816 53884 19880 53888
rect 19816 53828 19820 53884
rect 19820 53828 19876 53884
rect 19876 53828 19880 53884
rect 19816 53824 19880 53828
rect 4216 53340 4280 53344
rect 4216 53284 4220 53340
rect 4220 53284 4276 53340
rect 4276 53284 4280 53340
rect 4216 53280 4280 53284
rect 4296 53340 4360 53344
rect 4296 53284 4300 53340
rect 4300 53284 4356 53340
rect 4356 53284 4360 53340
rect 4296 53280 4360 53284
rect 4376 53340 4440 53344
rect 4376 53284 4380 53340
rect 4380 53284 4436 53340
rect 4436 53284 4440 53340
rect 4376 53280 4440 53284
rect 4456 53340 4520 53344
rect 4456 53284 4460 53340
rect 4460 53284 4516 53340
rect 4516 53284 4520 53340
rect 4456 53280 4520 53284
rect 34936 53340 35000 53344
rect 34936 53284 34940 53340
rect 34940 53284 34996 53340
rect 34996 53284 35000 53340
rect 34936 53280 35000 53284
rect 35016 53340 35080 53344
rect 35016 53284 35020 53340
rect 35020 53284 35076 53340
rect 35076 53284 35080 53340
rect 35016 53280 35080 53284
rect 35096 53340 35160 53344
rect 35096 53284 35100 53340
rect 35100 53284 35156 53340
rect 35156 53284 35160 53340
rect 35096 53280 35160 53284
rect 35176 53340 35240 53344
rect 35176 53284 35180 53340
rect 35180 53284 35236 53340
rect 35236 53284 35240 53340
rect 35176 53280 35240 53284
rect 19576 52796 19640 52800
rect 19576 52740 19580 52796
rect 19580 52740 19636 52796
rect 19636 52740 19640 52796
rect 19576 52736 19640 52740
rect 19656 52796 19720 52800
rect 19656 52740 19660 52796
rect 19660 52740 19716 52796
rect 19716 52740 19720 52796
rect 19656 52736 19720 52740
rect 19736 52796 19800 52800
rect 19736 52740 19740 52796
rect 19740 52740 19796 52796
rect 19796 52740 19800 52796
rect 19736 52736 19800 52740
rect 19816 52796 19880 52800
rect 19816 52740 19820 52796
rect 19820 52740 19876 52796
rect 19876 52740 19880 52796
rect 19816 52736 19880 52740
rect 4216 52252 4280 52256
rect 4216 52196 4220 52252
rect 4220 52196 4276 52252
rect 4276 52196 4280 52252
rect 4216 52192 4280 52196
rect 4296 52252 4360 52256
rect 4296 52196 4300 52252
rect 4300 52196 4356 52252
rect 4356 52196 4360 52252
rect 4296 52192 4360 52196
rect 4376 52252 4440 52256
rect 4376 52196 4380 52252
rect 4380 52196 4436 52252
rect 4436 52196 4440 52252
rect 4376 52192 4440 52196
rect 4456 52252 4520 52256
rect 4456 52196 4460 52252
rect 4460 52196 4516 52252
rect 4516 52196 4520 52252
rect 4456 52192 4520 52196
rect 34936 52252 35000 52256
rect 34936 52196 34940 52252
rect 34940 52196 34996 52252
rect 34996 52196 35000 52252
rect 34936 52192 35000 52196
rect 35016 52252 35080 52256
rect 35016 52196 35020 52252
rect 35020 52196 35076 52252
rect 35076 52196 35080 52252
rect 35016 52192 35080 52196
rect 35096 52252 35160 52256
rect 35096 52196 35100 52252
rect 35100 52196 35156 52252
rect 35156 52196 35160 52252
rect 35096 52192 35160 52196
rect 35176 52252 35240 52256
rect 35176 52196 35180 52252
rect 35180 52196 35236 52252
rect 35236 52196 35240 52252
rect 35176 52192 35240 52196
rect 19576 51708 19640 51712
rect 19576 51652 19580 51708
rect 19580 51652 19636 51708
rect 19636 51652 19640 51708
rect 19576 51648 19640 51652
rect 19656 51708 19720 51712
rect 19656 51652 19660 51708
rect 19660 51652 19716 51708
rect 19716 51652 19720 51708
rect 19656 51648 19720 51652
rect 19736 51708 19800 51712
rect 19736 51652 19740 51708
rect 19740 51652 19796 51708
rect 19796 51652 19800 51708
rect 19736 51648 19800 51652
rect 19816 51708 19880 51712
rect 19816 51652 19820 51708
rect 19820 51652 19876 51708
rect 19876 51652 19880 51708
rect 19816 51648 19880 51652
rect 4216 51164 4280 51168
rect 4216 51108 4220 51164
rect 4220 51108 4276 51164
rect 4276 51108 4280 51164
rect 4216 51104 4280 51108
rect 4296 51164 4360 51168
rect 4296 51108 4300 51164
rect 4300 51108 4356 51164
rect 4356 51108 4360 51164
rect 4296 51104 4360 51108
rect 4376 51164 4440 51168
rect 4376 51108 4380 51164
rect 4380 51108 4436 51164
rect 4436 51108 4440 51164
rect 4376 51104 4440 51108
rect 4456 51164 4520 51168
rect 4456 51108 4460 51164
rect 4460 51108 4516 51164
rect 4516 51108 4520 51164
rect 4456 51104 4520 51108
rect 34936 51164 35000 51168
rect 34936 51108 34940 51164
rect 34940 51108 34996 51164
rect 34996 51108 35000 51164
rect 34936 51104 35000 51108
rect 35016 51164 35080 51168
rect 35016 51108 35020 51164
rect 35020 51108 35076 51164
rect 35076 51108 35080 51164
rect 35016 51104 35080 51108
rect 35096 51164 35160 51168
rect 35096 51108 35100 51164
rect 35100 51108 35156 51164
rect 35156 51108 35160 51164
rect 35096 51104 35160 51108
rect 35176 51164 35240 51168
rect 35176 51108 35180 51164
rect 35180 51108 35236 51164
rect 35236 51108 35240 51164
rect 35176 51104 35240 51108
rect 19576 50620 19640 50624
rect 19576 50564 19580 50620
rect 19580 50564 19636 50620
rect 19636 50564 19640 50620
rect 19576 50560 19640 50564
rect 19656 50620 19720 50624
rect 19656 50564 19660 50620
rect 19660 50564 19716 50620
rect 19716 50564 19720 50620
rect 19656 50560 19720 50564
rect 19736 50620 19800 50624
rect 19736 50564 19740 50620
rect 19740 50564 19796 50620
rect 19796 50564 19800 50620
rect 19736 50560 19800 50564
rect 19816 50620 19880 50624
rect 19816 50564 19820 50620
rect 19820 50564 19876 50620
rect 19876 50564 19880 50620
rect 19816 50560 19880 50564
rect 4216 50076 4280 50080
rect 4216 50020 4220 50076
rect 4220 50020 4276 50076
rect 4276 50020 4280 50076
rect 4216 50016 4280 50020
rect 4296 50076 4360 50080
rect 4296 50020 4300 50076
rect 4300 50020 4356 50076
rect 4356 50020 4360 50076
rect 4296 50016 4360 50020
rect 4376 50076 4440 50080
rect 4376 50020 4380 50076
rect 4380 50020 4436 50076
rect 4436 50020 4440 50076
rect 4376 50016 4440 50020
rect 4456 50076 4520 50080
rect 4456 50020 4460 50076
rect 4460 50020 4516 50076
rect 4516 50020 4520 50076
rect 4456 50016 4520 50020
rect 34936 50076 35000 50080
rect 34936 50020 34940 50076
rect 34940 50020 34996 50076
rect 34996 50020 35000 50076
rect 34936 50016 35000 50020
rect 35016 50076 35080 50080
rect 35016 50020 35020 50076
rect 35020 50020 35076 50076
rect 35076 50020 35080 50076
rect 35016 50016 35080 50020
rect 35096 50076 35160 50080
rect 35096 50020 35100 50076
rect 35100 50020 35156 50076
rect 35156 50020 35160 50076
rect 35096 50016 35160 50020
rect 35176 50076 35240 50080
rect 35176 50020 35180 50076
rect 35180 50020 35236 50076
rect 35236 50020 35240 50076
rect 35176 50016 35240 50020
rect 19576 49532 19640 49536
rect 19576 49476 19580 49532
rect 19580 49476 19636 49532
rect 19636 49476 19640 49532
rect 19576 49472 19640 49476
rect 19656 49532 19720 49536
rect 19656 49476 19660 49532
rect 19660 49476 19716 49532
rect 19716 49476 19720 49532
rect 19656 49472 19720 49476
rect 19736 49532 19800 49536
rect 19736 49476 19740 49532
rect 19740 49476 19796 49532
rect 19796 49476 19800 49532
rect 19736 49472 19800 49476
rect 19816 49532 19880 49536
rect 19816 49476 19820 49532
rect 19820 49476 19876 49532
rect 19876 49476 19880 49532
rect 19816 49472 19880 49476
rect 4216 48988 4280 48992
rect 4216 48932 4220 48988
rect 4220 48932 4276 48988
rect 4276 48932 4280 48988
rect 4216 48928 4280 48932
rect 4296 48988 4360 48992
rect 4296 48932 4300 48988
rect 4300 48932 4356 48988
rect 4356 48932 4360 48988
rect 4296 48928 4360 48932
rect 4376 48988 4440 48992
rect 4376 48932 4380 48988
rect 4380 48932 4436 48988
rect 4436 48932 4440 48988
rect 4376 48928 4440 48932
rect 4456 48988 4520 48992
rect 4456 48932 4460 48988
rect 4460 48932 4516 48988
rect 4516 48932 4520 48988
rect 4456 48928 4520 48932
rect 34936 48988 35000 48992
rect 34936 48932 34940 48988
rect 34940 48932 34996 48988
rect 34996 48932 35000 48988
rect 34936 48928 35000 48932
rect 35016 48988 35080 48992
rect 35016 48932 35020 48988
rect 35020 48932 35076 48988
rect 35076 48932 35080 48988
rect 35016 48928 35080 48932
rect 35096 48988 35160 48992
rect 35096 48932 35100 48988
rect 35100 48932 35156 48988
rect 35156 48932 35160 48988
rect 35096 48928 35160 48932
rect 35176 48988 35240 48992
rect 35176 48932 35180 48988
rect 35180 48932 35236 48988
rect 35236 48932 35240 48988
rect 35176 48928 35240 48932
rect 19576 48444 19640 48448
rect 19576 48388 19580 48444
rect 19580 48388 19636 48444
rect 19636 48388 19640 48444
rect 19576 48384 19640 48388
rect 19656 48444 19720 48448
rect 19656 48388 19660 48444
rect 19660 48388 19716 48444
rect 19716 48388 19720 48444
rect 19656 48384 19720 48388
rect 19736 48444 19800 48448
rect 19736 48388 19740 48444
rect 19740 48388 19796 48444
rect 19796 48388 19800 48444
rect 19736 48384 19800 48388
rect 19816 48444 19880 48448
rect 19816 48388 19820 48444
rect 19820 48388 19876 48444
rect 19876 48388 19880 48444
rect 19816 48384 19880 48388
rect 4216 47900 4280 47904
rect 4216 47844 4220 47900
rect 4220 47844 4276 47900
rect 4276 47844 4280 47900
rect 4216 47840 4280 47844
rect 4296 47900 4360 47904
rect 4296 47844 4300 47900
rect 4300 47844 4356 47900
rect 4356 47844 4360 47900
rect 4296 47840 4360 47844
rect 4376 47900 4440 47904
rect 4376 47844 4380 47900
rect 4380 47844 4436 47900
rect 4436 47844 4440 47900
rect 4376 47840 4440 47844
rect 4456 47900 4520 47904
rect 4456 47844 4460 47900
rect 4460 47844 4516 47900
rect 4516 47844 4520 47900
rect 4456 47840 4520 47844
rect 34936 47900 35000 47904
rect 34936 47844 34940 47900
rect 34940 47844 34996 47900
rect 34996 47844 35000 47900
rect 34936 47840 35000 47844
rect 35016 47900 35080 47904
rect 35016 47844 35020 47900
rect 35020 47844 35076 47900
rect 35076 47844 35080 47900
rect 35016 47840 35080 47844
rect 35096 47900 35160 47904
rect 35096 47844 35100 47900
rect 35100 47844 35156 47900
rect 35156 47844 35160 47900
rect 35096 47840 35160 47844
rect 35176 47900 35240 47904
rect 35176 47844 35180 47900
rect 35180 47844 35236 47900
rect 35236 47844 35240 47900
rect 35176 47840 35240 47844
rect 19576 47356 19640 47360
rect 19576 47300 19580 47356
rect 19580 47300 19636 47356
rect 19636 47300 19640 47356
rect 19576 47296 19640 47300
rect 19656 47356 19720 47360
rect 19656 47300 19660 47356
rect 19660 47300 19716 47356
rect 19716 47300 19720 47356
rect 19656 47296 19720 47300
rect 19736 47356 19800 47360
rect 19736 47300 19740 47356
rect 19740 47300 19796 47356
rect 19796 47300 19800 47356
rect 19736 47296 19800 47300
rect 19816 47356 19880 47360
rect 19816 47300 19820 47356
rect 19820 47300 19876 47356
rect 19876 47300 19880 47356
rect 19816 47296 19880 47300
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 34936 46812 35000 46816
rect 34936 46756 34940 46812
rect 34940 46756 34996 46812
rect 34996 46756 35000 46812
rect 34936 46752 35000 46756
rect 35016 46812 35080 46816
rect 35016 46756 35020 46812
rect 35020 46756 35076 46812
rect 35076 46756 35080 46812
rect 35016 46752 35080 46756
rect 35096 46812 35160 46816
rect 35096 46756 35100 46812
rect 35100 46756 35156 46812
rect 35156 46756 35160 46812
rect 35096 46752 35160 46756
rect 35176 46812 35240 46816
rect 35176 46756 35180 46812
rect 35180 46756 35236 46812
rect 35236 46756 35240 46812
rect 35176 46752 35240 46756
rect 19576 46268 19640 46272
rect 19576 46212 19580 46268
rect 19580 46212 19636 46268
rect 19636 46212 19640 46268
rect 19576 46208 19640 46212
rect 19656 46268 19720 46272
rect 19656 46212 19660 46268
rect 19660 46212 19716 46268
rect 19716 46212 19720 46268
rect 19656 46208 19720 46212
rect 19736 46268 19800 46272
rect 19736 46212 19740 46268
rect 19740 46212 19796 46268
rect 19796 46212 19800 46268
rect 19736 46208 19800 46212
rect 19816 46268 19880 46272
rect 19816 46212 19820 46268
rect 19820 46212 19876 46268
rect 19876 46212 19880 46268
rect 19816 46208 19880 46212
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 34936 45724 35000 45728
rect 34936 45668 34940 45724
rect 34940 45668 34996 45724
rect 34996 45668 35000 45724
rect 34936 45664 35000 45668
rect 35016 45724 35080 45728
rect 35016 45668 35020 45724
rect 35020 45668 35076 45724
rect 35076 45668 35080 45724
rect 35016 45664 35080 45668
rect 35096 45724 35160 45728
rect 35096 45668 35100 45724
rect 35100 45668 35156 45724
rect 35156 45668 35160 45724
rect 35096 45664 35160 45668
rect 35176 45724 35240 45728
rect 35176 45668 35180 45724
rect 35180 45668 35236 45724
rect 35236 45668 35240 45724
rect 35176 45664 35240 45668
rect 19576 45180 19640 45184
rect 19576 45124 19580 45180
rect 19580 45124 19636 45180
rect 19636 45124 19640 45180
rect 19576 45120 19640 45124
rect 19656 45180 19720 45184
rect 19656 45124 19660 45180
rect 19660 45124 19716 45180
rect 19716 45124 19720 45180
rect 19656 45120 19720 45124
rect 19736 45180 19800 45184
rect 19736 45124 19740 45180
rect 19740 45124 19796 45180
rect 19796 45124 19800 45180
rect 19736 45120 19800 45124
rect 19816 45180 19880 45184
rect 19816 45124 19820 45180
rect 19820 45124 19876 45180
rect 19876 45124 19880 45180
rect 19816 45120 19880 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 34936 44636 35000 44640
rect 34936 44580 34940 44636
rect 34940 44580 34996 44636
rect 34996 44580 35000 44636
rect 34936 44576 35000 44580
rect 35016 44636 35080 44640
rect 35016 44580 35020 44636
rect 35020 44580 35076 44636
rect 35076 44580 35080 44636
rect 35016 44576 35080 44580
rect 35096 44636 35160 44640
rect 35096 44580 35100 44636
rect 35100 44580 35156 44636
rect 35156 44580 35160 44636
rect 35096 44576 35160 44580
rect 35176 44636 35240 44640
rect 35176 44580 35180 44636
rect 35180 44580 35236 44636
rect 35236 44580 35240 44636
rect 35176 44576 35240 44580
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 117536 4528 117552
rect 4208 117472 4216 117536
rect 4280 117472 4296 117536
rect 4360 117472 4376 117536
rect 4440 117472 4456 117536
rect 4520 117472 4528 117536
rect 4208 116448 4528 117472
rect 4208 116384 4216 116448
rect 4280 116384 4296 116448
rect 4360 116384 4376 116448
rect 4440 116384 4456 116448
rect 4520 116384 4528 116448
rect 4208 115360 4528 116384
rect 4208 115296 4216 115360
rect 4280 115296 4296 115360
rect 4360 115296 4376 115360
rect 4440 115296 4456 115360
rect 4520 115296 4528 115360
rect 4208 114272 4528 115296
rect 4208 114208 4216 114272
rect 4280 114208 4296 114272
rect 4360 114208 4376 114272
rect 4440 114208 4456 114272
rect 4520 114208 4528 114272
rect 4208 113184 4528 114208
rect 4208 113120 4216 113184
rect 4280 113120 4296 113184
rect 4360 113120 4376 113184
rect 4440 113120 4456 113184
rect 4520 113120 4528 113184
rect 4208 112096 4528 113120
rect 4208 112032 4216 112096
rect 4280 112032 4296 112096
rect 4360 112032 4376 112096
rect 4440 112032 4456 112096
rect 4520 112032 4528 112096
rect 4208 111008 4528 112032
rect 4208 110944 4216 111008
rect 4280 110944 4296 111008
rect 4360 110944 4376 111008
rect 4440 110944 4456 111008
rect 4520 110944 4528 111008
rect 4208 109920 4528 110944
rect 4208 109856 4216 109920
rect 4280 109856 4296 109920
rect 4360 109856 4376 109920
rect 4440 109856 4456 109920
rect 4520 109856 4528 109920
rect 4208 108832 4528 109856
rect 4208 108768 4216 108832
rect 4280 108768 4296 108832
rect 4360 108768 4376 108832
rect 4440 108768 4456 108832
rect 4520 108768 4528 108832
rect 4208 107744 4528 108768
rect 4208 107680 4216 107744
rect 4280 107680 4296 107744
rect 4360 107680 4376 107744
rect 4440 107680 4456 107744
rect 4520 107680 4528 107744
rect 4208 106656 4528 107680
rect 4208 106592 4216 106656
rect 4280 106592 4296 106656
rect 4360 106592 4376 106656
rect 4440 106592 4456 106656
rect 4520 106592 4528 106656
rect 4208 105568 4528 106592
rect 4208 105504 4216 105568
rect 4280 105504 4296 105568
rect 4360 105504 4376 105568
rect 4440 105504 4456 105568
rect 4520 105504 4528 105568
rect 4208 104480 4528 105504
rect 4208 104416 4216 104480
rect 4280 104416 4296 104480
rect 4360 104416 4376 104480
rect 4440 104416 4456 104480
rect 4520 104416 4528 104480
rect 4208 103392 4528 104416
rect 4208 103328 4216 103392
rect 4280 103328 4296 103392
rect 4360 103328 4376 103392
rect 4440 103328 4456 103392
rect 4520 103328 4528 103392
rect 4208 102304 4528 103328
rect 4208 102240 4216 102304
rect 4280 102240 4296 102304
rect 4360 102240 4376 102304
rect 4440 102240 4456 102304
rect 4520 102240 4528 102304
rect 4208 101216 4528 102240
rect 4208 101152 4216 101216
rect 4280 101152 4296 101216
rect 4360 101152 4376 101216
rect 4440 101152 4456 101216
rect 4520 101152 4528 101216
rect 4208 100128 4528 101152
rect 4208 100064 4216 100128
rect 4280 100064 4296 100128
rect 4360 100064 4376 100128
rect 4440 100064 4456 100128
rect 4520 100064 4528 100128
rect 4208 99040 4528 100064
rect 4208 98976 4216 99040
rect 4280 98976 4296 99040
rect 4360 98976 4376 99040
rect 4440 98976 4456 99040
rect 4520 98976 4528 99040
rect 4208 97952 4528 98976
rect 4208 97888 4216 97952
rect 4280 97888 4296 97952
rect 4360 97888 4376 97952
rect 4440 97888 4456 97952
rect 4520 97888 4528 97952
rect 4208 96864 4528 97888
rect 4208 96800 4216 96864
rect 4280 96800 4296 96864
rect 4360 96800 4376 96864
rect 4440 96800 4456 96864
rect 4520 96800 4528 96864
rect 4208 95776 4528 96800
rect 4208 95712 4216 95776
rect 4280 95712 4296 95776
rect 4360 95712 4376 95776
rect 4440 95712 4456 95776
rect 4520 95712 4528 95776
rect 4208 94688 4528 95712
rect 4208 94624 4216 94688
rect 4280 94624 4296 94688
rect 4360 94624 4376 94688
rect 4440 94624 4456 94688
rect 4520 94624 4528 94688
rect 4208 93600 4528 94624
rect 4208 93536 4216 93600
rect 4280 93536 4296 93600
rect 4360 93536 4376 93600
rect 4440 93536 4456 93600
rect 4520 93536 4528 93600
rect 4208 92512 4528 93536
rect 4208 92448 4216 92512
rect 4280 92448 4296 92512
rect 4360 92448 4376 92512
rect 4440 92448 4456 92512
rect 4520 92448 4528 92512
rect 4208 91424 4528 92448
rect 4208 91360 4216 91424
rect 4280 91360 4296 91424
rect 4360 91360 4376 91424
rect 4440 91360 4456 91424
rect 4520 91360 4528 91424
rect 4208 90336 4528 91360
rect 4208 90272 4216 90336
rect 4280 90272 4296 90336
rect 4360 90272 4376 90336
rect 4440 90272 4456 90336
rect 4520 90272 4528 90336
rect 4208 89248 4528 90272
rect 4208 89184 4216 89248
rect 4280 89184 4296 89248
rect 4360 89184 4376 89248
rect 4440 89184 4456 89248
rect 4520 89184 4528 89248
rect 4208 88160 4528 89184
rect 4208 88096 4216 88160
rect 4280 88096 4296 88160
rect 4360 88096 4376 88160
rect 4440 88096 4456 88160
rect 4520 88096 4528 88160
rect 4208 87072 4528 88096
rect 4208 87008 4216 87072
rect 4280 87008 4296 87072
rect 4360 87008 4376 87072
rect 4440 87008 4456 87072
rect 4520 87008 4528 87072
rect 4208 85984 4528 87008
rect 4208 85920 4216 85984
rect 4280 85920 4296 85984
rect 4360 85920 4376 85984
rect 4440 85920 4456 85984
rect 4520 85920 4528 85984
rect 4208 84896 4528 85920
rect 4208 84832 4216 84896
rect 4280 84832 4296 84896
rect 4360 84832 4376 84896
rect 4440 84832 4456 84896
rect 4520 84832 4528 84896
rect 4208 83808 4528 84832
rect 4208 83744 4216 83808
rect 4280 83744 4296 83808
rect 4360 83744 4376 83808
rect 4440 83744 4456 83808
rect 4520 83744 4528 83808
rect 4208 82720 4528 83744
rect 4208 82656 4216 82720
rect 4280 82656 4296 82720
rect 4360 82656 4376 82720
rect 4440 82656 4456 82720
rect 4520 82656 4528 82720
rect 4208 81632 4528 82656
rect 4208 81568 4216 81632
rect 4280 81568 4296 81632
rect 4360 81568 4376 81632
rect 4440 81568 4456 81632
rect 4520 81568 4528 81632
rect 4208 80544 4528 81568
rect 4208 80480 4216 80544
rect 4280 80480 4296 80544
rect 4360 80480 4376 80544
rect 4440 80480 4456 80544
rect 4520 80480 4528 80544
rect 4208 79456 4528 80480
rect 4208 79392 4216 79456
rect 4280 79392 4296 79456
rect 4360 79392 4376 79456
rect 4440 79392 4456 79456
rect 4520 79392 4528 79456
rect 4208 78368 4528 79392
rect 4208 78304 4216 78368
rect 4280 78304 4296 78368
rect 4360 78304 4376 78368
rect 4440 78304 4456 78368
rect 4520 78304 4528 78368
rect 4208 77280 4528 78304
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 76192 4528 77216
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 75104 4528 76128
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 4208 74016 4528 75040
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 72928 4528 73952
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 71840 4528 72864
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 70752 4528 71776
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 69664 4528 70688
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 68576 4528 69600
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 67488 4528 68512
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 66400 4528 67424
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 65312 4528 66336
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 64224 4528 65248
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 63136 4528 64160
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 62048 4528 63072
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 60960 4528 61984
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 59872 4528 60896
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 58784 4528 59808
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 57696 4528 58720
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 56608 4528 57632
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 55520 4528 56544
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 54432 4528 55456
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 53344 4528 54368
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 52256 4528 53280
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 51168 4528 52192
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 50080 4528 51104
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 48992 4528 50016
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 47904 4528 48928
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 46816 4528 47840
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 116992 19888 117552
rect 19568 116928 19576 116992
rect 19640 116928 19656 116992
rect 19720 116928 19736 116992
rect 19800 116928 19816 116992
rect 19880 116928 19888 116992
rect 19568 115904 19888 116928
rect 19568 115840 19576 115904
rect 19640 115840 19656 115904
rect 19720 115840 19736 115904
rect 19800 115840 19816 115904
rect 19880 115840 19888 115904
rect 19568 114816 19888 115840
rect 19568 114752 19576 114816
rect 19640 114752 19656 114816
rect 19720 114752 19736 114816
rect 19800 114752 19816 114816
rect 19880 114752 19888 114816
rect 19568 113728 19888 114752
rect 19568 113664 19576 113728
rect 19640 113664 19656 113728
rect 19720 113664 19736 113728
rect 19800 113664 19816 113728
rect 19880 113664 19888 113728
rect 19568 112640 19888 113664
rect 19568 112576 19576 112640
rect 19640 112576 19656 112640
rect 19720 112576 19736 112640
rect 19800 112576 19816 112640
rect 19880 112576 19888 112640
rect 19568 111552 19888 112576
rect 19568 111488 19576 111552
rect 19640 111488 19656 111552
rect 19720 111488 19736 111552
rect 19800 111488 19816 111552
rect 19880 111488 19888 111552
rect 19568 110464 19888 111488
rect 19568 110400 19576 110464
rect 19640 110400 19656 110464
rect 19720 110400 19736 110464
rect 19800 110400 19816 110464
rect 19880 110400 19888 110464
rect 19568 109376 19888 110400
rect 19568 109312 19576 109376
rect 19640 109312 19656 109376
rect 19720 109312 19736 109376
rect 19800 109312 19816 109376
rect 19880 109312 19888 109376
rect 19568 108288 19888 109312
rect 19568 108224 19576 108288
rect 19640 108224 19656 108288
rect 19720 108224 19736 108288
rect 19800 108224 19816 108288
rect 19880 108224 19888 108288
rect 19568 107200 19888 108224
rect 19568 107136 19576 107200
rect 19640 107136 19656 107200
rect 19720 107136 19736 107200
rect 19800 107136 19816 107200
rect 19880 107136 19888 107200
rect 19568 106112 19888 107136
rect 19568 106048 19576 106112
rect 19640 106048 19656 106112
rect 19720 106048 19736 106112
rect 19800 106048 19816 106112
rect 19880 106048 19888 106112
rect 19568 105024 19888 106048
rect 19568 104960 19576 105024
rect 19640 104960 19656 105024
rect 19720 104960 19736 105024
rect 19800 104960 19816 105024
rect 19880 104960 19888 105024
rect 19568 103936 19888 104960
rect 19568 103872 19576 103936
rect 19640 103872 19656 103936
rect 19720 103872 19736 103936
rect 19800 103872 19816 103936
rect 19880 103872 19888 103936
rect 19568 102848 19888 103872
rect 19568 102784 19576 102848
rect 19640 102784 19656 102848
rect 19720 102784 19736 102848
rect 19800 102784 19816 102848
rect 19880 102784 19888 102848
rect 19568 101760 19888 102784
rect 19568 101696 19576 101760
rect 19640 101696 19656 101760
rect 19720 101696 19736 101760
rect 19800 101696 19816 101760
rect 19880 101696 19888 101760
rect 19568 100672 19888 101696
rect 19568 100608 19576 100672
rect 19640 100608 19656 100672
rect 19720 100608 19736 100672
rect 19800 100608 19816 100672
rect 19880 100608 19888 100672
rect 19568 99584 19888 100608
rect 19568 99520 19576 99584
rect 19640 99520 19656 99584
rect 19720 99520 19736 99584
rect 19800 99520 19816 99584
rect 19880 99520 19888 99584
rect 19568 98496 19888 99520
rect 19568 98432 19576 98496
rect 19640 98432 19656 98496
rect 19720 98432 19736 98496
rect 19800 98432 19816 98496
rect 19880 98432 19888 98496
rect 19568 97408 19888 98432
rect 19568 97344 19576 97408
rect 19640 97344 19656 97408
rect 19720 97344 19736 97408
rect 19800 97344 19816 97408
rect 19880 97344 19888 97408
rect 19568 96320 19888 97344
rect 19568 96256 19576 96320
rect 19640 96256 19656 96320
rect 19720 96256 19736 96320
rect 19800 96256 19816 96320
rect 19880 96256 19888 96320
rect 19568 95232 19888 96256
rect 19568 95168 19576 95232
rect 19640 95168 19656 95232
rect 19720 95168 19736 95232
rect 19800 95168 19816 95232
rect 19880 95168 19888 95232
rect 19568 94144 19888 95168
rect 19568 94080 19576 94144
rect 19640 94080 19656 94144
rect 19720 94080 19736 94144
rect 19800 94080 19816 94144
rect 19880 94080 19888 94144
rect 19568 93056 19888 94080
rect 19568 92992 19576 93056
rect 19640 92992 19656 93056
rect 19720 92992 19736 93056
rect 19800 92992 19816 93056
rect 19880 92992 19888 93056
rect 19568 91968 19888 92992
rect 19568 91904 19576 91968
rect 19640 91904 19656 91968
rect 19720 91904 19736 91968
rect 19800 91904 19816 91968
rect 19880 91904 19888 91968
rect 19568 90880 19888 91904
rect 19568 90816 19576 90880
rect 19640 90816 19656 90880
rect 19720 90816 19736 90880
rect 19800 90816 19816 90880
rect 19880 90816 19888 90880
rect 19568 89792 19888 90816
rect 19568 89728 19576 89792
rect 19640 89728 19656 89792
rect 19720 89728 19736 89792
rect 19800 89728 19816 89792
rect 19880 89728 19888 89792
rect 19568 88704 19888 89728
rect 19568 88640 19576 88704
rect 19640 88640 19656 88704
rect 19720 88640 19736 88704
rect 19800 88640 19816 88704
rect 19880 88640 19888 88704
rect 19568 87616 19888 88640
rect 19568 87552 19576 87616
rect 19640 87552 19656 87616
rect 19720 87552 19736 87616
rect 19800 87552 19816 87616
rect 19880 87552 19888 87616
rect 19568 86528 19888 87552
rect 19568 86464 19576 86528
rect 19640 86464 19656 86528
rect 19720 86464 19736 86528
rect 19800 86464 19816 86528
rect 19880 86464 19888 86528
rect 19568 85440 19888 86464
rect 19568 85376 19576 85440
rect 19640 85376 19656 85440
rect 19720 85376 19736 85440
rect 19800 85376 19816 85440
rect 19880 85376 19888 85440
rect 19568 84352 19888 85376
rect 19568 84288 19576 84352
rect 19640 84288 19656 84352
rect 19720 84288 19736 84352
rect 19800 84288 19816 84352
rect 19880 84288 19888 84352
rect 19568 83264 19888 84288
rect 19568 83200 19576 83264
rect 19640 83200 19656 83264
rect 19720 83200 19736 83264
rect 19800 83200 19816 83264
rect 19880 83200 19888 83264
rect 19568 82176 19888 83200
rect 19568 82112 19576 82176
rect 19640 82112 19656 82176
rect 19720 82112 19736 82176
rect 19800 82112 19816 82176
rect 19880 82112 19888 82176
rect 19568 81088 19888 82112
rect 19568 81024 19576 81088
rect 19640 81024 19656 81088
rect 19720 81024 19736 81088
rect 19800 81024 19816 81088
rect 19880 81024 19888 81088
rect 19568 80000 19888 81024
rect 19568 79936 19576 80000
rect 19640 79936 19656 80000
rect 19720 79936 19736 80000
rect 19800 79936 19816 80000
rect 19880 79936 19888 80000
rect 19568 78912 19888 79936
rect 19568 78848 19576 78912
rect 19640 78848 19656 78912
rect 19720 78848 19736 78912
rect 19800 78848 19816 78912
rect 19880 78848 19888 78912
rect 19568 77824 19888 78848
rect 19568 77760 19576 77824
rect 19640 77760 19656 77824
rect 19720 77760 19736 77824
rect 19800 77760 19816 77824
rect 19880 77760 19888 77824
rect 19568 76736 19888 77760
rect 19568 76672 19576 76736
rect 19640 76672 19656 76736
rect 19720 76672 19736 76736
rect 19800 76672 19816 76736
rect 19880 76672 19888 76736
rect 19568 75648 19888 76672
rect 19568 75584 19576 75648
rect 19640 75584 19656 75648
rect 19720 75584 19736 75648
rect 19800 75584 19816 75648
rect 19880 75584 19888 75648
rect 19568 74560 19888 75584
rect 19568 74496 19576 74560
rect 19640 74496 19656 74560
rect 19720 74496 19736 74560
rect 19800 74496 19816 74560
rect 19880 74496 19888 74560
rect 19568 73472 19888 74496
rect 19568 73408 19576 73472
rect 19640 73408 19656 73472
rect 19720 73408 19736 73472
rect 19800 73408 19816 73472
rect 19880 73408 19888 73472
rect 19568 72384 19888 73408
rect 19568 72320 19576 72384
rect 19640 72320 19656 72384
rect 19720 72320 19736 72384
rect 19800 72320 19816 72384
rect 19880 72320 19888 72384
rect 19568 71296 19888 72320
rect 19568 71232 19576 71296
rect 19640 71232 19656 71296
rect 19720 71232 19736 71296
rect 19800 71232 19816 71296
rect 19880 71232 19888 71296
rect 19568 70208 19888 71232
rect 19568 70144 19576 70208
rect 19640 70144 19656 70208
rect 19720 70144 19736 70208
rect 19800 70144 19816 70208
rect 19880 70144 19888 70208
rect 19568 69120 19888 70144
rect 19568 69056 19576 69120
rect 19640 69056 19656 69120
rect 19720 69056 19736 69120
rect 19800 69056 19816 69120
rect 19880 69056 19888 69120
rect 19568 68032 19888 69056
rect 19568 67968 19576 68032
rect 19640 67968 19656 68032
rect 19720 67968 19736 68032
rect 19800 67968 19816 68032
rect 19880 67968 19888 68032
rect 19568 66944 19888 67968
rect 19568 66880 19576 66944
rect 19640 66880 19656 66944
rect 19720 66880 19736 66944
rect 19800 66880 19816 66944
rect 19880 66880 19888 66944
rect 19568 65856 19888 66880
rect 19568 65792 19576 65856
rect 19640 65792 19656 65856
rect 19720 65792 19736 65856
rect 19800 65792 19816 65856
rect 19880 65792 19888 65856
rect 19568 64768 19888 65792
rect 19568 64704 19576 64768
rect 19640 64704 19656 64768
rect 19720 64704 19736 64768
rect 19800 64704 19816 64768
rect 19880 64704 19888 64768
rect 19568 63680 19888 64704
rect 19568 63616 19576 63680
rect 19640 63616 19656 63680
rect 19720 63616 19736 63680
rect 19800 63616 19816 63680
rect 19880 63616 19888 63680
rect 19568 62592 19888 63616
rect 19568 62528 19576 62592
rect 19640 62528 19656 62592
rect 19720 62528 19736 62592
rect 19800 62528 19816 62592
rect 19880 62528 19888 62592
rect 19568 61504 19888 62528
rect 19568 61440 19576 61504
rect 19640 61440 19656 61504
rect 19720 61440 19736 61504
rect 19800 61440 19816 61504
rect 19880 61440 19888 61504
rect 19568 60416 19888 61440
rect 19568 60352 19576 60416
rect 19640 60352 19656 60416
rect 19720 60352 19736 60416
rect 19800 60352 19816 60416
rect 19880 60352 19888 60416
rect 19568 59328 19888 60352
rect 19568 59264 19576 59328
rect 19640 59264 19656 59328
rect 19720 59264 19736 59328
rect 19800 59264 19816 59328
rect 19880 59264 19888 59328
rect 19568 58240 19888 59264
rect 19568 58176 19576 58240
rect 19640 58176 19656 58240
rect 19720 58176 19736 58240
rect 19800 58176 19816 58240
rect 19880 58176 19888 58240
rect 19568 57152 19888 58176
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 19568 56064 19888 57088
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 19568 54976 19888 56000
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 19568 53888 19888 54912
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 52800 19888 53824
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 19568 51712 19888 52736
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 50624 19888 51648
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 19568 49536 19888 50560
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 48448 19888 49472
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 19568 47360 19888 48384
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 46272 19888 47296
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 45184 19888 46208
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 44096 19888 45120
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
rect 34928 117536 35248 117552
rect 34928 117472 34936 117536
rect 35000 117472 35016 117536
rect 35080 117472 35096 117536
rect 35160 117472 35176 117536
rect 35240 117472 35248 117536
rect 34928 116448 35248 117472
rect 34928 116384 34936 116448
rect 35000 116384 35016 116448
rect 35080 116384 35096 116448
rect 35160 116384 35176 116448
rect 35240 116384 35248 116448
rect 34928 115360 35248 116384
rect 34928 115296 34936 115360
rect 35000 115296 35016 115360
rect 35080 115296 35096 115360
rect 35160 115296 35176 115360
rect 35240 115296 35248 115360
rect 34928 114272 35248 115296
rect 34928 114208 34936 114272
rect 35000 114208 35016 114272
rect 35080 114208 35096 114272
rect 35160 114208 35176 114272
rect 35240 114208 35248 114272
rect 34928 113184 35248 114208
rect 34928 113120 34936 113184
rect 35000 113120 35016 113184
rect 35080 113120 35096 113184
rect 35160 113120 35176 113184
rect 35240 113120 35248 113184
rect 34928 112096 35248 113120
rect 34928 112032 34936 112096
rect 35000 112032 35016 112096
rect 35080 112032 35096 112096
rect 35160 112032 35176 112096
rect 35240 112032 35248 112096
rect 34928 111008 35248 112032
rect 34928 110944 34936 111008
rect 35000 110944 35016 111008
rect 35080 110944 35096 111008
rect 35160 110944 35176 111008
rect 35240 110944 35248 111008
rect 34928 109920 35248 110944
rect 34928 109856 34936 109920
rect 35000 109856 35016 109920
rect 35080 109856 35096 109920
rect 35160 109856 35176 109920
rect 35240 109856 35248 109920
rect 34928 108832 35248 109856
rect 34928 108768 34936 108832
rect 35000 108768 35016 108832
rect 35080 108768 35096 108832
rect 35160 108768 35176 108832
rect 35240 108768 35248 108832
rect 34928 107744 35248 108768
rect 34928 107680 34936 107744
rect 35000 107680 35016 107744
rect 35080 107680 35096 107744
rect 35160 107680 35176 107744
rect 35240 107680 35248 107744
rect 34928 106656 35248 107680
rect 34928 106592 34936 106656
rect 35000 106592 35016 106656
rect 35080 106592 35096 106656
rect 35160 106592 35176 106656
rect 35240 106592 35248 106656
rect 34928 105568 35248 106592
rect 34928 105504 34936 105568
rect 35000 105504 35016 105568
rect 35080 105504 35096 105568
rect 35160 105504 35176 105568
rect 35240 105504 35248 105568
rect 34928 104480 35248 105504
rect 34928 104416 34936 104480
rect 35000 104416 35016 104480
rect 35080 104416 35096 104480
rect 35160 104416 35176 104480
rect 35240 104416 35248 104480
rect 34928 103392 35248 104416
rect 34928 103328 34936 103392
rect 35000 103328 35016 103392
rect 35080 103328 35096 103392
rect 35160 103328 35176 103392
rect 35240 103328 35248 103392
rect 34928 102304 35248 103328
rect 34928 102240 34936 102304
rect 35000 102240 35016 102304
rect 35080 102240 35096 102304
rect 35160 102240 35176 102304
rect 35240 102240 35248 102304
rect 34928 101216 35248 102240
rect 34928 101152 34936 101216
rect 35000 101152 35016 101216
rect 35080 101152 35096 101216
rect 35160 101152 35176 101216
rect 35240 101152 35248 101216
rect 34928 100128 35248 101152
rect 34928 100064 34936 100128
rect 35000 100064 35016 100128
rect 35080 100064 35096 100128
rect 35160 100064 35176 100128
rect 35240 100064 35248 100128
rect 34928 99040 35248 100064
rect 34928 98976 34936 99040
rect 35000 98976 35016 99040
rect 35080 98976 35096 99040
rect 35160 98976 35176 99040
rect 35240 98976 35248 99040
rect 34928 97952 35248 98976
rect 34928 97888 34936 97952
rect 35000 97888 35016 97952
rect 35080 97888 35096 97952
rect 35160 97888 35176 97952
rect 35240 97888 35248 97952
rect 34928 96864 35248 97888
rect 34928 96800 34936 96864
rect 35000 96800 35016 96864
rect 35080 96800 35096 96864
rect 35160 96800 35176 96864
rect 35240 96800 35248 96864
rect 34928 95776 35248 96800
rect 34928 95712 34936 95776
rect 35000 95712 35016 95776
rect 35080 95712 35096 95776
rect 35160 95712 35176 95776
rect 35240 95712 35248 95776
rect 34928 94688 35248 95712
rect 34928 94624 34936 94688
rect 35000 94624 35016 94688
rect 35080 94624 35096 94688
rect 35160 94624 35176 94688
rect 35240 94624 35248 94688
rect 34928 93600 35248 94624
rect 34928 93536 34936 93600
rect 35000 93536 35016 93600
rect 35080 93536 35096 93600
rect 35160 93536 35176 93600
rect 35240 93536 35248 93600
rect 34928 92512 35248 93536
rect 34928 92448 34936 92512
rect 35000 92448 35016 92512
rect 35080 92448 35096 92512
rect 35160 92448 35176 92512
rect 35240 92448 35248 92512
rect 34928 91424 35248 92448
rect 34928 91360 34936 91424
rect 35000 91360 35016 91424
rect 35080 91360 35096 91424
rect 35160 91360 35176 91424
rect 35240 91360 35248 91424
rect 34928 90336 35248 91360
rect 34928 90272 34936 90336
rect 35000 90272 35016 90336
rect 35080 90272 35096 90336
rect 35160 90272 35176 90336
rect 35240 90272 35248 90336
rect 34928 89248 35248 90272
rect 34928 89184 34936 89248
rect 35000 89184 35016 89248
rect 35080 89184 35096 89248
rect 35160 89184 35176 89248
rect 35240 89184 35248 89248
rect 34928 88160 35248 89184
rect 34928 88096 34936 88160
rect 35000 88096 35016 88160
rect 35080 88096 35096 88160
rect 35160 88096 35176 88160
rect 35240 88096 35248 88160
rect 34928 87072 35248 88096
rect 34928 87008 34936 87072
rect 35000 87008 35016 87072
rect 35080 87008 35096 87072
rect 35160 87008 35176 87072
rect 35240 87008 35248 87072
rect 34928 85984 35248 87008
rect 34928 85920 34936 85984
rect 35000 85920 35016 85984
rect 35080 85920 35096 85984
rect 35160 85920 35176 85984
rect 35240 85920 35248 85984
rect 34928 84896 35248 85920
rect 34928 84832 34936 84896
rect 35000 84832 35016 84896
rect 35080 84832 35096 84896
rect 35160 84832 35176 84896
rect 35240 84832 35248 84896
rect 34928 83808 35248 84832
rect 34928 83744 34936 83808
rect 35000 83744 35016 83808
rect 35080 83744 35096 83808
rect 35160 83744 35176 83808
rect 35240 83744 35248 83808
rect 34928 82720 35248 83744
rect 34928 82656 34936 82720
rect 35000 82656 35016 82720
rect 35080 82656 35096 82720
rect 35160 82656 35176 82720
rect 35240 82656 35248 82720
rect 34928 81632 35248 82656
rect 34928 81568 34936 81632
rect 35000 81568 35016 81632
rect 35080 81568 35096 81632
rect 35160 81568 35176 81632
rect 35240 81568 35248 81632
rect 34928 80544 35248 81568
rect 34928 80480 34936 80544
rect 35000 80480 35016 80544
rect 35080 80480 35096 80544
rect 35160 80480 35176 80544
rect 35240 80480 35248 80544
rect 34928 79456 35248 80480
rect 34928 79392 34936 79456
rect 35000 79392 35016 79456
rect 35080 79392 35096 79456
rect 35160 79392 35176 79456
rect 35240 79392 35248 79456
rect 34928 78368 35248 79392
rect 34928 78304 34936 78368
rect 35000 78304 35016 78368
rect 35080 78304 35096 78368
rect 35160 78304 35176 78368
rect 35240 78304 35248 78368
rect 34928 77280 35248 78304
rect 34928 77216 34936 77280
rect 35000 77216 35016 77280
rect 35080 77216 35096 77280
rect 35160 77216 35176 77280
rect 35240 77216 35248 77280
rect 34928 76192 35248 77216
rect 34928 76128 34936 76192
rect 35000 76128 35016 76192
rect 35080 76128 35096 76192
rect 35160 76128 35176 76192
rect 35240 76128 35248 76192
rect 34928 75104 35248 76128
rect 34928 75040 34936 75104
rect 35000 75040 35016 75104
rect 35080 75040 35096 75104
rect 35160 75040 35176 75104
rect 35240 75040 35248 75104
rect 34928 74016 35248 75040
rect 34928 73952 34936 74016
rect 35000 73952 35016 74016
rect 35080 73952 35096 74016
rect 35160 73952 35176 74016
rect 35240 73952 35248 74016
rect 34928 72928 35248 73952
rect 34928 72864 34936 72928
rect 35000 72864 35016 72928
rect 35080 72864 35096 72928
rect 35160 72864 35176 72928
rect 35240 72864 35248 72928
rect 34928 71840 35248 72864
rect 34928 71776 34936 71840
rect 35000 71776 35016 71840
rect 35080 71776 35096 71840
rect 35160 71776 35176 71840
rect 35240 71776 35248 71840
rect 34928 70752 35248 71776
rect 34928 70688 34936 70752
rect 35000 70688 35016 70752
rect 35080 70688 35096 70752
rect 35160 70688 35176 70752
rect 35240 70688 35248 70752
rect 34928 69664 35248 70688
rect 34928 69600 34936 69664
rect 35000 69600 35016 69664
rect 35080 69600 35096 69664
rect 35160 69600 35176 69664
rect 35240 69600 35248 69664
rect 34928 68576 35248 69600
rect 34928 68512 34936 68576
rect 35000 68512 35016 68576
rect 35080 68512 35096 68576
rect 35160 68512 35176 68576
rect 35240 68512 35248 68576
rect 34928 67488 35248 68512
rect 34928 67424 34936 67488
rect 35000 67424 35016 67488
rect 35080 67424 35096 67488
rect 35160 67424 35176 67488
rect 35240 67424 35248 67488
rect 34928 66400 35248 67424
rect 34928 66336 34936 66400
rect 35000 66336 35016 66400
rect 35080 66336 35096 66400
rect 35160 66336 35176 66400
rect 35240 66336 35248 66400
rect 34928 65312 35248 66336
rect 34928 65248 34936 65312
rect 35000 65248 35016 65312
rect 35080 65248 35096 65312
rect 35160 65248 35176 65312
rect 35240 65248 35248 65312
rect 34928 64224 35248 65248
rect 34928 64160 34936 64224
rect 35000 64160 35016 64224
rect 35080 64160 35096 64224
rect 35160 64160 35176 64224
rect 35240 64160 35248 64224
rect 34928 63136 35248 64160
rect 34928 63072 34936 63136
rect 35000 63072 35016 63136
rect 35080 63072 35096 63136
rect 35160 63072 35176 63136
rect 35240 63072 35248 63136
rect 34928 62048 35248 63072
rect 34928 61984 34936 62048
rect 35000 61984 35016 62048
rect 35080 61984 35096 62048
rect 35160 61984 35176 62048
rect 35240 61984 35248 62048
rect 34928 60960 35248 61984
rect 34928 60896 34936 60960
rect 35000 60896 35016 60960
rect 35080 60896 35096 60960
rect 35160 60896 35176 60960
rect 35240 60896 35248 60960
rect 34928 59872 35248 60896
rect 34928 59808 34936 59872
rect 35000 59808 35016 59872
rect 35080 59808 35096 59872
rect 35160 59808 35176 59872
rect 35240 59808 35248 59872
rect 34928 58784 35248 59808
rect 34928 58720 34936 58784
rect 35000 58720 35016 58784
rect 35080 58720 35096 58784
rect 35160 58720 35176 58784
rect 35240 58720 35248 58784
rect 34928 57696 35248 58720
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 56608 35248 57632
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 34928 55520 35248 56544
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 54432 35248 55456
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 34928 53344 35248 54368
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 34928 52256 35248 53280
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 34928 51168 35248 52192
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 34928 50080 35248 51104
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 48992 35248 50016
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 34928 47904 35248 48928
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 46816 35248 47840
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 45728 35248 46752
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 44640 35248 45664
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 43552 35248 44576
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 42464 35248 43488
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
use sky130_fd_sc_hd__decap_4  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3
timestamp 1623621585
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1623621585
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1623621585
transform 1 0 2300 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1623621585
transform 1 0 2300 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input330 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1748 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input319
timestamp 1623621585
transform 1 0 1748 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input455
timestamp 1623621585
transform 1 0 2668 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input341
timestamp 1623621585
transform 1 0 2668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1623621585
transform 1 0 3772 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input456 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 4232 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input500
timestamp 1623621585
transform 1 0 4600 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 3220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1623621585
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 4784 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_23
timestamp 1623621585
transform 1 0 3220 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_30
timestamp 1623621585
transform 1 0 3864 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1623621585
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input478
timestamp 1623621585
transform 1 0 5520 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input511
timestamp 1623621585
transform 1 0 5888 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1623621585
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1623621585
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_44
timestamp 1623621585
transform 1 0 5152 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_58
timestamp 1623621585
transform 1 0 6440 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  input481
timestamp 1623621585
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input482
timestamp 1623621585
transform 1 0 8188 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input514 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 7176 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output707 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69
timestamp 1623621585
transform 1 0 7452 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1623621585
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_70
timestamp 1623621585
transform 1 0 7544 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_78
timestamp 1623621585
transform 1 0 8280 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_87
timestamp 1623621585
transform 1 0 9108 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88
timestamp 1623621585
transform 1 0 9200 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input483
timestamp 1623621585
transform 1 0 9476 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1623621585
transform 1 0 9016 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1623621585
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_95
timestamp 1623621585
transform 1 0 9844 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_96 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 9936 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output709
timestamp 1623621585
transform 1 0 10212 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input484
timestamp 1623621585
transform 1 0 10120 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_103
timestamp 1623621585
transform 1 0 10580 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp 1623621585
transform 1 0 10672 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1623621585
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input485
timestamp 1623621585
transform 1 0 11132 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input486
timestamp 1623621585
transform 1 0 11040 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input517
timestamp 1623621585
transform 1 0 12236 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input518
timestamp 1623621585
transform 1 0 12052 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1623621585
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1623621585
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_115
timestamp 1623621585
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1623621585
transform 1 0 12604 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_129 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 12972 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1623621585
transform 1 0 13156 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127
timestamp 1623621585
transform 1 0 12788 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input520 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 13248 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input487
timestamp 1623621585
transform 1 0 13064 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_144
timestamp 1623621585
transform 1 0 14352 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_142
timestamp 1623621585
transform 1 0 14168 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_136
timestamp 1623621585
transform 1 0 13616 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1623621585
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1623621585
transform 1 0 14260 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1623621585
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_151
timestamp 1623621585
transform 1 0 14996 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1623621585
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input491
timestamp 1623621585
transform 1 0 15364 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input458 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 14720 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input457
timestamp 1623621585
transform 1 0 14904 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_161
timestamp 1623621585
transform 1 0 15916 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_160
timestamp 1623621585
transform 1 0 15824 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1623621585
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input492
timestamp 1623621585
transform 1 0 16284 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input459
timestamp 1623621585
transform 1 0 15916 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_175
timestamp 1623621585
transform 1 0 17204 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_169
timestamp 1623621585
transform 1 0 16652 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1623621585
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1623621585
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input493
timestamp 1623621585
transform 1 0 17296 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1623621585
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_186
timestamp 1623621585
transform 1 0 18216 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_182
timestamp 1623621585
transform 1 0 17848 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input460
timestamp 1623621585
transform 1 0 17572 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input494
timestamp 1623621585
transform 1 0 18308 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_193
timestamp 1623621585
transform 1 0 18860 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_192
timestamp 1623621585
transform 1 0 18768 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_188
timestamp 1623621585
transform 1 0 18400 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input462
timestamp 1623621585
transform 1 0 18860 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1623621585
transform 1 0 19596 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_199
timestamp 1623621585
transform 1 0 19412 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1623621585
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1623621585
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1623621585
transform 1 0 19504 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1623621585
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _614_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 19964 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input496
timestamp 1623621585
transform 1 0 20240 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input497
timestamp 1623621585
transform 1 0 21160 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output689
timestamp 1623621585
transform 1 0 21160 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output690
timestamp 1623621585
transform 1 0 21896 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_214
timestamp 1623621585
transform 1 0 20792 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_224
timestamp 1623621585
transform 1 0 21712 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_214
timestamp 1623621585
transform 1 0 20792 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_222
timestamp 1623621585
transform 1 0 21528 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_238
timestamp 1623621585
transform 1 0 23000 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_230
timestamp 1623621585
transform 1 0 22264 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1623621585
transform 1 0 22540 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output691
timestamp 1623621585
transform 1 0 22632 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input498
timestamp 1623621585
transform 1 0 22908 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1623621585
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_242
timestamp 1623621585
transform 1 0 23368 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_243
timestamp 1623621585
transform 1 0 23460 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output692
timestamp 1623621585
transform 1 0 23460 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_247
timestamp 1623621585
transform 1 0 23828 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_258
timestamp 1623621585
transform 1 0 24840 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_255
timestamp 1623621585
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1623621585
transform 1 0 24748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_251
timestamp 1623621585
transform 1 0 24196 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  input502
timestamp 1623621585
transform 1 0 24380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1623621585
transform 1 0 24748 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_262
timestamp 1623621585
transform 1 0 25208 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1623621585
transform 1 0 25116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _617_
timestamp 1623621585
transform 1 0 25208 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_270
timestamp 1623621585
transform 1 0 25944 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_279
timestamp 1623621585
transform 1 0 26772 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1623621585
transform 1 0 26036 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_277
timestamp 1623621585
transform 1 0 26588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output696
timestamp 1623621585
transform 1 0 26404 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input503
timestamp 1623621585
transform 1 0 26036 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1623621585
transform 1 0 27416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_281
timestamp 1623621585
transform 1 0 26956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input504
timestamp 1623621585
transform 1 0 27048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1623621585
transform 1 0 27784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _616_
timestamp 1623621585
transform 1 0 27508 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1623621585
transform 1 0 27876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input505
timestamp 1623621585
transform 1 0 28244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input507
timestamp 1623621585
transform 1 0 29532 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output698
timestamp 1623621585
transform 1 0 28704 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_299
timestamp 1623621585
transform 1 0 28612 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_307
timestamp 1623621585
transform 1 0 29348 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_296
timestamp 1623621585
transform 1 0 28336 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_304
timestamp 1623621585
transform 1 0 29072 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_312
timestamp 1623621585
transform 1 0 29808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__or4b_4  _620_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 30452 0 1 2720
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1623621585
transform 1 0 30452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1623621585
transform 1 0 29992 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input508
timestamp 1623621585
transform 1 0 30912 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_315
timestamp 1623621585
transform 1 0 30084 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp 1623621585
transform 1 0 30544 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_330
timestamp 1623621585
transform 1 0 31464 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_315
timestamp 1623621585
transform 1 0 30084 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_330
timestamp 1623621585
transform 1 0 31464 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_338
timestamp 1623621585
transform 1 0 32200 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_338
timestamp 1623621585
transform 1 0 32200 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output702
timestamp 1623621585
transform 1 0 32568 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output701
timestamp 1623621585
transform 1 0 31832 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output614
timestamp 1623621585
transform 1 0 32384 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_346
timestamp 1623621585
transform 1 0 32936 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1623621585
transform 1 0 33212 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_344
timestamp 1623621585
transform 1 0 32752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output703
timestamp 1623621585
transform 1 0 33304 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1623621585
transform 1 0 33120 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_354
timestamp 1623621585
transform 1 0 33672 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input510
timestamp 1623621585
transform 1 0 33580 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1623621585
transform 1 0 35236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input512
timestamp 1623621585
transform 1 0 34500 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output667
timestamp 1623621585
transform 1 0 34500 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1623621585
transform 1 0 34132 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_367
timestamp 1623621585
transform 1 0 34868 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_375
timestamp 1623621585
transform 1 0 35604 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_362
timestamp 1623621585
transform 1 0 34408 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_367
timestamp 1623621585
transform 1 0 34868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_372
timestamp 1623621585
transform 1 0 35328 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_380
timestamp 1623621585
transform 1 0 36064 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_378
timestamp 1623621585
transform 1 0 35880 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input513
timestamp 1623621585
transform 1 0 35696 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1623621585
transform 1 0 36248 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1623621585
transform 1 0 35788 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_389
timestamp 1623621585
transform 1 0 36892 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_384
timestamp 1623621585
transform 1 0 36432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_386
timestamp 1623621585
transform 1 0 36616 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output619
timestamp 1623621585
transform 1 0 36524 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_394
timestamp 1623621585
transform 1 0 37352 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input62
timestamp 1623621585
transform 1 0 37444 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1623621585
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1623621585
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1623621585
transform 1 0 38456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output618
timestamp 1623621585
transform 1 0 37812 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_401
timestamp 1623621585
transform 1 0 37996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_405
timestamp 1623621585
transform 1 0 38364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_397
timestamp 1623621585
transform 1 0 37628 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1623621585
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1623621585
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input344
timestamp 1623621585
transform 1 0 1748 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1623621585
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_13
timestamp 1623621585
transform 1 0 2300 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input489
timestamp 1623621585
transform 1 0 3312 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output681
timestamp 1623621585
transform 1 0 4232 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_21
timestamp 1623621585
transform 1 0 3036 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_30
timestamp 1623621585
transform 1 0 3864 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_38
timestamp 1623621585
transform 1 0 4600 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1623621585
transform 1 0 6348 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input521
timestamp 1623621585
transform 1 0 5704 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output693
timestamp 1623621585
transform 1 0 4968 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output704
timestamp 1623621585
transform 1 0 6808 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_46
timestamp 1623621585
transform 1 0 5336 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1623621585
transform 1 0 5980 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_58
timestamp 1623621585
transform 1 0 6440 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input515
timestamp 1623621585
transform 1 0 8188 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input524
timestamp 1623621585
transform 1 0 7544 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1623621585
transform 1 0 7176 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1623621585
transform 1 0 7820 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1623621585
transform 1 0 8464 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input516
timestamp 1623621585
transform 1 0 9568 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output708
timestamp 1623621585
transform 1 0 8832 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1623621585
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_95
timestamp 1623621585
transform 1 0 9844 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_103
timestamp 1623621585
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__and3b_1  _615_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 12052 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1623621585
transform 1 0 11592 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output710
timestamp 1623621585
transform 1 0 10764 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_109
timestamp 1623621585
transform 1 0 11132 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_113
timestamp 1623621585
transform 1 0 11500 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_115
timestamp 1623621585
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input519
timestamp 1623621585
transform 1 0 13064 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output713
timestamp 1623621585
transform 1 0 13984 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_126
timestamp 1623621585
transform 1 0 12696 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1623621585
transform 1 0 13616 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1623621585
transform 1 0 14352 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output683
timestamp 1623621585
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output684
timestamp 1623621585
transform 1 0 15640 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_152
timestamp 1623621585
transform 1 0 15088 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_162
timestamp 1623621585
transform 1 0 16008 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1623621585
transform 1 0 16836 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input461
timestamp 1623621585
transform 1 0 17940 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_170
timestamp 1623621585
transform 1 0 16744 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_172
timestamp 1623621585
transform 1 0 16928 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_180
timestamp 1623621585
transform 1 0 17664 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1623621585
transform 1 0 18308 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input495
timestamp 1623621585
transform 1 0 19228 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output688
timestamp 1623621585
transform 1 0 19964 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_195
timestamp 1623621585
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_201
timestamp 1623621585
transform 1 0 19596 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _711_
timestamp 1623621585
transform 1 0 20700 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1623621585
transform 1 0 22080 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input464 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 21344 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1623621585
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_216
timestamp 1623621585
transform 1 0 20976 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_223
timestamp 1623621585
transform 1 0 21620 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_227
timestamp 1623621585
transform 1 0 21988 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_229
timestamp 1623621585
transform 1 0 22172 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _726_
timestamp 1623621585
transform 1 0 22540 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _727_
timestamp 1623621585
transform 1 0 23184 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input468
timestamp 1623621585
transform 1 0 23828 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_236
timestamp 1623621585
transform 1 0 22816 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_243
timestamp 1623621585
transform 1 0 23460 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_250
timestamp 1623621585
transform 1 0 24104 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output694
timestamp 1623621585
transform 1 0 24472 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output695
timestamp 1623621585
transform 1 0 25392 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_258
timestamp 1623621585
transform 1 0 24840 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_268
timestamp 1623621585
transform 1 0 25760 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _721_
timestamp 1623621585
transform 1 0 26404 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1623621585
transform 1 0 27324 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output697
timestamp 1623621585
transform 1 0 27784 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_274
timestamp 1623621585
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_278
timestamp 1623621585
transform 1 0 26680 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_284
timestamp 1623621585
transform 1 0 27232 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_286
timestamp 1623621585
transform 1 0 27416 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input472
timestamp 1623621585
transform 1 0 28520 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output699
timestamp 1623621585
transform 1 0 29348 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_294
timestamp 1623621585
transform 1 0 28152 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1623621585
transform 1 0 28796 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_311
timestamp 1623621585
transform 1 0 29716 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _741_
timestamp 1623621585
transform 1 0 31004 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _742_
timestamp 1623621585
transform 1 0 31648 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output700
timestamp 1623621585
transform 1 0 30268 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1623621585
transform 1 0 30636 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_328
timestamp 1623621585
transform 1 0 31280 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 33580 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1623621585
transform 1 0 32568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_335
timestamp 1623621585
transform 1 0 31924 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_341
timestamp 1623621585
transform 1 0 32476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_343
timestamp 1623621585
transform 1 0 32660 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_351
timestamp 1623621585
transform 1 0 33396 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output666
timestamp 1623621585
transform 1 0 35420 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output705
timestamp 1623621585
transform 1 0 34224 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_356
timestamp 1623621585
transform 1 0 33856 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_364
timestamp 1623621585
transform 1 0 34592 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_372
timestamp 1623621585
transform 1 0 35328 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output628
timestamp 1623621585
transform 1 0 36156 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output641
timestamp 1623621585
transform 1 0 37076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_377
timestamp 1623621585
transform 1 0 35788 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_385
timestamp 1623621585
transform 1 0 36524 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_395
timestamp 1623621585
transform 1 0 37444 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1623621585
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1623621585
transform 1 0 37812 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_400
timestamp 1623621585
transform 1 0 37904 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_406
timestamp 1623621585
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1623621585
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input345
timestamp 1623621585
transform 1 0 1748 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input526
timestamp 1623621585
transform 1 0 2668 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1623621585
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1623621585
transform 1 0 2300 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1623621585
transform 1 0 3772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output682
timestamp 1623621585
transform 1 0 4232 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_23
timestamp 1623621585
transform 1 0 3220 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1623621585
transform 1 0 3864 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_38
timestamp 1623621585
transform 1 0 4600 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input467
timestamp 1623621585
transform 1 0 4968 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input522
timestamp 1623621585
transform 1 0 5612 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input523
timestamp 1623621585
transform 1 0 6532 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_45
timestamp 1623621585
transform 1 0 5244 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_52
timestamp 1623621585
transform 1 0 5888 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_58
timestamp 1623621585
transform 1 0 6440 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1623621585
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1623621585
transform 1 0 9016 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_87
timestamp 1623621585
transform 1 0 9108 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_99
timestamp 1623621585
transform 1 0 10212 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output711
timestamp 1623621585
transform 1 0 11776 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_111
timestamp 1623621585
transform 1 0 11316 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_115
timestamp 1623621585
transform 1 0 11684 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_120
timestamp 1623621585
transform 1 0 12144 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1623621585
transform 1 0 14260 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output712
timestamp 1623621585
transform 1 0 12696 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_130
timestamp 1623621585
transform 1 0 13064 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_142
timestamp 1623621585
transform 1 0 14168 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_144
timestamp 1623621585
transform 1 0 14352 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input490
timestamp 1623621585
transform 1 0 14720 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_151
timestamp 1623621585
transform 1 0 14996 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_163
timestamp 1623621585
transform 1 0 16100 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output685
timestamp 1623621585
transform 1 0 16652 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output686
timestamp 1623621585
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_173
timestamp 1623621585
transform 1 0 17020 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_183
timestamp 1623621585
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1623621585
transform 1 0 19504 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input463
timestamp 1623621585
transform 1 0 19964 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output687
timestamp 1623621585
transform 1 0 18584 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1623621585
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_194
timestamp 1623621585
transform 1 0 18952 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_201
timestamp 1623621585
transform 1 0 19596 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1623621585
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input465
timestamp 1623621585
transform 1 0 21804 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1623621585
transform 1 0 21344 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_224
timestamp 1623621585
transform 1 0 21712 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_228
timestamp 1623621585
transform 1 0 22080 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input466
timestamp 1623621585
transform 1 0 22816 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input499
timestamp 1623621585
transform 1 0 23460 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input501
timestamp 1623621585
transform 1 0 24104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_239
timestamp 1623621585
transform 1 0 23092 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_246
timestamp 1623621585
transform 1 0 23736 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _732_
timestamp 1623621585
transform 1 0 25944 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1623621585
transform 1 0 24748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input469
timestamp 1623621585
transform 1 0 25208 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_253
timestamp 1623621585
transform 1 0 24380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_258
timestamp 1623621585
transform 1 0 24840 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_265
timestamp 1623621585
transform 1 0 25484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_269
timestamp 1623621585
transform 1 0 25852 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input470
timestamp 1623621585
transform 1 0 26588 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input471
timestamp 1623621585
transform 1 0 27232 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_273
timestamp 1623621585
transform 1 0 26220 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_280
timestamp 1623621585
transform 1 0 26864 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_287
timestamp 1623621585
transform 1 0 27508 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input473
timestamp 1623621585
transform 1 0 28704 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input506
timestamp 1623621585
transform 1 0 29348 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_299
timestamp 1623621585
transform 1 0 28612 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_303
timestamp 1623621585
transform 1 0 28980 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_310
timestamp 1623621585
transform 1 0 29624 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1623621585
transform 1 0 29992 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input474
timestamp 1623621585
transform 1 0 30452 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input475
timestamp 1623621585
transform 1 0 31096 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input476
timestamp 1623621585
transform 1 0 31740 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_315
timestamp 1623621585
transform 1 0 30084 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_322
timestamp 1623621585
transform 1 0 30728 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_329
timestamp 1623621585
transform 1 0 31372 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input90
timestamp 1623621585
transform 1 0 33396 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input477
timestamp 1623621585
transform 1 0 32568 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_336
timestamp 1623621585
transform 1 0 32016 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_345
timestamp 1623621585
transform 1 0 32844 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_354
timestamp 1623621585
transform 1 0 33672 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _747_
timestamp 1623621585
transform 1 0 34040 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1623621585
transform 1 0 35236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_361
timestamp 1623621585
transform 1 0 34316 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_369
timestamp 1623621585
transform 1 0 35052 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_372
timestamp 1623621585
transform 1 0 35328 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _750_
timestamp 1623621585
transform 1 0 35696 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output650
timestamp 1623621585
transform 1 0 37076 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output652
timestamp 1623621585
transform 1 0 36340 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_379
timestamp 1623621585
transform 1 0 35972 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1623621585
transform 1 0 36708 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_395
timestamp 1623621585
transform 1 0 37444 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1623621585
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output630
timestamp 1623621585
transform 1 0 37812 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1623621585
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1623621585
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input346
timestamp 1623621585
transform 1 0 1748 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output611
timestamp 1623621585
transform 1 0 2668 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1623621585
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1623621585
transform 1 0 2300 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _691_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 4140 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input488
timestamp 1623621585
transform 1 0 4784 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output613
timestamp 1623621585
transform 1 0 3404 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_21
timestamp 1623621585
transform 1 0 3036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1623621585
transform 1 0 3772 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_36
timestamp 1623621585
transform 1 0 4416 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1623621585
transform 1 0 6348 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_43
timestamp 1623621585
transform 1 0 5060 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_55
timestamp 1623621585
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_58
timestamp 1623621585
transform 1 0 6440 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_70
timestamp 1623621585
transform 1 0 7544 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_82
timestamp 1623621585
transform 1 0 8648 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_94
timestamp 1623621585
transform 1 0 9752 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1623621585
transform 1 0 11592 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_106
timestamp 1623621585
transform 1 0 10856 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_115
timestamp 1623621585
transform 1 0 11684 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_127
timestamp 1623621585
transform 1 0 12788 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_139
timestamp 1623621585
transform 1 0 13892 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_151
timestamp 1623621585
transform 1 0 14996 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_163
timestamp 1623621585
transform 1 0 16100 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1623621585
transform 1 0 16836 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_172
timestamp 1623621585
transform 1 0 16928 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_184
timestamp 1623621585
transform 1 0 18032 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_196
timestamp 1623621585
transform 1 0 19136 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_208
timestamp 1623621585
transform 1 0 20240 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1623621585
transform 1 0 22080 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_220
timestamp 1623621585
transform 1 0 21344 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_229
timestamp 1623621585
transform 1 0 22172 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_241
timestamp 1623621585
transform 1 0 23276 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1623621585
transform 1 0 24380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1623621585
transform 1 0 25484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1623621585
transform 1 0 27324 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_277
timestamp 1623621585
transform 1 0 26588 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_286
timestamp 1623621585
transform 1 0 27416 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_298
timestamp 1623621585
transform 1 0 28520 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_310
timestamp 1623621585
transform 1 0 29624 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_322
timestamp 1623621585
transform 1 0 30728 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1623621585
transform 1 0 32568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input479
timestamp 1623621585
transform 1 0 33580 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input509
timestamp 1623621585
transform 1 0 31924 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_334
timestamp 1623621585
transform 1 0 31832 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_338
timestamp 1623621585
transform 1 0 32200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_343
timestamp 1623621585
transform 1 0 32660 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_351
timestamp 1623621585
transform 1 0 33396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input89
timestamp 1623621585
transform 1 0 34500 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output706
timestamp 1623621585
transform 1 0 35144 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_356
timestamp 1623621585
transform 1 0 33856 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_362
timestamp 1623621585
transform 1 0 34408 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_366
timestamp 1623621585
transform 1 0 34776 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_374
timestamp 1623621585
transform 1 0 35512 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1623621585
transform 1 0 36432 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output660
timestamp 1623621585
transform 1 0 37076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_382
timestamp 1623621585
transform 1 0 36248 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_387
timestamp 1623621585
transform 1 0 36708 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_395
timestamp 1623621585
transform 1 0 37444 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1623621585
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1623621585
transform 1 0 37812 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_400
timestamp 1623621585
transform 1 0 37904 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1623621585
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1623621585
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input347
timestamp 1623621585
transform 1 0 1748 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output612
timestamp 1623621585
transform 1 0 2668 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1623621585
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1623621585
transform 1 0 2300 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1623621585
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_21
timestamp 1623621585
transform 1 0 3036 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_30
timestamp 1623621585
transform 1 0 3864 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_42
timestamp 1623621585
transform 1 0 4968 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_54
timestamp 1623621585
transform 1 0 6072 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_66
timestamp 1623621585
transform 1 0 7176 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_78
timestamp 1623621585
transform 1 0 8280 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1623621585
transform 1 0 9016 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_87
timestamp 1623621585
transform 1 0 9108 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_99
timestamp 1623621585
transform 1 0 10212 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_111
timestamp 1623621585
transform 1 0 11316 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1623621585
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1623621585
transform 1 0 14260 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_135
timestamp 1623621585
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_144
timestamp 1623621585
transform 1 0 14352 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_156
timestamp 1623621585
transform 1 0 15456 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_168
timestamp 1623621585
transform 1 0 16560 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_180
timestamp 1623621585
transform 1 0 17664 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1623621585
transform 1 0 19504 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_192
timestamp 1623621585
transform 1 0 18768 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_201
timestamp 1623621585
transform 1 0 19596 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_213
timestamp 1623621585
transform 1 0 20700 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1623621585
transform 1 0 21804 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1623621585
transform 1 0 22908 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_249
timestamp 1623621585
transform 1 0 24012 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1623621585
transform 1 0 24748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_258
timestamp 1623621585
transform 1 0 24840 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_270
timestamp 1623621585
transform 1 0 25944 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_282
timestamp 1623621585
transform 1 0 27048 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_294
timestamp 1623621585
transform 1 0 28152 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_306
timestamp 1623621585
transform 1 0 29256 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1623621585
transform 1 0 29992 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_315
timestamp 1623621585
transform 1 0 30084 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_327
timestamp 1623621585
transform 1 0 31188 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_339
timestamp 1623621585
transform 1 0 32292 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_351
timestamp 1623621585
transform 1 0 33396 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1623621585
transform 1 0 35236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input94
timestamp 1623621585
transform 1 0 34592 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_363
timestamp 1623621585
transform 1 0 34500 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_367
timestamp 1623621585
transform 1 0 34868 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_372
timestamp 1623621585
transform 1 0 35328 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1623621585
transform 1 0 37168 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input74
timestamp 1623621585
transform 1 0 36524 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input88
timestamp 1623621585
transform 1 0 35880 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_381
timestamp 1623621585
transform 1 0 36156 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1623621585
transform 1 0 36800 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_395
timestamp 1623621585
transform 1 0 37444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1623621585
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output657
timestamp 1623621585
transform 1 0 37812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1623621585
transform 1 0 38180 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1623621585
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1623621585
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input348
timestamp 1623621585
transform 1 0 1748 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1623621585
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_13
timestamp 1623621585
transform 1 0 2300 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1623621585
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1623621585
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _692_
timestamp 1623621585
transform 1 0 3036 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1623621585
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input525
timestamp 1623621585
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1623621585
transform 1 0 3312 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_31
timestamp 1623621585
transform 1 0 3956 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_27
timestamp 1623621585
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_30
timestamp 1623621585
transform 1 0 3864 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1623621585
transform 1 0 6348 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_43
timestamp 1623621585
transform 1 0 5060 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_55
timestamp 1623621585
transform 1 0 6164 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_58
timestamp 1623621585
transform 1 0 6440 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_42
timestamp 1623621585
transform 1 0 4968 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_54
timestamp 1623621585
transform 1 0 6072 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_70
timestamp 1623621585
transform 1 0 7544 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_82
timestamp 1623621585
transform 1 0 8648 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_66
timestamp 1623621585
transform 1 0 7176 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_78
timestamp 1623621585
transform 1 0 8280 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1623621585
transform 1 0 9016 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_94
timestamp 1623621585
transform 1 0 9752 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_87
timestamp 1623621585
transform 1 0 9108 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_99
timestamp 1623621585
transform 1 0 10212 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1623621585
transform 1 0 11592 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_106
timestamp 1623621585
transform 1 0 10856 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_115
timestamp 1623621585
transform 1 0 11684 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_111
timestamp 1623621585
transform 1 0 11316 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1623621585
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1623621585
transform 1 0 14260 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_127
timestamp 1623621585
transform 1 0 12788 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_139
timestamp 1623621585
transform 1 0 13892 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_135
timestamp 1623621585
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_144
timestamp 1623621585
transform 1 0 14352 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_151
timestamp 1623621585
transform 1 0 14996 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_163
timestamp 1623621585
transform 1 0 16100 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_156
timestamp 1623621585
transform 1 0 15456 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1623621585
transform 1 0 16836 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_172
timestamp 1623621585
transform 1 0 16928 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1623621585
transform 1 0 18032 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_168
timestamp 1623621585
transform 1 0 16560 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_180
timestamp 1623621585
transform 1 0 17664 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1623621585
transform 1 0 19504 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1623621585
transform 1 0 19136 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_208
timestamp 1623621585
transform 1 0 20240 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_192
timestamp 1623621585
transform 1 0 18768 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_201
timestamp 1623621585
transform 1 0 19596 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1623621585
transform 1 0 22080 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_220
timestamp 1623621585
transform 1 0 21344 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_229
timestamp 1623621585
transform 1 0 22172 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_213
timestamp 1623621585
transform 1 0 20700 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1623621585
transform 1 0 21804 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_241
timestamp 1623621585
transform 1 0 23276 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1623621585
transform 1 0 22908 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_249
timestamp 1623621585
transform 1 0 24012 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1623621585
transform 1 0 24748 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1623621585
transform 1 0 24380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1623621585
transform 1 0 25484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_258
timestamp 1623621585
transform 1 0 24840 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_270
timestamp 1623621585
transform 1 0 25944 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1623621585
transform 1 0 27324 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_277
timestamp 1623621585
transform 1 0 26588 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_286
timestamp 1623621585
transform 1 0 27416 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_282
timestamp 1623621585
transform 1 0 27048 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_298
timestamp 1623621585
transform 1 0 28520 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_310
timestamp 1623621585
transform 1 0 29624 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_294
timestamp 1623621585
transform 1 0 28152 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_306
timestamp 1623621585
transform 1 0 29256 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1623621585
transform 1 0 29992 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_322
timestamp 1623621585
transform 1 0 30728 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_315
timestamp 1623621585
transform 1 0 30084 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_327
timestamp 1623621585
transform 1 0 31188 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1623621585
transform 1 0 32568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_334
timestamp 1623621585
transform 1 0 31832 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_343
timestamp 1623621585
transform 1 0 32660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_339
timestamp 1623621585
transform 1 0 32292 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_351
timestamp 1623621585
transform 1 0 33396 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1623621585
transform 1 0 35236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input93
timestamp 1623621585
transform 1 0 35236 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input480
timestamp 1623621585
transform 1 0 34500 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_355
timestamp 1623621585
transform 1 0 33764 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_366
timestamp 1623621585
transform 1 0 34776 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_370
timestamp 1623621585
transform 1 0 35144 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_374
timestamp 1623621585
transform 1 0 35512 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_363
timestamp 1623621585
transform 1 0 34500 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_372
timestamp 1623621585
transform 1 0 35328 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input92
timestamp 1623621585
transform 1 0 35880 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_384
timestamp 1623621585
transform 1 0 36432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_381
timestamp 1623621585
transform 1 0 36156 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_389
timestamp 1623621585
transform 1 0 36892 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_388
timestamp 1623621585
transform 1 0 36800 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input91
timestamp 1623621585
transform 1 0 36616 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 1623621585
transform 1 0 36524 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1623621585
transform 1 0 37260 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1623621585
transform 1 0 37168 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_395
timestamp 1623621585
transform 1 0 37444 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1623621585
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1623621585
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1623621585
transform 1 0 37812 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1623621585
transform 1 0 37904 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_400
timestamp 1623621585
transform 1 0 37904 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_406
timestamp 1623621585
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_396
timestamp 1623621585
transform 1 0 37536 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1623621585
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1623621585
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input349
timestamp 1623621585
transform 1 0 1748 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1623621585
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_13
timestamp 1623621585
transform 1 0 2300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_25
timestamp 1623621585
transform 1 0 3404 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_37
timestamp 1623621585
transform 1 0 4508 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1623621585
transform 1 0 6348 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_49
timestamp 1623621585
transform 1 0 5612 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_58
timestamp 1623621585
transform 1 0 6440 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_70
timestamp 1623621585
transform 1 0 7544 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_82
timestamp 1623621585
transform 1 0 8648 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_94
timestamp 1623621585
transform 1 0 9752 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1623621585
transform 1 0 11592 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_106
timestamp 1623621585
transform 1 0 10856 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_115
timestamp 1623621585
transform 1 0 11684 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_127
timestamp 1623621585
transform 1 0 12788 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_139
timestamp 1623621585
transform 1 0 13892 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_151
timestamp 1623621585
transform 1 0 14996 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_163
timestamp 1623621585
transform 1 0 16100 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1623621585
transform 1 0 16836 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_172
timestamp 1623621585
transform 1 0 16928 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_184
timestamp 1623621585
transform 1 0 18032 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_196
timestamp 1623621585
transform 1 0 19136 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_208
timestamp 1623621585
transform 1 0 20240 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1623621585
transform 1 0 22080 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_220
timestamp 1623621585
transform 1 0 21344 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_229
timestamp 1623621585
transform 1 0 22172 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_8  _590_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 23552 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_8_241
timestamp 1623621585
transform 1 0 23276 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_257
timestamp 1623621585
transform 1 0 24748 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_269
timestamp 1623621585
transform 1 0 25852 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1623621585
transform 1 0 27324 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_281
timestamp 1623621585
transform 1 0 26956 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_286
timestamp 1623621585
transform 1 0 27416 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_298
timestamp 1623621585
transform 1 0 28520 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_310
timestamp 1623621585
transform 1 0 29624 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_322
timestamp 1623621585
transform 1 0 30728 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1623621585
transform 1 0 32568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_334
timestamp 1623621585
transform 1 0 31832 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_343
timestamp 1623621585
transform 1 0 32660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_355
timestamp 1623621585
transform 1 0 33764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_367
timestamp 1623621585
transform 1 0 34868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1623621585
transform 1 0 37168 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_379
timestamp 1623621585
transform 1 0 35972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_391
timestamp 1623621585
transform 1 0 37076 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_395
timestamp 1623621585
transform 1 0 37444 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1623621585
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1623621585
transform 1 0 37812 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_400
timestamp 1623621585
transform 1 0 37904 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_406
timestamp 1623621585
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1623621585
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input350
timestamp 1623621585
transform 1 0 1748 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1623621585
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_13
timestamp 1623621585
transform 1 0 2300 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1623621585
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_25
timestamp 1623621585
transform 1 0 3404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_30
timestamp 1623621585
transform 1 0 3864 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_42
timestamp 1623621585
transform 1 0 4968 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_54
timestamp 1623621585
transform 1 0 6072 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_66
timestamp 1623621585
transform 1 0 7176 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_78
timestamp 1623621585
transform 1 0 8280 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1623621585
transform 1 0 9016 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_87
timestamp 1623621585
transform 1 0 9108 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_99
timestamp 1623621585
transform 1 0 10212 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_111
timestamp 1623621585
transform 1 0 11316 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1623621585
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1623621585
transform 1 0 14260 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_135
timestamp 1623621585
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_144
timestamp 1623621585
transform 1 0 14352 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_156
timestamp 1623621585
transform 1 0 15456 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_168
timestamp 1623621585
transform 1 0 16560 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_180
timestamp 1623621585
transform 1 0 17664 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1623621585
transform 1 0 19504 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_192
timestamp 1623621585
transform 1 0 18768 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_201
timestamp 1623621585
transform 1 0 19596 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_213
timestamp 1623621585
transform 1 0 20700 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1623621585
transform 1 0 21804 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1623621585
transform 1 0 22908 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_249
timestamp 1623621585
transform 1 0 24012 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1623621585
transform 1 0 24748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_258
timestamp 1623621585
transform 1 0 24840 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_270
timestamp 1623621585
transform 1 0 25944 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_282
timestamp 1623621585
transform 1 0 27048 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_294
timestamp 1623621585
transform 1 0 28152 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_306
timestamp 1623621585
transform 1 0 29256 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1623621585
transform 1 0 29992 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_315
timestamp 1623621585
transform 1 0 30084 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_327
timestamp 1623621585
transform 1 0 31188 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_339
timestamp 1623621585
transform 1 0 32292 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_351
timestamp 1623621585
transform 1 0 33396 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1623621585
transform 1 0 35236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_363
timestamp 1623621585
transform 1 0 34500 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_372
timestamp 1623621585
transform 1 0 35328 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1623621585
transform 1 0 37260 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_384
timestamp 1623621585
transform 1 0 36432 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_392
timestamp 1623621585
transform 1 0 37168 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1623621585
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1623621585
transform 1 0 37904 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_396
timestamp 1623621585
transform 1 0 37536 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1623621585
transform 1 0 38180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1623621585
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1623621585
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1623621585
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_27
timestamp 1623621585
transform 1 0 3588 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1623621585
transform 1 0 4692 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1623621585
transform 1 0 6348 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_51
timestamp 1623621585
transform 1 0 5796 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_58
timestamp 1623621585
transform 1 0 6440 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_70
timestamp 1623621585
transform 1 0 7544 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_82
timestamp 1623621585
transform 1 0 8648 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_94
timestamp 1623621585
transform 1 0 9752 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1623621585
transform 1 0 11592 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_106
timestamp 1623621585
transform 1 0 10856 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_115
timestamp 1623621585
transform 1 0 11684 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_127
timestamp 1623621585
transform 1 0 12788 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_139
timestamp 1623621585
transform 1 0 13892 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_151
timestamp 1623621585
transform 1 0 14996 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_163
timestamp 1623621585
transform 1 0 16100 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1623621585
transform 1 0 16836 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_172
timestamp 1623621585
transform 1 0 16928 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_184
timestamp 1623621585
transform 1 0 18032 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_196
timestamp 1623621585
transform 1 0 19136 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_208
timestamp 1623621585
transform 1 0 20240 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1623621585
transform 1 0 22080 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_220
timestamp 1623621585
transform 1 0 21344 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_229
timestamp 1623621585
transform 1 0 22172 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_241
timestamp 1623621585
transform 1 0 23276 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1623621585
transform 1 0 24380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1623621585
transform 1 0 25484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1623621585
transform 1 0 27324 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_277
timestamp 1623621585
transform 1 0 26588 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_286
timestamp 1623621585
transform 1 0 27416 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__nor4_2  _621_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 29348 0 -1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_10_298
timestamp 1623621585
transform 1 0 28520 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_306
timestamp 1623621585
transform 1 0 29256 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_317
timestamp 1623621585
transform 1 0 30268 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_329
timestamp 1623621585
transform 1 0 31372 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1623621585
transform 1 0 32568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_341
timestamp 1623621585
transform 1 0 32476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_343
timestamp 1623621585
transform 1 0 32660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_355
timestamp 1623621585
transform 1 0 33764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_367
timestamp 1623621585
transform 1 0 34868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_379
timestamp 1623621585
transform 1 0 35972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_391
timestamp 1623621585
transform 1 0 37076 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1623621585
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1623621585
transform 1 0 37812 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_400
timestamp 1623621585
transform 1 0 37904 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_406
timestamp 1623621585
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1623621585
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input320
timestamp 1623621585
transform 1 0 1748 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1623621585
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_13
timestamp 1623621585
transform 1 0 2300 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1623621585
transform 1 0 3772 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_25
timestamp 1623621585
transform 1 0 3404 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_30
timestamp 1623621585
transform 1 0 3864 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_42
timestamp 1623621585
transform 1 0 4968 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_54
timestamp 1623621585
transform 1 0 6072 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_66
timestamp 1623621585
transform 1 0 7176 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_78
timestamp 1623621585
transform 1 0 8280 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1623621585
transform 1 0 9016 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_87
timestamp 1623621585
transform 1 0 9108 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_99
timestamp 1623621585
transform 1 0 10212 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_111
timestamp 1623621585
transform 1 0 11316 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1623621585
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1623621585
transform 1 0 14260 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_135
timestamp 1623621585
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_144
timestamp 1623621585
transform 1 0 14352 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_156
timestamp 1623621585
transform 1 0 15456 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_168
timestamp 1623621585
transform 1 0 16560 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_180
timestamp 1623621585
transform 1 0 17664 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1623621585
transform 1 0 19504 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_192
timestamp 1623621585
transform 1 0 18768 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_201
timestamp 1623621585
transform 1 0 19596 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_213
timestamp 1623621585
transform 1 0 20700 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1623621585
transform 1 0 21804 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1623621585
transform 1 0 22908 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_249
timestamp 1623621585
transform 1 0 24012 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1623621585
transform 1 0 24748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_258
timestamp 1623621585
transform 1 0 24840 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_270
timestamp 1623621585
transform 1 0 25944 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_282
timestamp 1623621585
transform 1 0 27048 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_294
timestamp 1623621585
transform 1 0 28152 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_306
timestamp 1623621585
transform 1 0 29256 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1623621585
transform 1 0 29992 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_315
timestamp 1623621585
transform 1 0 30084 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_327
timestamp 1623621585
transform 1 0 31188 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_339
timestamp 1623621585
transform 1 0 32292 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_351
timestamp 1623621585
transform 1 0 33396 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1623621585
transform 1 0 35236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_363
timestamp 1623621585
transform 1 0 34500 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_372
timestamp 1623621585
transform 1 0 35328 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1623621585
transform 1 0 37260 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_384
timestamp 1623621585
transform 1 0 36432 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_392
timestamp 1623621585
transform 1 0 37168 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1623621585
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1623621585
transform 1 0 37904 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_396
timestamp 1623621585
transform 1 0 37536 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1623621585
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1623621585
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input321
timestamp 1623621585
transform 1 0 1748 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1623621585
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_13
timestamp 1623621585
transform 1 0 2300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_25
timestamp 1623621585
transform 1 0 3404 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_37
timestamp 1623621585
transform 1 0 4508 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1623621585
transform 1 0 6348 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_49
timestamp 1623621585
transform 1 0 5612 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_58
timestamp 1623621585
transform 1 0 6440 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_70
timestamp 1623621585
transform 1 0 7544 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_82
timestamp 1623621585
transform 1 0 8648 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_94
timestamp 1623621585
transform 1 0 9752 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1623621585
transform 1 0 11592 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_106
timestamp 1623621585
transform 1 0 10856 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_115
timestamp 1623621585
transform 1 0 11684 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_127
timestamp 1623621585
transform 1 0 12788 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_139
timestamp 1623621585
transform 1 0 13892 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_151
timestamp 1623621585
transform 1 0 14996 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_163
timestamp 1623621585
transform 1 0 16100 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1623621585
transform 1 0 16836 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_172
timestamp 1623621585
transform 1 0 16928 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_184
timestamp 1623621585
transform 1 0 18032 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_196
timestamp 1623621585
transform 1 0 19136 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_208
timestamp 1623621585
transform 1 0 20240 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1623621585
transform 1 0 22080 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_220
timestamp 1623621585
transform 1 0 21344 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_229
timestamp 1623621585
transform 1 0 22172 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_241
timestamp 1623621585
transform 1 0 23276 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1623621585
transform 1 0 24380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1623621585
transform 1 0 25484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1623621585
transform 1 0 27324 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_277
timestamp 1623621585
transform 1 0 26588 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_286
timestamp 1623621585
transform 1 0 27416 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_298
timestamp 1623621585
transform 1 0 28520 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_310
timestamp 1623621585
transform 1 0 29624 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_322
timestamp 1623621585
transform 1 0 30728 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1623621585
transform 1 0 32568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_334
timestamp 1623621585
transform 1 0 31832 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_343
timestamp 1623621585
transform 1 0 32660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_355
timestamp 1623621585
transform 1 0 33764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_367
timestamp 1623621585
transform 1 0 34868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input75
timestamp 1623621585
transform 1 0 37168 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_379
timestamp 1623621585
transform 1 0 35972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_391
timestamp 1623621585
transform 1 0 37076 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_395
timestamp 1623621585
transform 1 0 37444 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1623621585
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1623621585
transform 1 0 37812 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_400
timestamp 1623621585
transform 1 0 37904 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_406
timestamp 1623621585
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1623621585
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1623621585
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input322
timestamp 1623621585
transform 1 0 1748 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1623621585
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1623621585
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1623621585
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_13
timestamp 1623621585
transform 1 0 2300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1623621585
transform 1 0 3772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_27
timestamp 1623621585
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_30
timestamp 1623621585
transform 1 0 3864 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_25
timestamp 1623621585
transform 1 0 3404 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_37
timestamp 1623621585
transform 1 0 4508 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1623621585
transform 1 0 6348 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_42
timestamp 1623621585
transform 1 0 4968 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_54
timestamp 1623621585
transform 1 0 6072 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_49
timestamp 1623621585
transform 1 0 5612 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_58
timestamp 1623621585
transform 1 0 6440 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_66
timestamp 1623621585
transform 1 0 7176 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_78
timestamp 1623621585
transform 1 0 8280 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_70
timestamp 1623621585
transform 1 0 7544 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_82
timestamp 1623621585
transform 1 0 8648 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1623621585
transform 1 0 9016 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_87
timestamp 1623621585
transform 1 0 9108 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_99
timestamp 1623621585
transform 1 0 10212 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_94
timestamp 1623621585
transform 1 0 9752 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1623621585
transform 1 0 11592 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_111
timestamp 1623621585
transform 1 0 11316 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1623621585
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_106
timestamp 1623621585
transform 1 0 10856 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_115
timestamp 1623621585
transform 1 0 11684 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1623621585
transform 1 0 14260 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_135
timestamp 1623621585
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_144
timestamp 1623621585
transform 1 0 14352 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_127
timestamp 1623621585
transform 1 0 12788 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_139
timestamp 1623621585
transform 1 0 13892 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_156
timestamp 1623621585
transform 1 0 15456 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_151
timestamp 1623621585
transform 1 0 14996 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_163
timestamp 1623621585
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1623621585
transform 1 0 16836 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_168
timestamp 1623621585
transform 1 0 16560 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_180
timestamp 1623621585
transform 1 0 17664 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_172
timestamp 1623621585
transform 1 0 16928 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_184
timestamp 1623621585
transform 1 0 18032 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1623621585
transform 1 0 19504 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_192
timestamp 1623621585
transform 1 0 18768 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_201
timestamp 1623621585
transform 1 0 19596 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_196
timestamp 1623621585
transform 1 0 19136 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_208
timestamp 1623621585
transform 1 0 20240 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1623621585
transform 1 0 22080 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_213
timestamp 1623621585
transform 1 0 20700 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1623621585
transform 1 0 21804 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_220
timestamp 1623621585
transform 1 0 21344 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_229
timestamp 1623621585
transform 1 0 22172 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1623621585
transform 1 0 22908 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_249
timestamp 1623621585
transform 1 0 24012 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_241
timestamp 1623621585
transform 1 0 23276 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1623621585
transform 1 0 24748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_258
timestamp 1623621585
transform 1 0 24840 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_270
timestamp 1623621585
transform 1 0 25944 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1623621585
transform 1 0 24380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1623621585
transform 1 0 25484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1623621585
transform 1 0 27324 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_282
timestamp 1623621585
transform 1 0 27048 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_277
timestamp 1623621585
transform 1 0 26588 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_286
timestamp 1623621585
transform 1 0 27416 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_294
timestamp 1623621585
transform 1 0 28152 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_306
timestamp 1623621585
transform 1 0 29256 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_298
timestamp 1623621585
transform 1 0 28520 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_310
timestamp 1623621585
transform 1 0 29624 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _709_
timestamp 1623621585
transform 1 0 30360 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1623621585
transform 1 0 29992 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_315
timestamp 1623621585
transform 1 0 30084 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_327
timestamp 1623621585
transform 1 0 31188 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1623621585
transform 1 0 30636 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_333
timestamp 1623621585
transform 1 0 31740 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1623621585
transform 1 0 32568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_339
timestamp 1623621585
transform 1 0 32292 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_351
timestamp 1623621585
transform 1 0 33396 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_341
timestamp 1623621585
transform 1 0 32476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_343
timestamp 1623621585
transform 1 0 32660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1623621585
transform 1 0 35236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_363
timestamp 1623621585
transform 1 0 34500 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_372
timestamp 1623621585
transform 1 0 35328 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_355
timestamp 1623621585
transform 1 0 33764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_367
timestamp 1623621585
transform 1 0 34868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input76
timestamp 1623621585
transform 1 0 37260 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_384
timestamp 1623621585
transform 1 0 36432 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_392
timestamp 1623621585
transform 1 0 37168 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_379
timestamp 1623621585
transform 1 0 35972 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_391
timestamp 1623621585
transform 1 0 37076 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1623621585
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1623621585
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1623621585
transform 1 0 37812 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1623621585
transform 1 0 37904 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_396
timestamp 1623621585
transform 1 0 37536 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1623621585
transform 1 0 38180 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_400
timestamp 1623621585
transform 1 0 37904 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1623621585
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1623621585
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input323
timestamp 1623621585
transform 1 0 1748 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1623621585
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_13
timestamp 1623621585
transform 1 0 2300 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1623621585
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_25
timestamp 1623621585
transform 1 0 3404 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_30
timestamp 1623621585
transform 1 0 3864 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_42
timestamp 1623621585
transform 1 0 4968 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_54
timestamp 1623621585
transform 1 0 6072 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_66
timestamp 1623621585
transform 1 0 7176 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_78
timestamp 1623621585
transform 1 0 8280 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1623621585
transform 1 0 9016 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_87
timestamp 1623621585
transform 1 0 9108 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_99
timestamp 1623621585
transform 1 0 10212 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_111
timestamp 1623621585
transform 1 0 11316 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1623621585
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1623621585
transform 1 0 14260 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_135
timestamp 1623621585
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_144
timestamp 1623621585
transform 1 0 14352 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_156
timestamp 1623621585
transform 1 0 15456 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_168
timestamp 1623621585
transform 1 0 16560 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_180
timestamp 1623621585
transform 1 0 17664 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1623621585
transform 1 0 19504 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_192
timestamp 1623621585
transform 1 0 18768 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_201
timestamp 1623621585
transform 1 0 19596 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_213
timestamp 1623621585
transform 1 0 20700 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1623621585
transform 1 0 21804 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1623621585
transform 1 0 22908 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_249
timestamp 1623621585
transform 1 0 24012 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1623621585
transform 1 0 24748 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_258
timestamp 1623621585
transform 1 0 24840 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_270
timestamp 1623621585
transform 1 0 25944 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_282
timestamp 1623621585
transform 1 0 27048 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_294
timestamp 1623621585
transform 1 0 28152 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_306
timestamp 1623621585
transform 1 0 29256 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1623621585
transform 1 0 29992 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_315
timestamp 1623621585
transform 1 0 30084 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_327
timestamp 1623621585
transform 1 0 31188 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_339
timestamp 1623621585
transform 1 0 32292 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_351
timestamp 1623621585
transform 1 0 33396 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1623621585
transform 1 0 35236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_363
timestamp 1623621585
transform 1 0 34500 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_372
timestamp 1623621585
transform 1 0 35328 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input78
timestamp 1623621585
transform 1 0 37260 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_384
timestamp 1623621585
transform 1 0 36432 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_392
timestamp 1623621585
transform 1 0 37168 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1623621585
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input77
timestamp 1623621585
transform 1 0 37904 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_396
timestamp 1623621585
transform 1 0 37536 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1623621585
transform 1 0 38180 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1623621585
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1623621585
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1623621585
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_27
timestamp 1623621585
transform 1 0 3588 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_39
timestamp 1623621585
transform 1 0 4692 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1623621585
transform 1 0 6348 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_51
timestamp 1623621585
transform 1 0 5796 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_58
timestamp 1623621585
transform 1 0 6440 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_70
timestamp 1623621585
transform 1 0 7544 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_82
timestamp 1623621585
transform 1 0 8648 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_94
timestamp 1623621585
transform 1 0 9752 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1623621585
transform 1 0 11592 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_106
timestamp 1623621585
transform 1 0 10856 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_115
timestamp 1623621585
transform 1 0 11684 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_127
timestamp 1623621585
transform 1 0 12788 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_139
timestamp 1623621585
transform 1 0 13892 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_151
timestamp 1623621585
transform 1 0 14996 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_163
timestamp 1623621585
transform 1 0 16100 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1623621585
transform 1 0 16836 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_172
timestamp 1623621585
transform 1 0 16928 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_184
timestamp 1623621585
transform 1 0 18032 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_196
timestamp 1623621585
transform 1 0 19136 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_208
timestamp 1623621585
transform 1 0 20240 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1623621585
transform 1 0 22080 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_220
timestamp 1623621585
transform 1 0 21344 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1623621585
transform 1 0 22172 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _776_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 22540 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_16_250
timestamp 1623621585
transform 1 0 24104 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_262
timestamp 1623621585
transform 1 0 25208 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1623621585
transform 1 0 27324 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_274
timestamp 1623621585
transform 1 0 26312 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_282
timestamp 1623621585
transform 1 0 27048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_286
timestamp 1623621585
transform 1 0 27416 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_298
timestamp 1623621585
transform 1 0 28520 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_310
timestamp 1623621585
transform 1 0 29624 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_1  _609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 30728 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_330
timestamp 1623621585
transform 1 0 31464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1623621585
transform 1 0 32568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_343
timestamp 1623621585
transform 1 0 32660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_355
timestamp 1623621585
transform 1 0 33764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_367
timestamp 1623621585
transform 1 0 34868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input80
timestamp 1623621585
transform 1 0 37168 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_379
timestamp 1623621585
transform 1 0 35972 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_391
timestamp 1623621585
transform 1 0 37076 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_395
timestamp 1623621585
transform 1 0 37444 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1623621585
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1623621585
transform 1 0 37812 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_400
timestamp 1623621585
transform 1 0 37904 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_406
timestamp 1623621585
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1623621585
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input324
timestamp 1623621585
transform 1 0 1748 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1623621585
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_13
timestamp 1623621585
transform 1 0 2300 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1623621585
transform 1 0 3772 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_25
timestamp 1623621585
transform 1 0 3404 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_30
timestamp 1623621585
transform 1 0 3864 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_42
timestamp 1623621585
transform 1 0 4968 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_54
timestamp 1623621585
transform 1 0 6072 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_66
timestamp 1623621585
transform 1 0 7176 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_78
timestamp 1623621585
transform 1 0 8280 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1623621585
transform 1 0 9016 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_87
timestamp 1623621585
transform 1 0 9108 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_99
timestamp 1623621585
transform 1 0 10212 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_111
timestamp 1623621585
transform 1 0 11316 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1623621585
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1623621585
transform 1 0 14260 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_135
timestamp 1623621585
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_144
timestamp 1623621585
transform 1 0 14352 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_156
timestamp 1623621585
transform 1 0 15456 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_168
timestamp 1623621585
transform 1 0 16560 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_180
timestamp 1623621585
transform 1 0 17664 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1623621585
transform 1 0 19504 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_192
timestamp 1623621585
transform 1 0 18768 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_201
timestamp 1623621585
transform 1 0 19596 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_213
timestamp 1623621585
transform 1 0 20700 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_225
timestamp 1623621585
transform 1 0 21804 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_229
timestamp 1623621585
transform 1 0 22172 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _775_
timestamp 1623621585
transform 1 0 22264 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_17_247
timestamp 1623621585
transform 1 0 23828 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1623621585
transform 1 0 24748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_255
timestamp 1623621585
transform 1 0 24564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_258
timestamp 1623621585
transform 1 0 24840 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_270
timestamp 1623621585
transform 1 0 25944 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_282
timestamp 1623621585
transform 1 0 27048 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_294
timestamp 1623621585
transform 1 0 28152 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_306
timestamp 1623621585
transform 1 0 29256 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1623621585
transform 1 0 29992 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_315
timestamp 1623621585
transform 1 0 30084 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_327
timestamp 1623621585
transform 1 0 31188 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_339
timestamp 1623621585
transform 1 0 32292 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_351
timestamp 1623621585
transform 1 0 33396 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1623621585
transform 1 0 35236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_363
timestamp 1623621585
transform 1 0 34500 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_372
timestamp 1623621585
transform 1 0 35328 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 1623621585
transform 1 0 37260 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_384
timestamp 1623621585
transform 1 0 36432 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_392
timestamp 1623621585
transform 1 0 37168 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1623621585
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input79
timestamp 1623621585
transform 1 0 37904 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_396
timestamp 1623621585
transform 1 0 37536 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_403
timestamp 1623621585
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1623621585
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input325
timestamp 1623621585
transform 1 0 1748 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1623621585
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_13
timestamp 1623621585
transform 1 0 2300 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_25
timestamp 1623621585
transform 1 0 3404 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_37
timestamp 1623621585
transform 1 0 4508 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1623621585
transform 1 0 6348 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_49
timestamp 1623621585
transform 1 0 5612 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_58
timestamp 1623621585
transform 1 0 6440 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_70
timestamp 1623621585
transform 1 0 7544 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_82
timestamp 1623621585
transform 1 0 8648 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_94
timestamp 1623621585
transform 1 0 9752 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1623621585
transform 1 0 11592 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_106
timestamp 1623621585
transform 1 0 10856 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_115
timestamp 1623621585
transform 1 0 11684 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_127
timestamp 1623621585
transform 1 0 12788 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_139
timestamp 1623621585
transform 1 0 13892 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_151
timestamp 1623621585
transform 1 0 14996 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_163
timestamp 1623621585
transform 1 0 16100 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1623621585
transform 1 0 16836 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_172
timestamp 1623621585
transform 1 0 16928 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_184
timestamp 1623621585
transform 1 0 18032 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_196
timestamp 1623621585
transform 1 0 19136 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_208
timestamp 1623621585
transform 1 0 20240 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1623621585
transform 1 0 22080 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_220
timestamp 1623621585
transform 1 0 21344 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_229
timestamp 1623621585
transform 1 0 22172 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _773_
timestamp 1623621585
transform 1 0 22540 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_18_250
timestamp 1623621585
transform 1 0 24104 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _777_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 24472 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_270
timestamp 1623621585
transform 1 0 25944 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1623621585
transform 1 0 27324 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_wb_clk_i
timestamp 1623621585
transform 1 0 26312 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_277
timestamp 1623621585
transform 1 0 26588 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_286
timestamp 1623621585
transform 1 0 27416 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_298
timestamp 1623621585
transform 1 0 28520 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_310
timestamp 1623621585
transform 1 0 29624 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_322
timestamp 1623621585
transform 1 0 30728 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1623621585
transform 1 0 32568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_334
timestamp 1623621585
transform 1 0 31832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_343
timestamp 1623621585
transform 1 0 32660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_355
timestamp 1623621585
transform 1 0 33764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_367
timestamp 1623621585
transform 1 0 34868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_379
timestamp 1623621585
transform 1 0 35972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_391
timestamp 1623621585
transform 1 0 37076 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1623621585
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1623621585
transform 1 0 37812 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_400
timestamp 1623621585
transform 1 0 37904 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1623621585
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1623621585
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1623621585
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input326
timestamp 1623621585
transform 1 0 1748 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1623621585
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1623621585
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1623621585
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_13
timestamp 1623621585
transform 1 0 2300 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1623621585
transform 1 0 3772 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_27
timestamp 1623621585
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_30
timestamp 1623621585
transform 1 0 3864 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_25
timestamp 1623621585
transform 1 0 3404 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_37
timestamp 1623621585
transform 1 0 4508 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1623621585
transform 1 0 6348 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_42
timestamp 1623621585
transform 1 0 4968 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_54
timestamp 1623621585
transform 1 0 6072 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_49
timestamp 1623621585
transform 1 0 5612 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_58
timestamp 1623621585
transform 1 0 6440 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_66
timestamp 1623621585
transform 1 0 7176 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_78
timestamp 1623621585
transform 1 0 8280 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_70
timestamp 1623621585
transform 1 0 7544 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_82
timestamp 1623621585
transform 1 0 8648 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1623621585
transform 1 0 9016 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_87
timestamp 1623621585
transform 1 0 9108 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_99
timestamp 1623621585
transform 1 0 10212 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_94
timestamp 1623621585
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1623621585
transform 1 0 11592 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_111
timestamp 1623621585
transform 1 0 11316 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1623621585
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_106
timestamp 1623621585
transform 1 0 10856 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_115
timestamp 1623621585
transform 1 0 11684 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1623621585
transform 1 0 14260 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_135
timestamp 1623621585
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_144
timestamp 1623621585
transform 1 0 14352 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_127
timestamp 1623621585
transform 1 0 12788 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_139
timestamp 1623621585
transform 1 0 13892 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_156
timestamp 1623621585
transform 1 0 15456 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_151
timestamp 1623621585
transform 1 0 14996 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_163
timestamp 1623621585
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1623621585
transform 1 0 16836 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_168
timestamp 1623621585
transform 1 0 16560 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_180
timestamp 1623621585
transform 1 0 17664 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_172
timestamp 1623621585
transform 1 0 16928 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_184
timestamp 1623621585
transform 1 0 18032 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1623621585
transform 1 0 19504 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_192
timestamp 1623621585
transform 1 0 18768 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_201
timestamp 1623621585
transform 1 0 19596 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_196
timestamp 1623621585
transform 1 0 19136 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_208
timestamp 1623621585
transform 1 0 20240 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_1  _622_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 20884 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _772_
timestamp 1623621585
transform 1 0 21988 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1623621585
transform 1 0 22080 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_213
timestamp 1623621585
transform 1 0 20700 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_223
timestamp 1623621585
transform 1 0 21620 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_220
timestamp 1623621585
transform 1 0 21344 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_229
timestamp 1623621585
transform 1 0 22172 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _774_
timestamp 1623621585
transform 1 0 22540 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_19_244
timestamp 1623621585
transform 1 0 23552 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_250
timestamp 1623621585
transform 1 0 24104 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _779_
timestamp 1623621585
transform 1 0 24472 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _780_
timestamp 1623621585
transform 1 0 25208 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1623621585
transform 1 0 24748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_256
timestamp 1623621585
transform 1 0 24656 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_258
timestamp 1623621585
transform 1 0 24840 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_270
timestamp 1623621585
transform 1 0 25944 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _552_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 26312 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _564_
timestamp 1623621585
transform 1 0 27048 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _789_
timestamp 1623621585
transform 1 0 27784 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1623621585
transform 1 0 27324 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_278
timestamp 1623621585
transform 1 0 26680 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_289
timestamp 1623621585
transform 1 0 27692 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_281
timestamp 1623621585
transform 1 0 26956 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_286
timestamp 1623621585
transform 1 0 27416 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _548_
timestamp 1623621585
transform 1 0 28612 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_297
timestamp 1623621585
transform 1 0 28428 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_303
timestamp 1623621585
transform 1 0 28980 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_311
timestamp 1623621585
transform 1 0 29716 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_306
timestamp 1623621585
transform 1 0 29256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1623621585
transform 1 0 29992 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_315
timestamp 1623621585
transform 1 0 30084 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_327
timestamp 1623621585
transform 1 0 31188 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_318
timestamp 1623621585
transform 1 0 30360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_330
timestamp 1623621585
transform 1 0 31464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1623621585
transform 1 0 32568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_339
timestamp 1623621585
transform 1 0 32292 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_351
timestamp 1623621585
transform 1 0 33396 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_343
timestamp 1623621585
transform 1 0 32660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1623621585
transform 1 0 35236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_363
timestamp 1623621585
transform 1 0 34500 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_372
timestamp 1623621585
transform 1 0 35328 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_355
timestamp 1623621585
transform 1 0 33764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_367
timestamp 1623621585
transform 1 0 34868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 1623621585
transform 1 0 37260 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1623621585
transform 1 0 37168 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_384
timestamp 1623621585
transform 1 0 36432 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_392
timestamp 1623621585
transform 1 0 37168 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_379
timestamp 1623621585
transform 1 0 35972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_391
timestamp 1623621585
transform 1 0 37076 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_395
timestamp 1623621585
transform 1 0 37444 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1623621585
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1623621585
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1623621585
transform 1 0 37812 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input82
timestamp 1623621585
transform 1 0 37904 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_396
timestamp 1623621585
transform 1 0 37536 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_403
timestamp 1623621585
transform 1 0 38180 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_400
timestamp 1623621585
transform 1 0 37904 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_406
timestamp 1623621585
transform 1 0 38456 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1623621585
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input327
timestamp 1623621585
transform 1 0 1748 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1623621585
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_13
timestamp 1623621585
transform 1 0 2300 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1623621585
transform 1 0 3772 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_25
timestamp 1623621585
transform 1 0 3404 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_30
timestamp 1623621585
transform 1 0 3864 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_42
timestamp 1623621585
transform 1 0 4968 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_54
timestamp 1623621585
transform 1 0 6072 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_66
timestamp 1623621585
transform 1 0 7176 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_78
timestamp 1623621585
transform 1 0 8280 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1623621585
transform 1 0 9016 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_87
timestamp 1623621585
transform 1 0 9108 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_99
timestamp 1623621585
transform 1 0 10212 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_111
timestamp 1623621585
transform 1 0 11316 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1623621585
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1623621585
transform 1 0 14260 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_135
timestamp 1623621585
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_144
timestamp 1623621585
transform 1 0 14352 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_156
timestamp 1623621585
transform 1 0 15456 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_168
timestamp 1623621585
transform 1 0 16560 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_180
timestamp 1623621585
transform 1 0 17664 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1623621585
transform 1 0 19504 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_192
timestamp 1623621585
transform 1 0 18768 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_201
timestamp 1623621585
transform 1 0 19596 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_213
timestamp 1623621585
transform 1 0 20700 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1623621585
transform 1 0 21804 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _778_
timestamp 1623621585
transform 1 0 22908 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _782_
timestamp 1623621585
transform 1 0 25208 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1623621585
transform 1 0 24748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_253
timestamp 1623621585
transform 1 0 24380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_258
timestamp 1623621585
transform 1 0 24840 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _784_
timestamp 1623621585
transform 1 0 27048 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_278
timestamp 1623621585
transform 1 0 26680 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _623_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 28888 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_21_298
timestamp 1623621585
transform 1 0 28520 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_307
timestamp 1623621585
transform 1 0 29348 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1623621585
transform 1 0 29992 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_313
timestamp 1623621585
transform 1 0 29900 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_315
timestamp 1623621585
transform 1 0 30084 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_327
timestamp 1623621585
transform 1 0 31188 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_1  _557_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 32844 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_21_339
timestamp 1623621585
transform 1 0 32292 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_352
timestamp 1623621585
transform 1 0 33488 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _491_
timestamp 1623621585
transform 1 0 33948 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _531_
timestamp 1623621585
transform 1 0 34592 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1623621585
transform 1 0 35236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_356
timestamp 1623621585
transform 1 0 33856 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_360
timestamp 1623621585
transform 1 0 34224 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_367
timestamp 1623621585
transform 1 0 34868 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_372
timestamp 1623621585
transform 1 0 35328 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input87
timestamp 1623621585
transform 1 0 37260 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_384
timestamp 1623621585
transform 1 0 36432 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_392
timestamp 1623621585
transform 1 0 37168 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1623621585
transform -1 0 38824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input84
timestamp 1623621585
transform 1 0 37904 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_396
timestamp 1623621585
transform 1 0 37536 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_403
timestamp 1623621585
transform 1 0 38180 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1623621585
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input328
timestamp 1623621585
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1623621585
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_11
timestamp 1623621585
transform 1 0 2116 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_23
timestamp 1623621585
transform 1 0 3220 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_35
timestamp 1623621585
transform 1 0 4324 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1623621585
transform 1 0 6348 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_47
timestamp 1623621585
transform 1 0 5428 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_55
timestamp 1623621585
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_58
timestamp 1623621585
transform 1 0 6440 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_70
timestamp 1623621585
transform 1 0 7544 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_82
timestamp 1623621585
transform 1 0 8648 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1623621585
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1623621585
transform 1 0 11592 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_106
timestamp 1623621585
transform 1 0 10856 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_115
timestamp 1623621585
transform 1 0 11684 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_127
timestamp 1623621585
transform 1 0 12788 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_139
timestamp 1623621585
transform 1 0 13892 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_151
timestamp 1623621585
transform 1 0 14996 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_163
timestamp 1623621585
transform 1 0 16100 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1623621585
transform 1 0 16836 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_172
timestamp 1623621585
transform 1 0 16928 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_184
timestamp 1623621585
transform 1 0 18032 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_196
timestamp 1623621585
transform 1 0 19136 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_208
timestamp 1623621585
transform 1 0 20240 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1623621585
transform 1 0 22080 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_220
timestamp 1623621585
transform 1 0 21344 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_229
timestamp 1623621585
transform 1 0 22172 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1623621585
transform 1 0 23368 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _781_
timestamp 1623621585
transform 1 0 24012 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_241
timestamp 1623621585
transform 1 0 23276 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_245
timestamp 1623621585
transform 1 0 23644 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_265
timestamp 1623621585
transform 1 0 25484 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _525_
timestamp 1623621585
transform 1 0 26312 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _786_
timestamp 1623621585
transform 1 0 27784 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1623621585
transform 1 0 27324 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_273
timestamp 1623621585
transform 1 0 26220 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_281
timestamp 1623621585
transform 1 0 26956 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_286
timestamp 1623621585
transform 1 0 27416 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _508_
timestamp 1623621585
transform 1 0 29624 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_306
timestamp 1623621585
transform 1 0 29256 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_314
timestamp 1623621585
transform 1 0 29992 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_326
timestamp 1623621585
transform 1 0 31096 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_1  _544_
timestamp 1623621585
transform 1 0 33028 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1623621585
transform 1 0 32568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_338
timestamp 1623621585
transform 1 0 32200 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_343
timestamp 1623621585
transform 1 0 32660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_354
timestamp 1623621585
transform 1 0 33672 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _563_
timestamp 1623621585
transform 1 0 34040 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1623621585
transform 1 0 34684 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input159
timestamp 1623621585
transform 1 0 37168 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1623621585
transform 1 0 35788 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_389
timestamp 1623621585
transform 1 0 36892 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_395
timestamp 1623621585
transform 1 0 37444 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1623621585
transform -1 0 38824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1623621585
transform 1 0 37812 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_400
timestamp 1623621585
transform 1 0 37904 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_406
timestamp 1623621585
transform 1 0 38456 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1623621585
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1623621585
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1623621585
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1623621585
transform 1 0 3772 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_27
timestamp 1623621585
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_30
timestamp 1623621585
transform 1 0 3864 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_42
timestamp 1623621585
transform 1 0 4968 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_54
timestamp 1623621585
transform 1 0 6072 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_66
timestamp 1623621585
transform 1 0 7176 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_78
timestamp 1623621585
transform 1 0 8280 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1623621585
transform 1 0 9016 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_87
timestamp 1623621585
transform 1 0 9108 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_99
timestamp 1623621585
transform 1 0 10212 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_111
timestamp 1623621585
transform 1 0 11316 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1623621585
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1623621585
transform 1 0 14260 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_135
timestamp 1623621585
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_144
timestamp 1623621585
transform 1 0 14352 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_156
timestamp 1623621585
transform 1 0 15456 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_168
timestamp 1623621585
transform 1 0 16560 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_180
timestamp 1623621585
transform 1 0 17664 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1623621585
transform 1 0 19504 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_192
timestamp 1623621585
transform 1 0 18768 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_201
timestamp 1623621585
transform 1 0 19596 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_213
timestamp 1623621585
transform 1 0 20700 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1623621585
transform 1 0 21804 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _558_
timestamp 1623621585
transform 1 0 23736 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _576_
timestamp 1623621585
transform 1 0 22724 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_23_233
timestamp 1623621585
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_242
timestamp 1623621585
transform 1 0 23368 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _783_
timestamp 1623621585
transform 1 0 25208 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1623621585
transform 1 0 24748 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_253
timestamp 1623621585
transform 1 0 24380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_258
timestamp 1623621585
transform 1 0 24840 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_8  _605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 27140 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_278
timestamp 1623621585
transform 1 0 26680 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_282
timestamp 1623621585
transform 1 0 27048 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _485_
timestamp 1623621585
transform 1 0 28980 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_299
timestamp 1623621585
transform 1 0 28612 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_310
timestamp 1623621585
transform 1 0 29624 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1623621585
transform 1 0 29992 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_315
timestamp 1623621585
transform 1 0 30084 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_327
timestamp 1623621585
transform 1 0 31188 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _538_
timestamp 1623621585
transform 1 0 32936 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _551_
timestamp 1623621585
transform 1 0 31924 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_342
timestamp 1623621585
transform 1 0 32568 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_353
timestamp 1623621585
transform 1 0 33580 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _569_
timestamp 1623621585
transform 1 0 33948 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1623621585
transform 1 0 35236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_364
timestamp 1623621585
transform 1 0 34592 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_370
timestamp 1623621585
transform 1 0 35144 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_372
timestamp 1623621585
transform 1 0 35328 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _366_
timestamp 1623621585
transform 1 0 35696 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_380
timestamp 1623621585
transform 1 0 36064 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_392
timestamp 1623621585
transform 1 0 37168 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1623621585
transform -1 0 38824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input95
timestamp 1623621585
transform 1 0 37904 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1623621585
transform 1 0 38180 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1623621585
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input329
timestamp 1623621585
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1623621585
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_11
timestamp 1623621585
transform 1 0 2116 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_23
timestamp 1623621585
transform 1 0 3220 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_35
timestamp 1623621585
transform 1 0 4324 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1623621585
transform 1 0 6348 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_47
timestamp 1623621585
transform 1 0 5428 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_55
timestamp 1623621585
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_58
timestamp 1623621585
transform 1 0 6440 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_70
timestamp 1623621585
transform 1 0 7544 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_82
timestamp 1623621585
transform 1 0 8648 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_94
timestamp 1623621585
transform 1 0 9752 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1623621585
transform 1 0 11592 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_106
timestamp 1623621585
transform 1 0 10856 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_115
timestamp 1623621585
transform 1 0 11684 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_127
timestamp 1623621585
transform 1 0 12788 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_139
timestamp 1623621585
transform 1 0 13892 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_151
timestamp 1623621585
transform 1 0 14996 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_163
timestamp 1623621585
transform 1 0 16100 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1623621585
transform 1 0 16836 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_172
timestamp 1623621585
transform 1 0 16928 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_184
timestamp 1623621585
transform 1 0 18032 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_196
timestamp 1623621585
transform 1 0 19136 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_208
timestamp 1623621585
transform 1 0 20240 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1623621585
transform 1 0 22080 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_220
timestamp 1623621585
transform 1 0 21344 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_229
timestamp 1623621585
transform 1 0 22172 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _545_
timestamp 1623621585
transform 1 0 23368 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_wb_clk_i
timestamp 1623621585
transform 1 0 22724 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_238
timestamp 1623621585
transform 1 0 23000 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_249
timestamp 1623621585
transform 1 0 24012 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _539_
timestamp 1623621585
transform 1 0 24380 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _785_
timestamp 1623621585
transform 1 0 25392 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_260
timestamp 1623621585
transform 1 0 25024 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _787_
timestamp 1623621585
transform 1 0 27784 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1623621585
transform 1 0 27324 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_280
timestamp 1623621585
transform 1 0 26864 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_284
timestamp 1623621585
transform 1 0 27232 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_286
timestamp 1623621585
transform 1 0 27416 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _499_
timestamp 1623621585
transform 1 0 29624 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_306
timestamp 1623621585
transform 1 0 29256 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _570_
timestamp 1623621585
transform 1 0 30636 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_317
timestamp 1623621585
transform 1 0 30268 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_328
timestamp 1623621585
transform 1 0 31280 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_1  _524_
timestamp 1623621585
transform 1 0 33120 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1623621585
transform 1 0 32568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_340
timestamp 1623621585
transform 1 0 32384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_343
timestamp 1623621585
transform 1 0 32660 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_347
timestamp 1623621585
transform 1 0 33028 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_1  _575_
timestamp 1623621585
transform 1 0 34132 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_355
timestamp 1623621585
transform 1 0 33764 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_366
timestamp 1623621585
transform 1 0 34776 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input127
timestamp 1623621585
transform 1 0 37168 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_378
timestamp 1623621585
transform 1 0 35880 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_390
timestamp 1623621585
transform 1 0 36984 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_395
timestamp 1623621585
transform 1 0 37444 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1623621585
transform -1 0 38824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1623621585
transform 1 0 37812 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_400
timestamp 1623621585
transform 1 0 37904 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_406
timestamp 1623621585
transform 1 0 38456 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1623621585
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input331
timestamp 1623621585
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1623621585
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_11
timestamp 1623621585
transform 1 0 2116 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1623621585
transform 1 0 3772 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_23
timestamp 1623621585
transform 1 0 3220 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_30
timestamp 1623621585
transform 1 0 3864 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_42
timestamp 1623621585
transform 1 0 4968 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_54
timestamp 1623621585
transform 1 0 6072 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_66
timestamp 1623621585
transform 1 0 7176 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_78
timestamp 1623621585
transform 1 0 8280 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1623621585
transform 1 0 9016 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_87
timestamp 1623621585
transform 1 0 9108 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_99
timestamp 1623621585
transform 1 0 10212 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_111
timestamp 1623621585
transform 1 0 11316 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1623621585
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1623621585
transform 1 0 14260 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1623621585
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_144
timestamp 1623621585
transform 1 0 14352 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_156
timestamp 1623621585
transform 1 0 15456 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_168
timestamp 1623621585
transform 1 0 16560 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_180
timestamp 1623621585
transform 1 0 17664 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1623621585
transform 1 0 19504 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_192
timestamp 1623621585
transform 1 0 18768 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_201
timestamp 1623621585
transform 1 0 19596 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_213
timestamp 1623621585
transform 1 0 20700 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1623621585
transform 1 0 21804 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _763_
timestamp 1623621585
transform 1 0 22540 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_25_249
timestamp 1623621585
transform 1 0 24012 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _808_
timestamp 1623621585
transform 1 0 25576 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1623621585
transform 1 0 24748 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_258
timestamp 1623621585
transform 1 0 24840 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _788_
timestamp 1623621585
transform 1 0 27508 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_283
timestamp 1623621585
transform 1 0 27140 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _306_
timestamp 1623621585
transform 1 0 29348 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_303
timestamp 1623621585
transform 1 0 28980 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_310
timestamp 1623621585
transform 1 0 29624 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _338_
timestamp 1623621585
transform 1 0 31464 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _505_
timestamp 1623621585
transform 1 0 30452 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1623621585
transform 1 0 29992 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_315
timestamp 1623621585
transform 1 0 30084 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_326
timestamp 1623621585
transform 1 0 31096 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _511_
timestamp 1623621585
transform 1 0 33212 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _581_
timestamp 1623621585
transform 1 0 32200 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_25_334
timestamp 1623621585
transform 1 0 31832 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_345
timestamp 1623621585
transform 1 0 32844 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _451_
timestamp 1623621585
transform 1 0 34224 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1623621585
transform 1 0 35236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_356
timestamp 1623621585
transform 1 0 33856 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_364
timestamp 1623621585
transform 1 0 34592 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_370
timestamp 1623621585
transform 1 0 35144 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_372
timestamp 1623621585
transform 1 0 35328 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input170
timestamp 1623621585
transform 1 0 37260 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_384
timestamp 1623621585
transform 1 0 36432 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_392
timestamp 1623621585
transform 1 0 37168 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1623621585
transform -1 0 38824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input106
timestamp 1623621585
transform 1 0 37904 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_396
timestamp 1623621585
transform 1 0 37536 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_403
timestamp 1623621585
transform 1 0 38180 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1623621585
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1623621585
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input332
timestamp 1623621585
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1623621585
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1623621585
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1623621585
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1623621585
transform 1 0 2116 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1623621585
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_27
timestamp 1623621585
transform 1 0 3588 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_39
timestamp 1623621585
transform 1 0 4692 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_23
timestamp 1623621585
transform 1 0 3220 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_30
timestamp 1623621585
transform 1 0 3864 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1623621585
transform 1 0 6348 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_51
timestamp 1623621585
transform 1 0 5796 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_58
timestamp 1623621585
transform 1 0 6440 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_42
timestamp 1623621585
transform 1 0 4968 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_54
timestamp 1623621585
transform 1 0 6072 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_70
timestamp 1623621585
transform 1 0 7544 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_82
timestamp 1623621585
transform 1 0 8648 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_66
timestamp 1623621585
transform 1 0 7176 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_78
timestamp 1623621585
transform 1 0 8280 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1623621585
transform 1 0 9016 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_94
timestamp 1623621585
transform 1 0 9752 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_87
timestamp 1623621585
transform 1 0 9108 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_99
timestamp 1623621585
transform 1 0 10212 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1623621585
transform 1 0 11592 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_106
timestamp 1623621585
transform 1 0 10856 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_115
timestamp 1623621585
transform 1 0 11684 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_111
timestamp 1623621585
transform 1 0 11316 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1623621585
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1623621585
transform 1 0 14260 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_127
timestamp 1623621585
transform 1 0 12788 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_139
timestamp 1623621585
transform 1 0 13892 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_135
timestamp 1623621585
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_144
timestamp 1623621585
transform 1 0 14352 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_151
timestamp 1623621585
transform 1 0 14996 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_163
timestamp 1623621585
transform 1 0 16100 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_156
timestamp 1623621585
transform 1 0 15456 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1623621585
transform 1 0 16836 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_172
timestamp 1623621585
transform 1 0 16928 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_184
timestamp 1623621585
transform 1 0 18032 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_168
timestamp 1623621585
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_180
timestamp 1623621585
transform 1 0 17664 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1623621585
transform 1 0 19504 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_196
timestamp 1623621585
transform 1 0 19136 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_208
timestamp 1623621585
transform 1 0 20240 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_192
timestamp 1623621585
transform 1 0 18768 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_201
timestamp 1623621585
transform 1 0 19596 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1623621585
transform 1 0 22080 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_220
timestamp 1623621585
transform 1 0 21344 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_229
timestamp 1623621585
transform 1 0 22172 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_213
timestamp 1623621585
transform 1 0 20700 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1623621585
transform 1 0 21804 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _350_
timestamp 1623621585
transform 1 0 24012 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _512_
timestamp 1623621585
transform 1 0 24012 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_wb_clk_i
timestamp 1623621585
transform 1 0 23368 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_241
timestamp 1623621585
transform 1 0 23276 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_245
timestamp 1623621585
transform 1 0 23644 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1623621585
transform 1 0 22908 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _766_
timestamp 1623621585
transform 1 0 25208 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _767_
timestamp 1623621585
transform 1 0 25024 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1623621585
transform 1 0 24748 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_256
timestamp 1623621585
transform 1 0 24656 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_253
timestamp 1623621585
transform 1 0 24380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_258
timestamp 1623621585
transform 1 0 24840 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _769_
timestamp 1623621585
transform 1 0 27048 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _771_
timestamp 1623621585
transform 1 0 27784 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1623621585
transform 1 0 27324 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_276
timestamp 1623621585
transform 1 0 26496 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_284
timestamp 1623621585
transform 1 0 27232 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_286
timestamp 1623621585
transform 1 0 27416 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_278
timestamp 1623621585
transform 1 0 26680 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _472_
timestamp 1623621585
transform 1 0 28980 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _791_
timestamp 1623621585
transform 1 0 29624 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_26_306
timestamp 1623621585
transform 1 0 29256 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_298
timestamp 1623621585
transform 1 0 28520 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_302
timestamp 1623621585
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_310
timestamp 1623621585
transform 1 0 29624 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _518_
timestamp 1623621585
transform 1 0 31464 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _793_
timestamp 1623621585
transform 1 0 30452 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1623621585
transform 1 0 29992 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_326
timestamp 1623621585
transform 1 0 31096 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_315
timestamp 1623621585
transform 1 0 30084 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_335
timestamp 1623621585
transform 1 0 31924 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_343
timestamp 1623621585
transform 1 0 32660 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_341
timestamp 1623621585
transform 1 0 32476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_337
timestamp 1623621585
transform 1 0 32108 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1623621585
transform 1 0 32568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _519_
timestamp 1623621585
transform 1 0 32292 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_354
timestamp 1623621585
transform 1 0 33672 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_351
timestamp 1623621585
transform 1 0 33396 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_1  _504_
timestamp 1623621585
transform 1 0 33488 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_27_342
timestamp 1623621585
transform 1 0 32568 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_1  _484_
timestamp 1623621585
transform 1 0 33764 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _517_
timestamp 1623621585
transform 1 0 34500 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1623621585
transform 1 0 35236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1623621585
transform 1 0 34132 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_370
timestamp 1623621585
transform 1 0 35144 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_362
timestamp 1623621585
transform 1 0 34408 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_370
timestamp 1623621585
transform 1 0 35144 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_372
timestamp 1623621585
transform 1 0 35328 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input181
timestamp 1623621585
transform 1 0 37260 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_382
timestamp 1623621585
transform 1 0 36248 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_394
timestamp 1623621585
transform 1 0 37352 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_384
timestamp 1623621585
transform 1 0 36432 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_392
timestamp 1623621585
transform 1 0 37168 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1623621585
transform -1 0 38824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1623621585
transform -1 0 38824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1623621585
transform 1 0 37812 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input138
timestamp 1623621585
transform 1 0 37904 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_398
timestamp 1623621585
transform 1 0 37720 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_400
timestamp 1623621585
transform 1 0 37904 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_406
timestamp 1623621585
transform 1 0 38456 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_396
timestamp 1623621585
transform 1 0 37536 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_403
timestamp 1623621585
transform 1 0 38180 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1623621585
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input333
timestamp 1623621585
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1623621585
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_11
timestamp 1623621585
transform 1 0 2116 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_23
timestamp 1623621585
transform 1 0 3220 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_35
timestamp 1623621585
transform 1 0 4324 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1623621585
transform 1 0 6348 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_47
timestamp 1623621585
transform 1 0 5428 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_55
timestamp 1623621585
transform 1 0 6164 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_58
timestamp 1623621585
transform 1 0 6440 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_70
timestamp 1623621585
transform 1 0 7544 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_82
timestamp 1623621585
transform 1 0 8648 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_94
timestamp 1623621585
transform 1 0 9752 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1623621585
transform 1 0 11592 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_106
timestamp 1623621585
transform 1 0 10856 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_115
timestamp 1623621585
transform 1 0 11684 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_127
timestamp 1623621585
transform 1 0 12788 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_139
timestamp 1623621585
transform 1 0 13892 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_151
timestamp 1623621585
transform 1 0 14996 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_163
timestamp 1623621585
transform 1 0 16100 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1623621585
transform 1 0 16836 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_172
timestamp 1623621585
transform 1 0 16928 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_184
timestamp 1623621585
transform 1 0 18032 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_196
timestamp 1623621585
transform 1 0 19136 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_208
timestamp 1623621585
transform 1 0 20240 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1623621585
transform 1 0 22080 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_220
timestamp 1623621585
transform 1 0 21344 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_229
timestamp 1623621585
transform 1 0 22172 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _764_
timestamp 1623621585
transform 1 0 23552 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_28_241
timestamp 1623621585
transform 1 0 23276 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _765_
timestamp 1623621585
transform 1 0 25392 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_260
timestamp 1623621585
transform 1 0 25024 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _790_
timestamp 1623621585
transform 1 0 27784 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1623621585
transform 1 0 27324 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_280
timestamp 1623621585
transform 1 0 26864 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_284
timestamp 1623621585
transform 1 0 27232 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_286
timestamp 1623621585
transform 1 0 27416 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _792_
timestamp 1623621585
transform 1 0 29624 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_306
timestamp 1623621585
transform 1 0 29256 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _478_
timestamp 1623621585
transform 1 0 31464 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_28_326
timestamp 1623621585
transform 1 0 31096 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _803_
timestamp 1623621585
transform 1 0 33028 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1623621585
transform 1 0 32568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_337
timestamp 1623621585
transform 1 0 32108 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_341
timestamp 1623621585
transform 1 0 32476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_343
timestamp 1623621585
transform 1 0 32660 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _498_
timestamp 1623621585
transform 1 0 34868 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_28_363
timestamp 1623621585
transform 1 0 34500 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_374
timestamp 1623621585
transform 1 0 35512 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_386
timestamp 1623621585
transform 1 0 36616 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1623621585
transform -1 0 38824 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1623621585
transform 1 0 37812 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_398
timestamp 1623621585
transform 1 0 37720 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_400
timestamp 1623621585
transform 1 0 37904 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_406
timestamp 1623621585
transform 1 0 38456 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1623621585
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1623621585
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1623621585
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1623621585
transform 1 0 3772 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_27
timestamp 1623621585
transform 1 0 3588 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_30
timestamp 1623621585
transform 1 0 3864 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_42
timestamp 1623621585
transform 1 0 4968 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_54
timestamp 1623621585
transform 1 0 6072 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_66
timestamp 1623621585
transform 1 0 7176 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_78
timestamp 1623621585
transform 1 0 8280 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1623621585
transform 1 0 9016 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_87
timestamp 1623621585
transform 1 0 9108 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_99
timestamp 1623621585
transform 1 0 10212 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_111
timestamp 1623621585
transform 1 0 11316 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1623621585
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1623621585
transform 1 0 14260 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_135
timestamp 1623621585
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_144
timestamp 1623621585
transform 1 0 14352 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_156
timestamp 1623621585
transform 1 0 15456 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_168
timestamp 1623621585
transform 1 0 16560 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_180
timestamp 1623621585
transform 1 0 17664 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1623621585
transform 1 0 19504 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_192
timestamp 1623621585
transform 1 0 18768 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_201
timestamp 1623621585
transform 1 0 19596 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_213
timestamp 1623621585
transform 1 0 20700 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1623621585
transform 1 0 21804 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1623621585
transform 1 0 22908 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_249
timestamp 1623621585
transform 1 0 24012 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _768_
timestamp 1623621585
transform 1 0 25208 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1623621585
transform 1 0 24748 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_258
timestamp 1623621585
transform 1 0 24840 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _770_
timestamp 1623621585
transform 1 0 27048 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_278
timestamp 1623621585
transform 1 0 26680 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _459_
timestamp 1623621585
transform 1 0 28980 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_29_298
timestamp 1623621585
transform 1 0 28520 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_302
timestamp 1623621585
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_310
timestamp 1623621585
transform 1 0 29624 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _795_
timestamp 1623621585
transform 1 0 30452 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1623621585
transform 1 0 29992 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_315
timestamp 1623621585
transform 1 0 30084 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _798_
timestamp 1623621585
transform 1 0 32292 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_335
timestamp 1623621585
transform 1 0 31924 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _471_
timestamp 1623621585
transform 1 0 34132 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1623621585
transform 1 0 35236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_355
timestamp 1623621585
transform 1 0 33764 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_366
timestamp 1623621585
transform 1 0 34776 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_370
timestamp 1623621585
transform 1 0 35144 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_372
timestamp 1623621585
transform 1 0 35328 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _468_
timestamp 1623621585
transform 1 0 35696 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input149
timestamp 1623621585
transform 1 0 37260 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_379
timestamp 1623621585
transform 1 0 35972 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_391
timestamp 1623621585
transform 1 0 37076 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1623621585
transform -1 0 38824 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input117
timestamp 1623621585
transform 1 0 37904 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_396
timestamp 1623621585
transform 1 0 37536 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1623621585
transform 1 0 38180 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1623621585
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input334
timestamp 1623621585
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1623621585
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_11
timestamp 1623621585
transform 1 0 2116 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_23
timestamp 1623621585
transform 1 0 3220 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_35
timestamp 1623621585
transform 1 0 4324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1623621585
transform 1 0 6348 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_47
timestamp 1623621585
transform 1 0 5428 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_55
timestamp 1623621585
transform 1 0 6164 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_58
timestamp 1623621585
transform 1 0 6440 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_70
timestamp 1623621585
transform 1 0 7544 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_82
timestamp 1623621585
transform 1 0 8648 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_94
timestamp 1623621585
transform 1 0 9752 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1623621585
transform 1 0 11592 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_106
timestamp 1623621585
transform 1 0 10856 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_115
timestamp 1623621585
transform 1 0 11684 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_127
timestamp 1623621585
transform 1 0 12788 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_139
timestamp 1623621585
transform 1 0 13892 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_151
timestamp 1623621585
transform 1 0 14996 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_163
timestamp 1623621585
transform 1 0 16100 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1623621585
transform 1 0 16836 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_172
timestamp 1623621585
transform 1 0 16928 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_184
timestamp 1623621585
transform 1 0 18032 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_196
timestamp 1623621585
transform 1 0 19136 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_208
timestamp 1623621585
transform 1 0 20240 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1623621585
transform 1 0 22080 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_220
timestamp 1623621585
transform 1 0 21344 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_229
timestamp 1623621585
transform 1 0 22172 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_241
timestamp 1623621585
transform 1 0 23276 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1623621585
transform 1 0 24012 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _318_
timestamp 1623621585
transform 1 0 24288 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_261
timestamp 1623621585
transform 1 0 25116 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_269
timestamp 1623621585
transform 1 0 25852 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_2  _320_
timestamp 1623621585
transform 1 0 27784 0 -1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _582_
timestamp 1623621585
transform 1 0 26128 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1623621585
transform 1 0 27324 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_279
timestamp 1623621585
transform 1 0 26772 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_286
timestamp 1623621585
transform 1 0 27416 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _794_
timestamp 1623621585
transform 1 0 29348 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_30_300
timestamp 1623621585
transform 1 0 28704 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_306
timestamp 1623621585
transform 1 0 29256 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _351_
timestamp 1623621585
transform 1 0 31188 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_323
timestamp 1623621585
transform 1 0 30820 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_331
timestamp 1623621585
transform 1 0 31556 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _801_
timestamp 1623621585
transform 1 0 33028 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1623621585
transform 1 0 32568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_wb_clk_i
timestamp 1623621585
transform 1 0 31924 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_338
timestamp 1623621585
transform 1 0 32200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_343
timestamp 1623621585
transform 1 0 32660 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _477_
timestamp 1623621585
transform 1 0 34868 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_30_363
timestamp 1623621585
transform 1 0 34500 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_374
timestamp 1623621585
transform 1 0 35512 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _411_
timestamp 1623621585
transform 1 0 35880 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input184
timestamp 1623621585
transform 1 0 37168 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_382
timestamp 1623621585
transform 1 0 36248 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_390
timestamp 1623621585
transform 1 0 36984 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_395
timestamp 1623621585
transform 1 0 37444 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1623621585
transform -1 0 38824 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1623621585
transform 1 0 37812 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_400
timestamp 1623621585
transform 1 0 37904 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1623621585
transform 1 0 38456 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1623621585
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input335
timestamp 1623621585
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1623621585
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_11
timestamp 1623621585
transform 1 0 2116 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1623621585
transform 1 0 3772 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_23
timestamp 1623621585
transform 1 0 3220 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_30
timestamp 1623621585
transform 1 0 3864 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_42
timestamp 1623621585
transform 1 0 4968 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_54
timestamp 1623621585
transform 1 0 6072 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_66
timestamp 1623621585
transform 1 0 7176 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_78
timestamp 1623621585
transform 1 0 8280 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1623621585
transform 1 0 9016 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_87
timestamp 1623621585
transform 1 0 9108 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_99
timestamp 1623621585
transform 1 0 10212 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_111
timestamp 1623621585
transform 1 0 11316 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1623621585
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1623621585
transform 1 0 14260 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_135
timestamp 1623621585
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_144
timestamp 1623621585
transform 1 0 14352 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_156
timestamp 1623621585
transform 1 0 15456 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_168
timestamp 1623621585
transform 1 0 16560 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_180
timestamp 1623621585
transform 1 0 17664 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1623621585
transform 1 0 19504 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_192
timestamp 1623621585
transform 1 0 18768 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_201
timestamp 1623621585
transform 1 0 19596 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_213
timestamp 1623621585
transform 1 0 20700 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1623621585
transform 1 0 21804 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_1  _319_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 23920 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_31_237
timestamp 1623621585
transform 1 0 22908 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_245
timestamp 1623621585
transform 1 0 23644 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _314_
timestamp 1623621585
transform 1 0 25852 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1623621585
transform 1 0 24748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_253
timestamp 1623621585
transform 1 0 24380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_258
timestamp 1623621585
transform 1 0 24840 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_266
timestamp 1623621585
transform 1 0 25576 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  _587_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 26588 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 27784 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_31_273
timestamp 1623621585
transform 1 0 26220 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_286
timestamp 1623621585
transform 1 0 27416 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_310
timestamp 1623621585
transform 1 0 29624 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _796_
timestamp 1623621585
transform 1 0 30452 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1623621585
transform 1 0 29992 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_315
timestamp 1623621585
transform 1 0 30084 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _797_
timestamp 1623621585
transform 1 0 32292 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_335
timestamp 1623621585
transform 1 0 31924 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _458_
timestamp 1623621585
transform 1 0 34132 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1623621585
transform 1 0 35236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_355
timestamp 1623621585
transform 1 0 33764 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_366
timestamp 1623621585
transform 1 0 34776 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_370
timestamp 1623621585
transform 1 0 35144 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_372
timestamp 1623621585
transform 1 0 35328 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _428_
timestamp 1623621585
transform 1 0 35696 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input152
timestamp 1623621585
transform 1 0 37260 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_379
timestamp 1623621585
transform 1 0 35972 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_391
timestamp 1623621585
transform 1 0 37076 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1623621585
transform -1 0 38824 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input120
timestamp 1623621585
transform 1 0 37904 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_396
timestamp 1623621585
transform 1 0 37536 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_403
timestamp 1623621585
transform 1 0 38180 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1623621585
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1623621585
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1623621585
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_27
timestamp 1623621585
transform 1 0 3588 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_39
timestamp 1623621585
transform 1 0 4692 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1623621585
transform 1 0 6348 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_51
timestamp 1623621585
transform 1 0 5796 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_58
timestamp 1623621585
transform 1 0 6440 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_70
timestamp 1623621585
transform 1 0 7544 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_82
timestamp 1623621585
transform 1 0 8648 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1623621585
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1623621585
transform 1 0 11592 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_106
timestamp 1623621585
transform 1 0 10856 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_115
timestamp 1623621585
transform 1 0 11684 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_127
timestamp 1623621585
transform 1 0 12788 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_139
timestamp 1623621585
transform 1 0 13892 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_151
timestamp 1623621585
transform 1 0 14996 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_163
timestamp 1623621585
transform 1 0 16100 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1623621585
transform 1 0 16836 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_172
timestamp 1623621585
transform 1 0 16928 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_184
timestamp 1623621585
transform 1 0 18032 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_196
timestamp 1623621585
transform 1 0 19136 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_208
timestamp 1623621585
transform 1 0 20240 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1623621585
transform 1 0 22080 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_220
timestamp 1623621585
transform 1 0 21344 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_229
timestamp 1623621585
transform 1 0 22172 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_241
timestamp 1623621585
transform 1 0 23276 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_4  _618_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 25668 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1623621585
transform 1 0 24380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_265
timestamp 1623621585
transform 1 0 25484 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _439_
timestamp 1623621585
transform 1 0 27876 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1623621585
transform 1 0 27324 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_276
timestamp 1623621585
transform 1 0 26496 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_284
timestamp 1623621585
transform 1 0 27232 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_286
timestamp 1623621585
transform 1 0 27416 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_290
timestamp 1623621585
transform 1 0 27784 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _445_
timestamp 1623621585
transform 1 0 29532 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _465_
timestamp 1623621585
transform 1 0 28520 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_32_294
timestamp 1623621585
transform 1 0 28152 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_305
timestamp 1623621585
transform 1 0 29164 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _399_
timestamp 1623621585
transform 1 0 31556 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _438_
timestamp 1623621585
transform 1 0 30544 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_32_316
timestamp 1623621585
transform 1 0 30176 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_327
timestamp 1623621585
transform 1 0 31188 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _800_
timestamp 1623621585
transform 1 0 33028 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1623621585
transform 1 0 32568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_334
timestamp 1623621585
transform 1 0 31832 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_343
timestamp 1623621585
transform 1 0 32660 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _464_
timestamp 1623621585
transform 1 0 34868 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_32_363
timestamp 1623621585
transform 1 0 34500 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_374
timestamp 1623621585
transform 1 0 35512 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _367_
timestamp 1623621585
transform 1 0 35880 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input185
timestamp 1623621585
transform 1 0 37168 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_382
timestamp 1623621585
transform 1 0 36248 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_390
timestamp 1623621585
transform 1 0 36984 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_395
timestamp 1623621585
transform 1 0 37444 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1623621585
transform -1 0 38824 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1623621585
transform 1 0 37812 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_400
timestamp 1623621585
transform 1 0 37904 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_406
timestamp 1623621585
transform 1 0 38456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1623621585
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1623621585
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input336
timestamp 1623621585
transform 1 0 1748 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input337
timestamp 1623621585
transform 1 0 1748 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1623621585
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_11
timestamp 1623621585
transform 1 0 2116 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1623621585
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_11
timestamp 1623621585
transform 1 0 2116 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1623621585
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_23
timestamp 1623621585
transform 1 0 3220 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_30
timestamp 1623621585
transform 1 0 3864 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_23
timestamp 1623621585
transform 1 0 3220 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_35
timestamp 1623621585
transform 1 0 4324 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1623621585
transform 1 0 6348 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_42
timestamp 1623621585
transform 1 0 4968 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_54
timestamp 1623621585
transform 1 0 6072 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_47
timestamp 1623621585
transform 1 0 5428 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_55
timestamp 1623621585
transform 1 0 6164 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_58
timestamp 1623621585
transform 1 0 6440 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_66
timestamp 1623621585
transform 1 0 7176 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_78
timestamp 1623621585
transform 1 0 8280 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_70
timestamp 1623621585
transform 1 0 7544 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_82
timestamp 1623621585
transform 1 0 8648 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1623621585
transform 1 0 9016 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_87
timestamp 1623621585
transform 1 0 9108 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_99
timestamp 1623621585
transform 1 0 10212 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_94
timestamp 1623621585
transform 1 0 9752 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1623621585
transform 1 0 11592 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_111
timestamp 1623621585
transform 1 0 11316 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1623621585
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_106
timestamp 1623621585
transform 1 0 10856 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_115
timestamp 1623621585
transform 1 0 11684 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1623621585
transform 1 0 14260 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_135
timestamp 1623621585
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_144
timestamp 1623621585
transform 1 0 14352 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_127
timestamp 1623621585
transform 1 0 12788 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_139
timestamp 1623621585
transform 1 0 13892 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_156
timestamp 1623621585
transform 1 0 15456 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_151
timestamp 1623621585
transform 1 0 14996 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_163
timestamp 1623621585
transform 1 0 16100 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1623621585
transform 1 0 16836 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_168
timestamp 1623621585
transform 1 0 16560 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_180
timestamp 1623621585
transform 1 0 17664 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_172
timestamp 1623621585
transform 1 0 16928 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_184
timestamp 1623621585
transform 1 0 18032 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1623621585
transform 1 0 19504 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_192
timestamp 1623621585
transform 1 0 18768 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_201
timestamp 1623621585
transform 1 0 19596 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_196
timestamp 1623621585
transform 1 0 19136 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_208
timestamp 1623621585
transform 1 0 20240 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1623621585
transform 1 0 22080 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_213
timestamp 1623621585
transform 1 0 20700 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1623621585
transform 1 0 21804 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_220
timestamp 1623621585
transform 1 0 21344 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_229
timestamp 1623621585
transform 1 0 22172 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1623621585
transform 1 0 22908 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_249
timestamp 1623621585
transform 1 0 24012 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_241
timestamp 1623621585
transform 1 0 23276 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1623621585
transform 1 0 24748 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_258
timestamp 1623621585
transform 1 0 24840 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_270
timestamp 1623621585
transform 1 0 25944 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1623621585
transform 1 0 24380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1623621585
transform 1 0 25484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _479_
timestamp 1623621585
transform 1 0 27876 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1623621585
transform 1 0 27324 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_wb_clk_i
timestamp 1623621585
transform 1 0 27232 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_282
timestamp 1623621585
transform 1 0 27048 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_287
timestamp 1623621585
transform 1 0 27508 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_277
timestamp 1623621585
transform 1 0 26588 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_286
timestamp 1623621585
transform 1 0 27416 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _307_
timestamp 1623621585
transform 1 0 28520 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_294
timestamp 1623621585
transform 1 0 28152 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_302
timestamp 1623621585
transform 1 0 28888 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_298
timestamp 1623621585
transform 1 0 28520 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_310
timestamp 1623621585
transform 1 0 29624 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _419_
timestamp 1623621585
transform 1 0 31280 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _425_
timestamp 1623621585
transform 1 0 30268 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _432_
timestamp 1623621585
transform 1 0 30636 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _799_
timestamp 1623621585
transform 1 0 31648 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1623621585
transform 1 0 29992 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_315
timestamp 1623621585
transform 1 0 30084 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_328
timestamp 1623621585
transform 1 0 31280 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_316
timestamp 1623621585
transform 1 0 30176 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_324
timestamp 1623621585
transform 1 0 30912 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _327_
timestamp 1623621585
transform 1 0 33488 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _802_
timestamp 1623621585
transform 1 0 33028 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1623621585
transform 1 0 32568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_348
timestamp 1623621585
transform 1 0 33120 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_335
timestamp 1623621585
transform 1 0 31924 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_341
timestamp 1623621585
transform 1 0 32476 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_343
timestamp 1623621585
transform 1 0 32660 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _431_
timestamp 1623621585
transform 1 0 34868 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _444_
timestamp 1623621585
transform 1 0 34224 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1623621585
transform 1 0 35236 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_356
timestamp 1623621585
transform 1 0 33856 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_367
timestamp 1623621585
transform 1 0 34868 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_372
timestamp 1623621585
transform 1 0 35328 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_363
timestamp 1623621585
transform 1 0 34500 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_374
timestamp 1623621585
transform 1 0 35512 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _388_
timestamp 1623621585
transform 1 0 35696 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _437_
timestamp 1623621585
transform 1 0 35880 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input153
timestamp 1623621585
transform 1 0 37168 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_380
timestamp 1623621585
transform 1 0 36064 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_392
timestamp 1623621585
transform 1 0 37168 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_385
timestamp 1623621585
transform 1 0 36524 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_391
timestamp 1623621585
transform 1 0 37076 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_395
timestamp 1623621585
transform 1 0 37444 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1623621585
transform -1 0 38824 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1623621585
transform -1 0 38824 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1623621585
transform 1 0 37812 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input121
timestamp 1623621585
transform 1 0 37904 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_403
timestamp 1623621585
transform 1 0 38180 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_400
timestamp 1623621585
transform 1 0 37904 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_406
timestamp 1623621585
transform 1 0 38456 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1623621585
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1623621585
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1623621585
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1623621585
transform 1 0 3772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_27
timestamp 1623621585
transform 1 0 3588 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_30
timestamp 1623621585
transform 1 0 3864 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_42
timestamp 1623621585
transform 1 0 4968 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_54
timestamp 1623621585
transform 1 0 6072 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_66
timestamp 1623621585
transform 1 0 7176 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_78
timestamp 1623621585
transform 1 0 8280 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1623621585
transform 1 0 9016 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_87
timestamp 1623621585
transform 1 0 9108 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_99
timestamp 1623621585
transform 1 0 10212 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_111
timestamp 1623621585
transform 1 0 11316 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1623621585
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1623621585
transform 1 0 14260 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_135
timestamp 1623621585
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_144
timestamp 1623621585
transform 1 0 14352 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1623621585
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1623621585
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_180
timestamp 1623621585
transform 1 0 17664 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1623621585
transform 1 0 19504 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_192
timestamp 1623621585
transform 1 0 18768 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_201
timestamp 1623621585
transform 1 0 19596 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_213
timestamp 1623621585
transform 1 0 20700 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1623621585
transform 1 0 21804 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1623621585
transform 1 0 22908 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_249
timestamp 1623621585
transform 1 0 24012 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1623621585
transform 1 0 24748 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_258
timestamp 1623621585
transform 1 0 24840 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_270
timestamp 1623621585
transform 1 0 25944 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_282
timestamp 1623621585
transform 1 0 27048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_294
timestamp 1623621585
transform 1 0 28152 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_306
timestamp 1623621585
transform 1 0 29256 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _405_
timestamp 1623621585
transform 1 0 31648 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1623621585
transform 1 0 29992 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_315
timestamp 1623621585
transform 1 0 30084 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_327
timestamp 1623621585
transform 1 0 31188 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_331
timestamp 1623621585
transform 1 0 31556 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_wb_clk_i
timestamp 1623621585
transform 1 0 32660 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_339
timestamp 1623621585
transform 1 0 32292 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_346
timestamp 1623621585
transform 1 0 32936 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _339_
timestamp 1623621585
transform 1 0 34040 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1623621585
transform 1 0 35236 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_362
timestamp 1623621585
transform 1 0 34408 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_370
timestamp 1623621585
transform 1 0 35144 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_372
timestamp 1623621585
transform 1 0 35328 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input186
timestamp 1623621585
transform 1 0 37260 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_384
timestamp 1623621585
transform 1 0 36432 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_392
timestamp 1623621585
transform 1 0 37168 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1623621585
transform -1 0 38824 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input122
timestamp 1623621585
transform 1 0 37904 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_396
timestamp 1623621585
transform 1 0 37536 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_403
timestamp 1623621585
transform 1 0 38180 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1623621585
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input338
timestamp 1623621585
transform 1 0 1748 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1623621585
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_11
timestamp 1623621585
transform 1 0 2116 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_23
timestamp 1623621585
transform 1 0 3220 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_35
timestamp 1623621585
transform 1 0 4324 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1623621585
transform 1 0 6348 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_47
timestamp 1623621585
transform 1 0 5428 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_55
timestamp 1623621585
transform 1 0 6164 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_58
timestamp 1623621585
transform 1 0 6440 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_70
timestamp 1623621585
transform 1 0 7544 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_82
timestamp 1623621585
transform 1 0 8648 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_94
timestamp 1623621585
transform 1 0 9752 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1623621585
transform 1 0 11592 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_106
timestamp 1623621585
transform 1 0 10856 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_115
timestamp 1623621585
transform 1 0 11684 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_127
timestamp 1623621585
transform 1 0 12788 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_139
timestamp 1623621585
transform 1 0 13892 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_151
timestamp 1623621585
transform 1 0 14996 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_163
timestamp 1623621585
transform 1 0 16100 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1623621585
transform 1 0 16836 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_172
timestamp 1623621585
transform 1 0 16928 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_184
timestamp 1623621585
transform 1 0 18032 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_196
timestamp 1623621585
transform 1 0 19136 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_208
timestamp 1623621585
transform 1 0 20240 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1623621585
transform 1 0 22080 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_220
timestamp 1623621585
transform 1 0 21344 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_229
timestamp 1623621585
transform 1 0 22172 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_241
timestamp 1623621585
transform 1 0 23276 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1623621585
transform 1 0 24380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1623621585
transform 1 0 25484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1623621585
transform 1 0 27324 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_277
timestamp 1623621585
transform 1 0 26588 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_286
timestamp 1623621585
transform 1 0 27416 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_298
timestamp 1623621585
transform 1 0 28520 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_310
timestamp 1623621585
transform 1 0 29624 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_322
timestamp 1623621585
transform 1 0 30728 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _392_
timestamp 1623621585
transform 1 0 33028 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1623621585
transform 1 0 32568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_334
timestamp 1623621585
transform 1 0 31832 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_343
timestamp 1623621585
transform 1 0 32660 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_354
timestamp 1623621585
transform 1 0 33672 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_1  _418_
timestamp 1623621585
transform 1 0 34868 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_36_366
timestamp 1623621585
transform 1 0 34776 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_374
timestamp 1623621585
transform 1 0 35512 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _424_
timestamp 1623621585
transform 1 0 35880 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_36_385
timestamp 1623621585
transform 1 0 36524 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1623621585
transform -1 0 38824 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1623621585
transform 1 0 37812 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_397
timestamp 1623621585
transform 1 0 37628 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_400
timestamp 1623621585
transform 1 0 37904 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_406
timestamp 1623621585
transform 1 0 38456 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1623621585
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input339
timestamp 1623621585
transform 1 0 1748 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1623621585
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_13
timestamp 1623621585
transform 1 0 2300 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1623621585
transform 1 0 3772 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_25
timestamp 1623621585
transform 1 0 3404 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_30
timestamp 1623621585
transform 1 0 3864 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_42
timestamp 1623621585
transform 1 0 4968 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_54
timestamp 1623621585
transform 1 0 6072 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_66
timestamp 1623621585
transform 1 0 7176 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_78
timestamp 1623621585
transform 1 0 8280 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1623621585
transform 1 0 9016 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_87
timestamp 1623621585
transform 1 0 9108 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_99
timestamp 1623621585
transform 1 0 10212 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_111
timestamp 1623621585
transform 1 0 11316 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1623621585
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1623621585
transform 1 0 14260 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_135
timestamp 1623621585
transform 1 0 13524 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_144
timestamp 1623621585
transform 1 0 14352 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_156
timestamp 1623621585
transform 1 0 15456 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_168
timestamp 1623621585
transform 1 0 16560 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_180
timestamp 1623621585
transform 1 0 17664 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1623621585
transform 1 0 19504 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_192
timestamp 1623621585
transform 1 0 18768 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_201
timestamp 1623621585
transform 1 0 19596 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_213
timestamp 1623621585
transform 1 0 20700 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1623621585
transform 1 0 21804 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1623621585
transform 1 0 22908 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_249
timestamp 1623621585
transform 1 0 24012 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1623621585
transform 1 0 24748 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_258
timestamp 1623621585
transform 1 0 24840 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_270
timestamp 1623621585
transform 1 0 25944 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _806_
timestamp 1623621585
transform 1 0 26404 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_37_274
timestamp 1623621585
transform 1 0 26312 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_291
timestamp 1623621585
transform 1 0 27876 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_303
timestamp 1623621585
transform 1 0 28980 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_311
timestamp 1623621585
transform 1 0 29716 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1623621585
transform 1 0 29992 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_315
timestamp 1623621585
transform 1 0 30084 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_327
timestamp 1623621585
transform 1 0 31188 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_333
timestamp 1623621585
transform 1 0 31740 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _349_
timestamp 1623621585
transform 1 0 32844 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _385_
timestamp 1623621585
transform 1 0 31832 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_37_341
timestamp 1623621585
transform 1 0 32476 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_352
timestamp 1623621585
transform 1 0 33488 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _398_
timestamp 1623621585
transform 1 0 33856 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1623621585
transform 1 0 35236 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_363
timestamp 1623621585
transform 1 0 34500 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_372
timestamp 1623621585
transform 1 0 35328 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _404_
timestamp 1623621585
transform 1 0 35696 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input187
timestamp 1623621585
transform 1 0 37260 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_383
timestamp 1623621585
transform 1 0 36340 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_391
timestamp 1623621585
transform 1 0 37076 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1623621585
transform -1 0 38824 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input154
timestamp 1623621585
transform 1 0 37904 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_396
timestamp 1623621585
transform 1 0 37536 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_403
timestamp 1623621585
transform 1 0 38180 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1623621585
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1623621585
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1623621585
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_27
timestamp 1623621585
transform 1 0 3588 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_39
timestamp 1623621585
transform 1 0 4692 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1623621585
transform 1 0 6348 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_51
timestamp 1623621585
transform 1 0 5796 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_58
timestamp 1623621585
transform 1 0 6440 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_70
timestamp 1623621585
transform 1 0 7544 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_82
timestamp 1623621585
transform 1 0 8648 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_94
timestamp 1623621585
transform 1 0 9752 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1623621585
transform 1 0 11592 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_106
timestamp 1623621585
transform 1 0 10856 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_115
timestamp 1623621585
transform 1 0 11684 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_127
timestamp 1623621585
transform 1 0 12788 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_139
timestamp 1623621585
transform 1 0 13892 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_151
timestamp 1623621585
transform 1 0 14996 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_163
timestamp 1623621585
transform 1 0 16100 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1623621585
transform 1 0 16836 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_172
timestamp 1623621585
transform 1 0 16928 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_184
timestamp 1623621585
transform 1 0 18032 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_196
timestamp 1623621585
transform 1 0 19136 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_208
timestamp 1623621585
transform 1 0 20240 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1623621585
transform 1 0 22080 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_220
timestamp 1623621585
transform 1 0 21344 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_229
timestamp 1623621585
transform 1 0 22172 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_241
timestamp 1623621585
transform 1 0 23276 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1623621585
transform 1 0 24380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1623621585
transform 1 0 25484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _805_
timestamp 1623621585
transform 1 0 27784 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1623621585
transform 1 0 27324 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_277
timestamp 1623621585
transform 1 0 26588 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_286
timestamp 1623621585
transform 1 0 27416 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_306
timestamp 1623621585
transform 1 0 29256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_318
timestamp 1623621585
transform 1 0 30360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_330
timestamp 1623621585
transform 1 0 31464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _335_
timestamp 1623621585
transform 1 0 33028 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1623621585
transform 1 0 32568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_343
timestamp 1623621585
transform 1 0 32660 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_354
timestamp 1623621585
transform 1 0 33672 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _357_
timestamp 1623621585
transform 1 0 34040 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _391_
timestamp 1623621585
transform 1 0 35236 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_38_365
timestamp 1623621585
transform 1 0 34684 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_378
timestamp 1623621585
transform 1 0 35880 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_390
timestamp 1623621585
transform 1 0 36984 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1623621585
transform -1 0 38824 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1623621585
transform 1 0 37812 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_398
timestamp 1623621585
transform 1 0 37720 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_400
timestamp 1623621585
transform 1 0 37904 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1623621585
transform 1 0 38456 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1623621585
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1623621585
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input340
timestamp 1623621585
transform 1 0 1748 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input342
timestamp 1623621585
transform 1 0 1748 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1623621585
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_13
timestamp 1623621585
transform 1 0 2300 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1623621585
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_13
timestamp 1623621585
transform 1 0 2300 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1623621585
transform 1 0 3772 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_25
timestamp 1623621585
transform 1 0 3404 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_30
timestamp 1623621585
transform 1 0 3864 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_25
timestamp 1623621585
transform 1 0 3404 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_37
timestamp 1623621585
transform 1 0 4508 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1623621585
transform 1 0 6348 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_42
timestamp 1623621585
transform 1 0 4968 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_54
timestamp 1623621585
transform 1 0 6072 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_49
timestamp 1623621585
transform 1 0 5612 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_58
timestamp 1623621585
transform 1 0 6440 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_66
timestamp 1623621585
transform 1 0 7176 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_78
timestamp 1623621585
transform 1 0 8280 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_70
timestamp 1623621585
transform 1 0 7544 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_82
timestamp 1623621585
transform 1 0 8648 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1623621585
transform 1 0 9016 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_87
timestamp 1623621585
transform 1 0 9108 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_99
timestamp 1623621585
transform 1 0 10212 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_94
timestamp 1623621585
transform 1 0 9752 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1623621585
transform 1 0 11592 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_111
timestamp 1623621585
transform 1 0 11316 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1623621585
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_106
timestamp 1623621585
transform 1 0 10856 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_115
timestamp 1623621585
transform 1 0 11684 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1623621585
transform 1 0 14260 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_135
timestamp 1623621585
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_144
timestamp 1623621585
transform 1 0 14352 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_127
timestamp 1623621585
transform 1 0 12788 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_139
timestamp 1623621585
transform 1 0 13892 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_156
timestamp 1623621585
transform 1 0 15456 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_151
timestamp 1623621585
transform 1 0 14996 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_163
timestamp 1623621585
transform 1 0 16100 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1623621585
transform 1 0 16836 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_168
timestamp 1623621585
transform 1 0 16560 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_180
timestamp 1623621585
transform 1 0 17664 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_172
timestamp 1623621585
transform 1 0 16928 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_184
timestamp 1623621585
transform 1 0 18032 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1623621585
transform 1 0 19504 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_192
timestamp 1623621585
transform 1 0 18768 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_201
timestamp 1623621585
transform 1 0 19596 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_196
timestamp 1623621585
transform 1 0 19136 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_208
timestamp 1623621585
transform 1 0 20240 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1623621585
transform 1 0 22080 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_213
timestamp 1623621585
transform 1 0 20700 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1623621585
transform 1 0 21804 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_220
timestamp 1623621585
transform 1 0 21344 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_229
timestamp 1623621585
transform 1 0 22172 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1623621585
transform 1 0 22908 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_249
timestamp 1623621585
transform 1 0 24012 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_241
timestamp 1623621585
transform 1 0 23276 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1623621585
transform 1 0 24748 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_258
timestamp 1623621585
transform 1 0 24840 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_270
timestamp 1623621585
transform 1 0 25944 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1623621585
transform 1 0 24380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1623621585
transform 1 0 25484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _315_
timestamp 1623621585
transform 1 0 27784 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 27232 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _317_
timestamp 1623621585
transform 1 0 27876 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1623621585
transform 1 0 27324 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_282
timestamp 1623621585
transform 1 0 27048 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_287
timestamp 1623621585
transform 1 0 27508 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_277
timestamp 1623621585
transform 1 0 26588 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_286
timestamp 1623621585
transform 1 0 27416 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _321_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 28888 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_294
timestamp 1623621585
transform 1 0 28152 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_306
timestamp 1623621585
transform 1 0 29256 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_297
timestamp 1623621585
transform 1 0 28428 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_301
timestamp 1623621585
transform 1 0 28796 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_310
timestamp 1623621585
transform 1 0 29624 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1623621585
transform 1 0 29992 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_315
timestamp 1623621585
transform 1 0 30084 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_327
timestamp 1623621585
transform 1 0 31188 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_322
timestamp 1623621585
transform 1 0 30728 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _343_
timestamp 1623621585
transform 1 0 33120 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _379_
timestamp 1623621585
transform 1 0 33028 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1623621585
transform 1 0 32568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_339
timestamp 1623621585
transform 1 0 32292 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_347
timestamp 1623621585
transform 1 0 33028 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_334
timestamp 1623621585
transform 1 0 31832 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_343
timestamp 1623621585
transform 1 0 32660 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_354
timestamp 1623621585
transform 1 0 33672 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_1  _378_
timestamp 1623621585
transform 1 0 35328 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1623621585
transform 1 0 35236 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_355
timestamp 1623621585
transform 1 0 33764 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_367
timestamp 1623621585
transform 1 0 34868 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_372
timestamp 1623621585
transform 1 0 35328 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_366
timestamp 1623621585
transform 1 0 34776 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _397_
timestamp 1623621585
transform 1 0 35696 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input155
timestamp 1623621585
transform 1 0 37260 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input188
timestamp 1623621585
transform 1 0 37168 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_383
timestamp 1623621585
transform 1 0 36340 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_391
timestamp 1623621585
transform 1 0 37076 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_379
timestamp 1623621585
transform 1 0 35972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_391
timestamp 1623621585
transform 1 0 37076 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_395
timestamp 1623621585
transform 1 0 37444 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1623621585
transform -1 0 38824 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1623621585
transform -1 0 38824 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1623621585
transform 1 0 37812 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input123
timestamp 1623621585
transform 1 0 37904 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_396
timestamp 1623621585
transform 1 0 37536 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_403
timestamp 1623621585
transform 1 0 38180 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_400
timestamp 1623621585
transform 1 0 37904 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_406
timestamp 1623621585
transform 1 0 38456 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1623621585
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1623621585
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1623621585
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1623621585
transform 1 0 3772 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_27
timestamp 1623621585
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_30
timestamp 1623621585
transform 1 0 3864 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_42
timestamp 1623621585
transform 1 0 4968 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_54
timestamp 1623621585
transform 1 0 6072 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_66
timestamp 1623621585
transform 1 0 7176 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_78
timestamp 1623621585
transform 1 0 8280 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1623621585
transform 1 0 9016 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_87
timestamp 1623621585
transform 1 0 9108 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_99
timestamp 1623621585
transform 1 0 10212 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_111
timestamp 1623621585
transform 1 0 11316 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1623621585
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1623621585
transform 1 0 14260 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_135
timestamp 1623621585
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_144
timestamp 1623621585
transform 1 0 14352 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_156
timestamp 1623621585
transform 1 0 15456 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_168
timestamp 1623621585
transform 1 0 16560 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_180
timestamp 1623621585
transform 1 0 17664 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1623621585
transform 1 0 19504 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_192
timestamp 1623621585
transform 1 0 18768 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_201
timestamp 1623621585
transform 1 0 19596 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_213
timestamp 1623621585
transform 1 0 20700 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1623621585
transform 1 0 21804 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1623621585
transform 1 0 22908 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_249
timestamp 1623621585
transform 1 0 24012 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1623621585
transform 1 0 24748 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_258
timestamp 1623621585
transform 1 0 24840 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_270
timestamp 1623621585
transform 1 0 25944 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1623621585
transform 1 0 27048 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1623621585
transform 1 0 27692 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_285
timestamp 1623621585
transform 1 0 27324 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_292
timestamp 1623621585
transform 1 0 27968 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_304
timestamp 1623621585
transform 1 0 29072 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_312
timestamp 1623621585
transform 1 0 29808 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1623621585
transform 1 0 29992 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_315
timestamp 1623621585
transform 1 0 30084 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_327
timestamp 1623621585
transform 1 0 31188 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _580_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 32844 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 32660 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_339
timestamp 1623621585
transform 1 0 32292 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_353
timestamp 1623621585
transform 1 0 33580 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1623621585
transform 1 0 35236 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_365
timestamp 1623621585
transform 1 0 34684 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_372
timestamp 1623621585
transform 1 0 35328 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _384_
timestamp 1623621585
transform 1 0 35696 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input156
timestamp 1623621585
transform 1 0 37260 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_383
timestamp 1623621585
transform 1 0 36340 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_391
timestamp 1623621585
transform 1 0 37076 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1623621585
transform -1 0 38824 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input124
timestamp 1623621585
transform 1 0 37904 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_396
timestamp 1623621585
transform 1 0 37536 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_403
timestamp 1623621585
transform 1 0 38180 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1623621585
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input343
timestamp 1623621585
transform 1 0 1748 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1623621585
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_13
timestamp 1623621585
transform 1 0 2300 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_25
timestamp 1623621585
transform 1 0 3404 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_37
timestamp 1623621585
transform 1 0 4508 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1623621585
transform 1 0 6348 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_49
timestamp 1623621585
transform 1 0 5612 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_58
timestamp 1623621585
transform 1 0 6440 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_70
timestamp 1623621585
transform 1 0 7544 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_82
timestamp 1623621585
transform 1 0 8648 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1623621585
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1623621585
transform 1 0 11592 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_106
timestamp 1623621585
transform 1 0 10856 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_115
timestamp 1623621585
transform 1 0 11684 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_127
timestamp 1623621585
transform 1 0 12788 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_139
timestamp 1623621585
transform 1 0 13892 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_151
timestamp 1623621585
transform 1 0 14996 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_163
timestamp 1623621585
transform 1 0 16100 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1623621585
transform 1 0 16836 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_172
timestamp 1623621585
transform 1 0 16928 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_184
timestamp 1623621585
transform 1 0 18032 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_196
timestamp 1623621585
transform 1 0 19136 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_208
timestamp 1623621585
transform 1 0 20240 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1623621585
transform 1 0 22080 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_220
timestamp 1623621585
transform 1 0 21344 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_229
timestamp 1623621585
transform 1 0 22172 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_241
timestamp 1623621585
transform 1 0 23276 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1623621585
transform 1 0 24380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1623621585
transform 1 0 25484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1623621585
transform 1 0 27324 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_277
timestamp 1623621585
transform 1 0 26588 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_286
timestamp 1623621585
transform 1 0 27416 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_298
timestamp 1623621585
transform 1 0 28520 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_310
timestamp 1623621585
transform 1 0 29624 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_322
timestamp 1623621585
transform 1 0 30728 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _574_
timestamp 1623621585
transform 1 0 33028 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1623621585
transform 1 0 32568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_13
timestamp 1623621585
transform 1 0 32844 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_334
timestamp 1623621585
transform 1 0 31832 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_343
timestamp 1623621585
transform 1 0 32660 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_1  _334_
timestamp 1623621585
transform 1 0 34132 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _348_
timestamp 1623621585
transform 1 0 35144 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_42_355
timestamp 1623621585
transform 1 0 33764 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_366
timestamp 1623621585
transform 1 0 34776 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _356_
timestamp 1623621585
transform 1 0 36156 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input189
timestamp 1623621585
transform 1 0 37168 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_377
timestamp 1623621585
transform 1 0 35788 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_388
timestamp 1623621585
transform 1 0 36800 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_395
timestamp 1623621585
transform 1 0 37444 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1623621585
transform -1 0 38824 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1623621585
transform 1 0 37812 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_400
timestamp 1623621585
transform 1 0 37904 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1623621585
transform 1 0 38456 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1623621585
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input351
timestamp 1623621585
transform 1 0 1748 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1623621585
transform 1 0 1380 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_11
timestamp 1623621585
transform 1 0 2116 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1623621585
transform 1 0 3772 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_23
timestamp 1623621585
transform 1 0 3220 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_30
timestamp 1623621585
transform 1 0 3864 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_42
timestamp 1623621585
transform 1 0 4968 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_54
timestamp 1623621585
transform 1 0 6072 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_66
timestamp 1623621585
transform 1 0 7176 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_78
timestamp 1623621585
transform 1 0 8280 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1623621585
transform 1 0 9016 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_87
timestamp 1623621585
transform 1 0 9108 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_99
timestamp 1623621585
transform 1 0 10212 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_111
timestamp 1623621585
transform 1 0 11316 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_123
timestamp 1623621585
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1623621585
transform 1 0 14260 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_135
timestamp 1623621585
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_144
timestamp 1623621585
transform 1 0 14352 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_156
timestamp 1623621585
transform 1 0 15456 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_168
timestamp 1623621585
transform 1 0 16560 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_180
timestamp 1623621585
transform 1 0 17664 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1623621585
transform 1 0 19504 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_192
timestamp 1623621585
transform 1 0 18768 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_201
timestamp 1623621585
transform 1 0 19596 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_213
timestamp 1623621585
transform 1 0 20700 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1623621585
transform 1 0 21804 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1623621585
transform 1 0 22908 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_249
timestamp 1623621585
transform 1 0 24012 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1623621585
transform 1 0 24748 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_258
timestamp 1623621585
transform 1 0 24840 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_270
timestamp 1623621585
transform 1 0 25944 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_282
timestamp 1623621585
transform 1 0 27048 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_294
timestamp 1623621585
transform 1 0 28152 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_306
timestamp 1623621585
transform 1 0 29256 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1623621585
transform 1 0 29992 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_315
timestamp 1623621585
transform 1 0 30084 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_327
timestamp 1623621585
transform 1 0 31188 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _562_
timestamp 1623621585
transform 1 0 32752 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_17
timestamp 1623621585
transform 1 0 32568 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_339
timestamp 1623621585
transform 1 0 32292 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_352
timestamp 1623621585
transform 1 0 33488 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1623621585
transform 1 0 35236 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_364
timestamp 1623621585
transform 1 0 34592 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_370
timestamp 1623621585
transform 1 0 35144 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_372
timestamp 1623621585
transform 1 0 35328 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _342_
timestamp 1623621585
transform 1 0 35696 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input157
timestamp 1623621585
transform 1 0 37260 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_383
timestamp 1623621585
transform 1 0 36340 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_391
timestamp 1623621585
transform 1 0 37076 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1623621585
transform -1 0 38824 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input125
timestamp 1623621585
transform 1 0 37904 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_396
timestamp 1623621585
transform 1 0 37536 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1623621585
transform 1 0 38180 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1623621585
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1623621585
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1623621585
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_27
timestamp 1623621585
transform 1 0 3588 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_39
timestamp 1623621585
transform 1 0 4692 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1623621585
transform 1 0 6348 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_51
timestamp 1623621585
transform 1 0 5796 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_58
timestamp 1623621585
transform 1 0 6440 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_70
timestamp 1623621585
transform 1 0 7544 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_82
timestamp 1623621585
transform 1 0 8648 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_94
timestamp 1623621585
transform 1 0 9752 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1623621585
transform 1 0 11592 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_106
timestamp 1623621585
transform 1 0 10856 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_115
timestamp 1623621585
transform 1 0 11684 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_127
timestamp 1623621585
transform 1 0 12788 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_139
timestamp 1623621585
transform 1 0 13892 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_151
timestamp 1623621585
transform 1 0 14996 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_163
timestamp 1623621585
transform 1 0 16100 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1623621585
transform 1 0 16836 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_172
timestamp 1623621585
transform 1 0 16928 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_184
timestamp 1623621585
transform 1 0 18032 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_196
timestamp 1623621585
transform 1 0 19136 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_208
timestamp 1623621585
transform 1 0 20240 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1623621585
transform 1 0 22080 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_220
timestamp 1623621585
transform 1 0 21344 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_229
timestamp 1623621585
transform 1 0 22172 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_241
timestamp 1623621585
transform 1 0 23276 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _807_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 25024 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_44_253
timestamp 1623621585
transform 1 0 24380 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_259
timestamp 1623621585
transform 1 0 24932 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1623621585
transform 1 0 27324 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_279
timestamp 1623621585
transform 1 0 26772 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_286
timestamp 1623621585
transform 1 0 27416 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_298
timestamp 1623621585
transform 1 0 28520 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_310
timestamp 1623621585
transform 1 0 29624 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_322
timestamp 1623621585
transform 1 0 30728 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _556_
timestamp 1623621585
transform 1 0 33028 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1623621585
transform 1 0 32568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE3_1
timestamp 1623621585
transform 1 0 32844 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_334
timestamp 1623621585
transform 1 0 31832 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_343
timestamp 1623621585
transform 1 0 32660 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__a221o_1  _568_
timestamp 1623621585
transform 1 0 34132 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_355
timestamp 1623621585
transform 1 0 33764 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_367
timestamp 1623621585
transform 1 0 34868 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input190
timestamp 1623621585
transform 1 0 37168 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_379
timestamp 1623621585
transform 1 0 35972 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_391
timestamp 1623621585
transform 1 0 37076 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_395
timestamp 1623621585
transform 1 0 37444 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1623621585
transform -1 0 38824 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1623621585
transform 1 0 37812 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_400
timestamp 1623621585
transform 1 0 37904 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_406
timestamp 1623621585
transform 1 0 38456 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1623621585
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input362
timestamp 1623621585
transform 1 0 1748 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1623621585
transform 1 0 1380 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_11
timestamp 1623621585
transform 1 0 2116 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1623621585
transform 1 0 3772 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_23
timestamp 1623621585
transform 1 0 3220 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_30
timestamp 1623621585
transform 1 0 3864 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_42
timestamp 1623621585
transform 1 0 4968 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_54
timestamp 1623621585
transform 1 0 6072 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_66
timestamp 1623621585
transform 1 0 7176 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_78
timestamp 1623621585
transform 1 0 8280 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1623621585
transform 1 0 9016 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_87
timestamp 1623621585
transform 1 0 9108 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_99
timestamp 1623621585
transform 1 0 10212 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_111
timestamp 1623621585
transform 1 0 11316 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1623621585
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1623621585
transform 1 0 14260 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_135
timestamp 1623621585
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_144
timestamp 1623621585
transform 1 0 14352 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_156
timestamp 1623621585
transform 1 0 15456 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_168
timestamp 1623621585
transform 1 0 16560 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_180
timestamp 1623621585
transform 1 0 17664 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1623621585
transform 1 0 19504 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_192
timestamp 1623621585
transform 1 0 18768 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_201
timestamp 1623621585
transform 1 0 19596 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_213
timestamp 1623621585
transform 1 0 20700 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1623621585
transform 1 0 21804 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1623621585
transform 1 0 22908 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_249
timestamp 1623621585
transform 1 0 24012 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1623621585
transform 1 0 25208 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1623621585
transform 1 0 24748 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_258
timestamp 1623621585
transform 1 0 24840 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_265
timestamp 1623621585
transform 1 0 25484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _312_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 26588 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1623621585
transform 1 0 26956 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1623621585
transform 1 0 28060 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_305
timestamp 1623621585
transform 1 0 29164 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _804_
timestamp 1623621585
transform 1 0 30452 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1623621585
transform 1 0 29992 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_313
timestamp 1623621585
transform 1 0 29900 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_315
timestamp 1623621585
transform 1 0 30084 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _550_
timestamp 1623621585
transform 1 0 32752 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_18
timestamp 1623621585
transform 1 0 32568 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_338
timestamp 1623621585
transform 1 0 32200 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_352
timestamp 1623621585
transform 1 0 33488 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1623621585
transform 1 0 35236 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_364
timestamp 1623621585
transform 1 0 34592 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_370
timestamp 1623621585
transform 1 0 35144 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_372
timestamp 1623621585
transform 1 0 35328 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_384
timestamp 1623621585
transform 1 0 36432 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1623621585
transform -1 0 38824 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input126
timestamp 1623621585
transform 1 0 37904 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_396
timestamp 1623621585
transform 1 0 37536 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_403
timestamp 1623621585
transform 1 0 38180 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1623621585
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1623621585
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input373
timestamp 1623621585
transform 1 0 1748 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input376
timestamp 1623621585
transform 1 0 1748 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1623621585
transform 1 0 1380 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_11
timestamp 1623621585
transform 1 0 2116 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1623621585
transform 1 0 1380 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_11
timestamp 1623621585
transform 1 0 2116 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1623621585
transform 1 0 3772 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_23
timestamp 1623621585
transform 1 0 3220 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_35
timestamp 1623621585
transform 1 0 4324 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_23
timestamp 1623621585
transform 1 0 3220 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_30
timestamp 1623621585
transform 1 0 3864 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1623621585
transform 1 0 6348 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_47
timestamp 1623621585
transform 1 0 5428 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_55
timestamp 1623621585
transform 1 0 6164 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_58
timestamp 1623621585
transform 1 0 6440 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_42
timestamp 1623621585
transform 1 0 4968 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_54
timestamp 1623621585
transform 1 0 6072 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_70
timestamp 1623621585
transform 1 0 7544 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_82
timestamp 1623621585
transform 1 0 8648 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_66
timestamp 1623621585
transform 1 0 7176 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_78
timestamp 1623621585
transform 1 0 8280 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1623621585
transform 1 0 9016 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_94
timestamp 1623621585
transform 1 0 9752 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_87
timestamp 1623621585
transform 1 0 9108 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_99
timestamp 1623621585
transform 1 0 10212 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1623621585
transform 1 0 11592 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_106
timestamp 1623621585
transform 1 0 10856 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_115
timestamp 1623621585
transform 1 0 11684 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_111
timestamp 1623621585
transform 1 0 11316 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1623621585
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1623621585
transform 1 0 14260 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_127
timestamp 1623621585
transform 1 0 12788 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_139
timestamp 1623621585
transform 1 0 13892 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_135
timestamp 1623621585
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_144
timestamp 1623621585
transform 1 0 14352 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_151
timestamp 1623621585
transform 1 0 14996 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_163
timestamp 1623621585
transform 1 0 16100 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_156
timestamp 1623621585
transform 1 0 15456 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1623621585
transform 1 0 16836 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_172
timestamp 1623621585
transform 1 0 16928 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_184
timestamp 1623621585
transform 1 0 18032 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_168
timestamp 1623621585
transform 1 0 16560 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_180
timestamp 1623621585
transform 1 0 17664 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1623621585
transform 1 0 19504 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_196
timestamp 1623621585
transform 1 0 19136 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_208
timestamp 1623621585
transform 1 0 20240 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_192
timestamp 1623621585
transform 1 0 18768 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_201
timestamp 1623621585
transform 1 0 19596 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1623621585
transform 1 0 22080 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_220
timestamp 1623621585
transform 1 0 21344 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_229
timestamp 1623621585
transform 1 0 22172 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_213
timestamp 1623621585
transform 1 0 20700 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1623621585
transform 1 0 21804 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_241
timestamp 1623621585
transform 1 0 23276 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1623621585
transform 1 0 22908 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_249
timestamp 1623621585
transform 1 0 24012 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1623621585
transform 1 0 24748 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1623621585
transform 1 0 24380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1623621585
transform 1 0 25484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_258
timestamp 1623621585
transform 1 0 24840 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_270
timestamp 1623621585
transform 1 0 25944 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _311_
timestamp 1623621585
transform 1 0 26772 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 27784 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1623621585
transform 1 0 27324 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_277
timestamp 1623621585
transform 1 0 26588 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_286
timestamp 1623621585
transform 1 0 27416 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_278
timestamp 1623621585
transform 1 0 26680 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_288
timestamp 1623621585
transform 1 0 27600 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_295
timestamp 1623621585
transform 1 0 28244 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_307
timestamp 1623621585
transform 1 0 29348 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_300
timestamp 1623621585
transform 1 0 28704 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_312
timestamp 1623621585
transform 1 0 29808 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1623621585
transform 1 0 29992 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_319
timestamp 1623621585
transform 1 0 30452 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_331
timestamp 1623621585
transform 1 0 31556 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_315
timestamp 1623621585
transform 1 0 30084 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_327
timestamp 1623621585
transform 1 0 31188 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _537_
timestamp 1623621585
transform 1 0 32752 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _543_
timestamp 1623621585
transform 1 0 33028 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1623621585
transform 1 0 32568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_19
timestamp 1623621585
transform 1 0 32844 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_20
timestamp 1623621585
transform 1 0 32568 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_339
timestamp 1623621585
transform 1 0 32292 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_343
timestamp 1623621585
transform 1 0 32660 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_339
timestamp 1623621585
transform 1 0 32292 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_352
timestamp 1623621585
transform 1 0 33488 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1623621585
transform 1 0 35236 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_355
timestamp 1623621585
transform 1 0 33764 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_367
timestamp 1623621585
transform 1 0 34868 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_364
timestamp 1623621585
transform 1 0 34592 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_370
timestamp 1623621585
transform 1 0 35144 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_372
timestamp 1623621585
transform 1 0 35328 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input158
timestamp 1623621585
transform 1 0 37168 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input160
timestamp 1623621585
transform 1 0 37260 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_379
timestamp 1623621585
transform 1 0 35972 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_391
timestamp 1623621585
transform 1 0 37076 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_395
timestamp 1623621585
transform 1 0 37444 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_384
timestamp 1623621585
transform 1 0 36432 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_392
timestamp 1623621585
transform 1 0 37168 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1623621585
transform -1 0 38824 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1623621585
transform -1 0 38824 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1623621585
transform 1 0 37812 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input128
timestamp 1623621585
transform 1 0 37904 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_400
timestamp 1623621585
transform 1 0 37904 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_406
timestamp 1623621585
transform 1 0 38456 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_396
timestamp 1623621585
transform 1 0 37536 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_403
timestamp 1623621585
transform 1 0 38180 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1623621585
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1623621585
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1623621585
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_27
timestamp 1623621585
transform 1 0 3588 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_39
timestamp 1623621585
transform 1 0 4692 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1623621585
transform 1 0 6348 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_51
timestamp 1623621585
transform 1 0 5796 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_58
timestamp 1623621585
transform 1 0 6440 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_70
timestamp 1623621585
transform 1 0 7544 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_82
timestamp 1623621585
transform 1 0 8648 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_94
timestamp 1623621585
transform 1 0 9752 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1623621585
transform 1 0 11592 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_106
timestamp 1623621585
transform 1 0 10856 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_115
timestamp 1623621585
transform 1 0 11684 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_127
timestamp 1623621585
transform 1 0 12788 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_139
timestamp 1623621585
transform 1 0 13892 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_151
timestamp 1623621585
transform 1 0 14996 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_163
timestamp 1623621585
transform 1 0 16100 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1623621585
transform 1 0 16836 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_172
timestamp 1623621585
transform 1 0 16928 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_184
timestamp 1623621585
transform 1 0 18032 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_196
timestamp 1623621585
transform 1 0 19136 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_208
timestamp 1623621585
transform 1 0 20240 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1623621585
transform 1 0 22080 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_220
timestamp 1623621585
transform 1 0 21344 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_229
timestamp 1623621585
transform 1 0 22172 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_241
timestamp 1623621585
transform 1 0 23276 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1623621585
transform 1 0 24380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1623621585
transform 1 0 25484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1623621585
transform 1 0 27324 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_277
timestamp 1623621585
transform 1 0 26588 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_286
timestamp 1623621585
transform 1 0 27416 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_298
timestamp 1623621585
transform 1 0 28520 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_310
timestamp 1623621585
transform 1 0 29624 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_322
timestamp 1623621585
transform 1 0 30728 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1623621585
transform 1 0 32568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_334
timestamp 1623621585
transform 1 0 31832 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_343
timestamp 1623621585
transform 1 0 32660 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_355
timestamp 1623621585
transform 1 0 33764 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_367
timestamp 1623621585
transform 1 0 34868 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_379
timestamp 1623621585
transform 1 0 35972 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_391
timestamp 1623621585
transform 1 0 37076 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1623621585
transform -1 0 38824 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1623621585
transform 1 0 37812 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_400
timestamp 1623621585
transform 1 0 37904 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_406
timestamp 1623621585
transform 1 0 38456 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1623621585
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input377
timestamp 1623621585
transform 1 0 1748 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1623621585
transform 1 0 1380 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_11
timestamp 1623621585
transform 1 0 2116 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1623621585
transform 1 0 3772 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_23
timestamp 1623621585
transform 1 0 3220 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_30
timestamp 1623621585
transform 1 0 3864 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_42
timestamp 1623621585
transform 1 0 4968 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_54
timestamp 1623621585
transform 1 0 6072 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_66
timestamp 1623621585
transform 1 0 7176 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_78
timestamp 1623621585
transform 1 0 8280 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1623621585
transform 1 0 9016 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_87
timestamp 1623621585
transform 1 0 9108 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_99
timestamp 1623621585
transform 1 0 10212 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_111
timestamp 1623621585
transform 1 0 11316 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_123
timestamp 1623621585
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1623621585
transform 1 0 14260 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_135
timestamp 1623621585
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_144
timestamp 1623621585
transform 1 0 14352 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_156
timestamp 1623621585
transform 1 0 15456 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_168
timestamp 1623621585
transform 1 0 16560 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_180
timestamp 1623621585
transform 1 0 17664 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1623621585
transform 1 0 19504 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_192
timestamp 1623621585
transform 1 0 18768 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_201
timestamp 1623621585
transform 1 0 19596 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_213
timestamp 1623621585
transform 1 0 20700 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1623621585
transform 1 0 21804 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1623621585
transform 1 0 22908 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_249
timestamp 1623621585
transform 1 0 24012 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1623621585
transform 1 0 24748 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_258
timestamp 1623621585
transform 1 0 24840 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_270
timestamp 1623621585
transform 1 0 25944 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_282
timestamp 1623621585
transform 1 0 27048 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_294
timestamp 1623621585
transform 1 0 28152 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_306
timestamp 1623621585
transform 1 0 29256 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1623621585
transform 1 0 29992 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_315
timestamp 1623621585
transform 1 0 30084 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_327
timestamp 1623621585
transform 1 0 31188 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_339
timestamp 1623621585
transform 1 0 32292 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_351
timestamp 1623621585
transform 1 0 33396 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1623621585
transform 1 0 35236 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_363
timestamp 1623621585
transform 1 0 34500 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_372
timestamp 1623621585
transform 1 0 35328 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input161
timestamp 1623621585
transform 1 0 37260 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 1623621585
transform 1 0 36432 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_392
timestamp 1623621585
transform 1 0 37168 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1623621585
transform -1 0 38824 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input96
timestamp 1623621585
transform 1 0 37904 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_396
timestamp 1623621585
transform 1 0 37536 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_403
timestamp 1623621585
transform 1 0 38180 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1623621585
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input378
timestamp 1623621585
transform 1 0 1748 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1623621585
transform 1 0 1380 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_11
timestamp 1623621585
transform 1 0 2116 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_23
timestamp 1623621585
transform 1 0 3220 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_35
timestamp 1623621585
transform 1 0 4324 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1623621585
transform 1 0 6348 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_47
timestamp 1623621585
transform 1 0 5428 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_55
timestamp 1623621585
transform 1 0 6164 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_58
timestamp 1623621585
transform 1 0 6440 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_70
timestamp 1623621585
transform 1 0 7544 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_82
timestamp 1623621585
transform 1 0 8648 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_94
timestamp 1623621585
transform 1 0 9752 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1623621585
transform 1 0 11592 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_106
timestamp 1623621585
transform 1 0 10856 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_115
timestamp 1623621585
transform 1 0 11684 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_127
timestamp 1623621585
transform 1 0 12788 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_139
timestamp 1623621585
transform 1 0 13892 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_151
timestamp 1623621585
transform 1 0 14996 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_163
timestamp 1623621585
transform 1 0 16100 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1623621585
transform 1 0 16836 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_172
timestamp 1623621585
transform 1 0 16928 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_184
timestamp 1623621585
transform 1 0 18032 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_196
timestamp 1623621585
transform 1 0 19136 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_208
timestamp 1623621585
transform 1 0 20240 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1623621585
transform 1 0 22080 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_220
timestamp 1623621585
transform 1 0 21344 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_229
timestamp 1623621585
transform 1 0 22172 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_241
timestamp 1623621585
transform 1 0 23276 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1623621585
transform 1 0 24380 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1623621585
transform 1 0 25484 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1623621585
transform 1 0 27324 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_277
timestamp 1623621585
transform 1 0 26588 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_286
timestamp 1623621585
transform 1 0 27416 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_298
timestamp 1623621585
transform 1 0 28520 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_310
timestamp 1623621585
transform 1 0 29624 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_322
timestamp 1623621585
transform 1 0 30728 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1623621585
transform 1 0 32568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_334
timestamp 1623621585
transform 1 0 31832 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_343
timestamp 1623621585
transform 1 0 32660 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_355
timestamp 1623621585
transform 1 0 33764 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_367
timestamp 1623621585
transform 1 0 34868 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_379
timestamp 1623621585
transform 1 0 35972 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_391
timestamp 1623621585
transform 1 0 37076 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1623621585
transform -1 0 38824 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1623621585
transform 1 0 37812 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_400
timestamp 1623621585
transform 1 0 37904 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_406
timestamp 1623621585
transform 1 0 38456 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1623621585
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1623621585
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1623621585
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1623621585
transform 1 0 3772 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_27
timestamp 1623621585
transform 1 0 3588 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_30
timestamp 1623621585
transform 1 0 3864 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_42
timestamp 1623621585
transform 1 0 4968 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_54
timestamp 1623621585
transform 1 0 6072 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_66
timestamp 1623621585
transform 1 0 7176 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_78
timestamp 1623621585
transform 1 0 8280 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1623621585
transform 1 0 9016 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_87
timestamp 1623621585
transform 1 0 9108 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_99
timestamp 1623621585
transform 1 0 10212 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_111
timestamp 1623621585
transform 1 0 11316 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_123
timestamp 1623621585
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1623621585
transform 1 0 14260 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_135
timestamp 1623621585
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_144
timestamp 1623621585
transform 1 0 14352 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_156
timestamp 1623621585
transform 1 0 15456 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_168
timestamp 1623621585
transform 1 0 16560 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_180
timestamp 1623621585
transform 1 0 17664 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1623621585
transform 1 0 19504 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_192
timestamp 1623621585
transform 1 0 18768 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_201
timestamp 1623621585
transform 1 0 19596 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_213
timestamp 1623621585
transform 1 0 20700 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1623621585
transform 1 0 21804 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1623621585
transform 1 0 22908 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_249
timestamp 1623621585
transform 1 0 24012 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1623621585
transform 1 0 24748 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_258
timestamp 1623621585
transform 1 0 24840 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_270
timestamp 1623621585
transform 1 0 25944 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_282
timestamp 1623621585
transform 1 0 27048 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_294
timestamp 1623621585
transform 1 0 28152 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_306
timestamp 1623621585
transform 1 0 29256 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_793
timestamp 1623621585
transform 1 0 29992 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_315
timestamp 1623621585
transform 1 0 30084 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_327
timestamp 1623621585
transform 1 0 31188 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _523_
timestamp 1623621585
transform 1 0 32844 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_21
timestamp 1623621585
transform 1 0 32660 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_339
timestamp 1623621585
transform 1 0 32292 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_353
timestamp 1623621585
transform 1 0 33580 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_794
timestamp 1623621585
transform 1 0 35236 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_365
timestamp 1623621585
transform 1 0 34684 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_372
timestamp 1623621585
transform 1 0 35328 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input129
timestamp 1623621585
transform 1 0 37260 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_384
timestamp 1623621585
transform 1 0 36432 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_392
timestamp 1623621585
transform 1 0 37168 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1623621585
transform -1 0 38824 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input97
timestamp 1623621585
transform 1 0 37904 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_396
timestamp 1623621585
transform 1 0 37536 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1623621585
transform 1 0 38180 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1623621585
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1623621585
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input379
timestamp 1623621585
transform 1 0 1748 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input380
timestamp 1623621585
transform 1 0 1748 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1623621585
transform 1 0 1380 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_11
timestamp 1623621585
transform 1 0 2116 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_3
timestamp 1623621585
transform 1 0 1380 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_11
timestamp 1623621585
transform 1 0 2116 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_802
timestamp 1623621585
transform 1 0 3772 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_23
timestamp 1623621585
transform 1 0 3220 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_35
timestamp 1623621585
transform 1 0 4324 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_23
timestamp 1623621585
transform 1 0 3220 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_30
timestamp 1623621585
transform 1 0 3864 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_795
timestamp 1623621585
transform 1 0 6348 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_47
timestamp 1623621585
transform 1 0 5428 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_55
timestamp 1623621585
transform 1 0 6164 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_58
timestamp 1623621585
transform 1 0 6440 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_42
timestamp 1623621585
transform 1 0 4968 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_54
timestamp 1623621585
transform 1 0 6072 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_70
timestamp 1623621585
transform 1 0 7544 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_82
timestamp 1623621585
transform 1 0 8648 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_66
timestamp 1623621585
transform 1 0 7176 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_78
timestamp 1623621585
transform 1 0 8280 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_803
timestamp 1623621585
transform 1 0 9016 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_94
timestamp 1623621585
transform 1 0 9752 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_87
timestamp 1623621585
transform 1 0 9108 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_99
timestamp 1623621585
transform 1 0 10212 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_796
timestamp 1623621585
transform 1 0 11592 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_106
timestamp 1623621585
transform 1 0 10856 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_115
timestamp 1623621585
transform 1 0 11684 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_111
timestamp 1623621585
transform 1 0 11316 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_123
timestamp 1623621585
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_804
timestamp 1623621585
transform 1 0 14260 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_127
timestamp 1623621585
transform 1 0 12788 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_139
timestamp 1623621585
transform 1 0 13892 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_135
timestamp 1623621585
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_144
timestamp 1623621585
transform 1 0 14352 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_151
timestamp 1623621585
transform 1 0 14996 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_163
timestamp 1623621585
transform 1 0 16100 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_156
timestamp 1623621585
transform 1 0 15456 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_797
timestamp 1623621585
transform 1 0 16836 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_172
timestamp 1623621585
transform 1 0 16928 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_184
timestamp 1623621585
transform 1 0 18032 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_168
timestamp 1623621585
transform 1 0 16560 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_180
timestamp 1623621585
transform 1 0 17664 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_805
timestamp 1623621585
transform 1 0 19504 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_196
timestamp 1623621585
transform 1 0 19136 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_208
timestamp 1623621585
transform 1 0 20240 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_192
timestamp 1623621585
transform 1 0 18768 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_201
timestamp 1623621585
transform 1 0 19596 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_798
timestamp 1623621585
transform 1 0 22080 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_220
timestamp 1623621585
transform 1 0 21344 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_229
timestamp 1623621585
transform 1 0 22172 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_213
timestamp 1623621585
transform 1 0 20700 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1623621585
transform 1 0 21804 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_241
timestamp 1623621585
transform 1 0 23276 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1623621585
transform 1 0 22908 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_249
timestamp 1623621585
transform 1 0 24012 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_806
timestamp 1623621585
transform 1 0 24748 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1623621585
transform 1 0 24380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1623621585
transform 1 0 25484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_258
timestamp 1623621585
transform 1 0 24840 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_270
timestamp 1623621585
transform 1 0 25944 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_799
timestamp 1623621585
transform 1 0 27324 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_277
timestamp 1623621585
transform 1 0 26588 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_286
timestamp 1623621585
transform 1 0 27416 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_282
timestamp 1623621585
transform 1 0 27048 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_298
timestamp 1623621585
transform 1 0 28520 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_310
timestamp 1623621585
transform 1 0 29624 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_294
timestamp 1623621585
transform 1 0 28152 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_306
timestamp 1623621585
transform 1 0 29256 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_807
timestamp 1623621585
transform 1 0 29992 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_322
timestamp 1623621585
transform 1 0 30728 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_315
timestamp 1623621585
transform 1 0 30084 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_327
timestamp 1623621585
transform 1 0 31188 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_343
timestamp 1623621585
transform 1 0 32660 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_339
timestamp 1623621585
transform 1 0 32292 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_343
timestamp 1623621585
transform 1 0 32660 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_334
timestamp 1623621585
transform 1 0 31832 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_800
timestamp 1623621585
transform 1 0 32568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_22
timestamp 1623621585
transform 1 0 32844 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_5
timestamp 1623621585
transform 1 0 32752 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__a221o_1  _516_
timestamp 1623621585
transform 1 0 33028 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _510_
timestamp 1623621585
transform 1 0 32936 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_354
timestamp 1623621585
transform 1 0 33672 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_808
timestamp 1623621585
transform 1 0 35236 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_355
timestamp 1623621585
transform 1 0 33764 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_367
timestamp 1623621585
transform 1 0 34868 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_366
timestamp 1623621585
transform 1 0 34776 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_370
timestamp 1623621585
transform 1 0 35144 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_372
timestamp 1623621585
transform 1 0 35328 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input130
timestamp 1623621585
transform 1 0 37260 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input162
timestamp 1623621585
transform 1 0 37168 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_379
timestamp 1623621585
transform 1 0 35972 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_391
timestamp 1623621585
transform 1 0 37076 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_395
timestamp 1623621585
transform 1 0 37444 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_384
timestamp 1623621585
transform 1 0 36432 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_392
timestamp 1623621585
transform 1 0 37168 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1623621585
transform -1 0 38824 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1623621585
transform -1 0 38824 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_801
timestamp 1623621585
transform 1 0 37812 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input98
timestamp 1623621585
transform 1 0 37904 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_400
timestamp 1623621585
transform 1 0 37904 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_406
timestamp 1623621585
transform 1 0 38456 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_396
timestamp 1623621585
transform 1 0 37536 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_403
timestamp 1623621585
transform 1 0 38180 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1623621585
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1623621585
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1623621585
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_27
timestamp 1623621585
transform 1 0 3588 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_39
timestamp 1623621585
transform 1 0 4692 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_809
timestamp 1623621585
transform 1 0 6348 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_51
timestamp 1623621585
transform 1 0 5796 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_58
timestamp 1623621585
transform 1 0 6440 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_70
timestamp 1623621585
transform 1 0 7544 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_82
timestamp 1623621585
transform 1 0 8648 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_94
timestamp 1623621585
transform 1 0 9752 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_810
timestamp 1623621585
transform 1 0 11592 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_106
timestamp 1623621585
transform 1 0 10856 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_115
timestamp 1623621585
transform 1 0 11684 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_127
timestamp 1623621585
transform 1 0 12788 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_139
timestamp 1623621585
transform 1 0 13892 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_151
timestamp 1623621585
transform 1 0 14996 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_163
timestamp 1623621585
transform 1 0 16100 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_811
timestamp 1623621585
transform 1 0 16836 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_172
timestamp 1623621585
transform 1 0 16928 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_184
timestamp 1623621585
transform 1 0 18032 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_196
timestamp 1623621585
transform 1 0 19136 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_208
timestamp 1623621585
transform 1 0 20240 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_812
timestamp 1623621585
transform 1 0 22080 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_220
timestamp 1623621585
transform 1 0 21344 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_229
timestamp 1623621585
transform 1 0 22172 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_241
timestamp 1623621585
transform 1 0 23276 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1623621585
transform 1 0 24380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1623621585
transform 1 0 25484 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_813
timestamp 1623621585
transform 1 0 27324 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_277
timestamp 1623621585
transform 1 0 26588 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_286
timestamp 1623621585
transform 1 0 27416 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_298
timestamp 1623621585
transform 1 0 28520 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_310
timestamp 1623621585
transform 1 0 29624 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_322
timestamp 1623621585
transform 1 0 30728 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _503_
timestamp 1623621585
transform 1 0 33028 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_814
timestamp 1623621585
transform 1 0 32568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_6
timestamp 1623621585
transform 1 0 32844 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_334
timestamp 1623621585
transform 1 0 31832 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_343
timestamp 1623621585
transform 1 0 32660 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_355
timestamp 1623621585
transform 1 0 33764 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_367
timestamp 1623621585
transform 1 0 34868 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input163
timestamp 1623621585
transform 1 0 37168 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_379
timestamp 1623621585
transform 1 0 35972 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_391
timestamp 1623621585
transform 1 0 37076 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_395
timestamp 1623621585
transform 1 0 37444 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1623621585
transform -1 0 38824 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_815
timestamp 1623621585
transform 1 0 37812 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_400
timestamp 1623621585
transform 1 0 37904 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_406
timestamp 1623621585
transform 1 0 38456 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1623621585
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input381
timestamp 1623621585
transform 1 0 1748 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1623621585
transform 1 0 1380 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_11
timestamp 1623621585
transform 1 0 2116 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_816
timestamp 1623621585
transform 1 0 3772 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_23
timestamp 1623621585
transform 1 0 3220 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_30
timestamp 1623621585
transform 1 0 3864 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_42
timestamp 1623621585
transform 1 0 4968 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_54
timestamp 1623621585
transform 1 0 6072 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_66
timestamp 1623621585
transform 1 0 7176 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_78
timestamp 1623621585
transform 1 0 8280 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_817
timestamp 1623621585
transform 1 0 9016 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_87
timestamp 1623621585
transform 1 0 9108 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_99
timestamp 1623621585
transform 1 0 10212 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_111
timestamp 1623621585
transform 1 0 11316 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_123
timestamp 1623621585
transform 1 0 12420 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_818
timestamp 1623621585
transform 1 0 14260 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_135
timestamp 1623621585
transform 1 0 13524 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_144
timestamp 1623621585
transform 1 0 14352 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_156
timestamp 1623621585
transform 1 0 15456 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_168
timestamp 1623621585
transform 1 0 16560 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_180
timestamp 1623621585
transform 1 0 17664 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_819
timestamp 1623621585
transform 1 0 19504 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_192
timestamp 1623621585
transform 1 0 18768 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_201
timestamp 1623621585
transform 1 0 19596 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_213
timestamp 1623621585
transform 1 0 20700 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1623621585
transform 1 0 21804 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1623621585
transform 1 0 22908 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_249
timestamp 1623621585
transform 1 0 24012 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_820
timestamp 1623621585
transform 1 0 24748 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_258
timestamp 1623621585
transform 1 0 24840 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_270
timestamp 1623621585
transform 1 0 25944 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_282
timestamp 1623621585
transform 1 0 27048 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_294
timestamp 1623621585
transform 1 0 28152 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_306
timestamp 1623621585
transform 1 0 29256 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_821
timestamp 1623621585
transform 1 0 29992 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_315
timestamp 1623621585
transform 1 0 30084 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_327
timestamp 1623621585
transform 1 0 31188 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _497_
timestamp 1623621585
transform 1 0 33028 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_7
timestamp 1623621585
transform 1 0 32844 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_339
timestamp 1623621585
transform 1 0 32292 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_822
timestamp 1623621585
transform 1 0 35236 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_355
timestamp 1623621585
transform 1 0 33764 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_367
timestamp 1623621585
transform 1 0 34868 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_372
timestamp 1623621585
transform 1 0 35328 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_384
timestamp 1623621585
transform 1 0 36432 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1623621585
transform -1 0 38824 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 1623621585
transform 1 0 37904 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_396
timestamp 1623621585
transform 1 0 37536 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1623621585
transform 1 0 38180 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1623621585
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input382
timestamp 1623621585
transform 1 0 1748 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_3
timestamp 1623621585
transform 1 0 1380 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_11
timestamp 1623621585
transform 1 0 2116 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_23
timestamp 1623621585
transform 1 0 3220 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_35
timestamp 1623621585
transform 1 0 4324 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_823
timestamp 1623621585
transform 1 0 6348 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_47
timestamp 1623621585
transform 1 0 5428 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_55
timestamp 1623621585
transform 1 0 6164 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_58
timestamp 1623621585
transform 1 0 6440 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_70
timestamp 1623621585
transform 1 0 7544 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_82
timestamp 1623621585
transform 1 0 8648 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_94
timestamp 1623621585
transform 1 0 9752 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_824
timestamp 1623621585
transform 1 0 11592 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_106
timestamp 1623621585
transform 1 0 10856 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_115
timestamp 1623621585
transform 1 0 11684 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_127
timestamp 1623621585
transform 1 0 12788 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_139
timestamp 1623621585
transform 1 0 13892 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_151
timestamp 1623621585
transform 1 0 14996 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_163
timestamp 1623621585
transform 1 0 16100 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_825
timestamp 1623621585
transform 1 0 16836 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_172
timestamp 1623621585
transform 1 0 16928 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_184
timestamp 1623621585
transform 1 0 18032 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_196
timestamp 1623621585
transform 1 0 19136 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_208
timestamp 1623621585
transform 1 0 20240 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_826
timestamp 1623621585
transform 1 0 22080 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_220
timestamp 1623621585
transform 1 0 21344 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_229
timestamp 1623621585
transform 1 0 22172 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_241
timestamp 1623621585
transform 1 0 23276 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1623621585
transform 1 0 24380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1623621585
transform 1 0 25484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_827
timestamp 1623621585
transform 1 0 27324 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_277
timestamp 1623621585
transform 1 0 26588 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_286
timestamp 1623621585
transform 1 0 27416 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_298
timestamp 1623621585
transform 1 0 28520 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_310
timestamp 1623621585
transform 1 0 29624 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_322
timestamp 1623621585
transform 1 0 30728 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_828
timestamp 1623621585
transform 1 0 32568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_334
timestamp 1623621585
transform 1 0 31832 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_343
timestamp 1623621585
transform 1 0 32660 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_355
timestamp 1623621585
transform 1 0 33764 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_367
timestamp 1623621585
transform 1 0 34868 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input131
timestamp 1623621585
transform 1 0 37168 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_379
timestamp 1623621585
transform 1 0 35972 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_391
timestamp 1623621585
transform 1 0 37076 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_395
timestamp 1623621585
transform 1 0 37444 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1623621585
transform -1 0 38824 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_829
timestamp 1623621585
transform 1 0 37812 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_400
timestamp 1623621585
transform 1 0 37904 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_406
timestamp 1623621585
transform 1 0 38456 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1623621585
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1623621585
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1623621585
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_830
timestamp 1623621585
transform 1 0 3772 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_27
timestamp 1623621585
transform 1 0 3588 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_30
timestamp 1623621585
transform 1 0 3864 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_42
timestamp 1623621585
transform 1 0 4968 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_54
timestamp 1623621585
transform 1 0 6072 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_66
timestamp 1623621585
transform 1 0 7176 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_78
timestamp 1623621585
transform 1 0 8280 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_831
timestamp 1623621585
transform 1 0 9016 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_87
timestamp 1623621585
transform 1 0 9108 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_99
timestamp 1623621585
transform 1 0 10212 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_111
timestamp 1623621585
transform 1 0 11316 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_123
timestamp 1623621585
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_832
timestamp 1623621585
transform 1 0 14260 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_135
timestamp 1623621585
transform 1 0 13524 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_144
timestamp 1623621585
transform 1 0 14352 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_156
timestamp 1623621585
transform 1 0 15456 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_168
timestamp 1623621585
transform 1 0 16560 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_180
timestamp 1623621585
transform 1 0 17664 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_833
timestamp 1623621585
transform 1 0 19504 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_192
timestamp 1623621585
transform 1 0 18768 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_201
timestamp 1623621585
transform 1 0 19596 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_213
timestamp 1623621585
transform 1 0 20700 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1623621585
transform 1 0 21804 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1623621585
transform 1 0 22908 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_249
timestamp 1623621585
transform 1 0 24012 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_834
timestamp 1623621585
transform 1 0 24748 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_258
timestamp 1623621585
transform 1 0 24840 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_270
timestamp 1623621585
transform 1 0 25944 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_282
timestamp 1623621585
transform 1 0 27048 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _532_
timestamp 1623621585
transform 1 0 28612 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_294
timestamp 1623621585
transform 1 0 28152 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_298
timestamp 1623621585
transform 1 0 28520 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_303
timestamp 1623621585
transform 1 0 28980 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_311
timestamp 1623621585
transform 1 0 29716 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_835
timestamp 1623621585
transform 1 0 29992 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_315
timestamp 1623621585
transform 1 0 30084 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_327
timestamp 1623621585
transform 1 0 31188 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _533_
timestamp 1623621585
transform 1 0 33580 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_339
timestamp 1623621585
transform 1 0 32292 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_351
timestamp 1623621585
transform 1 0 33396 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_836
timestamp 1623621585
transform 1 0 35236 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_357
timestamp 1623621585
transform 1 0 33948 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_369
timestamp 1623621585
transform 1 0 35052 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_372
timestamp 1623621585
transform 1 0 35328 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input164
timestamp 1623621585
transform 1 0 37260 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_384
timestamp 1623621585
transform 1 0 36432 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_392
timestamp 1623621585
transform 1 0 37168 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1623621585
transform -1 0 38824 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input100
timestamp 1623621585
transform 1 0 37904 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_396
timestamp 1623621585
transform 1 0 37536 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1623621585
transform 1 0 38180 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1623621585
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input352
timestamp 1623621585
transform 1 0 1748 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_3
timestamp 1623621585
transform 1 0 1380 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_11
timestamp 1623621585
transform 1 0 2116 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_23
timestamp 1623621585
transform 1 0 3220 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_35
timestamp 1623621585
transform 1 0 4324 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_837
timestamp 1623621585
transform 1 0 6348 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_47
timestamp 1623621585
transform 1 0 5428 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_55
timestamp 1623621585
transform 1 0 6164 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_58
timestamp 1623621585
transform 1 0 6440 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_70
timestamp 1623621585
transform 1 0 7544 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_82
timestamp 1623621585
transform 1 0 8648 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_94
timestamp 1623621585
transform 1 0 9752 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_838
timestamp 1623621585
transform 1 0 11592 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_106
timestamp 1623621585
transform 1 0 10856 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_115
timestamp 1623621585
transform 1 0 11684 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_127
timestamp 1623621585
transform 1 0 12788 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_139
timestamp 1623621585
transform 1 0 13892 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_151
timestamp 1623621585
transform 1 0 14996 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_163
timestamp 1623621585
transform 1 0 16100 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_839
timestamp 1623621585
transform 1 0 16836 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_172
timestamp 1623621585
transform 1 0 16928 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_184
timestamp 1623621585
transform 1 0 18032 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_196
timestamp 1623621585
transform 1 0 19136 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_208
timestamp 1623621585
transform 1 0 20240 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_840
timestamp 1623621585
transform 1 0 22080 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_220
timestamp 1623621585
transform 1 0 21344 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_229
timestamp 1623621585
transform 1 0 22172 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_241
timestamp 1623621585
transform 1 0 23276 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1623621585
transform 1 0 24380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1623621585
transform 1 0 25484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_841
timestamp 1623621585
transform 1 0 27324 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_277
timestamp 1623621585
transform 1 0 26588 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_286
timestamp 1623621585
transform 1 0 27416 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_298
timestamp 1623621585
transform 1 0 28520 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_310
timestamp 1623621585
transform 1 0 29624 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_322
timestamp 1623621585
transform 1 0 30728 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_842
timestamp 1623621585
transform 1 0 32568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_334
timestamp 1623621585
transform 1 0 31832 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_343
timestamp 1623621585
transform 1 0 32660 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_355
timestamp 1623621585
transform 1 0 33764 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_367
timestamp 1623621585
transform 1 0 34868 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_379
timestamp 1623621585
transform 1 0 35972 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_391
timestamp 1623621585
transform 1 0 37076 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1623621585
transform -1 0 38824 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_843
timestamp 1623621585
transform 1 0 37812 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_400
timestamp 1623621585
transform 1 0 37904 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1623621585
transform 1 0 38456 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1623621585
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1623621585
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input353
timestamp 1623621585
transform 1 0 1748 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1623621585
transform 1 0 1380 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_11
timestamp 1623621585
transform 1 0 2116 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1623621585
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1623621585
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_844
timestamp 1623621585
transform 1 0 3772 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_23
timestamp 1623621585
transform 1 0 3220 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_30
timestamp 1623621585
transform 1 0 3864 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_27
timestamp 1623621585
transform 1 0 3588 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_39
timestamp 1623621585
transform 1 0 4692 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_851
timestamp 1623621585
transform 1 0 6348 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_42
timestamp 1623621585
transform 1 0 4968 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_54
timestamp 1623621585
transform 1 0 6072 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_51
timestamp 1623621585
transform 1 0 5796 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_58
timestamp 1623621585
transform 1 0 6440 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_66
timestamp 1623621585
transform 1 0 7176 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_78
timestamp 1623621585
transform 1 0 8280 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_70
timestamp 1623621585
transform 1 0 7544 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_82
timestamp 1623621585
transform 1 0 8648 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_845
timestamp 1623621585
transform 1 0 9016 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_87
timestamp 1623621585
transform 1 0 9108 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_99
timestamp 1623621585
transform 1 0 10212 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_94
timestamp 1623621585
transform 1 0 9752 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_852
timestamp 1623621585
transform 1 0 11592 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_111
timestamp 1623621585
transform 1 0 11316 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_123
timestamp 1623621585
transform 1 0 12420 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_106
timestamp 1623621585
transform 1 0 10856 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_115
timestamp 1623621585
transform 1 0 11684 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_846
timestamp 1623621585
transform 1 0 14260 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_135
timestamp 1623621585
transform 1 0 13524 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_144
timestamp 1623621585
transform 1 0 14352 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_127
timestamp 1623621585
transform 1 0 12788 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_139
timestamp 1623621585
transform 1 0 13892 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_156
timestamp 1623621585
transform 1 0 15456 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_151
timestamp 1623621585
transform 1 0 14996 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_163
timestamp 1623621585
transform 1 0 16100 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_853
timestamp 1623621585
transform 1 0 16836 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_168
timestamp 1623621585
transform 1 0 16560 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_180
timestamp 1623621585
transform 1 0 17664 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_172
timestamp 1623621585
transform 1 0 16928 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_184
timestamp 1623621585
transform 1 0 18032 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_847
timestamp 1623621585
transform 1 0 19504 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_192
timestamp 1623621585
transform 1 0 18768 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_201
timestamp 1623621585
transform 1 0 19596 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_196
timestamp 1623621585
transform 1 0 19136 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_208
timestamp 1623621585
transform 1 0 20240 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_854
timestamp 1623621585
transform 1 0 22080 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_213
timestamp 1623621585
transform 1 0 20700 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1623621585
transform 1 0 21804 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_220
timestamp 1623621585
transform 1 0 21344 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_229
timestamp 1623621585
transform 1 0 22172 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1623621585
transform 1 0 22908 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_249
timestamp 1623621585
transform 1 0 24012 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_241
timestamp 1623621585
transform 1 0 23276 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_848
timestamp 1623621585
transform 1 0 24748 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_258
timestamp 1623621585
transform 1 0 24840 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_270
timestamp 1623621585
transform 1 0 25944 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1623621585
transform 1 0 24380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1623621585
transform 1 0 25484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_855
timestamp 1623621585
transform 1 0 27324 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_282
timestamp 1623621585
transform 1 0 27048 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_277
timestamp 1623621585
transform 1 0 26588 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_286
timestamp 1623621585
transform 1 0 27416 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_294
timestamp 1623621585
transform 1 0 28152 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_306
timestamp 1623621585
transform 1 0 29256 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_298
timestamp 1623621585
transform 1 0 28520 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_310
timestamp 1623621585
transform 1 0 29624 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_849
timestamp 1623621585
transform 1 0 29992 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_315
timestamp 1623621585
transform 1 0 30084 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_327
timestamp 1623621585
transform 1 0 31188 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_322
timestamp 1623621585
transform 1 0 30728 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _483_
timestamp 1623621585
transform 1 0 33120 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_856
timestamp 1623621585
transform 1 0 32568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_8
timestamp 1623621585
transform 1 0 32936 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_339
timestamp 1623621585
transform 1 0 32292 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_351
timestamp 1623621585
transform 1 0 33396 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_334
timestamp 1623621585
transform 1 0 31832 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_343
timestamp 1623621585
transform 1 0 32660 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _493_
timestamp 1623621585
transform 1 0 34224 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_850
timestamp 1623621585
transform 1 0 35236 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_363
timestamp 1623621585
transform 1 0 34500 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_372
timestamp 1623621585
transform 1 0 35328 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_356
timestamp 1623621585
transform 1 0 33856 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_364
timestamp 1623621585
transform 1 0 34592 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input165
timestamp 1623621585
transform 1 0 37260 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_384
timestamp 1623621585
transform 1 0 36432 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_392
timestamp 1623621585
transform 1 0 37168 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_376
timestamp 1623621585
transform 1 0 35696 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_388
timestamp 1623621585
transform 1 0 36800 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1623621585
transform -1 0 38824 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1623621585
transform -1 0 38824 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_857
timestamp 1623621585
transform 1 0 37812 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input132
timestamp 1623621585
transform 1 0 37904 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_396
timestamp 1623621585
transform 1 0 37536 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_403
timestamp 1623621585
transform 1 0 38180 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_396
timestamp 1623621585
transform 1 0 37536 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_400
timestamp 1623621585
transform 1 0 37904 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_406
timestamp 1623621585
transform 1 0 38456 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1623621585
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input354
timestamp 1623621585
transform 1 0 1748 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1623621585
transform 1 0 1380 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_11
timestamp 1623621585
transform 1 0 2116 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_858
timestamp 1623621585
transform 1 0 3772 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_23
timestamp 1623621585
transform 1 0 3220 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1623621585
transform 1 0 3864 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1623621585
transform 1 0 4968 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_54
timestamp 1623621585
transform 1 0 6072 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_66
timestamp 1623621585
transform 1 0 7176 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_78
timestamp 1623621585
transform 1 0 8280 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_859
timestamp 1623621585
transform 1 0 9016 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_87
timestamp 1623621585
transform 1 0 9108 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_99
timestamp 1623621585
transform 1 0 10212 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_111
timestamp 1623621585
transform 1 0 11316 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_123
timestamp 1623621585
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_860
timestamp 1623621585
transform 1 0 14260 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_135
timestamp 1623621585
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_144
timestamp 1623621585
transform 1 0 14352 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_156
timestamp 1623621585
transform 1 0 15456 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_168
timestamp 1623621585
transform 1 0 16560 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_180
timestamp 1623621585
transform 1 0 17664 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_861
timestamp 1623621585
transform 1 0 19504 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_192
timestamp 1623621585
transform 1 0 18768 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_201
timestamp 1623621585
transform 1 0 19596 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_213
timestamp 1623621585
transform 1 0 20700 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1623621585
transform 1 0 21804 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1623621585
transform 1 0 22908 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_249
timestamp 1623621585
transform 1 0 24012 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_862
timestamp 1623621585
transform 1 0 24748 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_258
timestamp 1623621585
transform 1 0 24840 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_270
timestamp 1623621585
transform 1 0 25944 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_282
timestamp 1623621585
transform 1 0 27048 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _492_
timestamp 1623621585
transform 1 0 28704 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_294
timestamp 1623621585
transform 1 0 28152 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_304
timestamp 1623621585
transform 1 0 29072 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_312
timestamp 1623621585
transform 1 0 29808 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_863
timestamp 1623621585
transform 1 0 29992 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_315
timestamp 1623621585
transform 1 0 30084 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_327
timestamp 1623621585
transform 1 0 31188 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _476_
timestamp 1623621585
transform 1 0 33212 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_9
timestamp 1623621585
transform 1 0 33028 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_339
timestamp 1623621585
transform 1 0 32292 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _370_
timestamp 1623621585
transform 1 0 34316 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_864
timestamp 1623621585
transform 1 0 35236 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_357
timestamp 1623621585
transform 1 0 33948 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_365
timestamp 1623621585
transform 1 0 34684 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_372
timestamp 1623621585
transform 1 0 35328 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input133
timestamp 1623621585
transform 1 0 37260 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_384
timestamp 1623621585
transform 1 0 36432 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_392
timestamp 1623621585
transform 1 0 37168 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1623621585
transform -1 0 38824 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input101
timestamp 1623621585
transform 1 0 37904 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_396
timestamp 1623621585
transform 1 0 37536 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_403
timestamp 1623621585
transform 1 0 38180 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1623621585
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input355
timestamp 1623621585
transform 1 0 1748 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_3
timestamp 1623621585
transform 1 0 1380 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_11
timestamp 1623621585
transform 1 0 2116 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_23
timestamp 1623621585
transform 1 0 3220 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_35
timestamp 1623621585
transform 1 0 4324 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_865
timestamp 1623621585
transform 1 0 6348 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_47
timestamp 1623621585
transform 1 0 5428 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_55
timestamp 1623621585
transform 1 0 6164 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_58
timestamp 1623621585
transform 1 0 6440 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_70
timestamp 1623621585
transform 1 0 7544 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_82
timestamp 1623621585
transform 1 0 8648 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_94
timestamp 1623621585
transform 1 0 9752 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_866
timestamp 1623621585
transform 1 0 11592 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_106
timestamp 1623621585
transform 1 0 10856 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_115
timestamp 1623621585
transform 1 0 11684 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_127
timestamp 1623621585
transform 1 0 12788 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_139
timestamp 1623621585
transform 1 0 13892 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_151
timestamp 1623621585
transform 1 0 14996 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_163
timestamp 1623621585
transform 1 0 16100 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_867
timestamp 1623621585
transform 1 0 16836 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_172
timestamp 1623621585
transform 1 0 16928 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_184
timestamp 1623621585
transform 1 0 18032 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_196
timestamp 1623621585
transform 1 0 19136 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_208
timestamp 1623621585
transform 1 0 20240 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_868
timestamp 1623621585
transform 1 0 22080 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_220
timestamp 1623621585
transform 1 0 21344 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_229
timestamp 1623621585
transform 1 0 22172 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_241
timestamp 1623621585
transform 1 0 23276 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1623621585
transform 1 0 24380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1623621585
transform 1 0 25484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_869
timestamp 1623621585
transform 1 0 27324 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_277
timestamp 1623621585
transform 1 0 26588 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_286
timestamp 1623621585
transform 1 0 27416 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _368_
timestamp 1623621585
transform 1 0 28612 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_298
timestamp 1623621585
transform 1 0 28520 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_303
timestamp 1623621585
transform 1 0 28980 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_315
timestamp 1623621585
transform 1 0 30084 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_327
timestamp 1623621585
transform 1 0 31188 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _470_
timestamp 1623621585
transform 1 0 33212 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_870
timestamp 1623621585
transform 1 0 32568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_10
timestamp 1623621585
transform 1 0 33028 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_339
timestamp 1623621585
transform 1 0 32292 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_343
timestamp 1623621585
transform 1 0 32660 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _412_
timestamp 1623621585
transform 1 0 34316 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_357
timestamp 1623621585
transform 1 0 33948 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1623621585
transform 1 0 34684 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input166
timestamp 1623621585
transform 1 0 37168 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1623621585
transform 1 0 35788 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_389
timestamp 1623621585
transform 1 0 36892 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_395
timestamp 1623621585
transform 1 0 37444 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1623621585
transform -1 0 38824 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_871
timestamp 1623621585
transform 1 0 37812 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_400
timestamp 1623621585
transform 1 0 37904 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_406
timestamp 1623621585
transform 1 0 38456 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1623621585
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1623621585
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1623621585
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_872
timestamp 1623621585
transform 1 0 3772 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_27
timestamp 1623621585
transform 1 0 3588 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_30
timestamp 1623621585
transform 1 0 3864 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_42
timestamp 1623621585
transform 1 0 4968 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_54
timestamp 1623621585
transform 1 0 6072 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_66
timestamp 1623621585
transform 1 0 7176 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_78
timestamp 1623621585
transform 1 0 8280 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_873
timestamp 1623621585
transform 1 0 9016 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_87
timestamp 1623621585
transform 1 0 9108 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_99
timestamp 1623621585
transform 1 0 10212 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_111
timestamp 1623621585
transform 1 0 11316 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1623621585
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_874
timestamp 1623621585
transform 1 0 14260 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_135
timestamp 1623621585
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_144
timestamp 1623621585
transform 1 0 14352 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_156
timestamp 1623621585
transform 1 0 15456 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_168
timestamp 1623621585
transform 1 0 16560 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_180
timestamp 1623621585
transform 1 0 17664 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_875
timestamp 1623621585
transform 1 0 19504 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_192
timestamp 1623621585
transform 1 0 18768 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_201
timestamp 1623621585
transform 1 0 19596 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_213
timestamp 1623621585
transform 1 0 20700 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1623621585
transform 1 0 21804 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1623621585
transform 1 0 22908 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_249
timestamp 1623621585
transform 1 0 24012 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_876
timestamp 1623621585
transform 1 0 24748 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_258
timestamp 1623621585
transform 1 0 24840 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_270
timestamp 1623621585
transform 1 0 25944 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_282
timestamp 1623621585
transform 1 0 27048 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_294
timestamp 1623621585
transform 1 0 28152 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_306
timestamp 1623621585
transform 1 0 29256 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_877
timestamp 1623621585
transform 1 0 29992 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_315
timestamp 1623621585
transform 1 0 30084 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_327
timestamp 1623621585
transform 1 0 31188 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _463_
timestamp 1623621585
transform 1 0 33212 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_11
timestamp 1623621585
transform 1 0 33028 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_339
timestamp 1623621585
transform 1 0 32292 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _413_
timestamp 1623621585
transform 1 0 34316 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_878
timestamp 1623621585
transform 1 0 35236 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_357
timestamp 1623621585
transform 1 0 33948 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_365
timestamp 1623621585
transform 1 0 34684 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_372
timestamp 1623621585
transform 1 0 35328 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input134
timestamp 1623621585
transform 1 0 37260 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_384
timestamp 1623621585
transform 1 0 36432 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_392
timestamp 1623621585
transform 1 0 37168 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1623621585
transform -1 0 38824 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input102
timestamp 1623621585
transform 1 0 37904 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_396
timestamp 1623621585
transform 1 0 37536 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1623621585
transform 1 0 38180 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1623621585
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input356
timestamp 1623621585
transform 1 0 1748 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1623621585
transform 1 0 1380 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_11
timestamp 1623621585
transform 1 0 2116 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_23
timestamp 1623621585
transform 1 0 3220 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_35
timestamp 1623621585
transform 1 0 4324 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_879
timestamp 1623621585
transform 1 0 6348 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_47
timestamp 1623621585
transform 1 0 5428 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_55
timestamp 1623621585
transform 1 0 6164 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_58
timestamp 1623621585
transform 1 0 6440 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_70
timestamp 1623621585
transform 1 0 7544 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_82
timestamp 1623621585
transform 1 0 8648 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_94
timestamp 1623621585
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_880
timestamp 1623621585
transform 1 0 11592 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_106
timestamp 1623621585
transform 1 0 10856 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_115
timestamp 1623621585
transform 1 0 11684 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_127
timestamp 1623621585
transform 1 0 12788 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_139
timestamp 1623621585
transform 1 0 13892 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_151
timestamp 1623621585
transform 1 0 14996 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_163
timestamp 1623621585
transform 1 0 16100 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_881
timestamp 1623621585
transform 1 0 16836 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_172
timestamp 1623621585
transform 1 0 16928 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_184
timestamp 1623621585
transform 1 0 18032 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_196
timestamp 1623621585
transform 1 0 19136 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_208
timestamp 1623621585
transform 1 0 20240 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_882
timestamp 1623621585
transform 1 0 22080 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_220
timestamp 1623621585
transform 1 0 21344 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_229
timestamp 1623621585
transform 1 0 22172 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_241
timestamp 1623621585
transform 1 0 23276 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1623621585
transform 1 0 24380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1623621585
transform 1 0 25484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_883
timestamp 1623621585
transform 1 0 27324 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_277
timestamp 1623621585
transform 1 0 26588 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_286
timestamp 1623621585
transform 1 0 27416 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_298
timestamp 1623621585
transform 1 0 28520 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_310
timestamp 1623621585
transform 1 0 29624 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_322
timestamp 1623621585
transform 1 0 30728 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_884
timestamp 1623621585
transform 1 0 32568 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_334
timestamp 1623621585
transform 1 0 31832 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_343
timestamp 1623621585
transform 1 0 32660 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_355
timestamp 1623621585
transform 1 0 33764 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_367
timestamp 1623621585
transform 1 0 34868 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input167
timestamp 1623621585
transform 1 0 37168 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_379
timestamp 1623621585
transform 1 0 35972 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1623621585
transform 1 0 37076 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_395
timestamp 1623621585
transform 1 0 37444 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1623621585
transform -1 0 38824 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_885
timestamp 1623621585
transform 1 0 37812 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_400
timestamp 1623621585
transform 1 0 37904 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_406
timestamp 1623621585
transform 1 0 38456 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1623621585
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input357
timestamp 1623621585
transform 1 0 1748 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_3
timestamp 1623621585
transform 1 0 1380 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_11
timestamp 1623621585
transform 1 0 2116 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_886
timestamp 1623621585
transform 1 0 3772 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_23
timestamp 1623621585
transform 1 0 3220 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_30
timestamp 1623621585
transform 1 0 3864 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_42
timestamp 1623621585
transform 1 0 4968 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_54
timestamp 1623621585
transform 1 0 6072 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_66
timestamp 1623621585
transform 1 0 7176 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_78
timestamp 1623621585
transform 1 0 8280 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_887
timestamp 1623621585
transform 1 0 9016 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_87
timestamp 1623621585
transform 1 0 9108 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_99
timestamp 1623621585
transform 1 0 10212 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_111
timestamp 1623621585
transform 1 0 11316 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_123
timestamp 1623621585
transform 1 0 12420 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_888
timestamp 1623621585
transform 1 0 14260 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_135
timestamp 1623621585
transform 1 0 13524 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_144
timestamp 1623621585
transform 1 0 14352 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_156
timestamp 1623621585
transform 1 0 15456 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_168
timestamp 1623621585
transform 1 0 16560 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_180
timestamp 1623621585
transform 1 0 17664 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_889
timestamp 1623621585
transform 1 0 19504 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_192
timestamp 1623621585
transform 1 0 18768 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_201
timestamp 1623621585
transform 1 0 19596 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_213
timestamp 1623621585
transform 1 0 20700 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1623621585
transform 1 0 21804 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1623621585
transform 1 0 22908 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_249
timestamp 1623621585
transform 1 0 24012 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_890
timestamp 1623621585
transform 1 0 24748 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_258
timestamp 1623621585
transform 1 0 24840 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_270
timestamp 1623621585
transform 1 0 25944 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_282
timestamp 1623621585
transform 1 0 27048 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_294
timestamp 1623621585
transform 1 0 28152 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_306
timestamp 1623621585
transform 1 0 29256 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_891
timestamp 1623621585
transform 1 0 29992 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_315
timestamp 1623621585
transform 1 0 30084 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_327
timestamp 1623621585
transform 1 0 31188 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _457_
timestamp 1623621585
transform 1 0 33304 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_12
timestamp 1623621585
transform 1 0 33120 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_339
timestamp 1623621585
transform 1 0 32292 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_347
timestamp 1623621585
transform 1 0 33028 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_892
timestamp 1623621585
transform 1 0 35236 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_358
timestamp 1623621585
transform 1 0 34040 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_370
timestamp 1623621585
transform 1 0 35144 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_372
timestamp 1623621585
transform 1 0 35328 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_384
timestamp 1623621585
transform 1 0 36432 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1623621585
transform -1 0 38824 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input103
timestamp 1623621585
transform 1 0 37904 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_396
timestamp 1623621585
transform 1 0 37536 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_403
timestamp 1623621585
transform 1 0 38180 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1623621585
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1623621585
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input358
timestamp 1623621585
transform 1 0 1748 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1623621585
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1623621585
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_3
timestamp 1623621585
transform 1 0 1380 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_11
timestamp 1623621585
transform 1 0 2116 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_900
timestamp 1623621585
transform 1 0 3772 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_27
timestamp 1623621585
transform 1 0 3588 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_39
timestamp 1623621585
transform 1 0 4692 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_23
timestamp 1623621585
transform 1 0 3220 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_30
timestamp 1623621585
transform 1 0 3864 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_893
timestamp 1623621585
transform 1 0 6348 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_51
timestamp 1623621585
transform 1 0 5796 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_58
timestamp 1623621585
transform 1 0 6440 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_42
timestamp 1623621585
transform 1 0 4968 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_54
timestamp 1623621585
transform 1 0 6072 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_70
timestamp 1623621585
transform 1 0 7544 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_82
timestamp 1623621585
transform 1 0 8648 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_66
timestamp 1623621585
transform 1 0 7176 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_78
timestamp 1623621585
transform 1 0 8280 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_901
timestamp 1623621585
transform 1 0 9016 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_94
timestamp 1623621585
transform 1 0 9752 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_87
timestamp 1623621585
transform 1 0 9108 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_99
timestamp 1623621585
transform 1 0 10212 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_894
timestamp 1623621585
transform 1 0 11592 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_106
timestamp 1623621585
transform 1 0 10856 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_115
timestamp 1623621585
transform 1 0 11684 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_111
timestamp 1623621585
transform 1 0 11316 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_123
timestamp 1623621585
transform 1 0 12420 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_902
timestamp 1623621585
transform 1 0 14260 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_127
timestamp 1623621585
transform 1 0 12788 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_139
timestamp 1623621585
transform 1 0 13892 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_135
timestamp 1623621585
transform 1 0 13524 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_144
timestamp 1623621585
transform 1 0 14352 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_151
timestamp 1623621585
transform 1 0 14996 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_163
timestamp 1623621585
transform 1 0 16100 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_156
timestamp 1623621585
transform 1 0 15456 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_895
timestamp 1623621585
transform 1 0 16836 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_172
timestamp 1623621585
transform 1 0 16928 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_184
timestamp 1623621585
transform 1 0 18032 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_168
timestamp 1623621585
transform 1 0 16560 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_180
timestamp 1623621585
transform 1 0 17664 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_903
timestamp 1623621585
transform 1 0 19504 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_196
timestamp 1623621585
transform 1 0 19136 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_208
timestamp 1623621585
transform 1 0 20240 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_192
timestamp 1623621585
transform 1 0 18768 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_201
timestamp 1623621585
transform 1 0 19596 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_896
timestamp 1623621585
transform 1 0 22080 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_220
timestamp 1623621585
transform 1 0 21344 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_229
timestamp 1623621585
transform 1 0 22172 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_213
timestamp 1623621585
transform 1 0 20700 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1623621585
transform 1 0 21804 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_241
timestamp 1623621585
transform 1 0 23276 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1623621585
transform 1 0 22908 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_249
timestamp 1623621585
transform 1 0 24012 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_904
timestamp 1623621585
transform 1 0 24748 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1623621585
transform 1 0 24380 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1623621585
transform 1 0 25484 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_258
timestamp 1623621585
transform 1 0 24840 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_270
timestamp 1623621585
transform 1 0 25944 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_897
timestamp 1623621585
transform 1 0 27324 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_277
timestamp 1623621585
transform 1 0 26588 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_286
timestamp 1623621585
transform 1 0 27416 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_282
timestamp 1623621585
transform 1 0 27048 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _452_
timestamp 1623621585
transform 1 0 28888 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_298
timestamp 1623621585
transform 1 0 28520 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_306
timestamp 1623621585
transform 1 0 29256 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_294
timestamp 1623621585
transform 1 0 28152 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_306
timestamp 1623621585
transform 1 0 29256 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_905
timestamp 1623621585
transform 1 0 29992 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_318
timestamp 1623621585
transform 1 0 30360 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_330
timestamp 1623621585
transform 1 0 31464 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_315
timestamp 1623621585
transform 1 0 30084 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_327
timestamp 1623621585
transform 1 0 31188 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _369_
timestamp 1623621585
transform 1 0 33120 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_898
timestamp 1623621585
transform 1 0 32568 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_343
timestamp 1623621585
transform 1 0 32660 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_347
timestamp 1623621585
transform 1 0 33028 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_352
timestamp 1623621585
transform 1 0 33488 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_339
timestamp 1623621585
transform 1 0 32292 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_351
timestamp 1623621585
transform 1 0 33396 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _371_
timestamp 1623621585
transform 1 0 33856 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _453_
timestamp 1623621585
transform 1 0 34592 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_906
timestamp 1623621585
transform 1 0 35236 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_360
timestamp 1623621585
transform 1 0 34224 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_367
timestamp 1623621585
transform 1 0 34868 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_363
timestamp 1623621585
transform 1 0 34500 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_372
timestamp 1623621585
transform 1 0 35328 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input135
timestamp 1623621585
transform 1 0 37168 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input168
timestamp 1623621585
transform 1 0 37260 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_379
timestamp 1623621585
transform 1 0 35972 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_391
timestamp 1623621585
transform 1 0 37076 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_395
timestamp 1623621585
transform 1 0 37444 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_384
timestamp 1623621585
transform 1 0 36432 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_392
timestamp 1623621585
transform 1 0 37168 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1623621585
transform -1 0 38824 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1623621585
transform -1 0 38824 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_899
timestamp 1623621585
transform 1 0 37812 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input104
timestamp 1623621585
transform 1 0 37904 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_400
timestamp 1623621585
transform 1 0 37904 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_406
timestamp 1623621585
transform 1 0 38456 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_396
timestamp 1623621585
transform 1 0 37536 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_403
timestamp 1623621585
transform 1 0 38180 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1623621585
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input359
timestamp 1623621585
transform 1 0 1748 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_3
timestamp 1623621585
transform 1 0 1380 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_11
timestamp 1623621585
transform 1 0 2116 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_23
timestamp 1623621585
transform 1 0 3220 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_35
timestamp 1623621585
transform 1 0 4324 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_907
timestamp 1623621585
transform 1 0 6348 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_47
timestamp 1623621585
transform 1 0 5428 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_55
timestamp 1623621585
transform 1 0 6164 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_58
timestamp 1623621585
transform 1 0 6440 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_70
timestamp 1623621585
transform 1 0 7544 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_82
timestamp 1623621585
transform 1 0 8648 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_94
timestamp 1623621585
transform 1 0 9752 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_908
timestamp 1623621585
transform 1 0 11592 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_106
timestamp 1623621585
transform 1 0 10856 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_115
timestamp 1623621585
transform 1 0 11684 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_127
timestamp 1623621585
transform 1 0 12788 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_139
timestamp 1623621585
transform 1 0 13892 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_151
timestamp 1623621585
transform 1 0 14996 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_163
timestamp 1623621585
transform 1 0 16100 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_909
timestamp 1623621585
transform 1 0 16836 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_172
timestamp 1623621585
transform 1 0 16928 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_184
timestamp 1623621585
transform 1 0 18032 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_196
timestamp 1623621585
transform 1 0 19136 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_208
timestamp 1623621585
transform 1 0 20240 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_910
timestamp 1623621585
transform 1 0 22080 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_220
timestamp 1623621585
transform 1 0 21344 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_229
timestamp 1623621585
transform 1 0 22172 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_241
timestamp 1623621585
transform 1 0 23276 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1623621585
transform 1 0 24380 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1623621585
transform 1 0 25484 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_911
timestamp 1623621585
transform 1 0 27324 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_277
timestamp 1623621585
transform 1 0 26588 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_286
timestamp 1623621585
transform 1 0 27416 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_298
timestamp 1623621585
transform 1 0 28520 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_310
timestamp 1623621585
transform 1 0 29624 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_322
timestamp 1623621585
transform 1 0 30728 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _443_
timestamp 1623621585
transform 1 0 33672 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_912
timestamp 1623621585
transform 1 0 32568 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_334
timestamp 1623621585
transform 1 0 31832 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_343
timestamp 1623621585
transform 1 0 32660 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_351
timestamp 1623621585
transform 1 0 33396 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_362
timestamp 1623621585
transform 1 0 34408 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_374
timestamp 1623621585
transform 1 0 35512 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_386
timestamp 1623621585
transform 1 0 36616 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1623621585
transform -1 0 38824 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_913
timestamp 1623621585
transform 1 0 37812 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_398
timestamp 1623621585
transform 1 0 37720 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_400
timestamp 1623621585
transform 1 0 37904 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_406
timestamp 1623621585
transform 1 0 38456 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1623621585
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1623621585
transform 1 0 1380 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1623621585
transform 1 0 2484 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_914
timestamp 1623621585
transform 1 0 3772 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_27
timestamp 1623621585
transform 1 0 3588 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_30
timestamp 1623621585
transform 1 0 3864 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_42
timestamp 1623621585
transform 1 0 4968 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_54
timestamp 1623621585
transform 1 0 6072 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_66
timestamp 1623621585
transform 1 0 7176 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_78
timestamp 1623621585
transform 1 0 8280 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_915
timestamp 1623621585
transform 1 0 9016 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_87
timestamp 1623621585
transform 1 0 9108 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_99
timestamp 1623621585
transform 1 0 10212 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_111
timestamp 1623621585
transform 1 0 11316 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_123
timestamp 1623621585
transform 1 0 12420 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_916
timestamp 1623621585
transform 1 0 14260 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_135
timestamp 1623621585
transform 1 0 13524 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_144
timestamp 1623621585
transform 1 0 14352 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _393_
timestamp 1623621585
transform 1 0 15640 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_69_156
timestamp 1623621585
transform 1 0 15456 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_163
timestamp 1623621585
transform 1 0 16100 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _364_
timestamp 1623621585
transform 1 0 16468 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _380_
timestamp 1623621585
transform 1 0 17296 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _400_
timestamp 1623621585
transform 1 0 18124 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_69_172
timestamp 1623621585
transform 1 0 16928 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_181
timestamp 1623621585
transform 1 0 17756 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_917
timestamp 1623621585
transform 1 0 19504 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_190
timestamp 1623621585
transform 1 0 18584 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_198
timestamp 1623621585
transform 1 0 19320 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_201
timestamp 1623621585
transform 1 0 19596 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_213
timestamp 1623621585
transform 1 0 20700 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1623621585
transform 1 0 21804 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1623621585
transform 1 0 22908 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_249
timestamp 1623621585
transform 1 0 24012 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_918
timestamp 1623621585
transform 1 0 24748 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_258
timestamp 1623621585
transform 1 0 24840 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_270
timestamp 1623621585
transform 1 0 25944 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_282
timestamp 1623621585
transform 1 0 27048 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_294
timestamp 1623621585
transform 1 0 28152 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_306
timestamp 1623621585
transform 1 0 29256 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_919
timestamp 1623621585
transform 1 0 29992 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_315
timestamp 1623621585
transform 1 0 30084 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_327
timestamp 1623621585
transform 1 0 31188 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _436_
timestamp 1623621585
transform 1 0 33672 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_339
timestamp 1623621585
transform 1 0 32292 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_351
timestamp 1623621585
transform 1 0 33396 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_920
timestamp 1623621585
transform 1 0 35236 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_362
timestamp 1623621585
transform 1 0 34408 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_370
timestamp 1623621585
transform 1 0 35144 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_372
timestamp 1623621585
transform 1 0 35328 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input169
timestamp 1623621585
transform 1 0 37260 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_384
timestamp 1623621585
transform 1 0 36432 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_392
timestamp 1623621585
transform 1 0 37168 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1623621585
transform -1 0 38824 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input136
timestamp 1623621585
transform 1 0 37904 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_396
timestamp 1623621585
transform 1 0 37536 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_403
timestamp 1623621585
transform 1 0 38180 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1623621585
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input360
timestamp 1623621585
transform 1 0 1748 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1623621585
transform 1 0 1380 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_11
timestamp 1623621585
transform 1 0 2116 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_23
timestamp 1623621585
transform 1 0 3220 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_35
timestamp 1623621585
transform 1 0 4324 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_921
timestamp 1623621585
transform 1 0 6348 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_47
timestamp 1623621585
transform 1 0 5428 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_55
timestamp 1623621585
transform 1 0 6164 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_58
timestamp 1623621585
transform 1 0 6440 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_70
timestamp 1623621585
transform 1 0 7544 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_82
timestamp 1623621585
transform 1 0 8648 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_94
timestamp 1623621585
transform 1 0 9752 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_922
timestamp 1623621585
transform 1 0 11592 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_106
timestamp 1623621585
transform 1 0 10856 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_115
timestamp 1623621585
transform 1 0 11684 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_127
timestamp 1623621585
transform 1 0 12788 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_139
timestamp 1623621585
transform 1 0 13892 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_151
timestamp 1623621585
transform 1 0 14996 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_163
timestamp 1623621585
transform 1 0 16100 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _386_
timestamp 1623621585
transform 1 0 17296 0 -1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_923
timestamp 1623621585
transform 1 0 16836 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_172
timestamp 1623621585
transform 1 0 16928 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_181
timestamp 1623621585
transform 1 0 17756 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_193
timestamp 1623621585
transform 1 0 18860 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_205
timestamp 1623621585
transform 1 0 19964 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_924
timestamp 1623621585
transform 1 0 22080 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_217
timestamp 1623621585
transform 1 0 21068 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_225
timestamp 1623621585
transform 1 0 21804 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_229
timestamp 1623621585
transform 1 0 22172 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_241
timestamp 1623621585
transform 1 0 23276 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1623621585
transform 1 0 24380 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1623621585
transform 1 0 25484 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_925
timestamp 1623621585
transform 1 0 27324 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_277
timestamp 1623621585
transform 1 0 26588 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_286
timestamp 1623621585
transform 1 0 27416 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_298
timestamp 1623621585
transform 1 0 28520 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_310
timestamp 1623621585
transform 1 0 29624 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_322
timestamp 1623621585
transform 1 0 30728 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_926
timestamp 1623621585
transform 1 0 32568 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_334
timestamp 1623621585
transform 1 0 31832 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_343
timestamp 1623621585
transform 1 0 32660 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_355
timestamp 1623621585
transform 1 0 33764 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_367
timestamp 1623621585
transform 1 0 34868 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_379
timestamp 1623621585
transform 1 0 35972 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_391
timestamp 1623621585
transform 1 0 37076 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1623621585
transform -1 0 38824 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_927
timestamp 1623621585
transform 1 0 37812 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_400
timestamp 1623621585
transform 1 0 37904 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_406
timestamp 1623621585
transform 1 0 38456 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1623621585
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input361
timestamp 1623621585
transform 1 0 1748 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_3
timestamp 1623621585
transform 1 0 1380 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_11
timestamp 1623621585
transform 1 0 2116 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_928
timestamp 1623621585
transform 1 0 3772 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_23
timestamp 1623621585
transform 1 0 3220 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_30
timestamp 1623621585
transform 1 0 3864 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_42
timestamp 1623621585
transform 1 0 4968 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_54
timestamp 1623621585
transform 1 0 6072 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_66
timestamp 1623621585
transform 1 0 7176 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_78
timestamp 1623621585
transform 1 0 8280 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_929
timestamp 1623621585
transform 1 0 9016 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_87
timestamp 1623621585
transform 1 0 9108 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_99
timestamp 1623621585
transform 1 0 10212 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_111
timestamp 1623621585
transform 1 0 11316 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_123
timestamp 1623621585
transform 1 0 12420 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_930
timestamp 1623621585
transform 1 0 14260 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_135
timestamp 1623621585
transform 1 0 13524 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_144
timestamp 1623621585
transform 1 0 14352 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_156
timestamp 1623621585
transform 1 0 15456 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_168
timestamp 1623621585
transform 1 0 16560 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_180
timestamp 1623621585
transform 1 0 17664 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_931
timestamp 1623621585
transform 1 0 19504 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_192
timestamp 1623621585
transform 1 0 18768 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_201
timestamp 1623621585
transform 1 0 19596 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_213
timestamp 1623621585
transform 1 0 20700 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1623621585
transform 1 0 21804 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1623621585
transform 1 0 22908 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_249
timestamp 1623621585
transform 1 0 24012 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_932
timestamp 1623621585
transform 1 0 24748 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_258
timestamp 1623621585
transform 1 0 24840 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_270
timestamp 1623621585
transform 1 0 25944 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_282
timestamp 1623621585
transform 1 0 27048 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_294
timestamp 1623621585
transform 1 0 28152 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_306
timestamp 1623621585
transform 1 0 29256 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_933
timestamp 1623621585
transform 1 0 29992 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_315
timestamp 1623621585
transform 1 0 30084 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_327
timestamp 1623621585
transform 1 0 31188 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _430_
timestamp 1623621585
transform 1 0 33672 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_339
timestamp 1623621585
transform 1 0 32292 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_351
timestamp 1623621585
transform 1 0 33396 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_934
timestamp 1623621585
transform 1 0 35236 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_362
timestamp 1623621585
transform 1 0 34408 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_370
timestamp 1623621585
transform 1 0 35144 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_372
timestamp 1623621585
transform 1 0 35328 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input137
timestamp 1623621585
transform 1 0 37260 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_384
timestamp 1623621585
transform 1 0 36432 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_392
timestamp 1623621585
transform 1 0 37168 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1623621585
transform -1 0 38824 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input105
timestamp 1623621585
transform 1 0 37904 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_396
timestamp 1623621585
transform 1 0 37536 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_403
timestamp 1623621585
transform 1 0 38180 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1623621585
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1623621585
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input363
timestamp 1623621585
transform 1 0 1748 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_3
timestamp 1623621585
transform 1 0 1380 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_11
timestamp 1623621585
transform 1 0 2116 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1623621585
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1623621585
transform 1 0 2484 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_942
timestamp 1623621585
transform 1 0 3772 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_23
timestamp 1623621585
transform 1 0 3220 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_35
timestamp 1623621585
transform 1 0 4324 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_27
timestamp 1623621585
transform 1 0 3588 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_30
timestamp 1623621585
transform 1 0 3864 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_935
timestamp 1623621585
transform 1 0 6348 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_47
timestamp 1623621585
transform 1 0 5428 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_55
timestamp 1623621585
transform 1 0 6164 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_58
timestamp 1623621585
transform 1 0 6440 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_42
timestamp 1623621585
transform 1 0 4968 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_54
timestamp 1623621585
transform 1 0 6072 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_70
timestamp 1623621585
transform 1 0 7544 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_82
timestamp 1623621585
transform 1 0 8648 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_66
timestamp 1623621585
transform 1 0 7176 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_78
timestamp 1623621585
transform 1 0 8280 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_943
timestamp 1623621585
transform 1 0 9016 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_94
timestamp 1623621585
transform 1 0 9752 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_87
timestamp 1623621585
transform 1 0 9108 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_99
timestamp 1623621585
transform 1 0 10212 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_936
timestamp 1623621585
transform 1 0 11592 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_106
timestamp 1623621585
transform 1 0 10856 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_115
timestamp 1623621585
transform 1 0 11684 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_111
timestamp 1623621585
transform 1 0 11316 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_123
timestamp 1623621585
transform 1 0 12420 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_944
timestamp 1623621585
transform 1 0 14260 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_127
timestamp 1623621585
transform 1 0 12788 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_139
timestamp 1623621585
transform 1 0 13892 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_135
timestamp 1623621585
transform 1 0 13524 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_144
timestamp 1623621585
transform 1 0 14352 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _409_
timestamp 1623621585
transform 1 0 16192 0 1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_72_151
timestamp 1623621585
transform 1 0 14996 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_163
timestamp 1623621585
transform 1 0 16100 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_156
timestamp 1623621585
transform 1 0 15456 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_937
timestamp 1623621585
transform 1 0 16836 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_172
timestamp 1623621585
transform 1 0 16928 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_184
timestamp 1623621585
transform 1 0 18032 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1623621585
transform 1 0 16652 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1623621585
transform 1 0 17756 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_945
timestamp 1623621585
transform 1 0 19504 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_196
timestamp 1623621585
transform 1 0 19136 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_208
timestamp 1623621585
transform 1 0 20240 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_193
timestamp 1623621585
transform 1 0 18860 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_199
timestamp 1623621585
transform 1 0 19412 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_201
timestamp 1623621585
transform 1 0 19596 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_938
timestamp 1623621585
transform 1 0 22080 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_220
timestamp 1623621585
transform 1 0 21344 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_229
timestamp 1623621585
transform 1 0 22172 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_213
timestamp 1623621585
transform 1 0 20700 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1623621585
transform 1 0 21804 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_241
timestamp 1623621585
transform 1 0 23276 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1623621585
transform 1 0 22908 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_249
timestamp 1623621585
transform 1 0 24012 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_946
timestamp 1623621585
transform 1 0 24748 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1623621585
transform 1 0 24380 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1623621585
transform 1 0 25484 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_258
timestamp 1623621585
transform 1 0 24840 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_270
timestamp 1623621585
transform 1 0 25944 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_939
timestamp 1623621585
transform 1 0 27324 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_277
timestamp 1623621585
transform 1 0 26588 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_286
timestamp 1623621585
transform 1 0 27416 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_282
timestamp 1623621585
transform 1 0 27048 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_298
timestamp 1623621585
transform 1 0 28520 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_310
timestamp 1623621585
transform 1 0 29624 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_294
timestamp 1623621585
transform 1 0 28152 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_306
timestamp 1623621585
transform 1 0 29256 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_947
timestamp 1623621585
transform 1 0 29992 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_322
timestamp 1623621585
transform 1 0 30728 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_315
timestamp 1623621585
transform 1 0 30084 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_327
timestamp 1623621585
transform 1 0 31188 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_940
timestamp 1623621585
transform 1 0 32568 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_334
timestamp 1623621585
transform 1 0 31832 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_343
timestamp 1623621585
transform 1 0 32660 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_339
timestamp 1623621585
transform 1 0 32292 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_351
timestamp 1623621585
transform 1 0 33396 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _417_
timestamp 1623621585
transform 1 0 33764 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _423_
timestamp 1623621585
transform 1 0 33764 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_948
timestamp 1623621585
transform 1 0 35236 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_363
timestamp 1623621585
transform 1 0 34500 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_375
timestamp 1623621585
transform 1 0 35604 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_363
timestamp 1623621585
transform 1 0 34500 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_372
timestamp 1623621585
transform 1 0 35328 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input139
timestamp 1623621585
transform 1 0 37260 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input171
timestamp 1623621585
transform 1 0 37168 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_387
timestamp 1623621585
transform 1 0 36708 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_391
timestamp 1623621585
transform 1 0 37076 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_395
timestamp 1623621585
transform 1 0 37444 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_384
timestamp 1623621585
transform 1 0 36432 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_392
timestamp 1623621585
transform 1 0 37168 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1623621585
transform -1 0 38824 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1623621585
transform -1 0 38824 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_941
timestamp 1623621585
transform 1 0 37812 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input107
timestamp 1623621585
transform 1 0 37904 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_72_400
timestamp 1623621585
transform 1 0 37904 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_406
timestamp 1623621585
transform 1 0 38456 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_396
timestamp 1623621585
transform 1 0 37536 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_403
timestamp 1623621585
transform 1 0 38180 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1623621585
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input364
timestamp 1623621585
transform 1 0 1748 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_3
timestamp 1623621585
transform 1 0 1380 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_11
timestamp 1623621585
transform 1 0 2116 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_23
timestamp 1623621585
transform 1 0 3220 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_35
timestamp 1623621585
transform 1 0 4324 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_949
timestamp 1623621585
transform 1 0 6348 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_47
timestamp 1623621585
transform 1 0 5428 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_55
timestamp 1623621585
transform 1 0 6164 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_58
timestamp 1623621585
transform 1 0 6440 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_70
timestamp 1623621585
transform 1 0 7544 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_82
timestamp 1623621585
transform 1 0 8648 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_94
timestamp 1623621585
transform 1 0 9752 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_950
timestamp 1623621585
transform 1 0 11592 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_106
timestamp 1623621585
transform 1 0 10856 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_115
timestamp 1623621585
transform 1 0 11684 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_127
timestamp 1623621585
transform 1 0 12788 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_139
timestamp 1623621585
transform 1 0 13892 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _433_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 15916 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_74_151
timestamp 1623621585
transform 1 0 14996 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_159
timestamp 1623621585
transform 1 0 15732 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__and2_1  _420_
timestamp 1623621585
transform 1 0 17296 0 -1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_951
timestamp 1623621585
transform 1 0 16836 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_167
timestamp 1623621585
transform 1 0 16468 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_172
timestamp 1623621585
transform 1 0 16928 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_181
timestamp 1623621585
transform 1 0 17756 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_193
timestamp 1623621585
transform 1 0 18860 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_205
timestamp 1623621585
transform 1 0 19964 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_952
timestamp 1623621585
transform 1 0 22080 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_217
timestamp 1623621585
transform 1 0 21068 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_225
timestamp 1623621585
transform 1 0 21804 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_229
timestamp 1623621585
transform 1 0 22172 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_241
timestamp 1623621585
transform 1 0 23276 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1623621585
transform 1 0 24380 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1623621585
transform 1 0 25484 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_953
timestamp 1623621585
transform 1 0 27324 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_277
timestamp 1623621585
transform 1 0 26588 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_286
timestamp 1623621585
transform 1 0 27416 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_298
timestamp 1623621585
transform 1 0 28520 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_310
timestamp 1623621585
transform 1 0 29624 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_322
timestamp 1623621585
transform 1 0 30728 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_954
timestamp 1623621585
transform 1 0 32568 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_334
timestamp 1623621585
transform 1 0 31832 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_343
timestamp 1623621585
transform 1 0 32660 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_355
timestamp 1623621585
transform 1 0 33764 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_367
timestamp 1623621585
transform 1 0 34868 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input172
timestamp 1623621585
transform 1 0 37168 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_379
timestamp 1623621585
transform 1 0 35972 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_391
timestamp 1623621585
transform 1 0 37076 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_395
timestamp 1623621585
transform 1 0 37444 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1623621585
transform -1 0 38824 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_955
timestamp 1623621585
transform 1 0 37812 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_400
timestamp 1623621585
transform 1 0 37904 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_406
timestamp 1623621585
transform 1 0 38456 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1623621585
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input365
timestamp 1623621585
transform 1 0 1748 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_3
timestamp 1623621585
transform 1 0 1380 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_11
timestamp 1623621585
transform 1 0 2116 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_956
timestamp 1623621585
transform 1 0 3772 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_23
timestamp 1623621585
transform 1 0 3220 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_30
timestamp 1623621585
transform 1 0 3864 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_42
timestamp 1623621585
transform 1 0 4968 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_54
timestamp 1623621585
transform 1 0 6072 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_66
timestamp 1623621585
transform 1 0 7176 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_78
timestamp 1623621585
transform 1 0 8280 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_957
timestamp 1623621585
transform 1 0 9016 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_87
timestamp 1623621585
transform 1 0 9108 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_99
timestamp 1623621585
transform 1 0 10212 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_111
timestamp 1623621585
transform 1 0 11316 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_123
timestamp 1623621585
transform 1 0 12420 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_958
timestamp 1623621585
transform 1 0 14260 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_135
timestamp 1623621585
transform 1 0 13524 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_75_144
timestamp 1623621585
transform 1 0 14352 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _426_
timestamp 1623621585
transform 1 0 16192 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _440_
timestamp 1623621585
transform 1 0 15272 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_75_152
timestamp 1623621585
transform 1 0 15088 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_160
timestamp 1623621585
transform 1 0 15824 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_170
timestamp 1623621585
transform 1 0 16744 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_182
timestamp 1623621585
transform 1 0 17848 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_959
timestamp 1623621585
transform 1 0 19504 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_194
timestamp 1623621585
transform 1 0 18952 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_201
timestamp 1623621585
transform 1 0 19596 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_213
timestamp 1623621585
transform 1 0 20700 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1623621585
transform 1 0 21804 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1623621585
transform 1 0 22908 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_249
timestamp 1623621585
transform 1 0 24012 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_960
timestamp 1623621585
transform 1 0 24748 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_258
timestamp 1623621585
transform 1 0 24840 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_270
timestamp 1623621585
transform 1 0 25944 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_282
timestamp 1623621585
transform 1 0 27048 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_294
timestamp 1623621585
transform 1 0 28152 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_306
timestamp 1623621585
transform 1 0 29256 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_961
timestamp 1623621585
transform 1 0 29992 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_315
timestamp 1623621585
transform 1 0 30084 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_327
timestamp 1623621585
transform 1 0 31188 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_339
timestamp 1623621585
transform 1 0 32292 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_351
timestamp 1623621585
transform 1 0 33396 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_962
timestamp 1623621585
transform 1 0 35236 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_363
timestamp 1623621585
transform 1 0 34500 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_372
timestamp 1623621585
transform 1 0 35328 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_384
timestamp 1623621585
transform 1 0 36432 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1623621585
transform -1 0 38824 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input108
timestamp 1623621585
transform 1 0 37904 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_396
timestamp 1623621585
transform 1 0 37536 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_403
timestamp 1623621585
transform 1 0 38180 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1623621585
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1623621585
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1623621585
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_27
timestamp 1623621585
transform 1 0 3588 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_39
timestamp 1623621585
transform 1 0 4692 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_963
timestamp 1623621585
transform 1 0 6348 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_51
timestamp 1623621585
transform 1 0 5796 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_58
timestamp 1623621585
transform 1 0 6440 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_70
timestamp 1623621585
transform 1 0 7544 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_82
timestamp 1623621585
transform 1 0 8648 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_94
timestamp 1623621585
transform 1 0 9752 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_964
timestamp 1623621585
transform 1 0 11592 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_106
timestamp 1623621585
transform 1 0 10856 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_115
timestamp 1623621585
transform 1 0 11684 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_127
timestamp 1623621585
transform 1 0 12788 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_139
timestamp 1623621585
transform 1 0 13892 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_151
timestamp 1623621585
transform 1 0 14996 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_163
timestamp 1623621585
transform 1 0 16100 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_965
timestamp 1623621585
transform 1 0 16836 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_172
timestamp 1623621585
transform 1 0 16928 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_184
timestamp 1623621585
transform 1 0 18032 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_196
timestamp 1623621585
transform 1 0 19136 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_208
timestamp 1623621585
transform 1 0 20240 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_966
timestamp 1623621585
transform 1 0 22080 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_220
timestamp 1623621585
transform 1 0 21344 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_229
timestamp 1623621585
transform 1 0 22172 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_241
timestamp 1623621585
transform 1 0 23276 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1623621585
transform 1 0 24380 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1623621585
transform 1 0 25484 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_967
timestamp 1623621585
transform 1 0 27324 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_277
timestamp 1623621585
transform 1 0 26588 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_286
timestamp 1623621585
transform 1 0 27416 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_298
timestamp 1623621585
transform 1 0 28520 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_310
timestamp 1623621585
transform 1 0 29624 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_322
timestamp 1623621585
transform 1 0 30728 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_968
timestamp 1623621585
transform 1 0 32568 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_334
timestamp 1623621585
transform 1 0 31832 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_343
timestamp 1623621585
transform 1 0 32660 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_355
timestamp 1623621585
transform 1 0 33764 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_367
timestamp 1623621585
transform 1 0 34868 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input140
timestamp 1623621585
transform 1 0 37168 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_379
timestamp 1623621585
transform 1 0 35972 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_391
timestamp 1623621585
transform 1 0 37076 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_395
timestamp 1623621585
transform 1 0 37444 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1623621585
transform -1 0 38824 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_969
timestamp 1623621585
transform 1 0 37812 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_400
timestamp 1623621585
transform 1 0 37904 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_406
timestamp 1623621585
transform 1 0 38456 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1623621585
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input366
timestamp 1623621585
transform 1 0 1748 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_3
timestamp 1623621585
transform 1 0 1380 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_11
timestamp 1623621585
transform 1 0 2116 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_970
timestamp 1623621585
transform 1 0 3772 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_23
timestamp 1623621585
transform 1 0 3220 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_30
timestamp 1623621585
transform 1 0 3864 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_42
timestamp 1623621585
transform 1 0 4968 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_54
timestamp 1623621585
transform 1 0 6072 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_66
timestamp 1623621585
transform 1 0 7176 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_78
timestamp 1623621585
transform 1 0 8280 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_971
timestamp 1623621585
transform 1 0 9016 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_87
timestamp 1623621585
transform 1 0 9108 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_99
timestamp 1623621585
transform 1 0 10212 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_111
timestamp 1623621585
transform 1 0 11316 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_123
timestamp 1623621585
transform 1 0 12420 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_972
timestamp 1623621585
transform 1 0 14260 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_135
timestamp 1623621585
transform 1 0 13524 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_144
timestamp 1623621585
transform 1 0 14352 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_156
timestamp 1623621585
transform 1 0 15456 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_168
timestamp 1623621585
transform 1 0 16560 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_180
timestamp 1623621585
transform 1 0 17664 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_973
timestamp 1623621585
transform 1 0 19504 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_192
timestamp 1623621585
transform 1 0 18768 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_201
timestamp 1623621585
transform 1 0 19596 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_213
timestamp 1623621585
transform 1 0 20700 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1623621585
transform 1 0 21804 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1623621585
transform 1 0 22908 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_249
timestamp 1623621585
transform 1 0 24012 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_974
timestamp 1623621585
transform 1 0 24748 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_258
timestamp 1623621585
transform 1 0 24840 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_270
timestamp 1623621585
transform 1 0 25944 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_282
timestamp 1623621585
transform 1 0 27048 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_294
timestamp 1623621585
transform 1 0 28152 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_306
timestamp 1623621585
transform 1 0 29256 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_975
timestamp 1623621585
transform 1 0 29992 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_315
timestamp 1623621585
transform 1 0 30084 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_327
timestamp 1623621585
transform 1 0 31188 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_339
timestamp 1623621585
transform 1 0 32292 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_351
timestamp 1623621585
transform 1 0 33396 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_2  _403_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 33856 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_976
timestamp 1623621585
transform 1 0 35236 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_355
timestamp 1623621585
transform 1 0 33764 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_365
timestamp 1623621585
transform 1 0 34684 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_372
timestamp 1623621585
transform 1 0 35328 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input173
timestamp 1623621585
transform 1 0 37260 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_384
timestamp 1623621585
transform 1 0 36432 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_392
timestamp 1623621585
transform 1 0 37168 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1623621585
transform -1 0 38824 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input109
timestamp 1623621585
transform 1 0 37904 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_396
timestamp 1623621585
transform 1 0 37536 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_403
timestamp 1623621585
transform 1 0 38180 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1623621585
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input367
timestamp 1623621585
transform 1 0 1748 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_3
timestamp 1623621585
transform 1 0 1380 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_11
timestamp 1623621585
transform 1 0 2116 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_23
timestamp 1623621585
transform 1 0 3220 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_35
timestamp 1623621585
transform 1 0 4324 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_977
timestamp 1623621585
transform 1 0 6348 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_47
timestamp 1623621585
transform 1 0 5428 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_55
timestamp 1623621585
transform 1 0 6164 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_58
timestamp 1623621585
transform 1 0 6440 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_70
timestamp 1623621585
transform 1 0 7544 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_82
timestamp 1623621585
transform 1 0 8648 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_94
timestamp 1623621585
transform 1 0 9752 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_978
timestamp 1623621585
transform 1 0 11592 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_106
timestamp 1623621585
transform 1 0 10856 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_115
timestamp 1623621585
transform 1 0 11684 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_127
timestamp 1623621585
transform 1 0 12788 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_139
timestamp 1623621585
transform 1 0 13892 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_151
timestamp 1623621585
transform 1 0 14996 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_163
timestamp 1623621585
transform 1 0 16100 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_979
timestamp 1623621585
transform 1 0 16836 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_172
timestamp 1623621585
transform 1 0 16928 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_184
timestamp 1623621585
transform 1 0 18032 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_196
timestamp 1623621585
transform 1 0 19136 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_208
timestamp 1623621585
transform 1 0 20240 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_980
timestamp 1623621585
transform 1 0 22080 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_220
timestamp 1623621585
transform 1 0 21344 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_229
timestamp 1623621585
transform 1 0 22172 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_241
timestamp 1623621585
transform 1 0 23276 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1623621585
transform 1 0 24380 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1623621585
transform 1 0 25484 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_981
timestamp 1623621585
transform 1 0 27324 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_277
timestamp 1623621585
transform 1 0 26588 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_286
timestamp 1623621585
transform 1 0 27416 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_298
timestamp 1623621585
transform 1 0 28520 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_310
timestamp 1623621585
transform 1 0 29624 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_322
timestamp 1623621585
transform 1 0 30728 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_982
timestamp 1623621585
transform 1 0 32568 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_334
timestamp 1623621585
transform 1 0 31832 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_343
timestamp 1623621585
transform 1 0 32660 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_355
timestamp 1623621585
transform 1 0 33764 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_367
timestamp 1623621585
transform 1 0 34868 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_379
timestamp 1623621585
transform 1 0 35972 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_391
timestamp 1623621585
transform 1 0 37076 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1623621585
transform -1 0 38824 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_983
timestamp 1623621585
transform 1 0 37812 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_400
timestamp 1623621585
transform 1 0 37904 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_406
timestamp 1623621585
transform 1 0 38456 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1623621585
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1623621585
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input368
timestamp 1623621585
transform 1 0 1748 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1623621585
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1623621585
transform 1 0 2484 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_3
timestamp 1623621585
transform 1 0 1380 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_11
timestamp 1623621585
transform 1 0 2116 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_984
timestamp 1623621585
transform 1 0 3772 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_27
timestamp 1623621585
transform 1 0 3588 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_30
timestamp 1623621585
transform 1 0 3864 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_23
timestamp 1623621585
transform 1 0 3220 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_35
timestamp 1623621585
transform 1 0 4324 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_991
timestamp 1623621585
transform 1 0 6348 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_42
timestamp 1623621585
transform 1 0 4968 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_54
timestamp 1623621585
transform 1 0 6072 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_47
timestamp 1623621585
transform 1 0 5428 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_55
timestamp 1623621585
transform 1 0 6164 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_58
timestamp 1623621585
transform 1 0 6440 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_66
timestamp 1623621585
transform 1 0 7176 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_78
timestamp 1623621585
transform 1 0 8280 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_70
timestamp 1623621585
transform 1 0 7544 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_82
timestamp 1623621585
transform 1 0 8648 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_985
timestamp 1623621585
transform 1 0 9016 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_87
timestamp 1623621585
transform 1 0 9108 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_99
timestamp 1623621585
transform 1 0 10212 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_94
timestamp 1623621585
transform 1 0 9752 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_992
timestamp 1623621585
transform 1 0 11592 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_111
timestamp 1623621585
transform 1 0 11316 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_123
timestamp 1623621585
transform 1 0 12420 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_106
timestamp 1623621585
transform 1 0 10856 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_115
timestamp 1623621585
transform 1 0 11684 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_986
timestamp 1623621585
transform 1 0 14260 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_135
timestamp 1623621585
transform 1 0 13524 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_144
timestamp 1623621585
transform 1 0 14352 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_127
timestamp 1623621585
transform 1 0 12788 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_139
timestamp 1623621585
transform 1 0 13892 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_156
timestamp 1623621585
transform 1 0 15456 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_151
timestamp 1623621585
transform 1 0 14996 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_163
timestamp 1623621585
transform 1 0 16100 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_993
timestamp 1623621585
transform 1 0 16836 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_168
timestamp 1623621585
transform 1 0 16560 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_180
timestamp 1623621585
transform 1 0 17664 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_172
timestamp 1623621585
transform 1 0 16928 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_184
timestamp 1623621585
transform 1 0 18032 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_987
timestamp 1623621585
transform 1 0 19504 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_192
timestamp 1623621585
transform 1 0 18768 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_201
timestamp 1623621585
transform 1 0 19596 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_196
timestamp 1623621585
transform 1 0 19136 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_208
timestamp 1623621585
transform 1 0 20240 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_994
timestamp 1623621585
transform 1 0 22080 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_213
timestamp 1623621585
transform 1 0 20700 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1623621585
transform 1 0 21804 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_220
timestamp 1623621585
transform 1 0 21344 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_229
timestamp 1623621585
transform 1 0 22172 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1623621585
transform 1 0 22908 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_249
timestamp 1623621585
transform 1 0 24012 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_241
timestamp 1623621585
transform 1 0 23276 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_988
timestamp 1623621585
transform 1 0 24748 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_258
timestamp 1623621585
transform 1 0 24840 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_270
timestamp 1623621585
transform 1 0 25944 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_253
timestamp 1623621585
transform 1 0 24380 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_265
timestamp 1623621585
transform 1 0 25484 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_995
timestamp 1623621585
transform 1 0 27324 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_282
timestamp 1623621585
transform 1 0 27048 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_277
timestamp 1623621585
transform 1 0 26588 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_286
timestamp 1623621585
transform 1 0 27416 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_294
timestamp 1623621585
transform 1 0 28152 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_306
timestamp 1623621585
transform 1 0 29256 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_298
timestamp 1623621585
transform 1 0 28520 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_310
timestamp 1623621585
transform 1 0 29624 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_989
timestamp 1623621585
transform 1 0 29992 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_315
timestamp 1623621585
transform 1 0 30084 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_327
timestamp 1623621585
transform 1 0 31188 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_322
timestamp 1623621585
transform 1 0 30728 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_996
timestamp 1623621585
transform 1 0 32568 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_339
timestamp 1623621585
transform 1 0 32292 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_351
timestamp 1623621585
transform 1 0 33396 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_80_334
timestamp 1623621585
transform 1 0 31832 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_343
timestamp 1623621585
transform 1 0 32660 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _390_
timestamp 1623621585
transform 1 0 33948 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _396_
timestamp 1623621585
transform 1 0 33948 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_990
timestamp 1623621585
transform 1 0 35236 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_366
timestamp 1623621585
transform 1 0 34776 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_370
timestamp 1623621585
transform 1 0 35144 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_372
timestamp 1623621585
transform 1 0 35328 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_355
timestamp 1623621585
transform 1 0 33764 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_366
timestamp 1623621585
transform 1 0 34776 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input142
timestamp 1623621585
transform 1 0 37168 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input174
timestamp 1623621585
transform 1 0 37260 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_384
timestamp 1623621585
transform 1 0 36432 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_392
timestamp 1623621585
transform 1 0 37168 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_378
timestamp 1623621585
transform 1 0 35880 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_390
timestamp 1623621585
transform 1 0 36984 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_395
timestamp 1623621585
transform 1 0 37444 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1623621585
transform -1 0 38824 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1623621585
transform -1 0 38824 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_997
timestamp 1623621585
transform 1 0 37812 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input141
timestamp 1623621585
transform 1 0 37904 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_396
timestamp 1623621585
transform 1 0 37536 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_403
timestamp 1623621585
transform 1 0 38180 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_400
timestamp 1623621585
transform 1 0 37904 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_406
timestamp 1623621585
transform 1 0 38456 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1623621585
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input369
timestamp 1623621585
transform 1 0 1748 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_3
timestamp 1623621585
transform 1 0 1380 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_11
timestamp 1623621585
transform 1 0 2116 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_998
timestamp 1623621585
transform 1 0 3772 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_23
timestamp 1623621585
transform 1 0 3220 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_30
timestamp 1623621585
transform 1 0 3864 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_42
timestamp 1623621585
transform 1 0 4968 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_54
timestamp 1623621585
transform 1 0 6072 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_66
timestamp 1623621585
transform 1 0 7176 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_78
timestamp 1623621585
transform 1 0 8280 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_999
timestamp 1623621585
transform 1 0 9016 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_87
timestamp 1623621585
transform 1 0 9108 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_99
timestamp 1623621585
transform 1 0 10212 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_111
timestamp 1623621585
transform 1 0 11316 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_123
timestamp 1623621585
transform 1 0 12420 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1000
timestamp 1623621585
transform 1 0 14260 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_135
timestamp 1623621585
transform 1 0 13524 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_144
timestamp 1623621585
transform 1 0 14352 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_156
timestamp 1623621585
transform 1 0 15456 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_168
timestamp 1623621585
transform 1 0 16560 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_180
timestamp 1623621585
transform 1 0 17664 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1001
timestamp 1623621585
transform 1 0 19504 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_192
timestamp 1623621585
transform 1 0 18768 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_201
timestamp 1623621585
transform 1 0 19596 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_213
timestamp 1623621585
transform 1 0 20700 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1623621585
transform 1 0 21804 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1623621585
transform 1 0 22908 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_249
timestamp 1623621585
transform 1 0 24012 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1002
timestamp 1623621585
transform 1 0 24748 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_258
timestamp 1623621585
transform 1 0 24840 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_270
timestamp 1623621585
transform 1 0 25944 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_282
timestamp 1623621585
transform 1 0 27048 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_294
timestamp 1623621585
transform 1 0 28152 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_306
timestamp 1623621585
transform 1 0 29256 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1003
timestamp 1623621585
transform 1 0 29992 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_315
timestamp 1623621585
transform 1 0 30084 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_327
timestamp 1623621585
transform 1 0 31188 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_339
timestamp 1623621585
transform 1 0 32292 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_351
timestamp 1623621585
transform 1 0 33396 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _383_
timestamp 1623621585
transform 1 0 33948 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1004
timestamp 1623621585
transform 1 0 35236 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_366
timestamp 1623621585
transform 1 0 34776 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_370
timestamp 1623621585
transform 1 0 35144 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_372
timestamp 1623621585
transform 1 0 35328 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input175
timestamp 1623621585
transform 1 0 37260 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_384
timestamp 1623621585
transform 1 0 36432 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_392
timestamp 1623621585
transform 1 0 37168 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1623621585
transform -1 0 38824 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input110
timestamp 1623621585
transform 1 0 37904 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_396
timestamp 1623621585
transform 1 0 37536 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_403
timestamp 1623621585
transform 1 0 38180 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1623621585
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1623621585
transform 1 0 1380 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1623621585
transform 1 0 2484 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_27
timestamp 1623621585
transform 1 0 3588 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_39
timestamp 1623621585
transform 1 0 4692 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1005
timestamp 1623621585
transform 1 0 6348 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_51
timestamp 1623621585
transform 1 0 5796 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_58
timestamp 1623621585
transform 1 0 6440 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_70
timestamp 1623621585
transform 1 0 7544 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_82
timestamp 1623621585
transform 1 0 8648 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_94
timestamp 1623621585
transform 1 0 9752 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1006
timestamp 1623621585
transform 1 0 11592 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_106
timestamp 1623621585
transform 1 0 10856 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_115
timestamp 1623621585
transform 1 0 11684 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_127
timestamp 1623621585
transform 1 0 12788 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_139
timestamp 1623621585
transform 1 0 13892 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_151
timestamp 1623621585
transform 1 0 14996 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_163
timestamp 1623621585
transform 1 0 16100 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1007
timestamp 1623621585
transform 1 0 16836 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_172
timestamp 1623621585
transform 1 0 16928 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_184
timestamp 1623621585
transform 1 0 18032 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_196
timestamp 1623621585
transform 1 0 19136 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_208
timestamp 1623621585
transform 1 0 20240 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1008
timestamp 1623621585
transform 1 0 22080 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_220
timestamp 1623621585
transform 1 0 21344 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_229
timestamp 1623621585
transform 1 0 22172 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_241
timestamp 1623621585
transform 1 0 23276 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_253
timestamp 1623621585
transform 1 0 24380 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_265
timestamp 1623621585
transform 1 0 25484 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1009
timestamp 1623621585
transform 1 0 27324 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_277
timestamp 1623621585
transform 1 0 26588 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_286
timestamp 1623621585
transform 1 0 27416 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_298
timestamp 1623621585
transform 1 0 28520 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_310
timestamp 1623621585
transform 1 0 29624 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_322
timestamp 1623621585
transform 1 0 30728 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1010
timestamp 1623621585
transform 1 0 32568 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_334
timestamp 1623621585
transform 1 0 31832 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_343
timestamp 1623621585
transform 1 0 32660 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _377_
timestamp 1623621585
transform 1 0 33948 0 -1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_82_355
timestamp 1623621585
transform 1 0 33764 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_366
timestamp 1623621585
transform 1 0 34776 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_378
timestamp 1623621585
transform 1 0 35880 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_390
timestamp 1623621585
transform 1 0 36984 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1623621585
transform -1 0 38824 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1011
timestamp 1623621585
transform 1 0 37812 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_398
timestamp 1623621585
transform 1 0 37720 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_400
timestamp 1623621585
transform 1 0 37904 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_406
timestamp 1623621585
transform 1 0 38456 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1623621585
transform 1 0 1104 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input370
timestamp 1623621585
transform 1 0 1748 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_3
timestamp 1623621585
transform 1 0 1380 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_11
timestamp 1623621585
transform 1 0 2116 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1012
timestamp 1623621585
transform 1 0 3772 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_23
timestamp 1623621585
transform 1 0 3220 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_30
timestamp 1623621585
transform 1 0 3864 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_42
timestamp 1623621585
transform 1 0 4968 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_54
timestamp 1623621585
transform 1 0 6072 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_66
timestamp 1623621585
transform 1 0 7176 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_78
timestamp 1623621585
transform 1 0 8280 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1013
timestamp 1623621585
transform 1 0 9016 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_87
timestamp 1623621585
transform 1 0 9108 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_99
timestamp 1623621585
transform 1 0 10212 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_111
timestamp 1623621585
transform 1 0 11316 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_123
timestamp 1623621585
transform 1 0 12420 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1014
timestamp 1623621585
transform 1 0 14260 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_135
timestamp 1623621585
transform 1 0 13524 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_144
timestamp 1623621585
transform 1 0 14352 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_156
timestamp 1623621585
transform 1 0 15456 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _363_
timestamp 1623621585
transform 1 0 16744 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_83_168
timestamp 1623621585
transform 1 0 16560 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_173
timestamp 1623621585
transform 1 0 17020 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_185
timestamp 1623621585
transform 1 0 18124 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1015
timestamp 1623621585
transform 1 0 19504 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_83_197
timestamp 1623621585
transform 1 0 19228 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_201
timestamp 1623621585
transform 1 0 19596 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_213
timestamp 1623621585
transform 1 0 20700 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_225
timestamp 1623621585
transform 1 0 21804 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_237
timestamp 1623621585
transform 1 0 22908 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_249
timestamp 1623621585
transform 1 0 24012 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1016
timestamp 1623621585
transform 1 0 24748 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_258
timestamp 1623621585
transform 1 0 24840 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_270
timestamp 1623621585
transform 1 0 25944 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_282
timestamp 1623621585
transform 1 0 27048 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_294
timestamp 1623621585
transform 1 0 28152 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_306
timestamp 1623621585
transform 1 0 29256 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1017
timestamp 1623621585
transform 1 0 29992 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_315
timestamp 1623621585
transform 1 0 30084 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_327
timestamp 1623621585
transform 1 0 31188 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_339
timestamp 1623621585
transform 1 0 32292 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_351
timestamp 1623621585
transform 1 0 33396 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1018
timestamp 1623621585
transform 1 0 35236 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_363
timestamp 1623621585
transform 1 0 34500 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_372
timestamp 1623621585
transform 1 0 35328 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input143
timestamp 1623621585
transform 1 0 37260 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_83_384
timestamp 1623621585
transform 1 0 36432 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_392
timestamp 1623621585
transform 1 0 37168 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1623621585
transform -1 0 38824 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input111
timestamp 1623621585
transform 1 0 37904 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_396
timestamp 1623621585
transform 1 0 37536 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_403
timestamp 1623621585
transform 1 0 38180 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1623621585
transform 1 0 1104 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input371
timestamp 1623621585
transform 1 0 1748 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_3
timestamp 1623621585
transform 1 0 1380 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_11
timestamp 1623621585
transform 1 0 2116 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_23
timestamp 1623621585
transform 1 0 3220 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_35
timestamp 1623621585
transform 1 0 4324 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1019
timestamp 1623621585
transform 1 0 6348 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_47
timestamp 1623621585
transform 1 0 5428 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_55
timestamp 1623621585
transform 1 0 6164 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_84_58
timestamp 1623621585
transform 1 0 6440 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_70
timestamp 1623621585
transform 1 0 7544 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_82
timestamp 1623621585
transform 1 0 8648 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_94
timestamp 1623621585
transform 1 0 9752 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1020
timestamp 1623621585
transform 1 0 11592 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_106
timestamp 1623621585
transform 1 0 10856 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_115
timestamp 1623621585
transform 1 0 11684 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_127
timestamp 1623621585
transform 1 0 12788 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_139
timestamp 1623621585
transform 1 0 13892 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_151
timestamp 1623621585
transform 1 0 14996 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_163
timestamp 1623621585
transform 1 0 16100 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1021
timestamp 1623621585
transform 1 0 16836 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_172
timestamp 1623621585
transform 1 0 16928 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_184
timestamp 1623621585
transform 1 0 18032 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_196
timestamp 1623621585
transform 1 0 19136 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_208
timestamp 1623621585
transform 1 0 20240 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1022
timestamp 1623621585
transform 1 0 22080 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_220
timestamp 1623621585
transform 1 0 21344 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_229
timestamp 1623621585
transform 1 0 22172 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_241
timestamp 1623621585
transform 1 0 23276 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_253
timestamp 1623621585
transform 1 0 24380 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_265
timestamp 1623621585
transform 1 0 25484 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1023
timestamp 1623621585
transform 1 0 27324 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_277
timestamp 1623621585
transform 1 0 26588 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_286
timestamp 1623621585
transform 1 0 27416 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_298
timestamp 1623621585
transform 1 0 28520 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_310
timestamp 1623621585
transform 1 0 29624 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_322
timestamp 1623621585
transform 1 0 30728 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1024
timestamp 1623621585
transform 1 0 32568 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_334
timestamp 1623621585
transform 1 0 31832 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_343
timestamp 1623621585
transform 1 0 32660 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_355
timestamp 1623621585
transform 1 0 33764 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_367
timestamp 1623621585
transform 1 0 34868 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input176
timestamp 1623621585
transform 1 0 37168 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_379
timestamp 1623621585
transform 1 0 35972 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_391
timestamp 1623621585
transform 1 0 37076 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_395
timestamp 1623621585
transform 1 0 37444 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1623621585
transform -1 0 38824 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1025
timestamp 1623621585
transform 1 0 37812 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_400
timestamp 1623621585
transform 1 0 37904 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_406
timestamp 1623621585
transform 1 0 38456 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1623621585
transform 1 0 1104 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1623621585
transform 1 0 1104 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input372
timestamp 1623621585
transform 1 0 1748 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1623621585
transform 1 0 1380 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1623621585
transform 1 0 2484 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_3
timestamp 1623621585
transform 1 0 1380 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_11
timestamp 1623621585
transform 1 0 2116 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1026
timestamp 1623621585
transform 1 0 3772 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_27
timestamp 1623621585
transform 1 0 3588 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_85_30
timestamp 1623621585
transform 1 0 3864 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_23
timestamp 1623621585
transform 1 0 3220 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_35
timestamp 1623621585
transform 1 0 4324 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1033
timestamp 1623621585
transform 1 0 6348 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_42
timestamp 1623621585
transform 1 0 4968 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_54
timestamp 1623621585
transform 1 0 6072 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_47
timestamp 1623621585
transform 1 0 5428 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_55
timestamp 1623621585
transform 1 0 6164 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_86_58
timestamp 1623621585
transform 1 0 6440 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_66
timestamp 1623621585
transform 1 0 7176 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_78
timestamp 1623621585
transform 1 0 8280 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_70
timestamp 1623621585
transform 1 0 7544 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_82
timestamp 1623621585
transform 1 0 8648 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1027
timestamp 1623621585
transform 1 0 9016 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_87
timestamp 1623621585
transform 1 0 9108 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_99
timestamp 1623621585
transform 1 0 10212 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_94
timestamp 1623621585
transform 1 0 9752 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1034
timestamp 1623621585
transform 1 0 11592 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_111
timestamp 1623621585
transform 1 0 11316 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_123
timestamp 1623621585
transform 1 0 12420 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_106
timestamp 1623621585
transform 1 0 10856 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_115
timestamp 1623621585
transform 1 0 11684 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1028
timestamp 1623621585
transform 1 0 14260 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_135
timestamp 1623621585
transform 1 0 13524 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_144
timestamp 1623621585
transform 1 0 14352 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_127
timestamp 1623621585
transform 1 0 12788 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_139
timestamp 1623621585
transform 1 0 13892 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_156
timestamp 1623621585
transform 1 0 15456 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_151
timestamp 1623621585
transform 1 0 14996 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_163
timestamp 1623621585
transform 1 0 16100 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _408_
timestamp 1623621585
transform 1 0 16652 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1035
timestamp 1623621585
transform 1 0 16836 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_168
timestamp 1623621585
transform 1 0 16560 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_172
timestamp 1623621585
transform 1 0 16928 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_184
timestamp 1623621585
transform 1 0 18032 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_172
timestamp 1623621585
transform 1 0 16928 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_184
timestamp 1623621585
transform 1 0 18032 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1029
timestamp 1623621585
transform 1 0 19504 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_196
timestamp 1623621585
transform 1 0 19136 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_201
timestamp 1623621585
transform 1 0 19596 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_196
timestamp 1623621585
transform 1 0 19136 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_208
timestamp 1623621585
transform 1 0 20240 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1036
timestamp 1623621585
transform 1 0 22080 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_213
timestamp 1623621585
transform 1 0 20700 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_225
timestamp 1623621585
transform 1 0 21804 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_220
timestamp 1623621585
transform 1 0 21344 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_229
timestamp 1623621585
transform 1 0 22172 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_237
timestamp 1623621585
transform 1 0 22908 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_249
timestamp 1623621585
transform 1 0 24012 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_241
timestamp 1623621585
transform 1 0 23276 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1030
timestamp 1623621585
transform 1 0 24748 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_258
timestamp 1623621585
transform 1 0 24840 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_270
timestamp 1623621585
transform 1 0 25944 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_253
timestamp 1623621585
transform 1 0 24380 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_265
timestamp 1623621585
transform 1 0 25484 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__a31oi_4  _586_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 27416 0 1 48416
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1037
timestamp 1623621585
transform 1 0 27324 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_282
timestamp 1623621585
transform 1 0 27048 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_277
timestamp 1623621585
transform 1 0 26588 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_286
timestamp 1623621585
transform 1 0 27416 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_303
timestamp 1623621585
transform 1 0 28980 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_311
timestamp 1623621585
transform 1 0 29716 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_298
timestamp 1623621585
transform 1 0 28520 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_310
timestamp 1623621585
transform 1 0 29624 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1031
timestamp 1623621585
transform 1 0 29992 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_315
timestamp 1623621585
transform 1 0 30084 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_327
timestamp 1623621585
transform 1 0 31188 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_322
timestamp 1623621585
transform 1 0 30728 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1038
timestamp 1623621585
transform 1 0 32568 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_339
timestamp 1623621585
transform 1 0 32292 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_351
timestamp 1623621585
transform 1 0 33396 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_334
timestamp 1623621585
transform 1 0 31832 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_343
timestamp 1623621585
transform 1 0 32660 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1032
timestamp 1623621585
transform 1 0 35236 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_363
timestamp 1623621585
transform 1 0 34500 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_372
timestamp 1623621585
transform 1 0 35328 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_355
timestamp 1623621585
transform 1 0 33764 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_367
timestamp 1623621585
transform 1 0 34868 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input144
timestamp 1623621585
transform 1 0 37260 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input177
timestamp 1623621585
transform 1 0 37168 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_85_384
timestamp 1623621585
transform 1 0 36432 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_392
timestamp 1623621585
transform 1 0 37168 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_379
timestamp 1623621585
transform 1 0 35972 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_391
timestamp 1623621585
transform 1 0 37076 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_395
timestamp 1623621585
transform 1 0 37444 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1623621585
transform -1 0 38824 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1623621585
transform -1 0 38824 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1039
timestamp 1623621585
transform 1 0 37812 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input112
timestamp 1623621585
transform 1 0 37904 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_396
timestamp 1623621585
transform 1 0 37536 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_403
timestamp 1623621585
transform 1 0 38180 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_400
timestamp 1623621585
transform 1 0 37904 0 -1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_406
timestamp 1623621585
transform 1 0 38456 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1623621585
transform 1 0 1104 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input374
timestamp 1623621585
transform 1 0 1748 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_3
timestamp 1623621585
transform 1 0 1380 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_11
timestamp 1623621585
transform 1 0 2116 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1040
timestamp 1623621585
transform 1 0 3772 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_23
timestamp 1623621585
transform 1 0 3220 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_87_30
timestamp 1623621585
transform 1 0 3864 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_42
timestamp 1623621585
transform 1 0 4968 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_54
timestamp 1623621585
transform 1 0 6072 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_66
timestamp 1623621585
transform 1 0 7176 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_78
timestamp 1623621585
transform 1 0 8280 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1041
timestamp 1623621585
transform 1 0 9016 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_87
timestamp 1623621585
transform 1 0 9108 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_99
timestamp 1623621585
transform 1 0 10212 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_111
timestamp 1623621585
transform 1 0 11316 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_123
timestamp 1623621585
transform 1 0 12420 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1042
timestamp 1623621585
transform 1 0 14260 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_135
timestamp 1623621585
transform 1 0 13524 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_144
timestamp 1623621585
transform 1 0 14352 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_156
timestamp 1623621585
transform 1 0 15456 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_168
timestamp 1623621585
transform 1 0 16560 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_180
timestamp 1623621585
transform 1 0 17664 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1043
timestamp 1623621585
transform 1 0 19504 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_192
timestamp 1623621585
transform 1 0 18768 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_201
timestamp 1623621585
transform 1 0 19596 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_213
timestamp 1623621585
transform 1 0 20700 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_225
timestamp 1623621585
transform 1 0 21804 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_237
timestamp 1623621585
transform 1 0 22908 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_249
timestamp 1623621585
transform 1 0 24012 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1044
timestamp 1623621585
transform 1 0 24748 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_258
timestamp 1623621585
transform 1 0 24840 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_270
timestamp 1623621585
transform 1 0 25944 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_282
timestamp 1623621585
transform 1 0 27048 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_294
timestamp 1623621585
transform 1 0 28152 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_306
timestamp 1623621585
transform 1 0 29256 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1045
timestamp 1623621585
transform 1 0 29992 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_315
timestamp 1623621585
transform 1 0 30084 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_327
timestamp 1623621585
transform 1 0 31188 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_2  _583_
timestamp 1623621585
transform 1 0 31924 0 1 49504
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_87_345
timestamp 1623621585
transform 1 0 32844 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1046
timestamp 1623621585
transform 1 0 35236 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_357
timestamp 1623621585
transform 1 0 33948 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_369
timestamp 1623621585
transform 1 0 35052 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_372
timestamp 1623621585
transform 1 0 35328 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_384
timestamp 1623621585
transform 1 0 36432 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1623621585
transform -1 0 38824 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 1623621585
transform 1 0 37904 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_87_396
timestamp 1623621585
transform 1 0 37536 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_403
timestamp 1623621585
transform 1 0 38180 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1623621585
transform 1 0 1104 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1623621585
transform 1 0 1380 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_15
timestamp 1623621585
transform 1 0 2484 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_27
timestamp 1623621585
transform 1 0 3588 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_39
timestamp 1623621585
transform 1 0 4692 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1047
timestamp 1623621585
transform 1 0 6348 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_51
timestamp 1623621585
transform 1 0 5796 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_88_58
timestamp 1623621585
transform 1 0 6440 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_70
timestamp 1623621585
transform 1 0 7544 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_82
timestamp 1623621585
transform 1 0 8648 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_94
timestamp 1623621585
transform 1 0 9752 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1048
timestamp 1623621585
transform 1 0 11592 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_106
timestamp 1623621585
transform 1 0 10856 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_115
timestamp 1623621585
transform 1 0 11684 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_127
timestamp 1623621585
transform 1 0 12788 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_139
timestamp 1623621585
transform 1 0 13892 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_151
timestamp 1623621585
transform 1 0 14996 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_163
timestamp 1623621585
transform 1 0 16100 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1049
timestamp 1623621585
transform 1 0 16836 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_172
timestamp 1623621585
transform 1 0 16928 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_184
timestamp 1623621585
transform 1 0 18032 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_196
timestamp 1623621585
transform 1 0 19136 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_208
timestamp 1623621585
transform 1 0 20240 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1050
timestamp 1623621585
transform 1 0 22080 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_220
timestamp 1623621585
transform 1 0 21344 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_229
timestamp 1623621585
transform 1 0 22172 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_241
timestamp 1623621585
transform 1 0 23276 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_253
timestamp 1623621585
transform 1 0 24380 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_265
timestamp 1623621585
transform 1 0 25484 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1051
timestamp 1623621585
transform 1 0 27324 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_277
timestamp 1623621585
transform 1 0 26588 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_286
timestamp 1623621585
transform 1 0 27416 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _328_
timestamp 1623621585
transform 1 0 28796 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_0
timestamp 1623621585
transform 1 0 28612 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_298
timestamp 1623621585
transform 1 0 28520 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_305
timestamp 1623621585
transform 1 0 29164 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_317
timestamp 1623621585
transform 1 0 30268 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_329
timestamp 1623621585
transform 1 0 31372 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _355_
timestamp 1623621585
transform 1 0 33304 0 -1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1052
timestamp 1623621585
transform 1 0 32568 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_341
timestamp 1623621585
transform 1 0 32476 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_343
timestamp 1623621585
transform 1 0 32660 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_349
timestamp 1623621585
transform 1 0 33212 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _329_
timestamp 1623621585
transform 1 0 34500 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_359
timestamp 1623621585
transform 1 0 34132 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_367
timestamp 1623621585
transform 1 0 34868 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_379
timestamp 1623621585
transform 1 0 35972 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_391
timestamp 1623621585
transform 1 0 37076 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1623621585
transform -1 0 38824 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1053
timestamp 1623621585
transform 1 0 37812 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_400
timestamp 1623621585
transform 1 0 37904 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_406
timestamp 1623621585
transform 1 0 38456 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1623621585
transform 1 0 1104 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input375
timestamp 1623621585
transform 1 0 1748 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_3
timestamp 1623621585
transform 1 0 1380 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_11
timestamp 1623621585
transform 1 0 2116 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1054
timestamp 1623621585
transform 1 0 3772 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_23
timestamp 1623621585
transform 1 0 3220 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_89_30
timestamp 1623621585
transform 1 0 3864 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_42
timestamp 1623621585
transform 1 0 4968 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_54
timestamp 1623621585
transform 1 0 6072 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_66
timestamp 1623621585
transform 1 0 7176 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_78
timestamp 1623621585
transform 1 0 8280 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1055
timestamp 1623621585
transform 1 0 9016 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_87
timestamp 1623621585
transform 1 0 9108 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_99
timestamp 1623621585
transform 1 0 10212 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_111
timestamp 1623621585
transform 1 0 11316 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_123
timestamp 1623621585
transform 1 0 12420 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1056
timestamp 1623621585
transform 1 0 14260 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_135
timestamp 1623621585
transform 1 0 13524 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_144
timestamp 1623621585
transform 1 0 14352 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_156
timestamp 1623621585
transform 1 0 15456 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_168
timestamp 1623621585
transform 1 0 16560 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_180
timestamp 1623621585
transform 1 0 17664 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1057
timestamp 1623621585
transform 1 0 19504 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_192
timestamp 1623621585
transform 1 0 18768 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_201
timestamp 1623621585
transform 1 0 19596 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_213
timestamp 1623621585
transform 1 0 20700 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_225
timestamp 1623621585
transform 1 0 21804 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_237
timestamp 1623621585
transform 1 0 22908 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_249
timestamp 1623621585
transform 1 0 24012 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1058
timestamp 1623621585
transform 1 0 24748 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_258
timestamp 1623621585
transform 1 0 24840 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_270
timestamp 1623621585
transform 1 0 25944 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_282
timestamp 1623621585
transform 1 0 27048 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_294
timestamp 1623621585
transform 1 0 28152 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_306
timestamp 1623621585
transform 1 0 29256 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1059
timestamp 1623621585
transform 1 0 29992 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_315
timestamp 1623621585
transform 1 0 30084 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_327
timestamp 1623621585
transform 1 0 31188 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _347_
timestamp 1623621585
transform 1 0 33304 0 1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_14
timestamp 1623621585
transform 1 0 33120 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_89_339
timestamp 1623621585
transform 1 0 32292 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_347
timestamp 1623621585
transform 1 0 33028 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1060
timestamp 1623621585
transform 1 0 35236 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_359
timestamp 1623621585
transform 1 0 34132 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_372
timestamp 1623621585
transform 1 0 35328 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input178
timestamp 1623621585
transform 1 0 37260 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_89_384
timestamp 1623621585
transform 1 0 36432 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_392
timestamp 1623621585
transform 1 0 37168 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1623621585
transform -1 0 38824 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input145
timestamp 1623621585
transform 1 0 37904 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_396
timestamp 1623621585
transform 1 0 37536 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_403
timestamp 1623621585
transform 1 0 38180 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1623621585
transform 1 0 1104 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input383
timestamp 1623621585
transform 1 0 1380 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_6
timestamp 1623621585
transform 1 0 1656 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_18
timestamp 1623621585
transform 1 0 2760 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_30
timestamp 1623621585
transform 1 0 3864 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1061
timestamp 1623621585
transform 1 0 6348 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_42
timestamp 1623621585
transform 1 0 4968 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_90_54
timestamp 1623621585
transform 1 0 6072 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_58
timestamp 1623621585
transform 1 0 6440 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_70
timestamp 1623621585
transform 1 0 7544 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_82
timestamp 1623621585
transform 1 0 8648 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_94
timestamp 1623621585
transform 1 0 9752 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1062
timestamp 1623621585
transform 1 0 11592 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_106
timestamp 1623621585
transform 1 0 10856 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_115
timestamp 1623621585
transform 1 0 11684 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_127
timestamp 1623621585
transform 1 0 12788 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_139
timestamp 1623621585
transform 1 0 13892 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_151
timestamp 1623621585
transform 1 0 14996 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_163
timestamp 1623621585
transform 1 0 16100 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1063
timestamp 1623621585
transform 1 0 16836 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_172
timestamp 1623621585
transform 1 0 16928 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_184
timestamp 1623621585
transform 1 0 18032 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_196
timestamp 1623621585
transform 1 0 19136 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_208
timestamp 1623621585
transform 1 0 20240 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1064
timestamp 1623621585
transform 1 0 22080 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_220
timestamp 1623621585
transform 1 0 21344 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_229
timestamp 1623621585
transform 1 0 22172 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_241
timestamp 1623621585
transform 1 0 23276 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_253
timestamp 1623621585
transform 1 0 24380 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_265
timestamp 1623621585
transform 1 0 25484 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1065
timestamp 1623621585
transform 1 0 27324 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_277
timestamp 1623621585
transform 1 0 26588 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_286
timestamp 1623621585
transform 1 0 27416 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_298
timestamp 1623621585
transform 1 0 28520 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_310
timestamp 1623621585
transform 1 0 29624 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_322
timestamp 1623621585
transform 1 0 30728 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _341_
timestamp 1623621585
transform 1 0 33304 0 -1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1066
timestamp 1623621585
transform 1 0 32568 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_15
timestamp 1623621585
transform 1 0 33120 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_90_334
timestamp 1623621585
transform 1 0 31832 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_90_343
timestamp 1623621585
transform 1 0 32660 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_347
timestamp 1623621585
transform 1 0 33028 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_359
timestamp 1623621585
transform 1 0 34132 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_371
timestamp 1623621585
transform 1 0 35236 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input146
timestamp 1623621585
transform 1 0 37168 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_90_383
timestamp 1623621585
transform 1 0 36340 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_391
timestamp 1623621585
transform 1 0 37076 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_395
timestamp 1623621585
transform 1 0 37444 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1623621585
transform -1 0 38824 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1067
timestamp 1623621585
transform 1 0 37812 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_400
timestamp 1623621585
transform 1 0 37904 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_406
timestamp 1623621585
transform 1 0 38456 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1623621585
transform 1 0 1104 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_3
timestamp 1623621585
transform 1 0 1380 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_15
timestamp 1623621585
transform 1 0 2484 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1068
timestamp 1623621585
transform 1 0 3772 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_27
timestamp 1623621585
transform 1 0 3588 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_91_30
timestamp 1623621585
transform 1 0 3864 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_42
timestamp 1623621585
transform 1 0 4968 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_54
timestamp 1623621585
transform 1 0 6072 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_66
timestamp 1623621585
transform 1 0 7176 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_78
timestamp 1623621585
transform 1 0 8280 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1069
timestamp 1623621585
transform 1 0 9016 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_87
timestamp 1623621585
transform 1 0 9108 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_99
timestamp 1623621585
transform 1 0 10212 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_111
timestamp 1623621585
transform 1 0 11316 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_123
timestamp 1623621585
transform 1 0 12420 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1070
timestamp 1623621585
transform 1 0 14260 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_135
timestamp 1623621585
transform 1 0 13524 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_144
timestamp 1623621585
transform 1 0 14352 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_156
timestamp 1623621585
transform 1 0 15456 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_168
timestamp 1623621585
transform 1 0 16560 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_180
timestamp 1623621585
transform 1 0 17664 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1071
timestamp 1623621585
transform 1 0 19504 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_192
timestamp 1623621585
transform 1 0 18768 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_201
timestamp 1623621585
transform 1 0 19596 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_213
timestamp 1623621585
transform 1 0 20700 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_225
timestamp 1623621585
transform 1 0 21804 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_237
timestamp 1623621585
transform 1 0 22908 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_249
timestamp 1623621585
transform 1 0 24012 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1072
timestamp 1623621585
transform 1 0 24748 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_258
timestamp 1623621585
transform 1 0 24840 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_270
timestamp 1623621585
transform 1 0 25944 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_282
timestamp 1623621585
transform 1 0 27048 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_294
timestamp 1623621585
transform 1 0 28152 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_306
timestamp 1623621585
transform 1 0 29256 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1073
timestamp 1623621585
transform 1 0 29992 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_315
timestamp 1623621585
transform 1 0 30084 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_327
timestamp 1623621585
transform 1 0 31188 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _333_
timestamp 1623621585
transform 1 0 33028 0 1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_16
timestamp 1623621585
transform 1 0 32844 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_91_339
timestamp 1623621585
transform 1 0 32292 0 1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1074
timestamp 1623621585
transform 1 0 35236 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_356
timestamp 1623621585
transform 1 0 33856 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_368
timestamp 1623621585
transform 1 0 34960 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_372
timestamp 1623621585
transform 1 0 35328 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input179
timestamp 1623621585
transform 1 0 37260 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_91_384
timestamp 1623621585
transform 1 0 36432 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_392
timestamp 1623621585
transform 1 0 37168 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1623621585
transform -1 0 38824 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input114
timestamp 1623621585
transform 1 0 37904 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_396
timestamp 1623621585
transform 1 0 37536 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_403
timestamp 1623621585
transform 1 0 38180 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1623621585
transform 1 0 1104 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1623621585
transform 1 0 1104 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input394
timestamp 1623621585
transform 1 0 1380 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input405
timestamp 1623621585
transform 1 0 1380 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_6
timestamp 1623621585
transform 1 0 1656 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_18
timestamp 1623621585
transform 1 0 2760 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_6
timestamp 1623621585
transform 1 0 1656 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_18
timestamp 1623621585
transform 1 0 2760 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1082
timestamp 1623621585
transform 1 0 3772 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_30
timestamp 1623621585
transform 1 0 3864 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_26
timestamp 1623621585
transform 1 0 3496 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_30
timestamp 1623621585
transform 1 0 3864 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1075
timestamp 1623621585
transform 1 0 6348 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_42
timestamp 1623621585
transform 1 0 4968 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_54
timestamp 1623621585
transform 1 0 6072 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_58
timestamp 1623621585
transform 1 0 6440 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_42
timestamp 1623621585
transform 1 0 4968 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_54
timestamp 1623621585
transform 1 0 6072 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_70
timestamp 1623621585
transform 1 0 7544 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_82
timestamp 1623621585
transform 1 0 8648 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_66
timestamp 1623621585
transform 1 0 7176 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_78
timestamp 1623621585
transform 1 0 8280 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1083
timestamp 1623621585
transform 1 0 9016 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_94
timestamp 1623621585
transform 1 0 9752 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_87
timestamp 1623621585
transform 1 0 9108 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_99
timestamp 1623621585
transform 1 0 10212 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1076
timestamp 1623621585
transform 1 0 11592 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_106
timestamp 1623621585
transform 1 0 10856 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_115
timestamp 1623621585
transform 1 0 11684 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_111
timestamp 1623621585
transform 1 0 11316 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_123
timestamp 1623621585
transform 1 0 12420 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1084
timestamp 1623621585
transform 1 0 14260 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_127
timestamp 1623621585
transform 1 0 12788 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_139
timestamp 1623621585
transform 1 0 13892 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_135
timestamp 1623621585
transform 1 0 13524 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_144
timestamp 1623621585
transform 1 0 14352 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_151
timestamp 1623621585
transform 1 0 14996 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_163
timestamp 1623621585
transform 1 0 16100 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_156
timestamp 1623621585
transform 1 0 15456 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1077
timestamp 1623621585
transform 1 0 16836 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_172
timestamp 1623621585
transform 1 0 16928 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_184
timestamp 1623621585
transform 1 0 18032 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_168
timestamp 1623621585
transform 1 0 16560 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_180
timestamp 1623621585
transform 1 0 17664 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1085
timestamp 1623621585
transform 1 0 19504 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_196
timestamp 1623621585
transform 1 0 19136 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_208
timestamp 1623621585
transform 1 0 20240 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_192
timestamp 1623621585
transform 1 0 18768 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_201
timestamp 1623621585
transform 1 0 19596 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1078
timestamp 1623621585
transform 1 0 22080 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_220
timestamp 1623621585
transform 1 0 21344 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_229
timestamp 1623621585
transform 1 0 22172 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_213
timestamp 1623621585
transform 1 0 20700 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_225
timestamp 1623621585
transform 1 0 21804 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_241
timestamp 1623621585
transform 1 0 23276 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_237
timestamp 1623621585
transform 1 0 22908 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_249
timestamp 1623621585
transform 1 0 24012 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1086
timestamp 1623621585
transform 1 0 24748 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_253
timestamp 1623621585
transform 1 0 24380 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_265
timestamp 1623621585
transform 1 0 25484 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_258
timestamp 1623621585
transform 1 0 24840 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_270
timestamp 1623621585
transform 1 0 25944 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1079
timestamp 1623621585
transform 1 0 27324 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_277
timestamp 1623621585
transform 1 0 26588 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_286
timestamp 1623621585
transform 1 0 27416 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_282
timestamp 1623621585
transform 1 0 27048 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_298
timestamp 1623621585
transform 1 0 28520 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_310
timestamp 1623621585
transform 1 0 29624 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_294
timestamp 1623621585
transform 1 0 28152 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_306
timestamp 1623621585
transform 1 0 29256 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1087
timestamp 1623621585
transform 1 0 29992 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_322
timestamp 1623621585
transform 1 0 30728 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_315
timestamp 1623621585
transform 1 0 30084 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_327
timestamp 1623621585
transform 1 0 31188 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1080
timestamp 1623621585
transform 1 0 32568 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_334
timestamp 1623621585
transform 1 0 31832 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_343
timestamp 1623621585
transform 1 0 32660 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_339
timestamp 1623621585
transform 1 0 32292 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_351
timestamp 1623621585
transform 1 0 33396 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1088
timestamp 1623621585
transform 1 0 35236 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_355
timestamp 1623621585
transform 1 0 33764 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_367
timestamp 1623621585
transform 1 0 34868 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_363
timestamp 1623621585
transform 1 0 34500 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_372
timestamp 1623621585
transform 1 0 35328 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input147
timestamp 1623621585
transform 1 0 37260 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_379
timestamp 1623621585
transform 1 0 35972 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_391
timestamp 1623621585
transform 1 0 37076 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_93_384
timestamp 1623621585
transform 1 0 36432 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_392
timestamp 1623621585
transform 1 0 37168 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1623621585
transform -1 0 38824 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1623621585
transform -1 0 38824 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1081
timestamp 1623621585
transform 1 0 37812 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input115
timestamp 1623621585
transform 1 0 37904 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_92_400
timestamp 1623621585
transform 1 0 37904 0 -1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_406
timestamp 1623621585
transform 1 0 38456 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_396
timestamp 1623621585
transform 1 0 37536 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_403
timestamp 1623621585
transform 1 0 38180 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1623621585
transform 1 0 1104 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input408
timestamp 1623621585
transform 1 0 1380 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_6
timestamp 1623621585
transform 1 0 1656 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_18
timestamp 1623621585
transform 1 0 2760 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_30
timestamp 1623621585
transform 1 0 3864 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1089
timestamp 1623621585
transform 1 0 6348 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_42
timestamp 1623621585
transform 1 0 4968 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_54
timestamp 1623621585
transform 1 0 6072 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_58
timestamp 1623621585
transform 1 0 6440 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_70
timestamp 1623621585
transform 1 0 7544 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_82
timestamp 1623621585
transform 1 0 8648 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_94
timestamp 1623621585
transform 1 0 9752 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1090
timestamp 1623621585
transform 1 0 11592 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_106
timestamp 1623621585
transform 1 0 10856 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_115
timestamp 1623621585
transform 1 0 11684 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_127
timestamp 1623621585
transform 1 0 12788 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_139
timestamp 1623621585
transform 1 0 13892 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_151
timestamp 1623621585
transform 1 0 14996 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_163
timestamp 1623621585
transform 1 0 16100 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1091
timestamp 1623621585
transform 1 0 16836 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_172
timestamp 1623621585
transform 1 0 16928 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_184
timestamp 1623621585
transform 1 0 18032 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _722_
timestamp 1623621585
transform 1 0 18952 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_94_192
timestamp 1623621585
transform 1 0 18768 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_94_200
timestamp 1623621585
transform 1 0 19504 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1092
timestamp 1623621585
transform 1 0 22080 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_212
timestamp 1623621585
transform 1 0 20608 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_224
timestamp 1623621585
transform 1 0 21712 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_229
timestamp 1623621585
transform 1 0 22172 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _715_
timestamp 1623621585
transform 1 0 22724 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_94_241
timestamp 1623621585
transform 1 0 23276 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _718_
timestamp 1623621585
transform 1 0 24840 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_94_253
timestamp 1623621585
transform 1 0 24380 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_257
timestamp 1623621585
transform 1 0 24748 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_264
timestamp 1623621585
transform 1 0 25392 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _734_
timestamp 1623621585
transform 1 0 27784 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1093
timestamp 1623621585
transform 1 0 27324 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_276
timestamp 1623621585
transform 1 0 26496 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_284
timestamp 1623621585
transform 1 0 27232 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_286
timestamp 1623621585
transform 1 0 27416 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _737_
timestamp 1623621585
transform 1 0 28888 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_94_296
timestamp 1623621585
transform 1 0 28336 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_94_308
timestamp 1623621585
transform 1 0 29440 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_320
timestamp 1623621585
transform 1 0 30544 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_332
timestamp 1623621585
transform 1 0 31648 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1094
timestamp 1623621585
transform 1 0 32568 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_340
timestamp 1623621585
transform 1 0 32384 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_94_343
timestamp 1623621585
transform 1 0 32660 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_355
timestamp 1623621585
transform 1 0 33764 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_367
timestamp 1623621585
transform 1 0 34868 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input116
timestamp 1623621585
transform 1 0 37168 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input180
timestamp 1623621585
transform 1 0 36524 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_94_379
timestamp 1623621585
transform 1 0 35972 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_94_388
timestamp 1623621585
transform 1 0 36800 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_395
timestamp 1623621585
transform 1 0 37444 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1623621585
transform -1 0 38824 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1095
timestamp 1623621585
transform 1 0 37812 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_400
timestamp 1623621585
transform 1 0 37904 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_406
timestamp 1623621585
transform 1 0 38456 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1623621585
transform 1 0 1104 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_3
timestamp 1623621585
transform 1 0 1380 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_15
timestamp 1623621585
transform 1 0 2484 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1096
timestamp 1623621585
transform 1 0 3772 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_27
timestamp 1623621585
transform 1 0 3588 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_95_30
timestamp 1623621585
transform 1 0 3864 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_42
timestamp 1623621585
transform 1 0 4968 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_54
timestamp 1623621585
transform 1 0 6072 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_66
timestamp 1623621585
transform 1 0 7176 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_78
timestamp 1623621585
transform 1 0 8280 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1097
timestamp 1623621585
transform 1 0 9016 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_87
timestamp 1623621585
transform 1 0 9108 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_99
timestamp 1623621585
transform 1 0 10212 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_111
timestamp 1623621585
transform 1 0 11316 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_123
timestamp 1623621585
transform 1 0 12420 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1098
timestamp 1623621585
transform 1 0 14260 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_135
timestamp 1623621585
transform 1 0 13524 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_144
timestamp 1623621585
transform 1 0 14352 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_156
timestamp 1623621585
transform 1 0 15456 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_168
timestamp 1623621585
transform 1 0 16560 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_180
timestamp 1623621585
transform 1 0 17664 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1099
timestamp 1623621585
transform 1 0 19504 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_192
timestamp 1623621585
transform 1 0 18768 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_201
timestamp 1623621585
transform 1 0 19596 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _725_
timestamp 1623621585
transform 1 0 21344 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_95_213
timestamp 1623621585
transform 1 0 20700 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_219
timestamp 1623621585
transform 1 0 21252 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_226
timestamp 1623621585
transform 1 0 21896 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_238
timestamp 1623621585
transform 1 0 23000 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_250
timestamp 1623621585
transform 1 0 24104 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1100
timestamp 1623621585
transform 1 0 24748 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_256
timestamp 1623621585
transform 1 0 24656 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_258
timestamp 1623621585
transform 1 0 24840 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_270
timestamp 1623621585
transform 1 0 25944 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_282
timestamp 1623621585
transform 1 0 27048 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_294
timestamp 1623621585
transform 1 0 28152 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_306
timestamp 1623621585
transform 1 0 29256 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1101
timestamp 1623621585
transform 1 0 29992 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_315
timestamp 1623621585
transform 1 0 30084 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_327
timestamp 1623621585
transform 1 0 31188 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _743_
timestamp 1623621585
transform 1 0 31924 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _745_
timestamp 1623621585
transform 1 0 33028 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_95_341
timestamp 1623621585
transform 1 0 32476 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_95_353
timestamp 1623621585
transform 1 0 33580 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _746_
timestamp 1623621585
transform 1 0 33948 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1102
timestamp 1623621585
transform 1 0 35236 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_363
timestamp 1623621585
transform 1 0 34500 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_372
timestamp 1623621585
transform 1 0 35328 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _753_
timestamp 1623621585
transform 1 0 37168 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_95_384
timestamp 1623621585
transform 1 0 36432 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1623621585
transform -1 0 38824 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_398
timestamp 1623621585
transform 1 0 37720 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_406
timestamp 1623621585
transform 1 0 38456 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1623621585
transform 1 0 1104 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input409
timestamp 1623621585
transform 1 0 1380 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_6
timestamp 1623621585
transform 1 0 1656 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_18
timestamp 1623621585
transform 1 0 2760 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_30
timestamp 1623621585
transform 1 0 3864 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1103
timestamp 1623621585
transform 1 0 6348 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_42
timestamp 1623621585
transform 1 0 4968 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_96_54
timestamp 1623621585
transform 1 0 6072 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_58
timestamp 1623621585
transform 1 0 6440 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_70
timestamp 1623621585
transform 1 0 7544 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_82
timestamp 1623621585
transform 1 0 8648 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_94
timestamp 1623621585
transform 1 0 9752 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1104
timestamp 1623621585
transform 1 0 11592 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_106
timestamp 1623621585
transform 1 0 10856 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_115
timestamp 1623621585
transform 1 0 11684 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_127
timestamp 1623621585
transform 1 0 12788 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_139
timestamp 1623621585
transform 1 0 13892 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_151
timestamp 1623621585
transform 1 0 14996 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_163
timestamp 1623621585
transform 1 0 16100 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1105
timestamp 1623621585
transform 1 0 16836 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_172
timestamp 1623621585
transform 1 0 16928 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_184
timestamp 1623621585
transform 1 0 18032 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_196
timestamp 1623621585
transform 1 0 19136 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_208
timestamp 1623621585
transform 1 0 20240 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1106
timestamp 1623621585
transform 1 0 22080 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_220
timestamp 1623621585
transform 1 0 21344 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_229
timestamp 1623621585
transform 1 0 22172 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_241
timestamp 1623621585
transform 1 0 23276 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_253
timestamp 1623621585
transform 1 0 24380 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_265
timestamp 1623621585
transform 1 0 25484 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1107
timestamp 1623621585
transform 1 0 27324 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_277
timestamp 1623621585
transform 1 0 26588 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_286
timestamp 1623621585
transform 1 0 27416 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_298
timestamp 1623621585
transform 1 0 28520 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_310
timestamp 1623621585
transform 1 0 29624 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_322
timestamp 1623621585
transform 1 0 30728 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _387_
timestamp 1623621585
transform 1 0 33120 0 -1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1108
timestamp 1623621585
transform 1 0 32568 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_334
timestamp 1623621585
transform 1 0 31832 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_96_343
timestamp 1623621585
transform 1 0 32660 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_347
timestamp 1623621585
transform 1 0 33028 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_357
timestamp 1623621585
transform 1 0 33948 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_369
timestamp 1623621585
transform 1 0 35052 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input148
timestamp 1623621585
transform 1 0 37168 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_96_381
timestamp 1623621585
transform 1 0 36156 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_96_389
timestamp 1623621585
transform 1 0 36892 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_395
timestamp 1623621585
transform 1 0 37444 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1623621585
transform -1 0 38824 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1109
timestamp 1623621585
transform 1 0 37812 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_400
timestamp 1623621585
transform 1 0 37904 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_406
timestamp 1623621585
transform 1 0 38456 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1623621585
transform 1 0 1104 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input410
timestamp 1623621585
transform 1 0 1380 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_6
timestamp 1623621585
transform 1 0 1656 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_18
timestamp 1623621585
transform 1 0 2760 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1110
timestamp 1623621585
transform 1 0 3772 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_97_26
timestamp 1623621585
transform 1 0 3496 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_30
timestamp 1623621585
transform 1 0 3864 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_42
timestamp 1623621585
transform 1 0 4968 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_54
timestamp 1623621585
transform 1 0 6072 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_66
timestamp 1623621585
transform 1 0 7176 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_78
timestamp 1623621585
transform 1 0 8280 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1111
timestamp 1623621585
transform 1 0 9016 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_87
timestamp 1623621585
transform 1 0 9108 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_99
timestamp 1623621585
transform 1 0 10212 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_111
timestamp 1623621585
transform 1 0 11316 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_123
timestamp 1623621585
transform 1 0 12420 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1112
timestamp 1623621585
transform 1 0 14260 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_135
timestamp 1623621585
transform 1 0 13524 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_144
timestamp 1623621585
transform 1 0 14352 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_156
timestamp 1623621585
transform 1 0 15456 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_168
timestamp 1623621585
transform 1 0 16560 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_180
timestamp 1623621585
transform 1 0 17664 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1113
timestamp 1623621585
transform 1 0 19504 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_192
timestamp 1623621585
transform 1 0 18768 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_201
timestamp 1623621585
transform 1 0 19596 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_213
timestamp 1623621585
transform 1 0 20700 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_225
timestamp 1623621585
transform 1 0 21804 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_237
timestamp 1623621585
transform 1 0 22908 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_249
timestamp 1623621585
transform 1 0 24012 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1114
timestamp 1623621585
transform 1 0 24748 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_258
timestamp 1623621585
transform 1 0 24840 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_270
timestamp 1623621585
transform 1 0 25944 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_282
timestamp 1623621585
transform 1 0 27048 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_294
timestamp 1623621585
transform 1 0 28152 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_306
timestamp 1623621585
transform 1 0 29256 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1115
timestamp 1623621585
transform 1 0 29992 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_315
timestamp 1623621585
transform 1 0 30084 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_327
timestamp 1623621585
transform 1 0 31188 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _365_
timestamp 1623621585
transform 1 0 33212 0 1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _401_
timestamp 1623621585
transform 1 0 32016 0 1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1623621585
transform 1 0 31924 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_345
timestamp 1623621585
transform 1 0 32844 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1116
timestamp 1623621585
transform 1 0 35236 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_358
timestamp 1623621585
transform 1 0 34040 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_370
timestamp 1623621585
transform 1 0 35144 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_372
timestamp 1623621585
transform 1 0 35328 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input182
timestamp 1623621585
transform 1 0 37260 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_97_384
timestamp 1623621585
transform 1 0 36432 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_392
timestamp 1623621585
transform 1 0 37168 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1623621585
transform -1 0 38824 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input118
timestamp 1623621585
transform 1 0 37904 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_396
timestamp 1623621585
transform 1 0 37536 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_403
timestamp 1623621585
transform 1 0 38180 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1623621585
transform 1 0 1104 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_3
timestamp 1623621585
transform 1 0 1380 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_15
timestamp 1623621585
transform 1 0 2484 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_27
timestamp 1623621585
transform 1 0 3588 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_39
timestamp 1623621585
transform 1 0 4692 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1117
timestamp 1623621585
transform 1 0 6348 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_51
timestamp 1623621585
transform 1 0 5796 0 -1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_98_58
timestamp 1623621585
transform 1 0 6440 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_70
timestamp 1623621585
transform 1 0 7544 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_82
timestamp 1623621585
transform 1 0 8648 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_94
timestamp 1623621585
transform 1 0 9752 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1118
timestamp 1623621585
transform 1 0 11592 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_106
timestamp 1623621585
transform 1 0 10856 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_115
timestamp 1623621585
transform 1 0 11684 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_127
timestamp 1623621585
transform 1 0 12788 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_139
timestamp 1623621585
transform 1 0 13892 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_151
timestamp 1623621585
transform 1 0 14996 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_163
timestamp 1623621585
transform 1 0 16100 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1119
timestamp 1623621585
transform 1 0 16836 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_172
timestamp 1623621585
transform 1 0 16928 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_184
timestamp 1623621585
transform 1 0 18032 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_196
timestamp 1623621585
transform 1 0 19136 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_208
timestamp 1623621585
transform 1 0 20240 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1120
timestamp 1623621585
transform 1 0 22080 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_220
timestamp 1623621585
transform 1 0 21344 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_229
timestamp 1623621585
transform 1 0 22172 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_241
timestamp 1623621585
transform 1 0 23276 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_253
timestamp 1623621585
transform 1 0 24380 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_265
timestamp 1623621585
transform 1 0 25484 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1121
timestamp 1623621585
transform 1 0 27324 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_277
timestamp 1623621585
transform 1 0 26588 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_286
timestamp 1623621585
transform 1 0 27416 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_298
timestamp 1623621585
transform 1 0 28520 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_310
timestamp 1623621585
transform 1 0 29624 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_322
timestamp 1623621585
transform 1 0 30728 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _381_
timestamp 1623621585
transform 1 0 33212 0 -1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1122
timestamp 1623621585
transform 1 0 32568 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_334
timestamp 1623621585
transform 1 0 31832 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_98_343
timestamp 1623621585
transform 1 0 32660 0 -1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_98_358
timestamp 1623621585
transform 1 0 34040 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_370
timestamp 1623621585
transform 1 0 35144 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input150
timestamp 1623621585
transform 1 0 37168 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_98_382
timestamp 1623621585
transform 1 0 36248 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_390
timestamp 1623621585
transform 1 0 36984 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_395
timestamp 1623621585
transform 1 0 37444 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1623621585
transform -1 0 38824 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1123
timestamp 1623621585
transform 1 0 37812 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_400
timestamp 1623621585
transform 1 0 37904 0 -1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_406
timestamp 1623621585
transform 1 0 38456 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1623621585
transform 1 0 1104 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1623621585
transform 1 0 1104 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input411
timestamp 1623621585
transform 1 0 1380 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input412
timestamp 1623621585
transform 1 0 1380 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_6
timestamp 1623621585
transform 1 0 1656 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_18
timestamp 1623621585
transform 1 0 2760 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_6
timestamp 1623621585
transform 1 0 1656 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_18
timestamp 1623621585
transform 1 0 2760 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1124
timestamp 1623621585
transform 1 0 3772 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_99_26
timestamp 1623621585
transform 1 0 3496 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_30
timestamp 1623621585
transform 1 0 3864 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_30
timestamp 1623621585
transform 1 0 3864 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1131
timestamp 1623621585
transform 1 0 6348 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_42
timestamp 1623621585
transform 1 0 4968 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_54
timestamp 1623621585
transform 1 0 6072 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_42
timestamp 1623621585
transform 1 0 4968 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_54
timestamp 1623621585
transform 1 0 6072 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_58
timestamp 1623621585
transform 1 0 6440 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_66
timestamp 1623621585
transform 1 0 7176 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_78
timestamp 1623621585
transform 1 0 8280 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_70
timestamp 1623621585
transform 1 0 7544 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_82
timestamp 1623621585
transform 1 0 8648 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1125
timestamp 1623621585
transform 1 0 9016 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_87
timestamp 1623621585
transform 1 0 9108 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_99
timestamp 1623621585
transform 1 0 10212 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_94
timestamp 1623621585
transform 1 0 9752 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1132
timestamp 1623621585
transform 1 0 11592 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_111
timestamp 1623621585
transform 1 0 11316 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_123
timestamp 1623621585
transform 1 0 12420 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_106
timestamp 1623621585
transform 1 0 10856 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_115
timestamp 1623621585
transform 1 0 11684 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1126
timestamp 1623621585
transform 1 0 14260 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_135
timestamp 1623621585
transform 1 0 13524 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_99_144
timestamp 1623621585
transform 1 0 14352 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_127
timestamp 1623621585
transform 1 0 12788 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_139
timestamp 1623621585
transform 1 0 13892 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _565_
timestamp 1623621585
transform 1 0 16284 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _577_
timestamp 1623621585
transform 1 0 15364 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_99_152
timestamp 1623621585
transform 1 0 15088 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_161
timestamp 1623621585
transform 1 0 15916 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_151
timestamp 1623621585
transform 1 0 14996 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_163
timestamp 1623621585
transform 1 0 16100 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _571_
timestamp 1623621585
transform 1 0 17204 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1133
timestamp 1623621585
transform 1 0 16836 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_2
timestamp 1623621585
transform 1 0 17020 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_171
timestamp 1623621585
transform 1 0 16836 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_99_181
timestamp 1623621585
transform 1 0 17756 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_172
timestamp 1623621585
transform 1 0 16928 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_184
timestamp 1623621585
transform 1 0 18032 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1127
timestamp 1623621585
transform 1 0 19504 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_193
timestamp 1623621585
transform 1 0 18860 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_199
timestamp 1623621585
transform 1 0 19412 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_201
timestamp 1623621585
transform 1 0 19596 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_196
timestamp 1623621585
transform 1 0 19136 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_208
timestamp 1623621585
transform 1 0 20240 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1134
timestamp 1623621585
transform 1 0 22080 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_213
timestamp 1623621585
transform 1 0 20700 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_225
timestamp 1623621585
transform 1 0 21804 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_220
timestamp 1623621585
transform 1 0 21344 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_229
timestamp 1623621585
transform 1 0 22172 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_237
timestamp 1623621585
transform 1 0 22908 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_249
timestamp 1623621585
transform 1 0 24012 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_241
timestamp 1623621585
transform 1 0 23276 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1128
timestamp 1623621585
transform 1 0 24748 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_258
timestamp 1623621585
transform 1 0 24840 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_270
timestamp 1623621585
transform 1 0 25944 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_253
timestamp 1623621585
transform 1 0 24380 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_265
timestamp 1623621585
transform 1 0 25484 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1135
timestamp 1623621585
transform 1 0 27324 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_282
timestamp 1623621585
transform 1 0 27048 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_277
timestamp 1623621585
transform 1 0 26588 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_286
timestamp 1623621585
transform 1 0 27416 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_294
timestamp 1623621585
transform 1 0 28152 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_306
timestamp 1623621585
transform 1 0 29256 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_298
timestamp 1623621585
transform 1 0 28520 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_310
timestamp 1623621585
transform 1 0 29624 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1129
timestamp 1623621585
transform 1 0 29992 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_315
timestamp 1623621585
transform 1 0 30084 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_327
timestamp 1623621585
transform 1 0 31188 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_322
timestamp 1623621585
transform 1 0 30728 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _394_
timestamp 1623621585
transform 1 0 33028 0 1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1136
timestamp 1623621585
transform 1 0 32568 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_339
timestamp 1623621585
transform 1 0 32292 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_100_334
timestamp 1623621585
transform 1 0 31832 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_343
timestamp 1623621585
transform 1 0 32660 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1130
timestamp 1623621585
transform 1 0 35236 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_356
timestamp 1623621585
transform 1 0 33856 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_368
timestamp 1623621585
transform 1 0 34960 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_372
timestamp 1623621585
transform 1 0 35328 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_355
timestamp 1623621585
transform 1 0 33764 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_367
timestamp 1623621585
transform 1 0 34868 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input183
timestamp 1623621585
transform 1 0 37260 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_99_384
timestamp 1623621585
transform 1 0 36432 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_392
timestamp 1623621585
transform 1 0 37168 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_379
timestamp 1623621585
transform 1 0 35972 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_391
timestamp 1623621585
transform 1 0 37076 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1623621585
transform -1 0 38824 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1623621585
transform -1 0 38824 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1137
timestamp 1623621585
transform 1 0 37812 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input119
timestamp 1623621585
transform 1 0 37904 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_396
timestamp 1623621585
transform 1 0 37536 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_403
timestamp 1623621585
transform 1 0 38180 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_400
timestamp 1623621585
transform 1 0 37904 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_406
timestamp 1623621585
transform 1 0 38456 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1623621585
transform 1 0 1104 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_3
timestamp 1623621585
transform 1 0 1380 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_15
timestamp 1623621585
transform 1 0 2484 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1138
timestamp 1623621585
transform 1 0 3772 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_27
timestamp 1623621585
transform 1 0 3588 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_101_30
timestamp 1623621585
transform 1 0 3864 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_42
timestamp 1623621585
transform 1 0 4968 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_54
timestamp 1623621585
transform 1 0 6072 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_66
timestamp 1623621585
transform 1 0 7176 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_78
timestamp 1623621585
transform 1 0 8280 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1139
timestamp 1623621585
transform 1 0 9016 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_87
timestamp 1623621585
transform 1 0 9108 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_99
timestamp 1623621585
transform 1 0 10212 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_111
timestamp 1623621585
transform 1 0 11316 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_123
timestamp 1623621585
transform 1 0 12420 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1140
timestamp 1623621585
transform 1 0 14260 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_135
timestamp 1623621585
transform 1 0 13524 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_144
timestamp 1623621585
transform 1 0 14352 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_156
timestamp 1623621585
transform 1 0 15456 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_168
timestamp 1623621585
transform 1 0 16560 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_180
timestamp 1623621585
transform 1 0 17664 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1141
timestamp 1623621585
transform 1 0 19504 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_192
timestamp 1623621585
transform 1 0 18768 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_201
timestamp 1623621585
transform 1 0 19596 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_213
timestamp 1623621585
transform 1 0 20700 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_225
timestamp 1623621585
transform 1 0 21804 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_237
timestamp 1623621585
transform 1 0 22908 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_249
timestamp 1623621585
transform 1 0 24012 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1142
timestamp 1623621585
transform 1 0 24748 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_258
timestamp 1623621585
transform 1 0 24840 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_270
timestamp 1623621585
transform 1 0 25944 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_282
timestamp 1623621585
transform 1 0 27048 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_294
timestamp 1623621585
transform 1 0 28152 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_306
timestamp 1623621585
transform 1 0 29256 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1143
timestamp 1623621585
transform 1 0 29992 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_315
timestamp 1623621585
transform 1 0 30084 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_327
timestamp 1623621585
transform 1 0 31188 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_339
timestamp 1623621585
transform 1 0 32292 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_351
timestamp 1623621585
transform 1 0 33396 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1144
timestamp 1623621585
transform 1 0 35236 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_363
timestamp 1623621585
transform 1 0 34500 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_372
timestamp 1623621585
transform 1 0 35328 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input191
timestamp 1623621585
transform 1 0 37260 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_384
timestamp 1623621585
transform 1 0 36432 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_392
timestamp 1623621585
transform 1 0 37168 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1623621585
transform -1 0 38824 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input151
timestamp 1623621585
transform 1 0 37904 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_396
timestamp 1623621585
transform 1 0 37536 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_403
timestamp 1623621585
transform 1 0 38180 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1623621585
transform 1 0 1104 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input413
timestamp 1623621585
transform 1 0 1380 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_102_6
timestamp 1623621585
transform 1 0 1656 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_18
timestamp 1623621585
transform 1 0 2760 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_30
timestamp 1623621585
transform 1 0 3864 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1145
timestamp 1623621585
transform 1 0 6348 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_42
timestamp 1623621585
transform 1 0 4968 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_102_54
timestamp 1623621585
transform 1 0 6072 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_102_58
timestamp 1623621585
transform 1 0 6440 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_70
timestamp 1623621585
transform 1 0 7544 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_82
timestamp 1623621585
transform 1 0 8648 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_94
timestamp 1623621585
transform 1 0 9752 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1146
timestamp 1623621585
transform 1 0 11592 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_106
timestamp 1623621585
transform 1 0 10856 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_115
timestamp 1623621585
transform 1 0 11684 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_127
timestamp 1623621585
transform 1 0 12788 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_139
timestamp 1623621585
transform 1 0 13892 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_151
timestamp 1623621585
transform 1 0 14996 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_163
timestamp 1623621585
transform 1 0 16100 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1147
timestamp 1623621585
transform 1 0 16836 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_172
timestamp 1623621585
transform 1 0 16928 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_184
timestamp 1623621585
transform 1 0 18032 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_196
timestamp 1623621585
transform 1 0 19136 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_208
timestamp 1623621585
transform 1 0 20240 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1148
timestamp 1623621585
transform 1 0 22080 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_220
timestamp 1623621585
transform 1 0 21344 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_229
timestamp 1623621585
transform 1 0 22172 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_241
timestamp 1623621585
transform 1 0 23276 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_253
timestamp 1623621585
transform 1 0 24380 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_265
timestamp 1623621585
transform 1 0 25484 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1149
timestamp 1623621585
transform 1 0 27324 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_277
timestamp 1623621585
transform 1 0 26588 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_286
timestamp 1623621585
transform 1 0 27416 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_298
timestamp 1623621585
transform 1 0 28520 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_310
timestamp 1623621585
transform 1 0 29624 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_322
timestamp 1623621585
transform 1 0 30728 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1150
timestamp 1623621585
transform 1 0 32568 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_334
timestamp 1623621585
transform 1 0 31832 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_343
timestamp 1623621585
transform 1 0 32660 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_355
timestamp 1623621585
transform 1 0 33764 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_367
timestamp 1623621585
transform 1 0 34868 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input202
timestamp 1623621585
transform 1 0 37168 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input216
timestamp 1623621585
transform 1 0 36524 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_102_379
timestamp 1623621585
transform 1 0 35972 0 -1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_102_388
timestamp 1623621585
transform 1 0 36800 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_395
timestamp 1623621585
transform 1 0 37444 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1623621585
transform -1 0 38824 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1151
timestamp 1623621585
transform 1 0 37812 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_102_400
timestamp 1623621585
transform 1 0 37904 0 -1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_406
timestamp 1623621585
transform 1 0 38456 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1623621585
transform 1 0 1104 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input414
timestamp 1623621585
transform 1 0 1380 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_6
timestamp 1623621585
transform 1 0 1656 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_18
timestamp 1623621585
transform 1 0 2760 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1152
timestamp 1623621585
transform 1 0 3772 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_103_26
timestamp 1623621585
transform 1 0 3496 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_30
timestamp 1623621585
transform 1 0 3864 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_42
timestamp 1623621585
transform 1 0 4968 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_54
timestamp 1623621585
transform 1 0 6072 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_66
timestamp 1623621585
transform 1 0 7176 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_78
timestamp 1623621585
transform 1 0 8280 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1153
timestamp 1623621585
transform 1 0 9016 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_87
timestamp 1623621585
transform 1 0 9108 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_99
timestamp 1623621585
transform 1 0 10212 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_111
timestamp 1623621585
transform 1 0 11316 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_123
timestamp 1623621585
transform 1 0 12420 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1154
timestamp 1623621585
transform 1 0 14260 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_103_135
timestamp 1623621585
transform 1 0 13524 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_103_144
timestamp 1623621585
transform 1 0 14352 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_156
timestamp 1623621585
transform 1 0 15456 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_168
timestamp 1623621585
transform 1 0 16560 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_180
timestamp 1623621585
transform 1 0 17664 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1155
timestamp 1623621585
transform 1 0 19504 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_103_192
timestamp 1623621585
transform 1 0 18768 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_103_201
timestamp 1623621585
transform 1 0 19596 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_213
timestamp 1623621585
transform 1 0 20700 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_225
timestamp 1623621585
transform 1 0 21804 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_237
timestamp 1623621585
transform 1 0 22908 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_249
timestamp 1623621585
transform 1 0 24012 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1156
timestamp 1623621585
transform 1 0 24748 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_258
timestamp 1623621585
transform 1 0 24840 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_270
timestamp 1623621585
transform 1 0 25944 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_282
timestamp 1623621585
transform 1 0 27048 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_294
timestamp 1623621585
transform 1 0 28152 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_306
timestamp 1623621585
transform 1 0 29256 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1157
timestamp 1623621585
transform 1 0 29992 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_315
timestamp 1623621585
transform 1 0 30084 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_327
timestamp 1623621585
transform 1 0 31188 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_4  _441_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 32384 0 1 58208
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_103_339
timestamp 1623621585
transform 1 0 32292 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1158
timestamp 1623621585
transform 1 0 35236 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_357
timestamp 1623621585
transform 1 0 33948 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_369
timestamp 1623621585
transform 1 0 35052 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_103_372
timestamp 1623621585
transform 1 0 35328 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 37076 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input213
timestamp 1623621585
transform 1 0 36432 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input217
timestamp 1623621585
transform 1 0 35788 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_103_376
timestamp 1623621585
transform 1 0 35696 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_380
timestamp 1623621585
transform 1 0 36064 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_387
timestamp 1623621585
transform 1 0 36708 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1623621585
transform -1 0 38824 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_103_399
timestamp 1623621585
transform 1 0 37812 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1623621585
transform 1 0 1104 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_104_3
timestamp 1623621585
transform 1 0 1380 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_15
timestamp 1623621585
transform 1 0 2484 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_27
timestamp 1623621585
transform 1 0 3588 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_39
timestamp 1623621585
transform 1 0 4692 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1159
timestamp 1623621585
transform 1 0 6348 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_104_51
timestamp 1623621585
transform 1 0 5796 0 -1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_104_58
timestamp 1623621585
transform 1 0 6440 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_70
timestamp 1623621585
transform 1 0 7544 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_82
timestamp 1623621585
transform 1 0 8648 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_94
timestamp 1623621585
transform 1 0 9752 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1160
timestamp 1623621585
transform 1 0 11592 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_106
timestamp 1623621585
transform 1 0 10856 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_115
timestamp 1623621585
transform 1 0 11684 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_127
timestamp 1623621585
transform 1 0 12788 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_139
timestamp 1623621585
transform 1 0 13892 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_151
timestamp 1623621585
transform 1 0 14996 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_163
timestamp 1623621585
transform 1 0 16100 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1161
timestamp 1623621585
transform 1 0 16836 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_172
timestamp 1623621585
transform 1 0 16928 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_184
timestamp 1623621585
transform 1 0 18032 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_196
timestamp 1623621585
transform 1 0 19136 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_208
timestamp 1623621585
transform 1 0 20240 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1162
timestamp 1623621585
transform 1 0 22080 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_220
timestamp 1623621585
transform 1 0 21344 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_229
timestamp 1623621585
transform 1 0 22172 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_241
timestamp 1623621585
transform 1 0 23276 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_253
timestamp 1623621585
transform 1 0 24380 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_265
timestamp 1623621585
transform 1 0 25484 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1163
timestamp 1623621585
transform 1 0 27324 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_277
timestamp 1623621585
transform 1 0 26588 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_286
timestamp 1623621585
transform 1 0 27416 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_298
timestamp 1623621585
transform 1 0 28520 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_310
timestamp 1623621585
transform 1 0 29624 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _421_
timestamp 1623621585
transform 1 0 31372 0 -1 59296
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_104_322
timestamp 1623621585
transform 1 0 30728 0 -1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_328
timestamp 1623621585
transform 1 0 31280 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_4  _427_
timestamp 1623621585
transform 1 0 33028 0 -1 59296
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1164
timestamp 1623621585
transform 1 0 32568 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_338
timestamp 1623621585
transform 1 0 32200 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_343
timestamp 1623621585
transform 1 0 32660 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _579_
timestamp 1623621585
transform 1 0 35604 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_104_364
timestamp 1623621585
transform 1 0 34592 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_104_372
timestamp 1623621585
transform 1 0 35328 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _555_
timestamp 1623621585
transform 1 0 36708 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_104_383
timestamp 1623621585
transform 1 0 36340 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_395
timestamp 1623621585
transform 1 0 37444 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1623621585
transform -1 0 38824 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1165
timestamp 1623621585
transform 1 0 37812 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_104_400
timestamp 1623621585
transform 1 0 37904 0 -1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_406
timestamp 1623621585
transform 1 0 38456 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1623621585
transform 1 0 1104 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1623621585
transform 1 0 1104 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input384
timestamp 1623621585
transform 1 0 1380 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input385
timestamp 1623621585
transform 1 0 1380 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_105_6
timestamp 1623621585
transform 1 0 1656 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_18
timestamp 1623621585
transform 1 0 2760 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_6
timestamp 1623621585
transform 1 0 1656 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_18
timestamp 1623621585
transform 1 0 2760 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1166
timestamp 1623621585
transform 1 0 3772 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_105_26
timestamp 1623621585
transform 1 0 3496 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_105_30
timestamp 1623621585
transform 1 0 3864 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_30
timestamp 1623621585
transform 1 0 3864 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1173
timestamp 1623621585
transform 1 0 6348 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_42
timestamp 1623621585
transform 1 0 4968 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_54
timestamp 1623621585
transform 1 0 6072 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_42
timestamp 1623621585
transform 1 0 4968 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_54
timestamp 1623621585
transform 1 0 6072 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_58
timestamp 1623621585
transform 1 0 6440 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_66
timestamp 1623621585
transform 1 0 7176 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_78
timestamp 1623621585
transform 1 0 8280 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_70
timestamp 1623621585
transform 1 0 7544 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_82
timestamp 1623621585
transform 1 0 8648 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1167
timestamp 1623621585
transform 1 0 9016 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_87
timestamp 1623621585
transform 1 0 9108 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_99
timestamp 1623621585
transform 1 0 10212 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_94
timestamp 1623621585
transform 1 0 9752 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1174
timestamp 1623621585
transform 1 0 11592 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_111
timestamp 1623621585
transform 1 0 11316 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_123
timestamp 1623621585
transform 1 0 12420 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_106
timestamp 1623621585
transform 1 0 10856 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_115
timestamp 1623621585
transform 1 0 11684 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1168
timestamp 1623621585
transform 1 0 14260 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_135
timestamp 1623621585
transform 1 0 13524 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_144
timestamp 1623621585
transform 1 0 14352 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_127
timestamp 1623621585
transform 1 0 12788 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_139
timestamp 1623621585
transform 1 0 13892 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_156
timestamp 1623621585
transform 1 0 15456 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_151
timestamp 1623621585
transform 1 0 14996 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_163
timestamp 1623621585
transform 1 0 16100 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1175
timestamp 1623621585
transform 1 0 16836 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_168
timestamp 1623621585
transform 1 0 16560 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_180
timestamp 1623621585
transform 1 0 17664 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_172
timestamp 1623621585
transform 1 0 16928 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_184
timestamp 1623621585
transform 1 0 18032 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1169
timestamp 1623621585
transform 1 0 19504 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_192
timestamp 1623621585
transform 1 0 18768 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_201
timestamp 1623621585
transform 1 0 19596 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_196
timestamp 1623621585
transform 1 0 19136 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_208
timestamp 1623621585
transform 1 0 20240 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1176
timestamp 1623621585
transform 1 0 22080 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_213
timestamp 1623621585
transform 1 0 20700 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_225
timestamp 1623621585
transform 1 0 21804 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_220
timestamp 1623621585
transform 1 0 21344 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_229
timestamp 1623621585
transform 1 0 22172 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_237
timestamp 1623621585
transform 1 0 22908 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_249
timestamp 1623621585
transform 1 0 24012 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_241
timestamp 1623621585
transform 1 0 23276 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1170
timestamp 1623621585
transform 1 0 24748 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_258
timestamp 1623621585
transform 1 0 24840 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_270
timestamp 1623621585
transform 1 0 25944 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_253
timestamp 1623621585
transform 1 0 24380 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_265
timestamp 1623621585
transform 1 0 25484 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1177
timestamp 1623621585
transform 1 0 27324 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_282
timestamp 1623621585
transform 1 0 27048 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_277
timestamp 1623621585
transform 1 0 26588 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_286
timestamp 1623621585
transform 1 0 27416 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_294
timestamp 1623621585
transform 1 0 28152 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_306
timestamp 1623621585
transform 1 0 29256 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_298
timestamp 1623621585
transform 1 0 28520 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_310
timestamp 1623621585
transform 1 0 29624 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1171
timestamp 1623621585
transform 1 0 29992 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_315
timestamp 1623621585
transform 1 0 30084 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_327
timestamp 1623621585
transform 1 0 31188 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_322
timestamp 1623621585
transform 1 0 30728 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _410_
timestamp 1623621585
transform 1 0 33028 0 -1 60384
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_4  _434_
timestamp 1623621585
transform 1 0 32476 0 1 59296
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1178
timestamp 1623621585
transform 1 0 32568 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_339
timestamp 1623621585
transform 1 0 32292 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_106_334
timestamp 1623621585
transform 1 0 31832 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_106_343
timestamp 1623621585
transform 1 0 32660 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _549_
timestamp 1623621585
transform 1 0 35604 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1172
timestamp 1623621585
transform 1 0 35236 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input218
timestamp 1623621585
transform 1 0 34592 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input219
timestamp 1623621585
transform 1 0 34960 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_105_358
timestamp 1623621585
transform 1 0 34040 0 1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_105_367
timestamp 1623621585
transform 1 0 34868 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_105_372
timestamp 1623621585
transform 1 0 35328 0 1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_106_356
timestamp 1623621585
transform 1 0 33856 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_371
timestamp 1623621585
transform 1 0 35236 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _536_
timestamp 1623621585
transform 1 0 36708 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _542_
timestamp 1623621585
transform 1 0 37076 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _573_
timestamp 1623621585
transform 1 0 35972 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_105_378
timestamp 1623621585
transform 1 0 35880 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_387
timestamp 1623621585
transform 1 0 36708 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_383
timestamp 1623621585
transform 1 0 36340 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_395
timestamp 1623621585
transform 1 0 37444 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1623621585
transform -1 0 38824 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1623621585
transform -1 0 38824 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1179
timestamp 1623621585
transform 1 0 37812 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_399
timestamp 1623621585
transform 1 0 37812 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_106_400
timestamp 1623621585
transform 1 0 37904 0 -1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_406
timestamp 1623621585
transform 1 0 38456 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1623621585
transform 1 0 1104 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_3
timestamp 1623621585
transform 1 0 1380 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_15
timestamp 1623621585
transform 1 0 2484 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1180
timestamp 1623621585
transform 1 0 3772 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_107_27
timestamp 1623621585
transform 1 0 3588 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_107_30
timestamp 1623621585
transform 1 0 3864 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_42
timestamp 1623621585
transform 1 0 4968 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_54
timestamp 1623621585
transform 1 0 6072 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_66
timestamp 1623621585
transform 1 0 7176 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_78
timestamp 1623621585
transform 1 0 8280 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1181
timestamp 1623621585
transform 1 0 9016 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_87
timestamp 1623621585
transform 1 0 9108 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_99
timestamp 1623621585
transform 1 0 10212 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_111
timestamp 1623621585
transform 1 0 11316 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_123
timestamp 1623621585
transform 1 0 12420 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1182
timestamp 1623621585
transform 1 0 14260 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_107_135
timestamp 1623621585
transform 1 0 13524 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_144
timestamp 1623621585
transform 1 0 14352 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_156
timestamp 1623621585
transform 1 0 15456 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_168
timestamp 1623621585
transform 1 0 16560 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_180
timestamp 1623621585
transform 1 0 17664 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1183
timestamp 1623621585
transform 1 0 19504 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_107_192
timestamp 1623621585
transform 1 0 18768 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_201
timestamp 1623621585
transform 1 0 19596 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_213
timestamp 1623621585
transform 1 0 20700 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_225
timestamp 1623621585
transform 1 0 21804 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_237
timestamp 1623621585
transform 1 0 22908 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_249
timestamp 1623621585
transform 1 0 24012 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1184
timestamp 1623621585
transform 1 0 24748 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_258
timestamp 1623621585
transform 1 0 24840 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_270
timestamp 1623621585
transform 1 0 25944 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_282
timestamp 1623621585
transform 1 0 27048 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_294
timestamp 1623621585
transform 1 0 28152 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_306
timestamp 1623621585
transform 1 0 29256 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1185
timestamp 1623621585
transform 1 0 29992 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_315
timestamp 1623621585
transform 1 0 30084 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_327
timestamp 1623621585
transform 1 0 31188 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_339
timestamp 1623621585
transform 1 0 32292 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_351
timestamp 1623621585
transform 1 0 33396 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1186
timestamp 1623621585
transform 1 0 35236 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_107_363
timestamp 1623621585
transform 1 0 34500 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_107_372
timestamp 1623621585
transform 1 0 35328 0 1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _522_
timestamp 1623621585
transform 1 0 37076 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _567_
timestamp 1623621585
transform 1 0 35972 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_378
timestamp 1623621585
transform 1 0 35880 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_387
timestamp 1623621585
transform 1 0 36708 0 1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1623621585
transform -1 0 38824 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_107_399
timestamp 1623621585
transform 1 0 37812 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1623621585
transform 1 0 1104 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input386
timestamp 1623621585
transform 1 0 1380 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_108_6
timestamp 1623621585
transform 1 0 1656 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_18
timestamp 1623621585
transform 1 0 2760 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_30
timestamp 1623621585
transform 1 0 3864 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1187
timestamp 1623621585
transform 1 0 6348 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_42
timestamp 1623621585
transform 1 0 4968 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_108_54
timestamp 1623621585
transform 1 0 6072 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_108_58
timestamp 1623621585
transform 1 0 6440 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_70
timestamp 1623621585
transform 1 0 7544 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_82
timestamp 1623621585
transform 1 0 8648 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_94
timestamp 1623621585
transform 1 0 9752 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1188
timestamp 1623621585
transform 1 0 11592 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_106
timestamp 1623621585
transform 1 0 10856 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_115
timestamp 1623621585
transform 1 0 11684 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_127
timestamp 1623621585
transform 1 0 12788 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_139
timestamp 1623621585
transform 1 0 13892 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_151
timestamp 1623621585
transform 1 0 14996 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_163
timestamp 1623621585
transform 1 0 16100 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1189
timestamp 1623621585
transform 1 0 16836 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_172
timestamp 1623621585
transform 1 0 16928 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_184
timestamp 1623621585
transform 1 0 18032 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_196
timestamp 1623621585
transform 1 0 19136 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_208
timestamp 1623621585
transform 1 0 20240 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1190
timestamp 1623621585
transform 1 0 22080 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_220
timestamp 1623621585
transform 1 0 21344 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_229
timestamp 1623621585
transform 1 0 22172 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_241
timestamp 1623621585
transform 1 0 23276 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_253
timestamp 1623621585
transform 1 0 24380 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_265
timestamp 1623621585
transform 1 0 25484 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1191
timestamp 1623621585
transform 1 0 27324 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_277
timestamp 1623621585
transform 1 0 26588 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_286
timestamp 1623621585
transform 1 0 27416 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_298
timestamp 1623621585
transform 1 0 28520 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_310
timestamp 1623621585
transform 1 0 29624 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_322
timestamp 1623621585
transform 1 0 30728 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1192
timestamp 1623621585
transform 1 0 32568 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_334
timestamp 1623621585
transform 1 0 31832 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_343
timestamp 1623621585
transform 1 0 32660 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input220
timestamp 1623621585
transform 1 0 35328 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input222
timestamp 1623621585
transform 1 0 34684 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_108_355
timestamp 1623621585
transform 1 0 33764 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_363
timestamp 1623621585
transform 1 0 34500 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_368
timestamp 1623621585
transform 1 0 34960 0 -1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_375
timestamp 1623621585
transform 1 0 35604 0 -1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _515_
timestamp 1623621585
transform 1 0 36708 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _752_
timestamp 1623621585
transform 1 0 35972 0 -1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_383
timestamp 1623621585
transform 1 0 36340 0 -1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_395
timestamp 1623621585
transform 1 0 37444 0 -1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1623621585
transform -1 0 38824 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1193
timestamp 1623621585
transform 1 0 37812 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_400
timestamp 1623621585
transform 1 0 37904 0 -1 61472
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_406
timestamp 1623621585
transform 1 0 38456 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1623621585
transform 1 0 1104 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input387
timestamp 1623621585
transform 1 0 1380 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_109_6
timestamp 1623621585
transform 1 0 1656 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_18
timestamp 1623621585
transform 1 0 2760 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1194
timestamp 1623621585
transform 1 0 3772 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_109_26
timestamp 1623621585
transform 1 0 3496 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_109_30
timestamp 1623621585
transform 1 0 3864 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_42
timestamp 1623621585
transform 1 0 4968 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_54
timestamp 1623621585
transform 1 0 6072 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_66
timestamp 1623621585
transform 1 0 7176 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_78
timestamp 1623621585
transform 1 0 8280 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1195
timestamp 1623621585
transform 1 0 9016 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_87
timestamp 1623621585
transform 1 0 9108 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_99
timestamp 1623621585
transform 1 0 10212 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_111
timestamp 1623621585
transform 1 0 11316 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_123
timestamp 1623621585
transform 1 0 12420 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1196
timestamp 1623621585
transform 1 0 14260 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_109_135
timestamp 1623621585
transform 1 0 13524 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_144
timestamp 1623621585
transform 1 0 14352 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_156
timestamp 1623621585
transform 1 0 15456 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_168
timestamp 1623621585
transform 1 0 16560 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_180
timestamp 1623621585
transform 1 0 17664 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1197
timestamp 1623621585
transform 1 0 19504 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_109_192
timestamp 1623621585
transform 1 0 18768 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_201
timestamp 1623621585
transform 1 0 19596 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_213
timestamp 1623621585
transform 1 0 20700 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_225
timestamp 1623621585
transform 1 0 21804 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_237
timestamp 1623621585
transform 1 0 22908 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_249
timestamp 1623621585
transform 1 0 24012 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1198
timestamp 1623621585
transform 1 0 24748 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_258
timestamp 1623621585
transform 1 0 24840 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_270
timestamp 1623621585
transform 1 0 25944 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_282
timestamp 1623621585
transform 1 0 27048 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_294
timestamp 1623621585
transform 1 0 28152 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_306
timestamp 1623621585
transform 1 0 29256 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1199
timestamp 1623621585
transform 1 0 29992 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_315
timestamp 1623621585
transform 1 0 30084 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_327
timestamp 1623621585
transform 1 0 31188 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_339
timestamp 1623621585
transform 1 0 32292 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_351
timestamp 1623621585
transform 1 0 33396 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1200
timestamp 1623621585
transform 1 0 35236 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_109_363
timestamp 1623621585
transform 1 0 34500 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_109_372
timestamp 1623621585
transform 1 0 35328 0 1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _509_
timestamp 1623621585
transform 1 0 37076 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input192
timestamp 1623621585
transform 1 0 36432 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input221
timestamp 1623621585
transform 1 0 35788 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_109_376
timestamp 1623621585
transform 1 0 35696 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_109_380
timestamp 1623621585
transform 1 0 36064 0 1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_387
timestamp 1623621585
transform 1 0 36708 0 1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1623621585
transform -1 0 38824 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_109_399
timestamp 1623621585
transform 1 0 37812 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1623621585
transform 1 0 1104 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_3
timestamp 1623621585
transform 1 0 1380 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_15
timestamp 1623621585
transform 1 0 2484 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_27
timestamp 1623621585
transform 1 0 3588 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_39
timestamp 1623621585
transform 1 0 4692 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1201
timestamp 1623621585
transform 1 0 6348 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_110_51
timestamp 1623621585
transform 1 0 5796 0 -1 62560
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_110_58
timestamp 1623621585
transform 1 0 6440 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_70
timestamp 1623621585
transform 1 0 7544 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_82
timestamp 1623621585
transform 1 0 8648 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_94
timestamp 1623621585
transform 1 0 9752 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1202
timestamp 1623621585
transform 1 0 11592 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_106
timestamp 1623621585
transform 1 0 10856 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_115
timestamp 1623621585
transform 1 0 11684 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_127
timestamp 1623621585
transform 1 0 12788 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_139
timestamp 1623621585
transform 1 0 13892 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _749_
timestamp 1623621585
transform 1 0 15272 0 -1 62560
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_110_151
timestamp 1623621585
transform 1 0 14996 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_110_160
timestamp 1623621585
transform 1 0 15824 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1203
timestamp 1623621585
transform 1 0 16836 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_110_168
timestamp 1623621585
transform 1 0 16560 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_172
timestamp 1623621585
transform 1 0 16928 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_184
timestamp 1623621585
transform 1 0 18032 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_196
timestamp 1623621585
transform 1 0 19136 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_208
timestamp 1623621585
transform 1 0 20240 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1204
timestamp 1623621585
transform 1 0 22080 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_220
timestamp 1623621585
transform 1 0 21344 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_229
timestamp 1623621585
transform 1 0 22172 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_241
timestamp 1623621585
transform 1 0 23276 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_253
timestamp 1623621585
transform 1 0 24380 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_265
timestamp 1623621585
transform 1 0 25484 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1205
timestamp 1623621585
transform 1 0 27324 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_277
timestamp 1623621585
transform 1 0 26588 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_286
timestamp 1623621585
transform 1 0 27416 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_298
timestamp 1623621585
transform 1 0 28520 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_310
timestamp 1623621585
transform 1 0 29624 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_322
timestamp 1623621585
transform 1 0 30728 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1206
timestamp 1623621585
transform 1 0 32568 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_334
timestamp 1623621585
transform 1 0 31832 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_343
timestamp 1623621585
transform 1 0 32660 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input194
timestamp 1623621585
transform 1 0 35420 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_355
timestamp 1623621585
transform 1 0 33764 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_367
timestamp 1623621585
transform 1 0 34868 0 -1 62560
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _502_
timestamp 1623621585
transform 1 0 36708 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input193
timestamp 1623621585
transform 1 0 36064 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_110_376
timestamp 1623621585
transform 1 0 35696 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_383
timestamp 1623621585
transform 1 0 36340 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_395
timestamp 1623621585
transform 1 0 37444 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1623621585
transform -1 0 38824 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1207
timestamp 1623621585
transform 1 0 37812 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_110_400
timestamp 1623621585
transform 1 0 37904 0 -1 62560
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_406
timestamp 1623621585
transform 1 0 38456 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1623621585
transform 1 0 1104 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input388
timestamp 1623621585
transform 1 0 1380 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_111_6
timestamp 1623621585
transform 1 0 1656 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_18
timestamp 1623621585
transform 1 0 2760 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1208
timestamp 1623621585
transform 1 0 3772 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_111_26
timestamp 1623621585
transform 1 0 3496 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_111_30
timestamp 1623621585
transform 1 0 3864 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_42
timestamp 1623621585
transform 1 0 4968 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_54
timestamp 1623621585
transform 1 0 6072 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_66
timestamp 1623621585
transform 1 0 7176 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_78
timestamp 1623621585
transform 1 0 8280 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1209
timestamp 1623621585
transform 1 0 9016 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_87
timestamp 1623621585
transform 1 0 9108 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_99
timestamp 1623621585
transform 1 0 10212 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_111
timestamp 1623621585
transform 1 0 11316 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_123
timestamp 1623621585
transform 1 0 12420 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1210
timestamp 1623621585
transform 1 0 14260 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_111_135
timestamp 1623621585
transform 1 0 13524 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_144
timestamp 1623621585
transform 1 0 14352 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_156
timestamp 1623621585
transform 1 0 15456 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_168
timestamp 1623621585
transform 1 0 16560 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_180
timestamp 1623621585
transform 1 0 17664 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1211
timestamp 1623621585
transform 1 0 19504 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_111_192
timestamp 1623621585
transform 1 0 18768 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_201
timestamp 1623621585
transform 1 0 19596 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_213
timestamp 1623621585
transform 1 0 20700 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_225
timestamp 1623621585
transform 1 0 21804 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_237
timestamp 1623621585
transform 1 0 22908 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_249
timestamp 1623621585
transform 1 0 24012 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1212
timestamp 1623621585
transform 1 0 24748 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_258
timestamp 1623621585
transform 1 0 24840 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_270
timestamp 1623621585
transform 1 0 25944 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_282
timestamp 1623621585
transform 1 0 27048 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_294
timestamp 1623621585
transform 1 0 28152 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_306
timestamp 1623621585
transform 1 0 29256 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _361_
timestamp 1623621585
transform 1 0 31740 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1213
timestamp 1623621585
transform 1 0 29992 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_315
timestamp 1623621585
transform 1 0 30084 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_327
timestamp 1623621585
transform 1 0 31188 0 1 62560
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _359_
timestamp 1623621585
transform 1 0 32568 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_111_337
timestamp 1623621585
transform 1 0 32108 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_341
timestamp 1623621585
transform 1 0 32476 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_346
timestamp 1623621585
transform 1 0 32936 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1214
timestamp 1623621585
transform 1 0 35236 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_358
timestamp 1623621585
transform 1 0 34040 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_111_370
timestamp 1623621585
transform 1 0 35144 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_111_372
timestamp 1623621585
transform 1 0 35328 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _482_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 36064 0 1 62560
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _496_
timestamp 1623621585
transform 1 0 37076 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_111_387
timestamp 1623621585
transform 1 0 36708 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1623621585
transform -1 0 38824 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_111_399
timestamp 1623621585
transform 1 0 37812 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1623621585
transform 1 0 1104 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1623621585
transform 1 0 1104 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input389
timestamp 1623621585
transform 1 0 1380 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_112_6
timestamp 1623621585
transform 1 0 1656 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_18
timestamp 1623621585
transform 1 0 2760 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_3
timestamp 1623621585
transform 1 0 1380 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_15
timestamp 1623621585
transform 1 0 2484 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1222
timestamp 1623621585
transform 1 0 3772 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_30
timestamp 1623621585
transform 1 0 3864 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_113_27
timestamp 1623621585
transform 1 0 3588 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_113_30
timestamp 1623621585
transform 1 0 3864 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1215
timestamp 1623621585
transform 1 0 6348 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_42
timestamp 1623621585
transform 1 0 4968 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_112_54
timestamp 1623621585
transform 1 0 6072 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_112_58
timestamp 1623621585
transform 1 0 6440 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_42
timestamp 1623621585
transform 1 0 4968 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_54
timestamp 1623621585
transform 1 0 6072 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_70
timestamp 1623621585
transform 1 0 7544 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_82
timestamp 1623621585
transform 1 0 8648 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_66
timestamp 1623621585
transform 1 0 7176 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_78
timestamp 1623621585
transform 1 0 8280 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1223
timestamp 1623621585
transform 1 0 9016 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_94
timestamp 1623621585
transform 1 0 9752 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_87
timestamp 1623621585
transform 1 0 9108 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_99
timestamp 1623621585
transform 1 0 10212 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1216
timestamp 1623621585
transform 1 0 11592 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_106
timestamp 1623621585
transform 1 0 10856 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_115
timestamp 1623621585
transform 1 0 11684 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_111
timestamp 1623621585
transform 1 0 11316 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_123
timestamp 1623621585
transform 1 0 12420 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1224
timestamp 1623621585
transform 1 0 14260 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_127
timestamp 1623621585
transform 1 0 12788 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_139
timestamp 1623621585
transform 1 0 13892 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_135
timestamp 1623621585
transform 1 0 13524 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_144
timestamp 1623621585
transform 1 0 14352 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_151
timestamp 1623621585
transform 1 0 14996 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_163
timestamp 1623621585
transform 1 0 16100 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_156
timestamp 1623621585
transform 1 0 15456 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1217
timestamp 1623621585
transform 1 0 16836 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_172
timestamp 1623621585
transform 1 0 16928 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_184
timestamp 1623621585
transform 1 0 18032 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_168
timestamp 1623621585
transform 1 0 16560 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_180
timestamp 1623621585
transform 1 0 17664 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1225
timestamp 1623621585
transform 1 0 19504 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_196
timestamp 1623621585
transform 1 0 19136 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_208
timestamp 1623621585
transform 1 0 20240 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_192
timestamp 1623621585
transform 1 0 18768 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_201
timestamp 1623621585
transform 1 0 19596 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1218
timestamp 1623621585
transform 1 0 22080 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_220
timestamp 1623621585
transform 1 0 21344 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_229
timestamp 1623621585
transform 1 0 22172 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_213
timestamp 1623621585
transform 1 0 20700 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_225
timestamp 1623621585
transform 1 0 21804 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_241
timestamp 1623621585
transform 1 0 23276 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_237
timestamp 1623621585
transform 1 0 22908 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_249
timestamp 1623621585
transform 1 0 24012 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1226
timestamp 1623621585
transform 1 0 24748 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_253
timestamp 1623621585
transform 1 0 24380 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_265
timestamp 1623621585
transform 1 0 25484 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_258
timestamp 1623621585
transform 1 0 24840 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_270
timestamp 1623621585
transform 1 0 25944 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1219
timestamp 1623621585
transform 1 0 27324 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_277
timestamp 1623621585
transform 1 0 26588 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_286
timestamp 1623621585
transform 1 0 27416 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_282
timestamp 1623621585
transform 1 0 27048 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_298
timestamp 1623621585
transform 1 0 28520 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_310
timestamp 1623621585
transform 1 0 29624 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_294
timestamp 1623621585
transform 1 0 28152 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_306
timestamp 1623621585
transform 1 0 29256 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1227
timestamp 1623621585
transform 1 0 29992 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_322
timestamp 1623621585
transform 1 0 30728 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_315
timestamp 1623621585
transform 1 0 30084 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_327
timestamp 1623621585
transform 1 0 31188 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1220
timestamp 1623621585
transform 1 0 32568 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_334
timestamp 1623621585
transform 1 0 31832 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_343
timestamp 1623621585
transform 1 0 32660 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_339
timestamp 1623621585
transform 1 0 32292 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_351
timestamp 1623621585
transform 1 0 33396 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_113_363
timestamp 1623621585
transform 1 0 34500 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_355
timestamp 1623621585
transform 1 0 33764 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _415_
timestamp 1623621585
transform 1 0 34500 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_113_367
timestamp 1623621585
transform 1 0 34868 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_366
timestamp 1623621585
transform 1 0 34776 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input195
timestamp 1623621585
transform 1 0 34592 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1228
timestamp 1623621585
transform 1 0 35236 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _414_
timestamp 1623621585
transform 1 0 35144 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_113_372
timestamp 1623621585
transform 1 0 35328 0 1 63648
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_112_373
timestamp 1623621585
transform 1 0 35420 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _375_
timestamp 1623621585
transform 1 0 35880 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _456_
timestamp 1623621585
transform 1 0 36524 0 1 63648
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _462_
timestamp 1623621585
transform 1 0 36800 0 -1 63648
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _475_
timestamp 1623621585
transform 1 0 35788 0 -1 63648
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_112_384
timestamp 1623621585
transform 1 0 36432 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_395
timestamp 1623621585
transform 1 0 37444 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_381
timestamp 1623621585
transform 1 0 36156 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_392
timestamp 1623621585
transform 1 0 37168 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _435_
timestamp 1623621585
transform 1 0 37536 0 1 63648
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1623621585
transform -1 0 38824 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1623621585
transform -1 0 38824 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1221
timestamp 1623621585
transform 1 0 37812 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_112_400
timestamp 1623621585
transform 1 0 37904 0 -1 63648
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_406
timestamp 1623621585
transform 1 0 38456 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_113_403
timestamp 1623621585
transform 1 0 38180 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1623621585
transform 1 0 1104 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input390
timestamp 1623621585
transform 1 0 1380 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_114_6
timestamp 1623621585
transform 1 0 1656 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_18
timestamp 1623621585
transform 1 0 2760 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_30
timestamp 1623621585
transform 1 0 3864 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1229
timestamp 1623621585
transform 1 0 6348 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_42
timestamp 1623621585
transform 1 0 4968 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_114_54
timestamp 1623621585
transform 1 0 6072 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_114_58
timestamp 1623621585
transform 1 0 6440 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_70
timestamp 1623621585
transform 1 0 7544 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_82
timestamp 1623621585
transform 1 0 8648 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_94
timestamp 1623621585
transform 1 0 9752 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1230
timestamp 1623621585
transform 1 0 11592 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_106
timestamp 1623621585
transform 1 0 10856 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_115
timestamp 1623621585
transform 1 0 11684 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_127
timestamp 1623621585
transform 1 0 12788 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_139
timestamp 1623621585
transform 1 0 13892 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_151
timestamp 1623621585
transform 1 0 14996 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_163
timestamp 1623621585
transform 1 0 16100 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1231
timestamp 1623621585
transform 1 0 16836 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_172
timestamp 1623621585
transform 1 0 16928 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_184
timestamp 1623621585
transform 1 0 18032 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _362_
timestamp 1623621585
transform 1 0 20056 0 -1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_114_196
timestamp 1623621585
transform 1 0 19136 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_114_204
timestamp 1623621585
transform 1 0 19872 0 -1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1232
timestamp 1623621585
transform 1 0 22080 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_210
timestamp 1623621585
transform 1 0 20424 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_222
timestamp 1623621585
transform 1 0 21528 0 -1 64736
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_114_229
timestamp 1623621585
transform 1 0 22172 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_241
timestamp 1623621585
transform 1 0 23276 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_253
timestamp 1623621585
transform 1 0 24380 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_265
timestamp 1623621585
transform 1 0 25484 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1233
timestamp 1623621585
transform 1 0 27324 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_277
timestamp 1623621585
transform 1 0 26588 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_286
timestamp 1623621585
transform 1 0 27416 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_298
timestamp 1623621585
transform 1 0 28520 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_310
timestamp 1623621585
transform 1 0 29624 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _407_
timestamp 1623621585
transform 1 0 31556 0 -1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_114_322
timestamp 1623621585
transform 1 0 30728 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_114_330
timestamp 1623621585
transform 1 0 31464 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _406_
timestamp 1623621585
transform 1 0 33028 0 -1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1234
timestamp 1623621585
transform 1 0 32568 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_114_335
timestamp 1623621585
transform 1 0 31924 0 -1 64736
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_341
timestamp 1623621585
transform 1 0 32476 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_114_343
timestamp 1623621585
transform 1 0 32660 0 -1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_114_351
timestamp 1623621585
transform 1 0 33396 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _373_
timestamp 1623621585
transform 1 0 35144 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input197
timestamp 1623621585
transform 1 0 34500 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_114_366
timestamp 1623621585
transform 1 0 34776 0 -1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_114_373
timestamp 1623621585
transform 1 0 35420 0 -1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _442_
timestamp 1623621585
transform 1 0 36800 0 -1 64736
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _469_
timestamp 1623621585
transform 1 0 35788 0 -1 64736
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_114_384
timestamp 1623621585
transform 1 0 36432 0 -1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_114_395
timestamp 1623621585
transform 1 0 37444 0 -1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1623621585
transform -1 0 38824 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1235
timestamp 1623621585
transform 1 0 37812 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_114_400
timestamp 1623621585
transform 1 0 37904 0 -1 64736
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_406
timestamp 1623621585
transform 1 0 38456 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1623621585
transform 1 0 1104 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input391
timestamp 1623621585
transform 1 0 1380 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_6
timestamp 1623621585
transform 1 0 1656 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_18
timestamp 1623621585
transform 1 0 2760 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1236
timestamp 1623621585
transform 1 0 3772 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_115_26
timestamp 1623621585
transform 1 0 3496 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_30
timestamp 1623621585
transform 1 0 3864 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_42
timestamp 1623621585
transform 1 0 4968 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_54
timestamp 1623621585
transform 1 0 6072 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_66
timestamp 1623621585
transform 1 0 7176 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_78
timestamp 1623621585
transform 1 0 8280 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1237
timestamp 1623621585
transform 1 0 9016 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_87
timestamp 1623621585
transform 1 0 9108 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_99
timestamp 1623621585
transform 1 0 10212 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_111
timestamp 1623621585
transform 1 0 11316 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_123
timestamp 1623621585
transform 1 0 12420 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1238
timestamp 1623621585
transform 1 0 14260 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_115_135
timestamp 1623621585
transform 1 0 13524 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_115_144
timestamp 1623621585
transform 1 0 14352 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_156
timestamp 1623621585
transform 1 0 15456 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_168
timestamp 1623621585
transform 1 0 16560 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_180
timestamp 1623621585
transform 1 0 17664 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1239
timestamp 1623621585
transform 1 0 19504 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_115_192
timestamp 1623621585
transform 1 0 18768 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_115_201
timestamp 1623621585
transform 1 0 19596 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_213
timestamp 1623621585
transform 1 0 20700 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_225
timestamp 1623621585
transform 1 0 21804 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_237
timestamp 1623621585
transform 1 0 22908 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_249
timestamp 1623621585
transform 1 0 24012 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1240
timestamp 1623621585
transform 1 0 24748 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_258
timestamp 1623621585
transform 1 0 24840 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_270
timestamp 1623621585
transform 1 0 25944 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_282
timestamp 1623621585
transform 1 0 27048 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_294
timestamp 1623621585
transform 1 0 28152 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_306
timestamp 1623621585
transform 1 0 29256 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1241
timestamp 1623621585
transform 1 0 29992 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_315
timestamp 1623621585
transform 1 0 30084 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_327
timestamp 1623621585
transform 1 0 31188 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _534_
timestamp 1623621585
transform 1 0 32752 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_339
timestamp 1623621585
transform 1 0 32292 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_343
timestamp 1623621585
transform 1 0 32660 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_348
timestamp 1623621585
transform 1 0 33120 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1242
timestamp 1623621585
transform 1 0 35236 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input199
timestamp 1623621585
transform 1 0 34592 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_115_360
timestamp 1623621585
transform 1 0 34224 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_367
timestamp 1623621585
transform 1 0 34868 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_372
timestamp 1623621585
transform 1 0 35328 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _429_
timestamp 1623621585
transform 1 0 36524 0 1 64736
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _535_
timestamp 1623621585
transform 1 0 35788 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_376
timestamp 1623621585
transform 1 0 35696 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_115_381
timestamp 1623621585
transform 1 0 36156 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_392
timestamp 1623621585
transform 1 0 37168 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _416_
timestamp 1623621585
transform 1 0 37536 0 1 64736
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1623621585
transform -1 0 38824 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_115_403
timestamp 1623621585
transform 1 0 38180 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1623621585
transform 1 0 1104 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_3
timestamp 1623621585
transform 1 0 1380 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_15
timestamp 1623621585
transform 1 0 2484 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_27
timestamp 1623621585
transform 1 0 3588 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_39
timestamp 1623621585
transform 1 0 4692 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1243
timestamp 1623621585
transform 1 0 6348 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_116_51
timestamp 1623621585
transform 1 0 5796 0 -1 65824
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_116_58
timestamp 1623621585
transform 1 0 6440 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_70
timestamp 1623621585
transform 1 0 7544 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_82
timestamp 1623621585
transform 1 0 8648 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_94
timestamp 1623621585
transform 1 0 9752 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1244
timestamp 1623621585
transform 1 0 11592 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_106
timestamp 1623621585
transform 1 0 10856 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_115
timestamp 1623621585
transform 1 0 11684 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_127
timestamp 1623621585
transform 1 0 12788 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_139
timestamp 1623621585
transform 1 0 13892 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_151
timestamp 1623621585
transform 1 0 14996 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_163
timestamp 1623621585
transform 1 0 16100 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1245
timestamp 1623621585
transform 1 0 16836 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_172
timestamp 1623621585
transform 1 0 16928 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_184
timestamp 1623621585
transform 1 0 18032 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_196
timestamp 1623621585
transform 1 0 19136 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_208
timestamp 1623621585
transform 1 0 20240 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1246
timestamp 1623621585
transform 1 0 22080 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_220
timestamp 1623621585
transform 1 0 21344 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_229
timestamp 1623621585
transform 1 0 22172 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_241
timestamp 1623621585
transform 1 0 23276 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_253
timestamp 1623621585
transform 1 0 24380 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_265
timestamp 1623621585
transform 1 0 25484 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1247
timestamp 1623621585
transform 1 0 27324 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_277
timestamp 1623621585
transform 1 0 26588 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_286
timestamp 1623621585
transform 1 0 27416 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_298
timestamp 1623621585
transform 1 0 28520 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_310
timestamp 1623621585
transform 1 0 29624 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_322
timestamp 1623621585
transform 1 0 30728 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _372_
timestamp 1623621585
transform 1 0 33028 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1248
timestamp 1623621585
transform 1 0 32568 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_334
timestamp 1623621585
transform 1 0 31832 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_116_343
timestamp 1623621585
transform 1 0 32660 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_116_351
timestamp 1623621585
transform 1 0 33396 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input198
timestamp 1623621585
transform 1 0 35512 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input200
timestamp 1623621585
transform 1 0 34868 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_116_363
timestamp 1623621585
transform 1 0 34500 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_370
timestamp 1623621585
transform 1 0 35144 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _422_
timestamp 1623621585
transform 1 0 36800 0 -1 65824
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input196
timestamp 1623621585
transform 1 0 36156 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_116_377
timestamp 1623621585
transform 1 0 35788 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_384
timestamp 1623621585
transform 1 0 36432 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_395
timestamp 1623621585
transform 1 0 37444 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1623621585
transform -1 0 38824 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1249
timestamp 1623621585
transform 1 0 37812 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_116_400
timestamp 1623621585
transform 1 0 37904 0 -1 65824
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_406
timestamp 1623621585
transform 1 0 38456 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1623621585
transform 1 0 1104 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input392
timestamp 1623621585
transform 1 0 1380 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_117_6
timestamp 1623621585
transform 1 0 1656 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_18
timestamp 1623621585
transform 1 0 2760 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1250
timestamp 1623621585
transform 1 0 3772 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_117_26
timestamp 1623621585
transform 1 0 3496 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_117_30
timestamp 1623621585
transform 1 0 3864 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_42
timestamp 1623621585
transform 1 0 4968 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_54
timestamp 1623621585
transform 1 0 6072 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_66
timestamp 1623621585
transform 1 0 7176 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_78
timestamp 1623621585
transform 1 0 8280 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1251
timestamp 1623621585
transform 1 0 9016 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_87
timestamp 1623621585
transform 1 0 9108 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_99
timestamp 1623621585
transform 1 0 10212 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_111
timestamp 1623621585
transform 1 0 11316 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_123
timestamp 1623621585
transform 1 0 12420 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1252
timestamp 1623621585
transform 1 0 14260 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_117_135
timestamp 1623621585
transform 1 0 13524 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_144
timestamp 1623621585
transform 1 0 14352 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_156
timestamp 1623621585
transform 1 0 15456 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_168
timestamp 1623621585
transform 1 0 16560 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_180
timestamp 1623621585
transform 1 0 17664 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1253
timestamp 1623621585
transform 1 0 19504 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_117_192
timestamp 1623621585
transform 1 0 18768 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_201
timestamp 1623621585
transform 1 0 19596 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_213
timestamp 1623621585
transform 1 0 20700 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_225
timestamp 1623621585
transform 1 0 21804 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_237
timestamp 1623621585
transform 1 0 22908 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_249
timestamp 1623621585
transform 1 0 24012 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1254
timestamp 1623621585
transform 1 0 24748 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_258
timestamp 1623621585
transform 1 0 24840 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_270
timestamp 1623621585
transform 1 0 25944 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_282
timestamp 1623621585
transform 1 0 27048 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_294
timestamp 1623621585
transform 1 0 28152 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_306
timestamp 1623621585
transform 1 0 29256 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1255
timestamp 1623621585
transform 1 0 29992 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_315
timestamp 1623621585
transform 1 0 30084 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_327
timestamp 1623621585
transform 1 0 31188 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _494_
timestamp 1623621585
transform 1 0 32844 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_117_339
timestamp 1623621585
transform 1 0 32292 0 1 65824
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_117_349
timestamp 1623621585
transform 1 0 33212 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1256
timestamp 1623621585
transform 1 0 35236 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_117_361
timestamp 1623621585
transform 1 0 34316 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_117_369
timestamp 1623621585
transform 1 0 35052 0 1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_117_372
timestamp 1623621585
transform 1 0 35328 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _374_
timestamp 1623621585
transform 1 0 36524 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _495_
timestamp 1623621585
transform 1 0 35788 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_376
timestamp 1623621585
transform 1 0 35696 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_381
timestamp 1623621585
transform 1 0 36156 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_117_389
timestamp 1623621585
transform 1 0 36892 0 1 65824
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_395
timestamp 1623621585
transform 1 0 37444 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _389_
timestamp 1623621585
transform 1 0 37536 0 1 65824
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1623621585
transform -1 0 38824 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_117_403
timestamp 1623621585
transform 1 0 38180 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1623621585
transform 1 0 1104 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1623621585
transform 1 0 1104 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input393
timestamp 1623621585
transform 1 0 1380 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input395
timestamp 1623621585
transform 1 0 1380 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_6
timestamp 1623621585
transform 1 0 1656 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_18
timestamp 1623621585
transform 1 0 2760 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_6
timestamp 1623621585
transform 1 0 1656 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_18
timestamp 1623621585
transform 1 0 2760 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1264
timestamp 1623621585
transform 1 0 3772 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_30
timestamp 1623621585
transform 1 0 3864 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_119_26
timestamp 1623621585
transform 1 0 3496 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_119_30
timestamp 1623621585
transform 1 0 3864 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1257
timestamp 1623621585
transform 1 0 6348 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_42
timestamp 1623621585
transform 1 0 4968 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_118_54
timestamp 1623621585
transform 1 0 6072 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_58
timestamp 1623621585
transform 1 0 6440 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_42
timestamp 1623621585
transform 1 0 4968 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_54
timestamp 1623621585
transform 1 0 6072 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_70
timestamp 1623621585
transform 1 0 7544 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_82
timestamp 1623621585
transform 1 0 8648 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_66
timestamp 1623621585
transform 1 0 7176 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_78
timestamp 1623621585
transform 1 0 8280 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1265
timestamp 1623621585
transform 1 0 9016 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_94
timestamp 1623621585
transform 1 0 9752 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_87
timestamp 1623621585
transform 1 0 9108 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_99
timestamp 1623621585
transform 1 0 10212 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1258
timestamp 1623621585
transform 1 0 11592 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_106
timestamp 1623621585
transform 1 0 10856 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_115
timestamp 1623621585
transform 1 0 11684 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_111
timestamp 1623621585
transform 1 0 11316 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_123
timestamp 1623621585
transform 1 0 12420 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1266
timestamp 1623621585
transform 1 0 14260 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_127
timestamp 1623621585
transform 1 0 12788 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_139
timestamp 1623621585
transform 1 0 13892 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_135
timestamp 1623621585
transform 1 0 13524 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_119_144
timestamp 1623621585
transform 1 0 14352 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_151
timestamp 1623621585
transform 1 0 14996 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_163
timestamp 1623621585
transform 1 0 16100 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_119_156
timestamp 1623621585
transform 1 0 15456 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1259
timestamp 1623621585
transform 1 0 16836 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_172
timestamp 1623621585
transform 1 0 16928 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_184
timestamp 1623621585
transform 1 0 18032 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_168
timestamp 1623621585
transform 1 0 16560 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_180
timestamp 1623621585
transform 1 0 17664 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1267
timestamp 1623621585
transform 1 0 19504 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_196
timestamp 1623621585
transform 1 0 19136 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_208
timestamp 1623621585
transform 1 0 20240 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_192
timestamp 1623621585
transform 1 0 18768 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_119_201
timestamp 1623621585
transform 1 0 19596 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1260
timestamp 1623621585
transform 1 0 22080 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_220
timestamp 1623621585
transform 1 0 21344 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_229
timestamp 1623621585
transform 1 0 22172 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_213
timestamp 1623621585
transform 1 0 20700 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_225
timestamp 1623621585
transform 1 0 21804 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_241
timestamp 1623621585
transform 1 0 23276 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_237
timestamp 1623621585
transform 1 0 22908 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_249
timestamp 1623621585
transform 1 0 24012 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1268
timestamp 1623621585
transform 1 0 24748 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_253
timestamp 1623621585
transform 1 0 24380 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_265
timestamp 1623621585
transform 1 0 25484 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_258
timestamp 1623621585
transform 1 0 24840 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_270
timestamp 1623621585
transform 1 0 25944 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1261
timestamp 1623621585
transform 1 0 27324 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_277
timestamp 1623621585
transform 1 0 26588 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_286
timestamp 1623621585
transform 1 0 27416 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_282
timestamp 1623621585
transform 1 0 27048 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_298
timestamp 1623621585
transform 1 0 28520 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_310
timestamp 1623621585
transform 1 0 29624 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_294
timestamp 1623621585
transform 1 0 28152 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_306
timestamp 1623621585
transform 1 0 29256 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1269
timestamp 1623621585
transform 1 0 29992 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_322
timestamp 1623621585
transform 1 0 30728 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_315
timestamp 1623621585
transform 1 0 30084 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_327
timestamp 1623621585
transform 1 0 31188 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _454_
timestamp 1623621585
transform 1 0 32844 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1262
timestamp 1623621585
transform 1 0 32568 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_334
timestamp 1623621585
transform 1 0 31832 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_343
timestamp 1623621585
transform 1 0 32660 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_339
timestamp 1623621585
transform 1 0 32292 0 1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_119_349
timestamp 1623621585
transform 1 0 33212 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1270
timestamp 1623621585
transform 1 0 35236 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input203
timestamp 1623621585
transform 1 0 35144 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input204
timestamp 1623621585
transform 1 0 34500 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_118_355
timestamp 1623621585
transform 1 0 33764 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_118_366
timestamp 1623621585
transform 1 0 34776 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_373
timestamp 1623621585
transform 1 0 35420 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_119_361
timestamp 1623621585
transform 1 0 34316 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_119_369
timestamp 1623621585
transform 1 0 35052 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_119_372
timestamp 1623621585
transform 1 0 35328 0 1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _382_
timestamp 1623621585
transform 1 0 36524 0 1 66912
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _395_
timestamp 1623621585
transform 1 0 36800 0 -1 66912
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _402_
timestamp 1623621585
transform 1 0 35788 0 -1 66912
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _455_
timestamp 1623621585
transform 1 0 35880 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_118_384
timestamp 1623621585
transform 1 0 36432 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_395
timestamp 1623621585
transform 1 0 37444 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_381
timestamp 1623621585
transform 1 0 36156 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_392
timestamp 1623621585
transform 1 0 37168 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _376_
timestamp 1623621585
transform 1 0 37536 0 1 66912
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1623621585
transform -1 0 38824 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1623621585
transform -1 0 38824 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1263
timestamp 1623621585
transform 1 0 37812 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_118_400
timestamp 1623621585
transform 1 0 37904 0 -1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_406
timestamp 1623621585
transform 1 0 38456 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_403
timestamp 1623621585
transform 1 0 38180 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1623621585
transform 1 0 1104 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_120_3
timestamp 1623621585
transform 1 0 1380 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_15
timestamp 1623621585
transform 1 0 2484 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_27
timestamp 1623621585
transform 1 0 3588 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_39
timestamp 1623621585
transform 1 0 4692 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1271
timestamp 1623621585
transform 1 0 6348 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_120_51
timestamp 1623621585
transform 1 0 5796 0 -1 68000
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_120_58
timestamp 1623621585
transform 1 0 6440 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_70
timestamp 1623621585
transform 1 0 7544 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_82
timestamp 1623621585
transform 1 0 8648 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_94
timestamp 1623621585
transform 1 0 9752 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1272
timestamp 1623621585
transform 1 0 11592 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_106
timestamp 1623621585
transform 1 0 10856 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_120_115
timestamp 1623621585
transform 1 0 11684 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_127
timestamp 1623621585
transform 1 0 12788 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_139
timestamp 1623621585
transform 1 0 13892 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_151
timestamp 1623621585
transform 1 0 14996 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_163
timestamp 1623621585
transform 1 0 16100 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1273
timestamp 1623621585
transform 1 0 16836 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_172
timestamp 1623621585
transform 1 0 16928 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_184
timestamp 1623621585
transform 1 0 18032 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_196
timestamp 1623621585
transform 1 0 19136 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_208
timestamp 1623621585
transform 1 0 20240 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1274
timestamp 1623621585
transform 1 0 22080 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_220
timestamp 1623621585
transform 1 0 21344 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_120_229
timestamp 1623621585
transform 1 0 22172 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_241
timestamp 1623621585
transform 1 0 23276 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_253
timestamp 1623621585
transform 1 0 24380 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_265
timestamp 1623621585
transform 1 0 25484 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1275
timestamp 1623621585
transform 1 0 27324 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_277
timestamp 1623621585
transform 1 0 26588 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_120_286
timestamp 1623621585
transform 1 0 27416 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_298
timestamp 1623621585
transform 1 0 28520 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_310
timestamp 1623621585
transform 1 0 29624 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_322
timestamp 1623621585
transform 1 0 30728 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1276
timestamp 1623621585
transform 1 0 32568 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_334
timestamp 1623621585
transform 1 0 31832 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_120_343
timestamp 1623621585
transform 1 0 32660 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_355
timestamp 1623621585
transform 1 0 33764 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_367
timestamp 1623621585
transform 1 0 34868 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _354_
timestamp 1623621585
transform 1 0 36708 0 -1 68000
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _751_
timestamp 1623621585
transform 1 0 35972 0 -1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_120_383
timestamp 1623621585
transform 1 0 36340 0 -1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_120_394
timestamp 1623621585
transform 1 0 37352 0 -1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1623621585
transform -1 0 38824 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1277
timestamp 1623621585
transform 1 0 37812 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_120_398
timestamp 1623621585
transform 1 0 37720 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_120_400
timestamp 1623621585
transform 1 0 37904 0 -1 68000
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_406
timestamp 1623621585
transform 1 0 38456 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1623621585
transform 1 0 1104 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input396
timestamp 1623621585
transform 1 0 1380 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_121_6
timestamp 1623621585
transform 1 0 1656 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_18
timestamp 1623621585
transform 1 0 2760 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1278
timestamp 1623621585
transform 1 0 3772 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_121_26
timestamp 1623621585
transform 1 0 3496 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_121_30
timestamp 1623621585
transform 1 0 3864 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_42
timestamp 1623621585
transform 1 0 4968 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_54
timestamp 1623621585
transform 1 0 6072 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_66
timestamp 1623621585
transform 1 0 7176 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_78
timestamp 1623621585
transform 1 0 8280 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1279
timestamp 1623621585
transform 1 0 9016 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_87
timestamp 1623621585
transform 1 0 9108 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_99
timestamp 1623621585
transform 1 0 10212 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_111
timestamp 1623621585
transform 1 0 11316 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_123
timestamp 1623621585
transform 1 0 12420 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1280
timestamp 1623621585
transform 1 0 14260 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_121_135
timestamp 1623621585
transform 1 0 13524 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_121_144
timestamp 1623621585
transform 1 0 14352 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_156
timestamp 1623621585
transform 1 0 15456 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_168
timestamp 1623621585
transform 1 0 16560 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_180
timestamp 1623621585
transform 1 0 17664 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1281
timestamp 1623621585
transform 1 0 19504 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_121_192
timestamp 1623621585
transform 1 0 18768 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_121_201
timestamp 1623621585
transform 1 0 19596 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_213
timestamp 1623621585
transform 1 0 20700 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_225
timestamp 1623621585
transform 1 0 21804 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_237
timestamp 1623621585
transform 1 0 22908 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_249
timestamp 1623621585
transform 1 0 24012 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1282
timestamp 1623621585
transform 1 0 24748 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_258
timestamp 1623621585
transform 1 0 24840 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_270
timestamp 1623621585
transform 1 0 25944 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_282
timestamp 1623621585
transform 1 0 27048 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_294
timestamp 1623621585
transform 1 0 28152 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_306
timestamp 1623621585
transform 1 0 29256 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1283
timestamp 1623621585
transform 1 0 29992 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_1
timestamp 1623621585
transform 1 0 31740 0 1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_121_315
timestamp 1623621585
transform 1 0 30084 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_327
timestamp 1623621585
transform 1 0 31188 0 1 68000
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _330_
timestamp 1623621585
transform 1 0 31924 0 1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_121_339
timestamp 1623621585
transform 1 0 32292 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_351
timestamp 1623621585
transform 1 0 33396 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1284
timestamp 1623621585
transform 1 0 35236 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_121_363
timestamp 1623621585
transform 1 0 34500 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_121_372
timestamp 1623621585
transform 1 0 35328 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _346_
timestamp 1623621585
transform 1 0 36708 0 1 68000
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input206
timestamp 1623621585
transform 1 0 36064 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_121_383
timestamp 1623621585
transform 1 0 36340 0 1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_121_394
timestamp 1623621585
transform 1 0 37352 0 1 68000
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1623621585
transform -1 0 38824 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input201
timestamp 1623621585
transform 1 0 37904 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_121_403
timestamp 1623621585
transform 1 0 38180 0 1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1623621585
transform 1 0 1104 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input397
timestamp 1623621585
transform 1 0 1380 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_122_6
timestamp 1623621585
transform 1 0 1656 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_18
timestamp 1623621585
transform 1 0 2760 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_30
timestamp 1623621585
transform 1 0 3864 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1285
timestamp 1623621585
transform 1 0 6348 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_42
timestamp 1623621585
transform 1 0 4968 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_122_54
timestamp 1623621585
transform 1 0 6072 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_122_58
timestamp 1623621585
transform 1 0 6440 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_70
timestamp 1623621585
transform 1 0 7544 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_82
timestamp 1623621585
transform 1 0 8648 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_94
timestamp 1623621585
transform 1 0 9752 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1286
timestamp 1623621585
transform 1 0 11592 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_106
timestamp 1623621585
transform 1 0 10856 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_122_115
timestamp 1623621585
transform 1 0 11684 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_127
timestamp 1623621585
transform 1 0 12788 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_139
timestamp 1623621585
transform 1 0 13892 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_151
timestamp 1623621585
transform 1 0 14996 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_163
timestamp 1623621585
transform 1 0 16100 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1287
timestamp 1623621585
transform 1 0 16836 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_172
timestamp 1623621585
transform 1 0 16928 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_184
timestamp 1623621585
transform 1 0 18032 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_196
timestamp 1623621585
transform 1 0 19136 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_208
timestamp 1623621585
transform 1 0 20240 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1288
timestamp 1623621585
transform 1 0 22080 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_220
timestamp 1623621585
transform 1 0 21344 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_122_229
timestamp 1623621585
transform 1 0 22172 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_241
timestamp 1623621585
transform 1 0 23276 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_253
timestamp 1623621585
transform 1 0 24380 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_265
timestamp 1623621585
transform 1 0 25484 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1289
timestamp 1623621585
transform 1 0 27324 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_277
timestamp 1623621585
transform 1 0 26588 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_122_286
timestamp 1623621585
transform 1 0 27416 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_298
timestamp 1623621585
transform 1 0 28520 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_310
timestamp 1623621585
transform 1 0 29624 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_322
timestamp 1623621585
transform 1 0 30728 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1290
timestamp 1623621585
transform 1 0 32568 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_334
timestamp 1623621585
transform 1 0 31832 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_122_343
timestamp 1623621585
transform 1 0 32660 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_355
timestamp 1623621585
transform 1 0 33764 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_367
timestamp 1623621585
transform 1 0 34868 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _340_
timestamp 1623621585
transform 1 0 36708 0 -1 69088
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input207
timestamp 1623621585
transform 1 0 36064 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_122_379
timestamp 1623621585
transform 1 0 35972 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_383
timestamp 1623621585
transform 1 0 36340 0 -1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_122_394
timestamp 1623621585
transform 1 0 37352 0 -1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1623621585
transform -1 0 38824 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1291
timestamp 1623621585
transform 1 0 37812 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_122_398
timestamp 1623621585
transform 1 0 37720 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_122_400
timestamp 1623621585
transform 1 0 37904 0 -1 69088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_406
timestamp 1623621585
transform 1 0 38456 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1623621585
transform 1 0 1104 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_3
timestamp 1623621585
transform 1 0 1380 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_15
timestamp 1623621585
transform 1 0 2484 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1292
timestamp 1623621585
transform 1 0 3772 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_123_27
timestamp 1623621585
transform 1 0 3588 0 1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_123_30
timestamp 1623621585
transform 1 0 3864 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_42
timestamp 1623621585
transform 1 0 4968 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_54
timestamp 1623621585
transform 1 0 6072 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_66
timestamp 1623621585
transform 1 0 7176 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_78
timestamp 1623621585
transform 1 0 8280 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1293
timestamp 1623621585
transform 1 0 9016 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_87
timestamp 1623621585
transform 1 0 9108 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_99
timestamp 1623621585
transform 1 0 10212 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_111
timestamp 1623621585
transform 1 0 11316 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_123
timestamp 1623621585
transform 1 0 12420 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1294
timestamp 1623621585
transform 1 0 14260 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_123_135
timestamp 1623621585
transform 1 0 13524 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_123_144
timestamp 1623621585
transform 1 0 14352 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _553_
timestamp 1623621585
transform 1 0 16100 0 1 69088
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_123_156
timestamp 1623621585
transform 1 0 15456 0 1 69088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_162
timestamp 1623621585
transform 1 0 16008 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_168
timestamp 1623621585
transform 1 0 16560 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_180
timestamp 1623621585
transform 1 0 17664 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1295
timestamp 1623621585
transform 1 0 19504 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_123_192
timestamp 1623621585
transform 1 0 18768 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_123_201
timestamp 1623621585
transform 1 0 19596 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_213
timestamp 1623621585
transform 1 0 20700 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_225
timestamp 1623621585
transform 1 0 21804 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_237
timestamp 1623621585
transform 1 0 22908 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_249
timestamp 1623621585
transform 1 0 24012 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1296
timestamp 1623621585
transform 1 0 24748 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_258
timestamp 1623621585
transform 1 0 24840 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_270
timestamp 1623621585
transform 1 0 25944 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_282
timestamp 1623621585
transform 1 0 27048 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_294
timestamp 1623621585
transform 1 0 28152 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_306
timestamp 1623621585
transform 1 0 29256 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1297
timestamp 1623621585
transform 1 0 29992 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_315
timestamp 1623621585
transform 1 0 30084 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_327
timestamp 1623621585
transform 1 0 31188 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_339
timestamp 1623621585
transform 1 0 32292 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_351
timestamp 1623621585
transform 1 0 33396 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1298
timestamp 1623621585
transform 1 0 35236 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_123_363
timestamp 1623621585
transform 1 0 34500 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_123_372
timestamp 1623621585
transform 1 0 35328 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _332_
timestamp 1623621585
transform 1 0 36616 0 1 69088
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_123_384
timestamp 1623621585
transform 1 0 36432 0 1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_123_393
timestamp 1623621585
transform 1 0 37260 0 1 69088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1623621585
transform -1 0 38824 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input205
timestamp 1623621585
transform 1 0 37904 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_123_399
timestamp 1623621585
transform 1 0 37812 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_123_403
timestamp 1623621585
transform 1 0 38180 0 1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1623621585
transform 1 0 1104 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input398
timestamp 1623621585
transform 1 0 1380 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_124_6
timestamp 1623621585
transform 1 0 1656 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_18
timestamp 1623621585
transform 1 0 2760 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_30
timestamp 1623621585
transform 1 0 3864 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1299
timestamp 1623621585
transform 1 0 6348 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_42
timestamp 1623621585
transform 1 0 4968 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_124_54
timestamp 1623621585
transform 1 0 6072 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_124_58
timestamp 1623621585
transform 1 0 6440 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_70
timestamp 1623621585
transform 1 0 7544 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_82
timestamp 1623621585
transform 1 0 8648 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_94
timestamp 1623621585
transform 1 0 9752 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1300
timestamp 1623621585
transform 1 0 11592 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_106
timestamp 1623621585
transform 1 0 10856 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_124_115
timestamp 1623621585
transform 1 0 11684 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_127
timestamp 1623621585
transform 1 0 12788 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_139
timestamp 1623621585
transform 1 0 13892 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _546_
timestamp 1623621585
transform 1 0 16008 0 -1 70176
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_124_151
timestamp 1623621585
transform 1 0 14996 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_124_159
timestamp 1623621585
transform 1 0 15732 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1301
timestamp 1623621585
transform 1 0 16836 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_124_167
timestamp 1623621585
transform 1 0 16468 0 -1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_124_172
timestamp 1623621585
transform 1 0 16928 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_184
timestamp 1623621585
transform 1 0 18032 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_196
timestamp 1623621585
transform 1 0 19136 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_208
timestamp 1623621585
transform 1 0 20240 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1302
timestamp 1623621585
transform 1 0 22080 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_220
timestamp 1623621585
transform 1 0 21344 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_124_229
timestamp 1623621585
transform 1 0 22172 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_241
timestamp 1623621585
transform 1 0 23276 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_253
timestamp 1623621585
transform 1 0 24380 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_265
timestamp 1623621585
transform 1 0 25484 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1303
timestamp 1623621585
transform 1 0 27324 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_277
timestamp 1623621585
transform 1 0 26588 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_124_286
timestamp 1623621585
transform 1 0 27416 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_298
timestamp 1623621585
transform 1 0 28520 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_310
timestamp 1623621585
transform 1 0 29624 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_322
timestamp 1623621585
transform 1 0 30728 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1304
timestamp 1623621585
transform 1 0 32568 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_334
timestamp 1623621585
transform 1 0 31832 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_124_343
timestamp 1623621585
transform 1 0 32660 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_355
timestamp 1623621585
transform 1 0 33764 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_367
timestamp 1623621585
transform 1 0 34868 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input209
timestamp 1623621585
transform 1 0 37168 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input211
timestamp 1623621585
transform 1 0 36524 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_124_379
timestamp 1623621585
transform 1 0 35972 0 -1 70176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_124_388
timestamp 1623621585
transform 1 0 36800 0 -1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_124_395
timestamp 1623621585
transform 1 0 37444 0 -1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1623621585
transform -1 0 38824 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1305
timestamp 1623621585
transform 1 0 37812 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_124_400
timestamp 1623621585
transform 1 0 37904 0 -1 70176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_406
timestamp 1623621585
transform 1 0 38456 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1623621585
transform 1 0 1104 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1623621585
transform 1 0 1104 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input399
timestamp 1623621585
transform 1 0 1380 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_6
timestamp 1623621585
transform 1 0 1656 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_18
timestamp 1623621585
transform 1 0 2760 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_3
timestamp 1623621585
transform 1 0 1380 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_15
timestamp 1623621585
transform 1 0 2484 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1306
timestamp 1623621585
transform 1 0 3772 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_125_26
timestamp 1623621585
transform 1 0 3496 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_30
timestamp 1623621585
transform 1 0 3864 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_27
timestamp 1623621585
transform 1 0 3588 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_39
timestamp 1623621585
transform 1 0 4692 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1313
timestamp 1623621585
transform 1 0 6348 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_42
timestamp 1623621585
transform 1 0 4968 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_54
timestamp 1623621585
transform 1 0 6072 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_51
timestamp 1623621585
transform 1 0 5796 0 -1 71264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_126_58
timestamp 1623621585
transform 1 0 6440 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_66
timestamp 1623621585
transform 1 0 7176 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_78
timestamp 1623621585
transform 1 0 8280 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_70
timestamp 1623621585
transform 1 0 7544 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_82
timestamp 1623621585
transform 1 0 8648 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1307
timestamp 1623621585
transform 1 0 9016 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_87
timestamp 1623621585
transform 1 0 9108 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_99
timestamp 1623621585
transform 1 0 10212 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_94
timestamp 1623621585
transform 1 0 9752 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1314
timestamp 1623621585
transform 1 0 11592 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_111
timestamp 1623621585
transform 1 0 11316 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_123
timestamp 1623621585
transform 1 0 12420 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_106
timestamp 1623621585
transform 1 0 10856 0 -1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_115
timestamp 1623621585
transform 1 0 11684 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1308
timestamp 1623621585
transform 1 0 14260 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_125_135
timestamp 1623621585
transform 1 0 13524 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_125_144
timestamp 1623621585
transform 1 0 14352 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_127
timestamp 1623621585
transform 1 0 12788 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_139
timestamp 1623621585
transform 1 0 13892 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _513_
timestamp 1623621585
transform 1 0 16008 0 -1 71264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _520_
timestamp 1623621585
transform 1 0 16284 0 1 70176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _529_
timestamp 1623621585
transform 1 0 15456 0 1 70176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _559_
timestamp 1623621585
transform 1 0 15180 0 -1 71264
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_125_161
timestamp 1623621585
transform 1 0 15916 0 1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_126_151
timestamp 1623621585
transform 1 0 14996 0 -1 71264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_126_158
timestamp 1623621585
transform 1 0 15640 0 -1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _540_
timestamp 1623621585
transform 1 0 17112 0 1 70176
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1315
timestamp 1623621585
transform 1 0 16836 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_3
timestamp 1623621585
transform 1 0 16928 0 1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_125_170
timestamp 1623621585
transform 1 0 16744 0 1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_125_179
timestamp 1623621585
transform 1 0 17572 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_126_167
timestamp 1623621585
transform 1 0 16468 0 -1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_126_172
timestamp 1623621585
transform 1 0 16928 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_184
timestamp 1623621585
transform 1 0 18032 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1309
timestamp 1623621585
transform 1 0 19504 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_125_191
timestamp 1623621585
transform 1 0 18676 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_125_199
timestamp 1623621585
transform 1 0 19412 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_201
timestamp 1623621585
transform 1 0 19596 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_196
timestamp 1623621585
transform 1 0 19136 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_208
timestamp 1623621585
transform 1 0 20240 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1316
timestamp 1623621585
transform 1 0 22080 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_213
timestamp 1623621585
transform 1 0 20700 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_225
timestamp 1623621585
transform 1 0 21804 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_220
timestamp 1623621585
transform 1 0 21344 0 -1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_229
timestamp 1623621585
transform 1 0 22172 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_237
timestamp 1623621585
transform 1 0 22908 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_249
timestamp 1623621585
transform 1 0 24012 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_241
timestamp 1623621585
transform 1 0 23276 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1310
timestamp 1623621585
transform 1 0 24748 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_258
timestamp 1623621585
transform 1 0 24840 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_270
timestamp 1623621585
transform 1 0 25944 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_253
timestamp 1623621585
transform 1 0 24380 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_265
timestamp 1623621585
transform 1 0 25484 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1317
timestamp 1623621585
transform 1 0 27324 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_282
timestamp 1623621585
transform 1 0 27048 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_277
timestamp 1623621585
transform 1 0 26588 0 -1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_286
timestamp 1623621585
transform 1 0 27416 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_294
timestamp 1623621585
transform 1 0 28152 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_306
timestamp 1623621585
transform 1 0 29256 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_298
timestamp 1623621585
transform 1 0 28520 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_310
timestamp 1623621585
transform 1 0 29624 0 -1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _572_
timestamp 1623621585
transform 1 0 30636 0 -1 71264
box -38 -48 1602 592
use sky130_fd_sc_hd__a221o_4  _578_
timestamp 1623621585
transform 1 0 30912 0 1 70176
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1311
timestamp 1623621585
transform 1 0 29992 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_125_315
timestamp 1623621585
transform 1 0 30084 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_125_323
timestamp 1623621585
transform 1 0 30820 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_126_318
timestamp 1623621585
transform 1 0 30360 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1318
timestamp 1623621585
transform 1 0 32568 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_341
timestamp 1623621585
transform 1 0 32476 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_353
timestamp 1623621585
transform 1 0 33580 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_126_338
timestamp 1623621585
transform 1 0 32200 0 -1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_126_343
timestamp 1623621585
transform 1 0 32660 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1312
timestamp 1623621585
transform 1 0 35236 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_125_365
timestamp 1623621585
transform 1 0 34684 0 1 70176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_125_372
timestamp 1623621585
transform 1 0 35328 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_355
timestamp 1623621585
transform 1 0 33764 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_367
timestamp 1623621585
transform 1 0 34868 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input210
timestamp 1623621585
transform 1 0 37260 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input214
timestamp 1623621585
transform 1 0 37168 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_125_384
timestamp 1623621585
transform 1 0 36432 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_125_392
timestamp 1623621585
transform 1 0 37168 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_379
timestamp 1623621585
transform 1 0 35972 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_391
timestamp 1623621585
transform 1 0 37076 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_126_395
timestamp 1623621585
transform 1 0 37444 0 -1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1623621585
transform -1 0 38824 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1623621585
transform -1 0 38824 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1319
timestamp 1623621585
transform 1 0 37812 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input208
timestamp 1623621585
transform 1 0 37904 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_125_396
timestamp 1623621585
transform 1 0 37536 0 1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_125_403
timestamp 1623621585
transform 1 0 38180 0 1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_126_400
timestamp 1623621585
transform 1 0 37904 0 -1 71264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_406
timestamp 1623621585
transform 1 0 38456 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1623621585
transform 1 0 1104 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input400
timestamp 1623621585
transform 1 0 1380 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_127_6
timestamp 1623621585
transform 1 0 1656 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_18
timestamp 1623621585
transform 1 0 2760 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1320
timestamp 1623621585
transform 1 0 3772 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_127_26
timestamp 1623621585
transform 1 0 3496 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_127_30
timestamp 1623621585
transform 1 0 3864 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_42
timestamp 1623621585
transform 1 0 4968 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_54
timestamp 1623621585
transform 1 0 6072 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_66
timestamp 1623621585
transform 1 0 7176 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_78
timestamp 1623621585
transform 1 0 8280 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1321
timestamp 1623621585
transform 1 0 9016 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_87
timestamp 1623621585
transform 1 0 9108 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_99
timestamp 1623621585
transform 1 0 10212 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_111
timestamp 1623621585
transform 1 0 11316 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_123
timestamp 1623621585
transform 1 0 12420 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1322
timestamp 1623621585
transform 1 0 14260 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_127_135
timestamp 1623621585
transform 1 0 13524 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_127_144
timestamp 1623621585
transform 1 0 14352 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _500_
timestamp 1623621585
transform 1 0 15732 0 1 71264
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_127_156
timestamp 1623621585
transform 1 0 15456 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_127_164
timestamp 1623621585
transform 1 0 16192 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _473_
timestamp 1623621585
transform 1 0 16560 0 1 71264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _506_
timestamp 1623621585
transform 1 0 17388 0 1 71264
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_127_173
timestamp 1623621585
transform 1 0 17020 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_127_182
timestamp 1623621585
transform 1 0 17848 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1323
timestamp 1623621585
transform 1 0 19504 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_127_194
timestamp 1623621585
transform 1 0 18952 0 1 71264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_127_201
timestamp 1623621585
transform 1 0 19596 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_213
timestamp 1623621585
transform 1 0 20700 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_225
timestamp 1623621585
transform 1 0 21804 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_237
timestamp 1623621585
transform 1 0 22908 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_249
timestamp 1623621585
transform 1 0 24012 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1324
timestamp 1623621585
transform 1 0 24748 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_258
timestamp 1623621585
transform 1 0 24840 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_270
timestamp 1623621585
transform 1 0 25944 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_282
timestamp 1623621585
transform 1 0 27048 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_294
timestamp 1623621585
transform 1 0 28152 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_306
timestamp 1623621585
transform 1 0 29256 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _566_
timestamp 1623621585
transform 1 0 31004 0 1 71264
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1325
timestamp 1623621585
transform 1 0 29992 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_127_315
timestamp 1623621585
transform 1 0 30084 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_127_323
timestamp 1623621585
transform 1 0 30820 0 1 71264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_127_342
timestamp 1623621585
transform 1 0 32568 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_354
timestamp 1623621585
transform 1 0 33672 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1326
timestamp 1623621585
transform 1 0 35236 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_127_366
timestamp 1623621585
transform 1 0 34776 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_370
timestamp 1623621585
transform 1 0 35144 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_127_372
timestamp 1623621585
transform 1 0 35328 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _331_
timestamp 1623621585
transform 1 0 35696 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input215
timestamp 1623621585
transform 1 0 37260 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_127_380
timestamp 1623621585
transform 1 0 36064 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_127_392
timestamp 1623621585
transform 1 0 37168 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1623621585
transform -1 0 38824 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input212
timestamp 1623621585
transform 1 0 37904 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_127_396
timestamp 1623621585
transform 1 0 37536 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_127_403
timestamp 1623621585
transform 1 0 38180 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1623621585
transform 1 0 1104 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input401
timestamp 1623621585
transform 1 0 1380 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_128_6
timestamp 1623621585
transform 1 0 1656 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_18
timestamp 1623621585
transform 1 0 2760 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_30
timestamp 1623621585
transform 1 0 3864 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1327
timestamp 1623621585
transform 1 0 6348 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_42
timestamp 1623621585
transform 1 0 4968 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_128_54
timestamp 1623621585
transform 1 0 6072 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_128_58
timestamp 1623621585
transform 1 0 6440 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_70
timestamp 1623621585
transform 1 0 7544 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_82
timestamp 1623621585
transform 1 0 8648 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_94
timestamp 1623621585
transform 1 0 9752 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1328
timestamp 1623621585
transform 1 0 11592 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_106
timestamp 1623621585
transform 1 0 10856 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_128_115
timestamp 1623621585
transform 1 0 11684 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_127
timestamp 1623621585
transform 1 0 12788 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_139
timestamp 1623621585
transform 1 0 13892 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _480_
timestamp 1623621585
transform 1 0 16008 0 -1 72352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_128_151
timestamp 1623621585
transform 1 0 14996 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_128_159
timestamp 1623621585
transform 1 0 15732 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _449_
timestamp 1623621585
transform 1 0 17296 0 -1 72352
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1329
timestamp 1623621585
transform 1 0 16836 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE3_0
timestamp 1623621585
transform 1 0 17112 0 -1 72352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_128_167
timestamp 1623621585
transform 1 0 16468 0 -1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_128_172
timestamp 1623621585
transform 1 0 16928 0 -1 72352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_128_181
timestamp 1623621585
transform 1 0 17756 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_193
timestamp 1623621585
transform 1 0 18860 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_205
timestamp 1623621585
transform 1 0 19964 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1330
timestamp 1623621585
transform 1 0 22080 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_217
timestamp 1623621585
transform 1 0 21068 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_128_225
timestamp 1623621585
transform 1 0 21804 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_128_229
timestamp 1623621585
transform 1 0 22172 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_241
timestamp 1623621585
transform 1 0 23276 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_253
timestamp 1623621585
transform 1 0 24380 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_265
timestamp 1623621585
transform 1 0 25484 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1331
timestamp 1623621585
transform 1 0 27324 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_277
timestamp 1623621585
transform 1 0 26588 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_128_286
timestamp 1623621585
transform 1 0 27416 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_298
timestamp 1623621585
transform 1 0 28520 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_310
timestamp 1623621585
transform 1 0 29624 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_322
timestamp 1623621585
transform 1 0 30728 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1332
timestamp 1623621585
transform 1 0 32568 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_334
timestamp 1623621585
transform 1 0 31832 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_128_343
timestamp 1623621585
transform 1 0 32660 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_355
timestamp 1623621585
transform 1 0 33764 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_367
timestamp 1623621585
transform 1 0 34868 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input234
timestamp 1623621585
transform 1 0 37168 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_128_379
timestamp 1623621585
transform 1 0 35972 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_391
timestamp 1623621585
transform 1 0 37076 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_128_395
timestamp 1623621585
transform 1 0 37444 0 -1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1623621585
transform -1 0 38824 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1333
timestamp 1623621585
transform 1 0 37812 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_128_400
timestamp 1623621585
transform 1 0 37904 0 -1 72352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_406
timestamp 1623621585
transform 1 0 38456 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1623621585
transform 1 0 1104 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_129_3
timestamp 1623621585
transform 1 0 1380 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_15
timestamp 1623621585
transform 1 0 2484 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1334
timestamp 1623621585
transform 1 0 3772 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_129_27
timestamp 1623621585
transform 1 0 3588 0 1 72352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_129_30
timestamp 1623621585
transform 1 0 3864 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_42
timestamp 1623621585
transform 1 0 4968 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_54
timestamp 1623621585
transform 1 0 6072 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_66
timestamp 1623621585
transform 1 0 7176 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_78
timestamp 1623621585
transform 1 0 8280 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1335
timestamp 1623621585
transform 1 0 9016 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_87
timestamp 1623621585
transform 1 0 9108 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_99
timestamp 1623621585
transform 1 0 10212 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_111
timestamp 1623621585
transform 1 0 11316 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_123
timestamp 1623621585
transform 1 0 12420 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1336
timestamp 1623621585
transform 1 0 14260 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_129_135
timestamp 1623621585
transform 1 0 13524 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_129_144
timestamp 1623621585
transform 1 0 14352 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _489_
timestamp 1623621585
transform 1 0 15732 0 1 72352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_129_156
timestamp 1623621585
transform 1 0 15456 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_129_164
timestamp 1623621585
transform 1 0 16192 0 1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _460_
timestamp 1623621585
transform 1 0 16560 0 1 72352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _466_
timestamp 1623621585
transform 1 0 17388 0 1 72352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_129_173
timestamp 1623621585
transform 1 0 17020 0 1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_129_182
timestamp 1623621585
transform 1 0 17848 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _528_
timestamp 1623621585
transform 1 0 19964 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1337
timestamp 1623621585
transform 1 0 19504 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_129_194
timestamp 1623621585
transform 1 0 18952 0 1 72352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_129_201
timestamp 1623621585
transform 1 0 19596 0 1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_129_208
timestamp 1623621585
transform 1 0 20240 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_220
timestamp 1623621585
transform 1 0 21344 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_232
timestamp 1623621585
transform 1 0 22448 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_244
timestamp 1623621585
transform 1 0 23552 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1338
timestamp 1623621585
transform 1 0 24748 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_129_256
timestamp 1623621585
transform 1 0 24656 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_258
timestamp 1623621585
transform 1 0 24840 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_270
timestamp 1623621585
transform 1 0 25944 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_282
timestamp 1623621585
transform 1 0 27048 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_294
timestamp 1623621585
transform 1 0 28152 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_306
timestamp 1623621585
transform 1 0 29256 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1339
timestamp 1623621585
transform 1 0 29992 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_315
timestamp 1623621585
transform 1 0 30084 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_327
timestamp 1623621585
transform 1 0 31188 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_339
timestamp 1623621585
transform 1 0 32292 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_351
timestamp 1623621585
transform 1 0 33396 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1340
timestamp 1623621585
transform 1 0 35236 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_129_363
timestamp 1623621585
transform 1 0 34500 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_129_372
timestamp 1623621585
transform 1 0 35328 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input245
timestamp 1623621585
transform 1 0 37260 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_129_384
timestamp 1623621585
transform 1 0 36432 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_129_392
timestamp 1623621585
transform 1 0 37168 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1623621585
transform -1 0 38824 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input223
timestamp 1623621585
transform 1 0 37904 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_129_396
timestamp 1623621585
transform 1 0 37536 0 1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_129_403
timestamp 1623621585
transform 1 0 38180 0 1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1623621585
transform 1 0 1104 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input402
timestamp 1623621585
transform 1 0 1380 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_130_6
timestamp 1623621585
transform 1 0 1656 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_18
timestamp 1623621585
transform 1 0 2760 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_30
timestamp 1623621585
transform 1 0 3864 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1341
timestamp 1623621585
transform 1 0 6348 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_42
timestamp 1623621585
transform 1 0 4968 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_130_54
timestamp 1623621585
transform 1 0 6072 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_130_58
timestamp 1623621585
transform 1 0 6440 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_70
timestamp 1623621585
transform 1 0 7544 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_82
timestamp 1623621585
transform 1 0 8648 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_94
timestamp 1623621585
transform 1 0 9752 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1342
timestamp 1623621585
transform 1 0 11592 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_106
timestamp 1623621585
transform 1 0 10856 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_130_115
timestamp 1623621585
transform 1 0 11684 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_127
timestamp 1623621585
transform 1 0 12788 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_139
timestamp 1623621585
transform 1 0 13892 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_151
timestamp 1623621585
transform 1 0 14996 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_163
timestamp 1623621585
transform 1 0 16100 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1343
timestamp 1623621585
transform 1 0 16836 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_172
timestamp 1623621585
transform 1 0 16928 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_184
timestamp 1623621585
transform 1 0 18032 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_196
timestamp 1623621585
transform 1 0 19136 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_208
timestamp 1623621585
transform 1 0 20240 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1344
timestamp 1623621585
transform 1 0 22080 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_220
timestamp 1623621585
transform 1 0 21344 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_130_229
timestamp 1623621585
transform 1 0 22172 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_241
timestamp 1623621585
transform 1 0 23276 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_253
timestamp 1623621585
transform 1 0 24380 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_265
timestamp 1623621585
transform 1 0 25484 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1345
timestamp 1623621585
transform 1 0 27324 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_277
timestamp 1623621585
transform 1 0 26588 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_130_286
timestamp 1623621585
transform 1 0 27416 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_298
timestamp 1623621585
transform 1 0 28520 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_310
timestamp 1623621585
transform 1 0 29624 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_322
timestamp 1623621585
transform 1 0 30728 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1346
timestamp 1623621585
transform 1 0 32568 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_334
timestamp 1623621585
transform 1 0 31832 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_130_343
timestamp 1623621585
transform 1 0 32660 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_355
timestamp 1623621585
transform 1 0 33764 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_367
timestamp 1623621585
transform 1 0 34868 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_379
timestamp 1623621585
transform 1 0 35972 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_391
timestamp 1623621585
transform 1 0 37076 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1623621585
transform -1 0 38824 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1347
timestamp 1623621585
transform 1 0 37812 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_130_400
timestamp 1623621585
transform 1 0 37904 0 -1 73440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_406
timestamp 1623621585
transform 1 0 38456 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1623621585
transform 1 0 1104 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input403
timestamp 1623621585
transform 1 0 1380 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_131_6
timestamp 1623621585
transform 1 0 1656 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_131_18
timestamp 1623621585
transform 1 0 2760 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1348
timestamp 1623621585
transform 1 0 3772 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_131_26
timestamp 1623621585
transform 1 0 3496 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_131_30
timestamp 1623621585
transform 1 0 3864 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_42
timestamp 1623621585
transform 1 0 4968 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_54
timestamp 1623621585
transform 1 0 6072 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_66
timestamp 1623621585
transform 1 0 7176 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_131_78
timestamp 1623621585
transform 1 0 8280 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1349
timestamp 1623621585
transform 1 0 9016 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_87
timestamp 1623621585
transform 1 0 9108 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_99
timestamp 1623621585
transform 1 0 10212 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_111
timestamp 1623621585
transform 1 0 11316 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_123
timestamp 1623621585
transform 1 0 12420 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1350
timestamp 1623621585
transform 1 0 14260 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_131_135
timestamp 1623621585
transform 1 0 13524 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_131_144
timestamp 1623621585
transform 1 0 14352 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_156
timestamp 1623621585
transform 1 0 15456 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_168
timestamp 1623621585
transform 1 0 16560 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_180
timestamp 1623621585
transform 1 0 17664 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _448_
timestamp 1623621585
transform 1 0 20056 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1351
timestamp 1623621585
transform 1 0 19504 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_131_192
timestamp 1623621585
transform 1 0 18768 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_131_201
timestamp 1623621585
transform 1 0 19596 0 1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_205
timestamp 1623621585
transform 1 0 19964 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _488_
timestamp 1623621585
transform 1 0 20700 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_131_209
timestamp 1623621585
transform 1 0 20332 0 1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_131_216
timestamp 1623621585
transform 1 0 20976 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_228
timestamp 1623621585
transform 1 0 22080 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_240
timestamp 1623621585
transform 1 0 23184 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1352
timestamp 1623621585
transform 1 0 24748 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_131_252
timestamp 1623621585
transform 1 0 24288 0 1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_256
timestamp 1623621585
transform 1 0 24656 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_258
timestamp 1623621585
transform 1 0 24840 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_270
timestamp 1623621585
transform 1 0 25944 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_282
timestamp 1623621585
transform 1 0 27048 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_294
timestamp 1623621585
transform 1 0 28152 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_131_306
timestamp 1623621585
transform 1 0 29256 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1353
timestamp 1623621585
transform 1 0 29992 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_315
timestamp 1623621585
transform 1 0 30084 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_327
timestamp 1623621585
transform 1 0 31188 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_339
timestamp 1623621585
transform 1 0 32292 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_351
timestamp 1623621585
transform 1 0 33396 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1354
timestamp 1623621585
transform 1 0 35236 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_131_363
timestamp 1623621585
transform 1 0 34500 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_131_372
timestamp 1623621585
transform 1 0 35328 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input249
timestamp 1623621585
transform 1 0 37260 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_131_384
timestamp 1623621585
transform 1 0 36432 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_131_392
timestamp 1623621585
transform 1 0 37168 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1623621585
transform -1 0 38824 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input248
timestamp 1623621585
transform 1 0 37904 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_131_396
timestamp 1623621585
transform 1 0 37536 0 1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_131_403
timestamp 1623621585
transform 1 0 38180 0 1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1623621585
transform 1 0 1104 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1623621585
transform 1 0 1104 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input404
timestamp 1623621585
transform 1 0 1380 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_132_3
timestamp 1623621585
transform 1 0 1380 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_15
timestamp 1623621585
transform 1 0 2484 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_6
timestamp 1623621585
transform 1 0 1656 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_18
timestamp 1623621585
transform 1 0 2760 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1362
timestamp 1623621585
transform 1 0 3772 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_27
timestamp 1623621585
transform 1 0 3588 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_39
timestamp 1623621585
transform 1 0 4692 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_133_26
timestamp 1623621585
transform 1 0 3496 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_133_30
timestamp 1623621585
transform 1 0 3864 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1355
timestamp 1623621585
transform 1 0 6348 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_132_51
timestamp 1623621585
transform 1 0 5796 0 -1 74528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_132_58
timestamp 1623621585
transform 1 0 6440 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_42
timestamp 1623621585
transform 1 0 4968 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_54
timestamp 1623621585
transform 1 0 6072 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_70
timestamp 1623621585
transform 1 0 7544 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_82
timestamp 1623621585
transform 1 0 8648 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_66
timestamp 1623621585
transform 1 0 7176 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_78
timestamp 1623621585
transform 1 0 8280 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1363
timestamp 1623621585
transform 1 0 9016 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_94
timestamp 1623621585
transform 1 0 9752 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_87
timestamp 1623621585
transform 1 0 9108 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_99
timestamp 1623621585
transform 1 0 10212 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1356
timestamp 1623621585
transform 1 0 11592 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_106
timestamp 1623621585
transform 1 0 10856 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_132_115
timestamp 1623621585
transform 1 0 11684 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_111
timestamp 1623621585
transform 1 0 11316 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_123
timestamp 1623621585
transform 1 0 12420 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1364
timestamp 1623621585
transform 1 0 14260 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_127
timestamp 1623621585
transform 1 0 12788 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_139
timestamp 1623621585
transform 1 0 13892 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_135
timestamp 1623621585
transform 1 0 13524 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_133_144
timestamp 1623621585
transform 1 0 14352 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_151
timestamp 1623621585
transform 1 0 14996 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_163
timestamp 1623621585
transform 1 0 16100 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_133_156
timestamp 1623621585
transform 1 0 15456 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1357
timestamp 1623621585
transform 1 0 16836 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_172
timestamp 1623621585
transform 1 0 16928 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_184
timestamp 1623621585
transform 1 0 18032 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_168
timestamp 1623621585
transform 1 0 16560 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_180
timestamp 1623621585
transform 1 0 17664 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _352_
timestamp 1623621585
transform 1 0 19964 0 1 74528
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1365
timestamp 1623621585
transform 1 0 19504 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_196
timestamp 1623621585
transform 1 0 19136 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_208
timestamp 1623621585
transform 1 0 20240 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_192
timestamp 1623621585
transform 1 0 18768 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_133_201
timestamp 1623621585
transform 1 0 19596 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1358
timestamp 1623621585
transform 1 0 22080 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_220
timestamp 1623621585
transform 1 0 21344 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_132_229
timestamp 1623621585
transform 1 0 22172 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_210
timestamp 1623621585
transform 1 0 20424 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_222
timestamp 1623621585
transform 1 0 21528 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_241
timestamp 1623621585
transform 1 0 23276 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_234
timestamp 1623621585
transform 1 0 22632 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_246
timestamp 1623621585
transform 1 0 23736 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1366
timestamp 1623621585
transform 1 0 24748 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_253
timestamp 1623621585
transform 1 0 24380 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_265
timestamp 1623621585
transform 1 0 25484 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_133_254
timestamp 1623621585
transform 1 0 24472 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_133_258
timestamp 1623621585
transform 1 0 24840 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_270
timestamp 1623621585
transform 1 0 25944 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1359
timestamp 1623621585
transform 1 0 27324 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_277
timestamp 1623621585
transform 1 0 26588 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_132_286
timestamp 1623621585
transform 1 0 27416 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_282
timestamp 1623621585
transform 1 0 27048 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_298
timestamp 1623621585
transform 1 0 28520 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_310
timestamp 1623621585
transform 1 0 29624 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_294
timestamp 1623621585
transform 1 0 28152 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_306
timestamp 1623621585
transform 1 0 29256 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1367
timestamp 1623621585
transform 1 0 29992 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_322
timestamp 1623621585
transform 1 0 30728 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_315
timestamp 1623621585
transform 1 0 30084 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_327
timestamp 1623621585
transform 1 0 31188 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1360
timestamp 1623621585
transform 1 0 32568 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_334
timestamp 1623621585
transform 1 0 31832 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_132_343
timestamp 1623621585
transform 1 0 32660 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_339
timestamp 1623621585
transform 1 0 32292 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_351
timestamp 1623621585
transform 1 0 33396 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1368
timestamp 1623621585
transform 1 0 35236 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_355
timestamp 1623621585
transform 1 0 33764 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_367
timestamp 1623621585
transform 1 0 34868 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_363
timestamp 1623621585
transform 1 0 34500 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_133_372
timestamp 1623621585
transform 1 0 35328 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input251
timestamp 1623621585
transform 1 0 37168 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input252
timestamp 1623621585
transform 1 0 37260 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_132_379
timestamp 1623621585
transform 1 0 35972 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_391
timestamp 1623621585
transform 1 0 37076 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_132_395
timestamp 1623621585
transform 1 0 37444 0 -1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_133_384
timestamp 1623621585
transform 1 0 36432 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_133_392
timestamp 1623621585
transform 1 0 37168 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1623621585
transform -1 0 38824 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1623621585
transform -1 0 38824 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1361
timestamp 1623621585
transform 1 0 37812 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input250
timestamp 1623621585
transform 1 0 37904 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_132_400
timestamp 1623621585
transform 1 0 37904 0 -1 74528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_406
timestamp 1623621585
transform 1 0 38456 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_133_396
timestamp 1623621585
transform 1 0 37536 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_133_403
timestamp 1623621585
transform 1 0 38180 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1623621585
transform 1 0 1104 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input406
timestamp 1623621585
transform 1 0 1380 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_134_6
timestamp 1623621585
transform 1 0 1656 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_18
timestamp 1623621585
transform 1 0 2760 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_30
timestamp 1623621585
transform 1 0 3864 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1369
timestamp 1623621585
transform 1 0 6348 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_42
timestamp 1623621585
transform 1 0 4968 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_134_54
timestamp 1623621585
transform 1 0 6072 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_134_58
timestamp 1623621585
transform 1 0 6440 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_70
timestamp 1623621585
transform 1 0 7544 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_82
timestamp 1623621585
transform 1 0 8648 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_94
timestamp 1623621585
transform 1 0 9752 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1370
timestamp 1623621585
transform 1 0 11592 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_106
timestamp 1623621585
transform 1 0 10856 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_134_115
timestamp 1623621585
transform 1 0 11684 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_127
timestamp 1623621585
transform 1 0 12788 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_139
timestamp 1623621585
transform 1 0 13892 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_151
timestamp 1623621585
transform 1 0 14996 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_163
timestamp 1623621585
transform 1 0 16100 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1371
timestamp 1623621585
transform 1 0 16836 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_172
timestamp 1623621585
transform 1 0 16928 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_184
timestamp 1623621585
transform 1 0 18032 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _325_
timestamp 1623621585
transform 1 0 19964 0 -1 75616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_134_196
timestamp 1623621585
transform 1 0 19136 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_134_204
timestamp 1623621585
transform 1 0 19872 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _336_
timestamp 1623621585
transform 1 0 20792 0 -1 75616
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1372
timestamp 1623621585
transform 1 0 22080 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_134_210
timestamp 1623621585
transform 1 0 20424 0 -1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_134_219
timestamp 1623621585
transform 1 0 21252 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_134_227
timestamp 1623621585
transform 1 0 21988 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_229
timestamp 1623621585
transform 1 0 22172 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_241
timestamp 1623621585
transform 1 0 23276 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_253
timestamp 1623621585
transform 1 0 24380 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_265
timestamp 1623621585
transform 1 0 25484 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1373
timestamp 1623621585
transform 1 0 27324 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_277
timestamp 1623621585
transform 1 0 26588 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_134_286
timestamp 1623621585
transform 1 0 27416 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__nor4_2  _584_
timestamp 1623621585
transform 1 0 29348 0 -1 75616
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_134_298
timestamp 1623621585
transform 1 0 28520 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_134_306
timestamp 1623621585
transform 1 0 29256 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_317
timestamp 1623621585
transform 1 0 30268 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_329
timestamp 1623621585
transform 1 0 31372 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1374
timestamp 1623621585
transform 1 0 32568 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_134_341
timestamp 1623621585
transform 1 0 32476 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_343
timestamp 1623621585
transform 1 0 32660 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_355
timestamp 1623621585
transform 1 0 33764 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_367
timestamp 1623621585
transform 1 0 34868 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input253
timestamp 1623621585
transform 1 0 37168 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_134_379
timestamp 1623621585
transform 1 0 35972 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_391
timestamp 1623621585
transform 1 0 37076 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_134_395
timestamp 1623621585
transform 1 0 37444 0 -1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1623621585
transform -1 0 38824 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1375
timestamp 1623621585
transform 1 0 37812 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_134_400
timestamp 1623621585
transform 1 0 37904 0 -1 75616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_406
timestamp 1623621585
transform 1 0 38456 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1623621585
transform 1 0 1104 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_3
timestamp 1623621585
transform 1 0 1380 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_15
timestamp 1623621585
transform 1 0 2484 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1376
timestamp 1623621585
transform 1 0 3772 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_135_27
timestamp 1623621585
transform 1 0 3588 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_135_30
timestamp 1623621585
transform 1 0 3864 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_42
timestamp 1623621585
transform 1 0 4968 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_54
timestamp 1623621585
transform 1 0 6072 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_66
timestamp 1623621585
transform 1 0 7176 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_78
timestamp 1623621585
transform 1 0 8280 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1377
timestamp 1623621585
transform 1 0 9016 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_87
timestamp 1623621585
transform 1 0 9108 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_99
timestamp 1623621585
transform 1 0 10212 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_111
timestamp 1623621585
transform 1 0 11316 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_123
timestamp 1623621585
transform 1 0 12420 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1378
timestamp 1623621585
transform 1 0 14260 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_135_135
timestamp 1623621585
transform 1 0 13524 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_135_144
timestamp 1623621585
transform 1 0 14352 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_156
timestamp 1623621585
transform 1 0 15456 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_168
timestamp 1623621585
transform 1 0 16560 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_180
timestamp 1623621585
transform 1 0 17664 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _344_
timestamp 1623621585
transform 1 0 19964 0 1 75616
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1379
timestamp 1623621585
transform 1 0 19504 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_135_192
timestamp 1623621585
transform 1 0 18768 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_135_201
timestamp 1623621585
transform 1 0 19596 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_135_210
timestamp 1623621585
transform 1 0 20424 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_222
timestamp 1623621585
transform 1 0 21528 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_234
timestamp 1623621585
transform 1 0 22632 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_246
timestamp 1623621585
transform 1 0 23736 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1380
timestamp 1623621585
transform 1 0 24748 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_135_254
timestamp 1623621585
transform 1 0 24472 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_258
timestamp 1623621585
transform 1 0 24840 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_270
timestamp 1623621585
transform 1 0 25944 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_282
timestamp 1623621585
transform 1 0 27048 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_294
timestamp 1623621585
transform 1 0 28152 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_306
timestamp 1623621585
transform 1 0 29256 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1381
timestamp 1623621585
transform 1 0 29992 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_315
timestamp 1623621585
transform 1 0 30084 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_327
timestamp 1623621585
transform 1 0 31188 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_339
timestamp 1623621585
transform 1 0 32292 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_351
timestamp 1623621585
transform 1 0 33396 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1382
timestamp 1623621585
transform 1 0 35236 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_135_363
timestamp 1623621585
transform 1 0 34500 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_135_372
timestamp 1623621585
transform 1 0 35328 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input254
timestamp 1623621585
transform 1 0 37260 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_135_384
timestamp 1623621585
transform 1 0 36432 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_135_392
timestamp 1623621585
transform 1 0 37168 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1623621585
transform -1 0 38824 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input225
timestamp 1623621585
transform 1 0 37904 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_135_396
timestamp 1623621585
transform 1 0 37536 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_135_403
timestamp 1623621585
transform 1 0 38180 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1623621585
transform 1 0 1104 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input407
timestamp 1623621585
transform 1 0 1380 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_136_6
timestamp 1623621585
transform 1 0 1656 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_18
timestamp 1623621585
transform 1 0 2760 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_30
timestamp 1623621585
transform 1 0 3864 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1383
timestamp 1623621585
transform 1 0 6348 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_42
timestamp 1623621585
transform 1 0 4968 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_136_54
timestamp 1623621585
transform 1 0 6072 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_136_58
timestamp 1623621585
transform 1 0 6440 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_70
timestamp 1623621585
transform 1 0 7544 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_82
timestamp 1623621585
transform 1 0 8648 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_94
timestamp 1623621585
transform 1 0 9752 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1384
timestamp 1623621585
transform 1 0 11592 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_136_106
timestamp 1623621585
transform 1 0 10856 0 -1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_136_115
timestamp 1623621585
transform 1 0 11684 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_127
timestamp 1623621585
transform 1 0 12788 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_139
timestamp 1623621585
transform 1 0 13892 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_151
timestamp 1623621585
transform 1 0 14996 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_163
timestamp 1623621585
transform 1 0 16100 0 -1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1385
timestamp 1623621585
transform 1 0 16836 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_172
timestamp 1623621585
transform 1 0 16928 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_184
timestamp 1623621585
transform 1 0 18032 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_196
timestamp 1623621585
transform 1 0 19136 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_208
timestamp 1623621585
transform 1 0 20240 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1386
timestamp 1623621585
transform 1 0 22080 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_136_220
timestamp 1623621585
transform 1 0 21344 0 -1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_136_229
timestamp 1623621585
transform 1 0 22172 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _324_
timestamp 1623621585
transform 1 0 23368 0 -1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_241
timestamp 1623621585
transform 1 0 23276 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_246
timestamp 1623621585
transform 1 0 23736 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_258
timestamp 1623621585
transform 1 0 24840 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_270
timestamp 1623621585
transform 1 0 25944 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1387
timestamp 1623621585
transform 1 0 27324 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_136_282
timestamp 1623621585
transform 1 0 27048 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_136_286
timestamp 1623621585
transform 1 0 27416 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_298
timestamp 1623621585
transform 1 0 28520 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_310
timestamp 1623621585
transform 1 0 29624 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _740_
timestamp 1623621585
transform 1 0 30912 0 -1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_136_322
timestamp 1623621585
transform 1 0 30728 0 -1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_136_328
timestamp 1623621585
transform 1 0 31280 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1388
timestamp 1623621585
transform 1 0 32568 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_136_340
timestamp 1623621585
transform 1 0 32384 0 -1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_136_343
timestamp 1623621585
transform 1 0 32660 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_355
timestamp 1623621585
transform 1 0 33764 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_367
timestamp 1623621585
transform 1 0 34868 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_379
timestamp 1623621585
transform 1 0 35972 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_391
timestamp 1623621585
transform 1 0 37076 0 -1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1623621585
transform -1 0 38824 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1389
timestamp 1623621585
transform 1 0 37812 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_136_400
timestamp 1623621585
transform 1 0 37904 0 -1 76704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_406
timestamp 1623621585
transform 1 0 38456 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1623621585
transform 1 0 1104 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input415
timestamp 1623621585
transform 1 0 1380 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_137_6
timestamp 1623621585
transform 1 0 1656 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_18
timestamp 1623621585
transform 1 0 2760 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1390
timestamp 1623621585
transform 1 0 3772 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_137_26
timestamp 1623621585
transform 1 0 3496 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_137_30
timestamp 1623621585
transform 1 0 3864 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_42
timestamp 1623621585
transform 1 0 4968 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_54
timestamp 1623621585
transform 1 0 6072 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_66
timestamp 1623621585
transform 1 0 7176 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_78
timestamp 1623621585
transform 1 0 8280 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1391
timestamp 1623621585
transform 1 0 9016 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_87
timestamp 1623621585
transform 1 0 9108 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_99
timestamp 1623621585
transform 1 0 10212 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_111
timestamp 1623621585
transform 1 0 11316 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_123
timestamp 1623621585
transform 1 0 12420 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1392
timestamp 1623621585
transform 1 0 14260 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_137_135
timestamp 1623621585
transform 1 0 13524 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_137_144
timestamp 1623621585
transform 1 0 14352 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_156
timestamp 1623621585
transform 1 0 15456 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_168
timestamp 1623621585
transform 1 0 16560 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_180
timestamp 1623621585
transform 1 0 17664 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1393
timestamp 1623621585
transform 1 0 19504 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_137_192
timestamp 1623621585
transform 1 0 18768 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_137_201
timestamp 1623621585
transform 1 0 19596 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_213
timestamp 1623621585
transform 1 0 20700 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_225
timestamp 1623621585
transform 1 0 21804 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_237
timestamp 1623621585
transform 1 0 22908 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_249
timestamp 1623621585
transform 1 0 24012 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1394
timestamp 1623621585
transform 1 0 24748 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_258
timestamp 1623621585
transform 1 0 24840 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_270
timestamp 1623621585
transform 1 0 25944 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_282
timestamp 1623621585
transform 1 0 27048 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_294
timestamp 1623621585
transform 1 0 28152 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_306
timestamp 1623621585
transform 1 0 29256 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1395
timestamp 1623621585
transform 1 0 29992 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_315
timestamp 1623621585
transform 1 0 30084 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_327
timestamp 1623621585
transform 1 0 31188 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_339
timestamp 1623621585
transform 1 0 32292 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_351
timestamp 1623621585
transform 1 0 33396 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1396
timestamp 1623621585
transform 1 0 35236 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_137_363
timestamp 1623621585
transform 1 0 34500 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_137_372
timestamp 1623621585
transform 1 0 35328 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input226
timestamp 1623621585
transform 1 0 37260 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_137_384
timestamp 1623621585
transform 1 0 36432 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_137_392
timestamp 1623621585
transform 1 0 37168 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1623621585
transform -1 0 38824 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input224
timestamp 1623621585
transform 1 0 37904 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_396
timestamp 1623621585
transform 1 0 37536 0 1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_403
timestamp 1623621585
transform 1 0 38180 0 1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1623621585
transform 1 0 1104 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_278
timestamp 1623621585
transform 1 0 1104 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input426
timestamp 1623621585
transform 1 0 1380 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_3
timestamp 1623621585
transform 1 0 1380 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_15
timestamp 1623621585
transform 1 0 2484 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_6
timestamp 1623621585
transform 1 0 1656 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_18
timestamp 1623621585
transform 1 0 2760 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1404
timestamp 1623621585
transform 1 0 3772 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_27
timestamp 1623621585
transform 1 0 3588 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_39
timestamp 1623621585
transform 1 0 4692 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_139_26
timestamp 1623621585
transform 1 0 3496 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_139_30
timestamp 1623621585
transform 1 0 3864 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1397
timestamp 1623621585
transform 1 0 6348 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_138_51
timestamp 1623621585
transform 1 0 5796 0 -1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_138_58
timestamp 1623621585
transform 1 0 6440 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_42
timestamp 1623621585
transform 1 0 4968 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_54
timestamp 1623621585
transform 1 0 6072 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_70
timestamp 1623621585
transform 1 0 7544 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_82
timestamp 1623621585
transform 1 0 8648 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_66
timestamp 1623621585
transform 1 0 7176 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_78
timestamp 1623621585
transform 1 0 8280 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1405
timestamp 1623621585
transform 1 0 9016 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_94
timestamp 1623621585
transform 1 0 9752 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_87
timestamp 1623621585
transform 1 0 9108 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_99
timestamp 1623621585
transform 1 0 10212 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1398
timestamp 1623621585
transform 1 0 11592 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_106
timestamp 1623621585
transform 1 0 10856 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_138_115
timestamp 1623621585
transform 1 0 11684 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_111
timestamp 1623621585
transform 1 0 11316 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_123
timestamp 1623621585
transform 1 0 12420 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1406
timestamp 1623621585
transform 1 0 14260 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_127
timestamp 1623621585
transform 1 0 12788 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_139
timestamp 1623621585
transform 1 0 13892 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_135
timestamp 1623621585
transform 1 0 13524 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_139_144
timestamp 1623621585
transform 1 0 14352 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_151
timestamp 1623621585
transform 1 0 14996 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_163
timestamp 1623621585
transform 1 0 16100 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_139_156
timestamp 1623621585
transform 1 0 15456 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1399
timestamp 1623621585
transform 1 0 16836 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_172
timestamp 1623621585
transform 1 0 16928 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_184
timestamp 1623621585
transform 1 0 18032 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_168
timestamp 1623621585
transform 1 0 16560 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_180
timestamp 1623621585
transform 1 0 17664 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1407
timestamp 1623621585
transform 1 0 19504 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_196
timestamp 1623621585
transform 1 0 19136 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_208
timestamp 1623621585
transform 1 0 20240 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_192
timestamp 1623621585
transform 1 0 18768 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_139_201
timestamp 1623621585
transform 1 0 19596 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1400
timestamp 1623621585
transform 1 0 22080 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_220
timestamp 1623621585
transform 1 0 21344 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_138_229
timestamp 1623621585
transform 1 0 22172 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_213
timestamp 1623621585
transform 1 0 20700 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_225
timestamp 1623621585
transform 1 0 21804 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_241
timestamp 1623621585
transform 1 0 23276 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_237
timestamp 1623621585
transform 1 0 22908 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_249
timestamp 1623621585
transform 1 0 24012 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1408
timestamp 1623621585
transform 1 0 24748 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_253
timestamp 1623621585
transform 1 0 24380 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_265
timestamp 1623621585
transform 1 0 25484 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_258
timestamp 1623621585
transform 1 0 24840 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_270
timestamp 1623621585
transform 1 0 25944 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1401
timestamp 1623621585
transform 1 0 27324 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_277
timestamp 1623621585
transform 1 0 26588 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_138_286
timestamp 1623621585
transform 1 0 27416 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_282
timestamp 1623621585
transform 1 0 27048 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_298
timestamp 1623621585
transform 1 0 28520 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_310
timestamp 1623621585
transform 1 0 29624 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_294
timestamp 1623621585
transform 1 0 28152 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_306
timestamp 1623621585
transform 1 0 29256 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1409
timestamp 1623621585
transform 1 0 29992 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_322
timestamp 1623621585
transform 1 0 30728 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_315
timestamp 1623621585
transform 1 0 30084 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_327
timestamp 1623621585
transform 1 0 31188 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _358_
timestamp 1623621585
transform 1 0 32384 0 1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1402
timestamp 1623621585
transform 1 0 32568 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_334
timestamp 1623621585
transform 1 0 31832 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_138_343
timestamp 1623621585
transform 1 0 32660 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_139_339
timestamp 1623621585
transform 1 0 32292 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_344
timestamp 1623621585
transform 1 0 32752 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1410
timestamp 1623621585
transform 1 0 35236 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_355
timestamp 1623621585
transform 1 0 33764 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_367
timestamp 1623621585
transform 1 0 34868 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_356
timestamp 1623621585
transform 1 0 33856 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_139_368
timestamp 1623621585
transform 1 0 34960 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_139_372
timestamp 1623621585
transform 1 0 35328 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input228
timestamp 1623621585
transform 1 0 37260 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_379
timestamp 1623621585
transform 1 0 35972 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_391
timestamp 1623621585
transform 1 0 37076 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_139_384
timestamp 1623621585
transform 1 0 36432 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_139_392
timestamp 1623621585
transform 1 0 37168 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1623621585
transform -1 0 38824 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_279
timestamp 1623621585
transform -1 0 38824 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1403
timestamp 1623621585
transform 1 0 37812 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input227
timestamp 1623621585
transform 1 0 37904 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_138_400
timestamp 1623621585
transform 1 0 37904 0 -1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_406
timestamp 1623621585
transform 1 0 38456 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_139_396
timestamp 1623621585
transform 1 0 37536 0 1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_139_403
timestamp 1623621585
transform 1 0 38180 0 1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_280
timestamp 1623621585
transform 1 0 1104 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input437
timestamp 1623621585
transform 1 0 1380 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_140_6
timestamp 1623621585
transform 1 0 1656 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_18
timestamp 1623621585
transform 1 0 2760 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_30
timestamp 1623621585
transform 1 0 3864 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1411
timestamp 1623621585
transform 1 0 6348 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_42
timestamp 1623621585
transform 1 0 4968 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_140_54
timestamp 1623621585
transform 1 0 6072 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_140_58
timestamp 1623621585
transform 1 0 6440 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_70
timestamp 1623621585
transform 1 0 7544 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_82
timestamp 1623621585
transform 1 0 8648 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_94
timestamp 1623621585
transform 1 0 9752 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1412
timestamp 1623621585
transform 1 0 11592 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_140_106
timestamp 1623621585
transform 1 0 10856 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_140_115
timestamp 1623621585
transform 1 0 11684 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_127
timestamp 1623621585
transform 1 0 12788 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_139
timestamp 1623621585
transform 1 0 13892 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_151
timestamp 1623621585
transform 1 0 14996 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_140_163
timestamp 1623621585
transform 1 0 16100 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1413
timestamp 1623621585
transform 1 0 16836 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_172
timestamp 1623621585
transform 1 0 16928 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_184
timestamp 1623621585
transform 1 0 18032 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_196
timestamp 1623621585
transform 1 0 19136 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_208
timestamp 1623621585
transform 1 0 20240 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1414
timestamp 1623621585
transform 1 0 22080 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_140_220
timestamp 1623621585
transform 1 0 21344 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_140_229
timestamp 1623621585
transform 1 0 22172 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_241
timestamp 1623621585
transform 1 0 23276 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_253
timestamp 1623621585
transform 1 0 24380 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_265
timestamp 1623621585
transform 1 0 25484 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _360_
timestamp 1623621585
transform 1 0 27784 0 -1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1415
timestamp 1623621585
transform 1 0 27324 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_140_277
timestamp 1623621585
transform 1 0 26588 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_140_286
timestamp 1623621585
transform 1 0 27416 0 -1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_140_294
timestamp 1623621585
transform 1 0 28152 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_306
timestamp 1623621585
transform 1 0 29256 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_318
timestamp 1623621585
transform 1 0 30360 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_330
timestamp 1623621585
transform 1 0 31464 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1416
timestamp 1623621585
transform 1 0 32568 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_343
timestamp 1623621585
transform 1 0 32660 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_355
timestamp 1623621585
transform 1 0 33764 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_367
timestamp 1623621585
transform 1 0 34868 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_379
timestamp 1623621585
transform 1 0 35972 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_140_391
timestamp 1623621585
transform 1 0 37076 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_281
timestamp 1623621585
transform -1 0 38824 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1417
timestamp 1623621585
transform 1 0 37812 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_140_400
timestamp 1623621585
transform 1 0 37904 0 -1 78880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_406
timestamp 1623621585
transform 1 0 38456 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_282
timestamp 1623621585
transform 1 0 1104 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_141_3
timestamp 1623621585
transform 1 0 1380 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_15
timestamp 1623621585
transform 1 0 2484 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1418
timestamp 1623621585
transform 1 0 3772 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_141_27
timestamp 1623621585
transform 1 0 3588 0 1 78880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_141_30
timestamp 1623621585
transform 1 0 3864 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_42
timestamp 1623621585
transform 1 0 4968 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_54
timestamp 1623621585
transform 1 0 6072 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_66
timestamp 1623621585
transform 1 0 7176 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_141_78
timestamp 1623621585
transform 1 0 8280 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1419
timestamp 1623621585
transform 1 0 9016 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_87
timestamp 1623621585
transform 1 0 9108 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_99
timestamp 1623621585
transform 1 0 10212 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_111
timestamp 1623621585
transform 1 0 11316 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_123
timestamp 1623621585
transform 1 0 12420 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1420
timestamp 1623621585
transform 1 0 14260 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_141_135
timestamp 1623621585
transform 1 0 13524 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_141_144
timestamp 1623621585
transform 1 0 14352 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_156
timestamp 1623621585
transform 1 0 15456 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_168
timestamp 1623621585
transform 1 0 16560 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_180
timestamp 1623621585
transform 1 0 17664 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1421
timestamp 1623621585
transform 1 0 19504 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_141_192
timestamp 1623621585
transform 1 0 18768 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_141_201
timestamp 1623621585
transform 1 0 19596 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_213
timestamp 1623621585
transform 1 0 20700 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_225
timestamp 1623621585
transform 1 0 21804 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_237
timestamp 1623621585
transform 1 0 22908 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_141_249
timestamp 1623621585
transform 1 0 24012 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1422
timestamp 1623621585
transform 1 0 24748 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_258
timestamp 1623621585
transform 1 0 24840 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_270
timestamp 1623621585
transform 1 0 25944 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_282
timestamp 1623621585
transform 1 0 27048 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_294
timestamp 1623621585
transform 1 0 28152 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_141_306
timestamp 1623621585
transform 1 0 29256 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1423
timestamp 1623621585
transform 1 0 29992 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_315
timestamp 1623621585
transform 1 0 30084 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_327
timestamp 1623621585
transform 1 0 31188 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_339
timestamp 1623621585
transform 1 0 32292 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_351
timestamp 1623621585
transform 1 0 33396 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1424
timestamp 1623621585
transform 1 0 35236 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_141_363
timestamp 1623621585
transform 1 0 34500 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_141_372
timestamp 1623621585
transform 1 0 35328 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input230
timestamp 1623621585
transform 1 0 37260 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_141_384
timestamp 1623621585
transform 1 0 36432 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_141_392
timestamp 1623621585
transform 1 0 37168 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_283
timestamp 1623621585
transform -1 0 38824 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input229
timestamp 1623621585
transform 1 0 37904 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_141_396
timestamp 1623621585
transform 1 0 37536 0 1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_141_403
timestamp 1623621585
transform 1 0 38180 0 1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_284
timestamp 1623621585
transform 1 0 1104 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input440
timestamp 1623621585
transform 1 0 1380 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_142_6
timestamp 1623621585
transform 1 0 1656 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_18
timestamp 1623621585
transform 1 0 2760 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_30
timestamp 1623621585
transform 1 0 3864 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1425
timestamp 1623621585
transform 1 0 6348 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_42
timestamp 1623621585
transform 1 0 4968 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_142_54
timestamp 1623621585
transform 1 0 6072 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_142_58
timestamp 1623621585
transform 1 0 6440 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_70
timestamp 1623621585
transform 1 0 7544 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_82
timestamp 1623621585
transform 1 0 8648 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_94
timestamp 1623621585
transform 1 0 9752 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1426
timestamp 1623621585
transform 1 0 11592 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_142_106
timestamp 1623621585
transform 1 0 10856 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_142_115
timestamp 1623621585
transform 1 0 11684 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_127
timestamp 1623621585
transform 1 0 12788 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_142_139
timestamp 1623621585
transform 1 0 13892 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _748_
timestamp 1623621585
transform 1 0 14812 0 -1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_142_147
timestamp 1623621585
transform 1 0 14628 0 -1 79968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_142_153
timestamp 1623621585
transform 1 0 15180 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_165
timestamp 1623621585
transform 1 0 16284 0 -1 79968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1427
timestamp 1623621585
transform 1 0 16836 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_172
timestamp 1623621585
transform 1 0 16928 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_184
timestamp 1623621585
transform 1 0 18032 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_196
timestamp 1623621585
transform 1 0 19136 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_208
timestamp 1623621585
transform 1 0 20240 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1428
timestamp 1623621585
transform 1 0 22080 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_142_220
timestamp 1623621585
transform 1 0 21344 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_142_229
timestamp 1623621585
transform 1 0 22172 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_241
timestamp 1623621585
transform 1 0 23276 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_253
timestamp 1623621585
transform 1 0 24380 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_265
timestamp 1623621585
transform 1 0 25484 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1429
timestamp 1623621585
transform 1 0 27324 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_142_277
timestamp 1623621585
transform 1 0 26588 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_142_286
timestamp 1623621585
transform 1 0 27416 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_298
timestamp 1623621585
transform 1 0 28520 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_310
timestamp 1623621585
transform 1 0 29624 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_322
timestamp 1623621585
transform 1 0 30728 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1430
timestamp 1623621585
transform 1 0 32568 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_142_334
timestamp 1623621585
transform 1 0 31832 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_142_343
timestamp 1623621585
transform 1 0 32660 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_355
timestamp 1623621585
transform 1 0 33764 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_367
timestamp 1623621585
transform 1 0 34868 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input232
timestamp 1623621585
transform 1 0 37168 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_142_379
timestamp 1623621585
transform 1 0 35972 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_391
timestamp 1623621585
transform 1 0 37076 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_142_395
timestamp 1623621585
transform 1 0 37444 0 -1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_285
timestamp 1623621585
transform -1 0 38824 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1431
timestamp 1623621585
transform 1 0 37812 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_142_400
timestamp 1623621585
transform 1 0 37904 0 -1 79968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_406
timestamp 1623621585
transform 1 0 38456 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_286
timestamp 1623621585
transform 1 0 1104 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input441
timestamp 1623621585
transform 1 0 1380 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_143_6
timestamp 1623621585
transform 1 0 1656 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_143_18
timestamp 1623621585
transform 1 0 2760 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1432
timestamp 1623621585
transform 1 0 3772 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_143_26
timestamp 1623621585
transform 1 0 3496 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_143_30
timestamp 1623621585
transform 1 0 3864 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_42
timestamp 1623621585
transform 1 0 4968 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_54
timestamp 1623621585
transform 1 0 6072 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_66
timestamp 1623621585
transform 1 0 7176 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_143_78
timestamp 1623621585
transform 1 0 8280 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1433
timestamp 1623621585
transform 1 0 9016 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_87
timestamp 1623621585
transform 1 0 9108 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_99
timestamp 1623621585
transform 1 0 10212 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_111
timestamp 1623621585
transform 1 0 11316 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_123
timestamp 1623621585
transform 1 0 12420 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1434
timestamp 1623621585
transform 1 0 14260 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_143_135
timestamp 1623621585
transform 1 0 13524 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_143_144
timestamp 1623621585
transform 1 0 14352 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_156
timestamp 1623621585
transform 1 0 15456 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_168
timestamp 1623621585
transform 1 0 16560 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_180
timestamp 1623621585
transform 1 0 17664 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1435
timestamp 1623621585
transform 1 0 19504 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_143_192
timestamp 1623621585
transform 1 0 18768 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_143_201
timestamp 1623621585
transform 1 0 19596 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_213
timestamp 1623621585
transform 1 0 20700 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_225
timestamp 1623621585
transform 1 0 21804 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_237
timestamp 1623621585
transform 1 0 22908 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_143_249
timestamp 1623621585
transform 1 0 24012 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1436
timestamp 1623621585
transform 1 0 24748 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_258
timestamp 1623621585
transform 1 0 24840 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_270
timestamp 1623621585
transform 1 0 25944 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_282
timestamp 1623621585
transform 1 0 27048 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_294
timestamp 1623621585
transform 1 0 28152 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_143_306
timestamp 1623621585
transform 1 0 29256 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _547_
timestamp 1623621585
transform 1 0 30912 0 1 79968
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1437
timestamp 1623621585
transform 1 0 29992 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_143_315
timestamp 1623621585
transform 1 0 30084 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_143_323
timestamp 1623621585
transform 1 0 30820 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_341
timestamp 1623621585
transform 1 0 32476 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_353
timestamp 1623621585
transform 1 0 33580 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1438
timestamp 1623621585
transform 1 0 35236 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_143_365
timestamp 1623621585
transform 1 0 34684 0 1 79968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_143_372
timestamp 1623621585
transform 1 0 35328 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input233
timestamp 1623621585
transform 1 0 37260 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_143_384
timestamp 1623621585
transform 1 0 36432 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_143_392
timestamp 1623621585
transform 1 0 37168 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_287
timestamp 1623621585
transform -1 0 38824 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input231
timestamp 1623621585
transform 1 0 37904 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_143_396
timestamp 1623621585
transform 1 0 37536 0 1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_143_403
timestamp 1623621585
transform 1 0 38180 0 1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_288
timestamp 1623621585
transform 1 0 1104 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input442
timestamp 1623621585
transform 1 0 1380 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_144_6
timestamp 1623621585
transform 1 0 1656 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_18
timestamp 1623621585
transform 1 0 2760 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_30
timestamp 1623621585
transform 1 0 3864 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1439
timestamp 1623621585
transform 1 0 6348 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_42
timestamp 1623621585
transform 1 0 4968 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_144_54
timestamp 1623621585
transform 1 0 6072 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_144_58
timestamp 1623621585
transform 1 0 6440 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_70
timestamp 1623621585
transform 1 0 7544 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_82
timestamp 1623621585
transform 1 0 8648 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_94
timestamp 1623621585
transform 1 0 9752 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1440
timestamp 1623621585
transform 1 0 11592 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_144_106
timestamp 1623621585
transform 1 0 10856 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_144_115
timestamp 1623621585
transform 1 0 11684 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_127
timestamp 1623621585
transform 1 0 12788 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_139
timestamp 1623621585
transform 1 0 13892 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_151
timestamp 1623621585
transform 1 0 14996 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_144_163
timestamp 1623621585
transform 1 0 16100 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1441
timestamp 1623621585
transform 1 0 16836 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_172
timestamp 1623621585
transform 1 0 16928 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_184
timestamp 1623621585
transform 1 0 18032 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_196
timestamp 1623621585
transform 1 0 19136 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_208
timestamp 1623621585
transform 1 0 20240 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1442
timestamp 1623621585
transform 1 0 22080 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_144_220
timestamp 1623621585
transform 1 0 21344 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_144_229
timestamp 1623621585
transform 1 0 22172 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_241
timestamp 1623621585
transform 1 0 23276 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_253
timestamp 1623621585
transform 1 0 24380 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_265
timestamp 1623621585
transform 1 0 25484 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1443
timestamp 1623621585
transform 1 0 27324 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_144_277
timestamp 1623621585
transform 1 0 26588 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_144_286
timestamp 1623621585
transform 1 0 27416 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_298
timestamp 1623621585
transform 1 0 28520 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_144_310
timestamp 1623621585
transform 1 0 29624 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _541_
timestamp 1623621585
transform 1 0 30636 0 -1 81056
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_144_318
timestamp 1623621585
transform 1 0 30360 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_4  _560_
timestamp 1623621585
transform 1 0 33028 0 -1 81056
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1444
timestamp 1623621585
transform 1 0 32568 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_144_338
timestamp 1623621585
transform 1 0 32200 0 -1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_144_343
timestamp 1623621585
transform 1 0 32660 0 -1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_144_364
timestamp 1623621585
transform 1 0 34592 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_376
timestamp 1623621585
transform 1 0 35696 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_144_388
timestamp 1623621585
transform 1 0 36800 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_289
timestamp 1623621585
transform -1 0 38824 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1445
timestamp 1623621585
transform 1 0 37812 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_144_396
timestamp 1623621585
transform 1 0 37536 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_144_400
timestamp 1623621585
transform 1 0 37904 0 -1 81056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_406
timestamp 1623621585
transform 1 0 38456 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_290
timestamp 1623621585
transform 1 0 1104 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_292
timestamp 1623621585
transform 1 0 1104 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input443
timestamp 1623621585
transform 1 0 1380 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_145_3
timestamp 1623621585
transform 1 0 1380 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_15
timestamp 1623621585
transform 1 0 2484 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_6
timestamp 1623621585
transform 1 0 1656 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_18
timestamp 1623621585
transform 1 0 2760 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1446
timestamp 1623621585
transform 1 0 3772 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_145_27
timestamp 1623621585
transform 1 0 3588 0 1 81056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_145_30
timestamp 1623621585
transform 1 0 3864 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_30
timestamp 1623621585
transform 1 0 3864 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1453
timestamp 1623621585
transform 1 0 6348 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_42
timestamp 1623621585
transform 1 0 4968 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_54
timestamp 1623621585
transform 1 0 6072 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_42
timestamp 1623621585
transform 1 0 4968 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_146_54
timestamp 1623621585
transform 1 0 6072 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_146_58
timestamp 1623621585
transform 1 0 6440 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_66
timestamp 1623621585
transform 1 0 7176 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_145_78
timestamp 1623621585
transform 1 0 8280 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_146_70
timestamp 1623621585
transform 1 0 7544 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_82
timestamp 1623621585
transform 1 0 8648 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1447
timestamp 1623621585
transform 1 0 9016 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_87
timestamp 1623621585
transform 1 0 9108 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_99
timestamp 1623621585
transform 1 0 10212 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_94
timestamp 1623621585
transform 1 0 9752 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1454
timestamp 1623621585
transform 1 0 11592 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_111
timestamp 1623621585
transform 1 0 11316 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_123
timestamp 1623621585
transform 1 0 12420 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_106
timestamp 1623621585
transform 1 0 10856 0 -1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_146_115
timestamp 1623621585
transform 1 0 11684 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1448
timestamp 1623621585
transform 1 0 14260 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_145_135
timestamp 1623621585
transform 1 0 13524 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_145_144
timestamp 1623621585
transform 1 0 14352 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_127
timestamp 1623621585
transform 1 0 12788 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_139
timestamp 1623621585
transform 1 0 13892 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_156
timestamp 1623621585
transform 1 0 15456 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_151
timestamp 1623621585
transform 1 0 14996 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_163
timestamp 1623621585
transform 1 0 16100 0 -1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1455
timestamp 1623621585
transform 1 0 16836 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_168
timestamp 1623621585
transform 1 0 16560 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_180
timestamp 1623621585
transform 1 0 17664 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_172
timestamp 1623621585
transform 1 0 16928 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_184
timestamp 1623621585
transform 1 0 18032 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1449
timestamp 1623621585
transform 1 0 19504 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_145_192
timestamp 1623621585
transform 1 0 18768 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_145_201
timestamp 1623621585
transform 1 0 19596 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_196
timestamp 1623621585
transform 1 0 19136 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_208
timestamp 1623621585
transform 1 0 20240 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1456
timestamp 1623621585
transform 1 0 22080 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_213
timestamp 1623621585
transform 1 0 20700 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_225
timestamp 1623621585
transform 1 0 21804 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_220
timestamp 1623621585
transform 1 0 21344 0 -1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_146_229
timestamp 1623621585
transform 1 0 22172 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_237
timestamp 1623621585
transform 1 0 22908 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_145_249
timestamp 1623621585
transform 1 0 24012 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_146_241
timestamp 1623621585
transform 1 0 23276 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1450
timestamp 1623621585
transform 1 0 24748 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_258
timestamp 1623621585
transform 1 0 24840 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_270
timestamp 1623621585
transform 1 0 25944 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_253
timestamp 1623621585
transform 1 0 24380 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_265
timestamp 1623621585
transform 1 0 25484 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1457
timestamp 1623621585
transform 1 0 27324 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_282
timestamp 1623621585
transform 1 0 27048 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_277
timestamp 1623621585
transform 1 0 26588 0 -1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_146_286
timestamp 1623621585
transform 1 0 27416 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_294
timestamp 1623621585
transform 1 0 28152 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_145_306
timestamp 1623621585
transform 1 0 29256 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_146_298
timestamp 1623621585
transform 1 0 28520 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_310
timestamp 1623621585
transform 1 0 29624 0 -1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _514_
timestamp 1623621585
transform 1 0 31280 0 1 81056
box -38 -48 1602 592
use sky130_fd_sc_hd__a221o_4  _521_
timestamp 1623621585
transform 1 0 30636 0 -1 82144
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1451
timestamp 1623621585
transform 1 0 29992 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_315
timestamp 1623621585
transform 1 0 30084 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_145_327
timestamp 1623621585
transform 1 0 31188 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_146_318
timestamp 1623621585
transform 1 0 30360 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_4  _530_
timestamp 1623621585
transform 1 0 33028 0 -1 82144
box -38 -48 1602 592
use sky130_fd_sc_hd__a221o_4  _554_
timestamp 1623621585
transform 1 0 33212 0 1 81056
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1458
timestamp 1623621585
transform 1 0 32568 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_145_345
timestamp 1623621585
transform 1 0 32844 0 1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_146_338
timestamp 1623621585
transform 1 0 32200 0 -1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_146_343
timestamp 1623621585
transform 1 0 32660 0 -1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1452
timestamp 1623621585
transform 1 0 35236 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_145_366
timestamp 1623621585
transform 1 0 34776 0 1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_145_370
timestamp 1623621585
transform 1 0 35144 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_372
timestamp 1623621585
transform 1 0 35328 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_364
timestamp 1623621585
transform 1 0 34592 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input236
timestamp 1623621585
transform 1 0 37260 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input238
timestamp 1623621585
transform 1 0 37168 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_145_384
timestamp 1623621585
transform 1 0 36432 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_145_392
timestamp 1623621585
transform 1 0 37168 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_376
timestamp 1623621585
transform 1 0 35696 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_146_388
timestamp 1623621585
transform 1 0 36800 0 -1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_146_395
timestamp 1623621585
transform 1 0 37444 0 -1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_291
timestamp 1623621585
transform -1 0 38824 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_293
timestamp 1623621585
transform -1 0 38824 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1459
timestamp 1623621585
transform 1 0 37812 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input235
timestamp 1623621585
transform 1 0 37904 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_145_396
timestamp 1623621585
transform 1 0 37536 0 1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_145_403
timestamp 1623621585
transform 1 0 38180 0 1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_146_400
timestamp 1623621585
transform 1 0 37904 0 -1 82144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_406
timestamp 1623621585
transform 1 0 38456 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_294
timestamp 1623621585
transform 1 0 1104 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input444
timestamp 1623621585
transform 1 0 1380 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_147_6
timestamp 1623621585
transform 1 0 1656 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_147_18
timestamp 1623621585
transform 1 0 2760 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1460
timestamp 1623621585
transform 1 0 3772 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_147_26
timestamp 1623621585
transform 1 0 3496 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_147_30
timestamp 1623621585
transform 1 0 3864 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_42
timestamp 1623621585
transform 1 0 4968 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_54
timestamp 1623621585
transform 1 0 6072 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_66
timestamp 1623621585
transform 1 0 7176 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_147_78
timestamp 1623621585
transform 1 0 8280 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1461
timestamp 1623621585
transform 1 0 9016 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_87
timestamp 1623621585
transform 1 0 9108 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_99
timestamp 1623621585
transform 1 0 10212 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_111
timestamp 1623621585
transform 1 0 11316 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_123
timestamp 1623621585
transform 1 0 12420 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1462
timestamp 1623621585
transform 1 0 14260 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_147_135
timestamp 1623621585
transform 1 0 13524 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_147_144
timestamp 1623621585
transform 1 0 14352 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_156
timestamp 1623621585
transform 1 0 15456 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_168
timestamp 1623621585
transform 1 0 16560 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_180
timestamp 1623621585
transform 1 0 17664 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1463
timestamp 1623621585
transform 1 0 19504 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_147_192
timestamp 1623621585
transform 1 0 18768 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_147_201
timestamp 1623621585
transform 1 0 19596 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_213
timestamp 1623621585
transform 1 0 20700 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_225
timestamp 1623621585
transform 1 0 21804 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_237
timestamp 1623621585
transform 1 0 22908 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_147_249
timestamp 1623621585
transform 1 0 24012 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1464
timestamp 1623621585
transform 1 0 24748 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_258
timestamp 1623621585
transform 1 0 24840 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_270
timestamp 1623621585
transform 1 0 25944 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_282
timestamp 1623621585
transform 1 0 27048 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_294
timestamp 1623621585
transform 1 0 28152 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_147_306
timestamp 1623621585
transform 1 0 29256 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _490_
timestamp 1623621585
transform 1 0 31464 0 1 82144
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1465
timestamp 1623621585
transform 1 0 29992 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_315
timestamp 1623621585
transform 1 0 30084 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_147_327
timestamp 1623621585
transform 1 0 31188 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_147_347
timestamp 1623621585
transform 1 0 33028 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1466
timestamp 1623621585
transform 1 0 35236 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_359
timestamp 1623621585
transform 1 0 34132 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_372
timestamp 1623621585
transform 1 0 35328 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input239
timestamp 1623621585
transform 1 0 37260 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_147_384
timestamp 1623621585
transform 1 0 36432 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_147_392
timestamp 1623621585
transform 1 0 37168 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_295
timestamp 1623621585
transform -1 0 38824 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input237
timestamp 1623621585
transform 1 0 37904 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_147_396
timestamp 1623621585
transform 1 0 37536 0 1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_147_403
timestamp 1623621585
transform 1 0 38180 0 1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_296
timestamp 1623621585
transform 1 0 1104 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_148_3
timestamp 1623621585
transform 1 0 1380 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_15
timestamp 1623621585
transform 1 0 2484 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_27
timestamp 1623621585
transform 1 0 3588 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_39
timestamp 1623621585
transform 1 0 4692 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1467
timestamp 1623621585
transform 1 0 6348 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_148_51
timestamp 1623621585
transform 1 0 5796 0 -1 83232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_148_58
timestamp 1623621585
transform 1 0 6440 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_70
timestamp 1623621585
transform 1 0 7544 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_82
timestamp 1623621585
transform 1 0 8648 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_94
timestamp 1623621585
transform 1 0 9752 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1468
timestamp 1623621585
transform 1 0 11592 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_148_106
timestamp 1623621585
transform 1 0 10856 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_148_115
timestamp 1623621585
transform 1 0 11684 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_127
timestamp 1623621585
transform 1 0 12788 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_139
timestamp 1623621585
transform 1 0 13892 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_151
timestamp 1623621585
transform 1 0 14996 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_148_163
timestamp 1623621585
transform 1 0 16100 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1469
timestamp 1623621585
transform 1 0 16836 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_172
timestamp 1623621585
transform 1 0 16928 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_184
timestamp 1623621585
transform 1 0 18032 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_196
timestamp 1623621585
transform 1 0 19136 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_208
timestamp 1623621585
transform 1 0 20240 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1470
timestamp 1623621585
transform 1 0 22080 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_148_220
timestamp 1623621585
transform 1 0 21344 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_148_229
timestamp 1623621585
transform 1 0 22172 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_241
timestamp 1623621585
transform 1 0 23276 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_253
timestamp 1623621585
transform 1 0 24380 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_265
timestamp 1623621585
transform 1 0 25484 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1471
timestamp 1623621585
transform 1 0 27324 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_148_277
timestamp 1623621585
transform 1 0 26588 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_148_286
timestamp 1623621585
transform 1 0 27416 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_298
timestamp 1623621585
transform 1 0 28520 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_148_310
timestamp 1623621585
transform 1 0 29624 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _501_
timestamp 1623621585
transform 1 0 30636 0 -1 83232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_148_318
timestamp 1623621585
transform 1 0 30360 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_4  _507_
timestamp 1623621585
transform 1 0 33028 0 -1 83232
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1472
timestamp 1623621585
transform 1 0 32568 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_148_338
timestamp 1623621585
transform 1 0 32200 0 -1 83232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_148_343
timestamp 1623621585
transform 1 0 32660 0 -1 83232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_148_364
timestamp 1623621585
transform 1 0 34592 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_376
timestamp 1623621585
transform 1 0 35696 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_148_388
timestamp 1623621585
transform 1 0 36800 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_297
timestamp 1623621585
transform -1 0 38824 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1473
timestamp 1623621585
transform 1 0 37812 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_148_396
timestamp 1623621585
transform 1 0 37536 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_148_400
timestamp 1623621585
transform 1 0 37904 0 -1 83232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_406
timestamp 1623621585
transform 1 0 38456 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_298
timestamp 1623621585
transform 1 0 1104 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input445
timestamp 1623621585
transform 1 0 1380 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_149_6
timestamp 1623621585
transform 1 0 1656 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_149_18
timestamp 1623621585
transform 1 0 2760 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1474
timestamp 1623621585
transform 1 0 3772 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_149_26
timestamp 1623621585
transform 1 0 3496 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_149_30
timestamp 1623621585
transform 1 0 3864 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_42
timestamp 1623621585
transform 1 0 4968 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_54
timestamp 1623621585
transform 1 0 6072 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_66
timestamp 1623621585
transform 1 0 7176 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_149_78
timestamp 1623621585
transform 1 0 8280 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1475
timestamp 1623621585
transform 1 0 9016 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_87
timestamp 1623621585
transform 1 0 9108 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_99
timestamp 1623621585
transform 1 0 10212 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_111
timestamp 1623621585
transform 1 0 11316 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_123
timestamp 1623621585
transform 1 0 12420 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1476
timestamp 1623621585
transform 1 0 14260 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_149_135
timestamp 1623621585
transform 1 0 13524 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_149_144
timestamp 1623621585
transform 1 0 14352 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_156
timestamp 1623621585
transform 1 0 15456 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_168
timestamp 1623621585
transform 1 0 16560 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_180
timestamp 1623621585
transform 1 0 17664 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1477
timestamp 1623621585
transform 1 0 19504 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_149_192
timestamp 1623621585
transform 1 0 18768 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_149_201
timestamp 1623621585
transform 1 0 19596 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_213
timestamp 1623621585
transform 1 0 20700 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_225
timestamp 1623621585
transform 1 0 21804 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_237
timestamp 1623621585
transform 1 0 22908 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_149_249
timestamp 1623621585
transform 1 0 24012 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1478
timestamp 1623621585
transform 1 0 24748 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_258
timestamp 1623621585
transform 1 0 24840 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_270
timestamp 1623621585
transform 1 0 25944 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_282
timestamp 1623621585
transform 1 0 27048 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_294
timestamp 1623621585
transform 1 0 28152 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_149_306
timestamp 1623621585
transform 1 0 29256 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1479
timestamp 1623621585
transform 1 0 29992 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_315
timestamp 1623621585
transform 1 0 30084 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_327
timestamp 1623621585
transform 1 0 31188 0 1 83232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_333
timestamp 1623621585
transform 1 0 31740 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_4  _467_
timestamp 1623621585
transform 1 0 31832 0 1 83232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_149_351
timestamp 1623621585
transform 1 0 33396 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1480
timestamp 1623621585
transform 1 0 35236 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_149_363
timestamp 1623621585
transform 1 0 34500 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_149_372
timestamp 1623621585
transform 1 0 35328 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input241
timestamp 1623621585
transform 1 0 37260 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_149_384
timestamp 1623621585
transform 1 0 36432 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_149_392
timestamp 1623621585
transform 1 0 37168 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_299
timestamp 1623621585
transform -1 0 38824 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input240
timestamp 1623621585
transform 1 0 37904 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_149_396
timestamp 1623621585
transform 1 0 37536 0 1 83232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_149_403
timestamp 1623621585
transform 1 0 38180 0 1 83232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_300
timestamp 1623621585
transform 1 0 1104 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input446
timestamp 1623621585
transform 1 0 1380 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_150_6
timestamp 1623621585
transform 1 0 1656 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_18
timestamp 1623621585
transform 1 0 2760 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_30
timestamp 1623621585
transform 1 0 3864 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1481
timestamp 1623621585
transform 1 0 6348 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_42
timestamp 1623621585
transform 1 0 4968 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_54
timestamp 1623621585
transform 1 0 6072 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_150_58
timestamp 1623621585
transform 1 0 6440 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_70
timestamp 1623621585
transform 1 0 7544 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_82
timestamp 1623621585
transform 1 0 8648 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_94
timestamp 1623621585
transform 1 0 9752 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1482
timestamp 1623621585
transform 1 0 11592 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_150_106
timestamp 1623621585
transform 1 0 10856 0 -1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_150_115
timestamp 1623621585
transform 1 0 11684 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_127
timestamp 1623621585
transform 1 0 12788 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_139
timestamp 1623621585
transform 1 0 13892 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_151
timestamp 1623621585
transform 1 0 14996 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_150_163
timestamp 1623621585
transform 1 0 16100 0 -1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1483
timestamp 1623621585
transform 1 0 16836 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_172
timestamp 1623621585
transform 1 0 16928 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_184
timestamp 1623621585
transform 1 0 18032 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_196
timestamp 1623621585
transform 1 0 19136 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_208
timestamp 1623621585
transform 1 0 20240 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1484
timestamp 1623621585
transform 1 0 22080 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_150_220
timestamp 1623621585
transform 1 0 21344 0 -1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_150_229
timestamp 1623621585
transform 1 0 22172 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_241
timestamp 1623621585
transform 1 0 23276 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_253
timestamp 1623621585
transform 1 0 24380 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_265
timestamp 1623621585
transform 1 0 25484 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1485
timestamp 1623621585
transform 1 0 27324 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_150_277
timestamp 1623621585
transform 1 0 26588 0 -1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_150_286
timestamp 1623621585
transform 1 0 27416 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_298
timestamp 1623621585
transform 1 0 28520 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_150_310
timestamp 1623621585
transform 1 0 29624 0 -1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _481_
timestamp 1623621585
transform 1 0 30636 0 -1 84320
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_150_318
timestamp 1623621585
transform 1 0 30360 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_4  _474_
timestamp 1623621585
transform 1 0 33028 0 -1 84320
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1486
timestamp 1623621585
transform 1 0 32568 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_150_338
timestamp 1623621585
transform 1 0 32200 0 -1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_150_343
timestamp 1623621585
transform 1 0 32660 0 -1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_150_364
timestamp 1623621585
transform 1 0 34592 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input243
timestamp 1623621585
transform 1 0 37168 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_150_376
timestamp 1623621585
transform 1 0 35696 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_150_388
timestamp 1623621585
transform 1 0 36800 0 -1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_150_395
timestamp 1623621585
transform 1 0 37444 0 -1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_301
timestamp 1623621585
transform -1 0 38824 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1487
timestamp 1623621585
transform 1 0 37812 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_150_400
timestamp 1623621585
transform 1 0 37904 0 -1 84320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_406
timestamp 1623621585
transform 1 0 38456 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_302
timestamp 1623621585
transform 1 0 1104 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_304
timestamp 1623621585
transform 1 0 1104 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input416
timestamp 1623621585
transform 1 0 1380 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_151_3
timestamp 1623621585
transform 1 0 1380 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_15
timestamp 1623621585
transform 1 0 2484 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_6
timestamp 1623621585
transform 1 0 1656 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_18
timestamp 1623621585
transform 1 0 2760 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1488
timestamp 1623621585
transform 1 0 3772 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_151_27
timestamp 1623621585
transform 1 0 3588 0 1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_151_30
timestamp 1623621585
transform 1 0 3864 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_30
timestamp 1623621585
transform 1 0 3864 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1495
timestamp 1623621585
transform 1 0 6348 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_42
timestamp 1623621585
transform 1 0 4968 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_54
timestamp 1623621585
transform 1 0 6072 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_42
timestamp 1623621585
transform 1 0 4968 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_152_54
timestamp 1623621585
transform 1 0 6072 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_152_58
timestamp 1623621585
transform 1 0 6440 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_66
timestamp 1623621585
transform 1 0 7176 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_78
timestamp 1623621585
transform 1 0 8280 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_152_70
timestamp 1623621585
transform 1 0 7544 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_82
timestamp 1623621585
transform 1 0 8648 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1489
timestamp 1623621585
transform 1 0 9016 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_87
timestamp 1623621585
transform 1 0 9108 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_99
timestamp 1623621585
transform 1 0 10212 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_94
timestamp 1623621585
transform 1 0 9752 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1496
timestamp 1623621585
transform 1 0 11592 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_111
timestamp 1623621585
transform 1 0 11316 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_123
timestamp 1623621585
transform 1 0 12420 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_106
timestamp 1623621585
transform 1 0 10856 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_152_115
timestamp 1623621585
transform 1 0 11684 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1490
timestamp 1623621585
transform 1 0 14260 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_135
timestamp 1623621585
transform 1 0 13524 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_151_144
timestamp 1623621585
transform 1 0 14352 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_127
timestamp 1623621585
transform 1 0 12788 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_139
timestamp 1623621585
transform 1 0 13892 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_156
timestamp 1623621585
transform 1 0 15456 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_151
timestamp 1623621585
transform 1 0 14996 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_163
timestamp 1623621585
transform 1 0 16100 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1497
timestamp 1623621585
transform 1 0 16836 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_168
timestamp 1623621585
transform 1 0 16560 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_180
timestamp 1623621585
transform 1 0 17664 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_172
timestamp 1623621585
transform 1 0 16928 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_184
timestamp 1623621585
transform 1 0 18032 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1491
timestamp 1623621585
transform 1 0 19504 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_192
timestamp 1623621585
transform 1 0 18768 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_151_201
timestamp 1623621585
transform 1 0 19596 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_196
timestamp 1623621585
transform 1 0 19136 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_208
timestamp 1623621585
transform 1 0 20240 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1498
timestamp 1623621585
transform 1 0 22080 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_213
timestamp 1623621585
transform 1 0 20700 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_225
timestamp 1623621585
transform 1 0 21804 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_220
timestamp 1623621585
transform 1 0 21344 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_152_229
timestamp 1623621585
transform 1 0 22172 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_237
timestamp 1623621585
transform 1 0 22908 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_249
timestamp 1623621585
transform 1 0 24012 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_152_241
timestamp 1623621585
transform 1 0 23276 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1492
timestamp 1623621585
transform 1 0 24748 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_258
timestamp 1623621585
transform 1 0 24840 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_270
timestamp 1623621585
transform 1 0 25944 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_152_253
timestamp 1623621585
transform 1 0 24380 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_265
timestamp 1623621585
transform 1 0 25484 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _527_
timestamp 1623621585
transform 1 0 26956 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1499
timestamp 1623621585
transform 1 0 27324 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_151_278
timestamp 1623621585
transform 1 0 26680 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_151_285
timestamp 1623621585
transform 1 0 27324 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_277
timestamp 1623621585
transform 1 0 26588 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_152_286
timestamp 1623621585
transform 1 0 27416 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_297
timestamp 1623621585
transform 1 0 28428 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_151_309
timestamp 1623621585
transform 1 0 29532 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_152_298
timestamp 1623621585
transform 1 0 28520 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_310
timestamp 1623621585
transform 1 0 29624 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _526_
timestamp 1623621585
transform 1 0 31280 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1493
timestamp 1623621585
transform 1 0 29992 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_151_313
timestamp 1623621585
transform 1 0 29900 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_315
timestamp 1623621585
transform 1 0 30084 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_151_327
timestamp 1623621585
transform 1 0 31188 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_151_332
timestamp 1623621585
transform 1 0 31648 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_152_322
timestamp 1623621585
transform 1 0 30728 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_4  _450_
timestamp 1623621585
transform 1 0 32016 0 1 84320
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _486_
timestamp 1623621585
transform 1 0 33028 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1500
timestamp 1623621585
transform 1 0 32568 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_353
timestamp 1623621585
transform 1 0 33580 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_334
timestamp 1623621585
transform 1 0 31832 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_152_343
timestamp 1623621585
transform 1 0 32660 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_152_351
timestamp 1623621585
transform 1 0 33396 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1494
timestamp 1623621585
transform 1 0 35236 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_151_365
timestamp 1623621585
transform 1 0 34684 0 1 84320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_151_372
timestamp 1623621585
transform 1 0 35328 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_363
timestamp 1623621585
transform 1 0 34500 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_375
timestamp 1623621585
transform 1 0 35604 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input244
timestamp 1623621585
transform 1 0 37260 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_151_384
timestamp 1623621585
transform 1 0 36432 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_392
timestamp 1623621585
transform 1 0 37168 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_387
timestamp 1623621585
transform 1 0 36708 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_303
timestamp 1623621585
transform -1 0 38824 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_305
timestamp 1623621585
transform -1 0 38824 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1501
timestamp 1623621585
transform 1 0 37812 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input242
timestamp 1623621585
transform 1 0 37904 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_151_396
timestamp 1623621585
transform 1 0 37536 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_403
timestamp 1623621585
transform 1 0 38180 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_152_400
timestamp 1623621585
transform 1 0 37904 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_406
timestamp 1623621585
transform 1 0 38456 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_306
timestamp 1623621585
transform 1 0 1104 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input417
timestamp 1623621585
transform 1 0 1380 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_153_6
timestamp 1623621585
transform 1 0 1656 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_153_18
timestamp 1623621585
transform 1 0 2760 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1502
timestamp 1623621585
transform 1 0 3772 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_153_26
timestamp 1623621585
transform 1 0 3496 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_153_30
timestamp 1623621585
transform 1 0 3864 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_42
timestamp 1623621585
transform 1 0 4968 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_54
timestamp 1623621585
transform 1 0 6072 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_66
timestamp 1623621585
transform 1 0 7176 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_153_78
timestamp 1623621585
transform 1 0 8280 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1503
timestamp 1623621585
transform 1 0 9016 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_87
timestamp 1623621585
transform 1 0 9108 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_99
timestamp 1623621585
transform 1 0 10212 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_111
timestamp 1623621585
transform 1 0 11316 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_123
timestamp 1623621585
transform 1 0 12420 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1504
timestamp 1623621585
transform 1 0 14260 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_153_135
timestamp 1623621585
transform 1 0 13524 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_153_144
timestamp 1623621585
transform 1 0 14352 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_156
timestamp 1623621585
transform 1 0 15456 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_168
timestamp 1623621585
transform 1 0 16560 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_180
timestamp 1623621585
transform 1 0 17664 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1505
timestamp 1623621585
transform 1 0 19504 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_153_192
timestamp 1623621585
transform 1 0 18768 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_153_201
timestamp 1623621585
transform 1 0 19596 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_213
timestamp 1623621585
transform 1 0 20700 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_225
timestamp 1623621585
transform 1 0 21804 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_237
timestamp 1623621585
transform 1 0 22908 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_153_249
timestamp 1623621585
transform 1 0 24012 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1506
timestamp 1623621585
transform 1 0 24748 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_258
timestamp 1623621585
transform 1 0 24840 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_270
timestamp 1623621585
transform 1 0 25944 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _487_
timestamp 1623621585
transform 1 0 27140 0 1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_153_282
timestamp 1623621585
transform 1 0 27048 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_287
timestamp 1623621585
transform 1 0 27508 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_299
timestamp 1623621585
transform 1 0 28612 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_153_311
timestamp 1623621585
transform 1 0 29716 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1507
timestamp 1623621585
transform 1 0 29992 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_315
timestamp 1623621585
transform 1 0 30084 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_153_327
timestamp 1623621585
transform 1 0 31188 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _461_
timestamp 1623621585
transform 1 0 31924 0 1 85408
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_153_352
timestamp 1623621585
transform 1 0 33488 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1508
timestamp 1623621585
transform 1 0 35236 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_153_364
timestamp 1623621585
transform 1 0 34592 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_370
timestamp 1623621585
transform 1 0 35144 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_372
timestamp 1623621585
transform 1 0 35328 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input247
timestamp 1623621585
transform 1 0 37260 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_153_384
timestamp 1623621585
transform 1 0 36432 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_153_392
timestamp 1623621585
transform 1 0 37168 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_307
timestamp 1623621585
transform -1 0 38824 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input246
timestamp 1623621585
transform 1 0 37904 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_153_396
timestamp 1623621585
transform 1 0 37536 0 1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_153_403
timestamp 1623621585
transform 1 0 38180 0 1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_308
timestamp 1623621585
transform 1 0 1104 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_154_3
timestamp 1623621585
transform 1 0 1380 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_15
timestamp 1623621585
transform 1 0 2484 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_27
timestamp 1623621585
transform 1 0 3588 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_39
timestamp 1623621585
transform 1 0 4692 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1509
timestamp 1623621585
transform 1 0 6348 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_154_51
timestamp 1623621585
transform 1 0 5796 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_154_58
timestamp 1623621585
transform 1 0 6440 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_70
timestamp 1623621585
transform 1 0 7544 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_82
timestamp 1623621585
transform 1 0 8648 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_94
timestamp 1623621585
transform 1 0 9752 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1510
timestamp 1623621585
transform 1 0 11592 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_154_106
timestamp 1623621585
transform 1 0 10856 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_154_115
timestamp 1623621585
transform 1 0 11684 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_127
timestamp 1623621585
transform 1 0 12788 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_139
timestamp 1623621585
transform 1 0 13892 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_151
timestamp 1623621585
transform 1 0 14996 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_154_163
timestamp 1623621585
transform 1 0 16100 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1511
timestamp 1623621585
transform 1 0 16836 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_172
timestamp 1623621585
transform 1 0 16928 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_184
timestamp 1623621585
transform 1 0 18032 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_196
timestamp 1623621585
transform 1 0 19136 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_208
timestamp 1623621585
transform 1 0 20240 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1512
timestamp 1623621585
transform 1 0 22080 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_154_220
timestamp 1623621585
transform 1 0 21344 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_154_229
timestamp 1623621585
transform 1 0 22172 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_241
timestamp 1623621585
transform 1 0 23276 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_253
timestamp 1623621585
transform 1 0 24380 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_265
timestamp 1623621585
transform 1 0 25484 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1513
timestamp 1623621585
transform 1 0 27324 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_154_277
timestamp 1623621585
transform 1 0 26588 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_154_286
timestamp 1623621585
transform 1 0 27416 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_298
timestamp 1623621585
transform 1 0 28520 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_310
timestamp 1623621585
transform 1 0 29624 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_322
timestamp 1623621585
transform 1 0 30728 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_4  _345_
timestamp 1623621585
transform 1 0 33212 0 -1 86496
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1514
timestamp 1623621585
transform 1 0 32568 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_154_334
timestamp 1623621585
transform 1 0 31832 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_154_343
timestamp 1623621585
transform 1 0 32660 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_154_366
timestamp 1623621585
transform 1 0 34776 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_378
timestamp 1623621585
transform 1 0 35880 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_154_390
timestamp 1623621585
transform 1 0 36984 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_309
timestamp 1623621585
transform -1 0 38824 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1515
timestamp 1623621585
transform 1 0 37812 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_154_398
timestamp 1623621585
transform 1 0 37720 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_154_400
timestamp 1623621585
transform 1 0 37904 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_406
timestamp 1623621585
transform 1 0 38456 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_310
timestamp 1623621585
transform 1 0 1104 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input418
timestamp 1623621585
transform 1 0 1380 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_155_6
timestamp 1623621585
transform 1 0 1656 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_155_18
timestamp 1623621585
transform 1 0 2760 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1516
timestamp 1623621585
transform 1 0 3772 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_155_26
timestamp 1623621585
transform 1 0 3496 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_155_30
timestamp 1623621585
transform 1 0 3864 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_42
timestamp 1623621585
transform 1 0 4968 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_54
timestamp 1623621585
transform 1 0 6072 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_66
timestamp 1623621585
transform 1 0 7176 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_155_78
timestamp 1623621585
transform 1 0 8280 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1517
timestamp 1623621585
transform 1 0 9016 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_87
timestamp 1623621585
transform 1 0 9108 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_99
timestamp 1623621585
transform 1 0 10212 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_111
timestamp 1623621585
transform 1 0 11316 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_123
timestamp 1623621585
transform 1 0 12420 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1518
timestamp 1623621585
transform 1 0 14260 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_155_135
timestamp 1623621585
transform 1 0 13524 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_155_144
timestamp 1623621585
transform 1 0 14352 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_156
timestamp 1623621585
transform 1 0 15456 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_168
timestamp 1623621585
transform 1 0 16560 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_180
timestamp 1623621585
transform 1 0 17664 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1519
timestamp 1623621585
transform 1 0 19504 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_155_192
timestamp 1623621585
transform 1 0 18768 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_155_201
timestamp 1623621585
transform 1 0 19596 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_213
timestamp 1623621585
transform 1 0 20700 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_225
timestamp 1623621585
transform 1 0 21804 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_237
timestamp 1623621585
transform 1 0 22908 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_155_249
timestamp 1623621585
transform 1 0 24012 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1520
timestamp 1623621585
transform 1 0 24748 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_258
timestamp 1623621585
transform 1 0 24840 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_270
timestamp 1623621585
transform 1 0 25944 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _323_
timestamp 1623621585
transform 1 0 27784 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _447_
timestamp 1623621585
transform 1 0 27048 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_155_286
timestamp 1623621585
transform 1 0 27416 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_155_294
timestamp 1623621585
transform 1 0 28152 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_155_306
timestamp 1623621585
transform 1 0 29256 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _446_
timestamp 1623621585
transform 1 0 31740 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1521
timestamp 1623621585
transform 1 0 29992 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_315
timestamp 1623621585
transform 1 0 30084 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_327
timestamp 1623621585
transform 1 0 31188 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _322_
timestamp 1623621585
transform 1 0 32476 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_4  _326_
timestamp 1623621585
transform 1 0 33212 0 1 86496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_155_337
timestamp 1623621585
transform 1 0 32108 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_155_345
timestamp 1623621585
transform 1 0 32844 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1522
timestamp 1623621585
transform 1 0 35236 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_155_366
timestamp 1623621585
transform 1 0 34776 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_155_370
timestamp 1623621585
transform 1 0 35144 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_372
timestamp 1623621585
transform 1 0 35328 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input266
timestamp 1623621585
transform 1 0 37260 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_155_384
timestamp 1623621585
transform 1 0 36432 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_155_392
timestamp 1623621585
transform 1 0 37168 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_311
timestamp 1623621585
transform -1 0 38824 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input255
timestamp 1623621585
transform 1 0 37904 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_155_396
timestamp 1623621585
transform 1 0 37536 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_155_403
timestamp 1623621585
transform 1 0 38180 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_312
timestamp 1623621585
transform 1 0 1104 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input419
timestamp 1623621585
transform 1 0 1380 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_156_6
timestamp 1623621585
transform 1 0 1656 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_18
timestamp 1623621585
transform 1 0 2760 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_30
timestamp 1623621585
transform 1 0 3864 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1523
timestamp 1623621585
transform 1 0 6348 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_42
timestamp 1623621585
transform 1 0 4968 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_156_54
timestamp 1623621585
transform 1 0 6072 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_156_58
timestamp 1623621585
transform 1 0 6440 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_70
timestamp 1623621585
transform 1 0 7544 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_82
timestamp 1623621585
transform 1 0 8648 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_94
timestamp 1623621585
transform 1 0 9752 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1524
timestamp 1623621585
transform 1 0 11592 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_156_106
timestamp 1623621585
transform 1 0 10856 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_156_115
timestamp 1623621585
transform 1 0 11684 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_127
timestamp 1623621585
transform 1 0 12788 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_139
timestamp 1623621585
transform 1 0 13892 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_151
timestamp 1623621585
transform 1 0 14996 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_156_163
timestamp 1623621585
transform 1 0 16100 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1525
timestamp 1623621585
transform 1 0 16836 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_172
timestamp 1623621585
transform 1 0 16928 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_184
timestamp 1623621585
transform 1 0 18032 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_196
timestamp 1623621585
transform 1 0 19136 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_208
timestamp 1623621585
transform 1 0 20240 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1526
timestamp 1623621585
transform 1 0 22080 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_156_220
timestamp 1623621585
transform 1 0 21344 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_156_229
timestamp 1623621585
transform 1 0 22172 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_241
timestamp 1623621585
transform 1 0 23276 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_253
timestamp 1623621585
transform 1 0 24380 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_265
timestamp 1623621585
transform 1 0 25484 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1527
timestamp 1623621585
transform 1 0 27324 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_156_277
timestamp 1623621585
transform 1 0 26588 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_156_286
timestamp 1623621585
transform 1 0 27416 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_298
timestamp 1623621585
transform 1 0 28520 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_310
timestamp 1623621585
transform 1 0 29624 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_322
timestamp 1623621585
transform 1 0 30728 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_4  _337_
timestamp 1623621585
transform 1 0 33212 0 -1 87584
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1528
timestamp 1623621585
transform 1 0 32568 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_156_334
timestamp 1623621585
transform 1 0 31832 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_156_343
timestamp 1623621585
transform 1 0 32660 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_156_366
timestamp 1623621585
transform 1 0 34776 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input280
timestamp 1623621585
transform 1 0 37168 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_156_378
timestamp 1623621585
transform 1 0 35880 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_156_390
timestamp 1623621585
transform 1 0 36984 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_156_395
timestamp 1623621585
transform 1 0 37444 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_313
timestamp 1623621585
transform -1 0 38824 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1529
timestamp 1623621585
transform 1 0 37812 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_156_400
timestamp 1623621585
transform 1 0 37904 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_406
timestamp 1623621585
transform 1 0 38456 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_314
timestamp 1623621585
transform 1 0 1104 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_157_3
timestamp 1623621585
transform 1 0 1380 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_15
timestamp 1623621585
transform 1 0 2484 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1530
timestamp 1623621585
transform 1 0 3772 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_157_27
timestamp 1623621585
transform 1 0 3588 0 1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_157_30
timestamp 1623621585
transform 1 0 3864 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_42
timestamp 1623621585
transform 1 0 4968 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_54
timestamp 1623621585
transform 1 0 6072 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_66
timestamp 1623621585
transform 1 0 7176 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_157_78
timestamp 1623621585
transform 1 0 8280 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1531
timestamp 1623621585
transform 1 0 9016 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_87
timestamp 1623621585
transform 1 0 9108 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_99
timestamp 1623621585
transform 1 0 10212 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_111
timestamp 1623621585
transform 1 0 11316 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_123
timestamp 1623621585
transform 1 0 12420 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1532
timestamp 1623621585
transform 1 0 14260 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_157_135
timestamp 1623621585
transform 1 0 13524 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_157_144
timestamp 1623621585
transform 1 0 14352 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_156
timestamp 1623621585
transform 1 0 15456 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_168
timestamp 1623621585
transform 1 0 16560 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_180
timestamp 1623621585
transform 1 0 17664 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1533
timestamp 1623621585
transform 1 0 19504 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_157_192
timestamp 1623621585
transform 1 0 18768 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_157_201
timestamp 1623621585
transform 1 0 19596 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_213
timestamp 1623621585
transform 1 0 20700 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_225
timestamp 1623621585
transform 1 0 21804 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_237
timestamp 1623621585
transform 1 0 22908 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_157_249
timestamp 1623621585
transform 1 0 24012 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1534
timestamp 1623621585
transform 1 0 24748 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_258
timestamp 1623621585
transform 1 0 24840 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_270
timestamp 1623621585
transform 1 0 25944 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_282
timestamp 1623621585
transform 1 0 27048 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_294
timestamp 1623621585
transform 1 0 28152 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_157_306
timestamp 1623621585
transform 1 0 29256 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1535
timestamp 1623621585
transform 1 0 29992 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_315
timestamp 1623621585
transform 1 0 30084 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_327
timestamp 1623621585
transform 1 0 31188 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_4  _353_
timestamp 1623621585
transform 1 0 33212 0 1 87584
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_157_339
timestamp 1623621585
transform 1 0 32292 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_157_347
timestamp 1623621585
transform 1 0 33028 0 1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1536
timestamp 1623621585
transform 1 0 35236 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_157_366
timestamp 1623621585
transform 1 0 34776 0 1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_157_370
timestamp 1623621585
transform 1 0 35144 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_372
timestamp 1623621585
transform 1 0 35328 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input281
timestamp 1623621585
transform 1 0 37260 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_157_384
timestamp 1623621585
transform 1 0 36432 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_157_392
timestamp 1623621585
transform 1 0 37168 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_315
timestamp 1623621585
transform -1 0 38824 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input277
timestamp 1623621585
transform 1 0 37904 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_157_396
timestamp 1623621585
transform 1 0 37536 0 1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_157_403
timestamp 1623621585
transform 1 0 38180 0 1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_316
timestamp 1623621585
transform 1 0 1104 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_318
timestamp 1623621585
transform 1 0 1104 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input420
timestamp 1623621585
transform 1 0 1380 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input421
timestamp 1623621585
transform 1 0 1380 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_158_6
timestamp 1623621585
transform 1 0 1656 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_18
timestamp 1623621585
transform 1 0 2760 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_6
timestamp 1623621585
transform 1 0 1656 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_18
timestamp 1623621585
transform 1 0 2760 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1544
timestamp 1623621585
transform 1 0 3772 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_30
timestamp 1623621585
transform 1 0 3864 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_159_26
timestamp 1623621585
transform 1 0 3496 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_159_30
timestamp 1623621585
transform 1 0 3864 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1537
timestamp 1623621585
transform 1 0 6348 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_42
timestamp 1623621585
transform 1 0 4968 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_158_54
timestamp 1623621585
transform 1 0 6072 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_158_58
timestamp 1623621585
transform 1 0 6440 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_42
timestamp 1623621585
transform 1 0 4968 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_54
timestamp 1623621585
transform 1 0 6072 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_70
timestamp 1623621585
transform 1 0 7544 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_82
timestamp 1623621585
transform 1 0 8648 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_66
timestamp 1623621585
transform 1 0 7176 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_78
timestamp 1623621585
transform 1 0 8280 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1545
timestamp 1623621585
transform 1 0 9016 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_94
timestamp 1623621585
transform 1 0 9752 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_87
timestamp 1623621585
transform 1 0 9108 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_99
timestamp 1623621585
transform 1 0 10212 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1538
timestamp 1623621585
transform 1 0 11592 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_158_106
timestamp 1623621585
transform 1 0 10856 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_158_115
timestamp 1623621585
transform 1 0 11684 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_111
timestamp 1623621585
transform 1 0 11316 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_123
timestamp 1623621585
transform 1 0 12420 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1546
timestamp 1623621585
transform 1 0 14260 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_127
timestamp 1623621585
transform 1 0 12788 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_139
timestamp 1623621585
transform 1 0 13892 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_135
timestamp 1623621585
transform 1 0 13524 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_159_144
timestamp 1623621585
transform 1 0 14352 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_151
timestamp 1623621585
transform 1 0 14996 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_158_163
timestamp 1623621585
transform 1 0 16100 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_159_156
timestamp 1623621585
transform 1 0 15456 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1539
timestamp 1623621585
transform 1 0 16836 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_172
timestamp 1623621585
transform 1 0 16928 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_184
timestamp 1623621585
transform 1 0 18032 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_168
timestamp 1623621585
transform 1 0 16560 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_180
timestamp 1623621585
transform 1 0 17664 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1547
timestamp 1623621585
transform 1 0 19504 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_196
timestamp 1623621585
transform 1 0 19136 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_208
timestamp 1623621585
transform 1 0 20240 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_192
timestamp 1623621585
transform 1 0 18768 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_159_201
timestamp 1623621585
transform 1 0 19596 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1540
timestamp 1623621585
transform 1 0 22080 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_158_220
timestamp 1623621585
transform 1 0 21344 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_158_229
timestamp 1623621585
transform 1 0 22172 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_213
timestamp 1623621585
transform 1 0 20700 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_225
timestamp 1623621585
transform 1 0 21804 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_241
timestamp 1623621585
transform 1 0 23276 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_237
timestamp 1623621585
transform 1 0 22908 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_249
timestamp 1623621585
transform 1 0 24012 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1548
timestamp 1623621585
transform 1 0 24748 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_253
timestamp 1623621585
transform 1 0 24380 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_265
timestamp 1623621585
transform 1 0 25484 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_258
timestamp 1623621585
transform 1 0 24840 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_270
timestamp 1623621585
transform 1 0 25944 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1541
timestamp 1623621585
transform 1 0 27324 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_158_277
timestamp 1623621585
transform 1 0 26588 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_158_286
timestamp 1623621585
transform 1 0 27416 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_282
timestamp 1623621585
transform 1 0 27048 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_298
timestamp 1623621585
transform 1 0 28520 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_310
timestamp 1623621585
transform 1 0 29624 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_294
timestamp 1623621585
transform 1 0 28152 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_306
timestamp 1623621585
transform 1 0 29256 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1549
timestamp 1623621585
transform 1 0 29992 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_322
timestamp 1623621585
transform 1 0 30728 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_315
timestamp 1623621585
transform 1 0 30084 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_327
timestamp 1623621585
transform 1 0 31188 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1542
timestamp 1623621585
transform 1 0 32568 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_158_334
timestamp 1623621585
transform 1 0 31832 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_158_343
timestamp 1623621585
transform 1 0 32660 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_339
timestamp 1623621585
transform 1 0 32292 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_351
timestamp 1623621585
transform 1 0 33396 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1550
timestamp 1623621585
transform 1 0 35236 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_355
timestamp 1623621585
transform 1 0 33764 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_367
timestamp 1623621585
transform 1 0 34868 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_363
timestamp 1623621585
transform 1 0 34500 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_159_372
timestamp 1623621585
transform 1 0 35328 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input283
timestamp 1623621585
transform 1 0 37260 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_158_379
timestamp 1623621585
transform 1 0 35972 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_158_391
timestamp 1623621585
transform 1 0 37076 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_159_384
timestamp 1623621585
transform 1 0 36432 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_159_392
timestamp 1623621585
transform 1 0 37168 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_317
timestamp 1623621585
transform -1 0 38824 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_319
timestamp 1623621585
transform -1 0 38824 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1543
timestamp 1623621585
transform 1 0 37812 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input282
timestamp 1623621585
transform 1 0 37904 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_158_400
timestamp 1623621585
transform 1 0 37904 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_406
timestamp 1623621585
transform 1 0 38456 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_159_396
timestamp 1623621585
transform 1 0 37536 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_159_403
timestamp 1623621585
transform 1 0 38180 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_320
timestamp 1623621585
transform 1 0 1104 0 -1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_160_3
timestamp 1623621585
transform 1 0 1380 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_15
timestamp 1623621585
transform 1 0 2484 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_27
timestamp 1623621585
transform 1 0 3588 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_39
timestamp 1623621585
transform 1 0 4692 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1551
timestamp 1623621585
transform 1 0 6348 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_160_51
timestamp 1623621585
transform 1 0 5796 0 -1 89760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_160_58
timestamp 1623621585
transform 1 0 6440 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_70
timestamp 1623621585
transform 1 0 7544 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_82
timestamp 1623621585
transform 1 0 8648 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_94
timestamp 1623621585
transform 1 0 9752 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1552
timestamp 1623621585
transform 1 0 11592 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_160_106
timestamp 1623621585
transform 1 0 10856 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_160_115
timestamp 1623621585
transform 1 0 11684 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_127
timestamp 1623621585
transform 1 0 12788 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_139
timestamp 1623621585
transform 1 0 13892 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_151
timestamp 1623621585
transform 1 0 14996 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_160_163
timestamp 1623621585
transform 1 0 16100 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1553
timestamp 1623621585
transform 1 0 16836 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_172
timestamp 1623621585
transform 1 0 16928 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_184
timestamp 1623621585
transform 1 0 18032 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_196
timestamp 1623621585
transform 1 0 19136 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_208
timestamp 1623621585
transform 1 0 20240 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1554
timestamp 1623621585
transform 1 0 22080 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_160_220
timestamp 1623621585
transform 1 0 21344 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_160_229
timestamp 1623621585
transform 1 0 22172 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_241
timestamp 1623621585
transform 1 0 23276 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_253
timestamp 1623621585
transform 1 0 24380 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_265
timestamp 1623621585
transform 1 0 25484 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1555
timestamp 1623621585
transform 1 0 27324 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_160_277
timestamp 1623621585
transform 1 0 26588 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_160_286
timestamp 1623621585
transform 1 0 27416 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_298
timestamp 1623621585
transform 1 0 28520 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_310
timestamp 1623621585
transform 1 0 29624 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_322
timestamp 1623621585
transform 1 0 30728 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1556
timestamp 1623621585
transform 1 0 32568 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_160_334
timestamp 1623621585
transform 1 0 31832 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_160_343
timestamp 1623621585
transform 1 0 32660 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_355
timestamp 1623621585
transform 1 0 33764 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_367
timestamp 1623621585
transform 1 0 34868 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input285
timestamp 1623621585
transform 1 0 37168 0 -1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_160_379
timestamp 1623621585
transform 1 0 35972 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_391
timestamp 1623621585
transform 1 0 37076 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_160_395
timestamp 1623621585
transform 1 0 37444 0 -1 89760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_321
timestamp 1623621585
transform -1 0 38824 0 -1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1557
timestamp 1623621585
transform 1 0 37812 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_160_400
timestamp 1623621585
transform 1 0 37904 0 -1 89760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_406
timestamp 1623621585
transform 1 0 38456 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_322
timestamp 1623621585
transform 1 0 1104 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input422
timestamp 1623621585
transform 1 0 1380 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_161_6
timestamp 1623621585
transform 1 0 1656 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_18
timestamp 1623621585
transform 1 0 2760 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1558
timestamp 1623621585
transform 1 0 3772 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_161_26
timestamp 1623621585
transform 1 0 3496 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_161_30
timestamp 1623621585
transform 1 0 3864 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_42
timestamp 1623621585
transform 1 0 4968 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_54
timestamp 1623621585
transform 1 0 6072 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_66
timestamp 1623621585
transform 1 0 7176 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_78
timestamp 1623621585
transform 1 0 8280 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1559
timestamp 1623621585
transform 1 0 9016 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_87
timestamp 1623621585
transform 1 0 9108 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_99
timestamp 1623621585
transform 1 0 10212 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_111
timestamp 1623621585
transform 1 0 11316 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_123
timestamp 1623621585
transform 1 0 12420 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1560
timestamp 1623621585
transform 1 0 14260 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_161_135
timestamp 1623621585
transform 1 0 13524 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_161_144
timestamp 1623621585
transform 1 0 14352 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_156
timestamp 1623621585
transform 1 0 15456 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_168
timestamp 1623621585
transform 1 0 16560 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_180
timestamp 1623621585
transform 1 0 17664 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1561
timestamp 1623621585
transform 1 0 19504 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_161_192
timestamp 1623621585
transform 1 0 18768 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_161_201
timestamp 1623621585
transform 1 0 19596 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_213
timestamp 1623621585
transform 1 0 20700 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_225
timestamp 1623621585
transform 1 0 21804 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_237
timestamp 1623621585
transform 1 0 22908 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_249
timestamp 1623621585
transform 1 0 24012 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1562
timestamp 1623621585
transform 1 0 24748 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_258
timestamp 1623621585
transform 1 0 24840 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_270
timestamp 1623621585
transform 1 0 25944 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_282
timestamp 1623621585
transform 1 0 27048 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_294
timestamp 1623621585
transform 1 0 28152 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_306
timestamp 1623621585
transform 1 0 29256 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1563
timestamp 1623621585
transform 1 0 29992 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_315
timestamp 1623621585
transform 1 0 30084 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_327
timestamp 1623621585
transform 1 0 31188 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_339
timestamp 1623621585
transform 1 0 32292 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_351
timestamp 1623621585
transform 1 0 33396 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1564
timestamp 1623621585
transform 1 0 35236 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_161_363
timestamp 1623621585
transform 1 0 34500 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_161_372
timestamp 1623621585
transform 1 0 35328 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input286
timestamp 1623621585
transform 1 0 37260 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_161_384
timestamp 1623621585
transform 1 0 36432 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_161_392
timestamp 1623621585
transform 1 0 37168 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_323
timestamp 1623621585
transform -1 0 38824 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input284
timestamp 1623621585
transform 1 0 37904 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_161_396
timestamp 1623621585
transform 1 0 37536 0 1 89760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_161_403
timestamp 1623621585
transform 1 0 38180 0 1 89760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _754_
timestamp 1623621585
transform 1 0 1380 0 -1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_324
timestamp 1623621585
transform 1 0 1104 0 -1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input423
timestamp 1623621585
transform 1 0 2024 0 -1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_162_6
timestamp 1623621585
transform 1 0 1656 0 -1 90848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_162_13
timestamp 1623621585
transform 1 0 2300 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_25
timestamp 1623621585
transform 1 0 3404 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_37
timestamp 1623621585
transform 1 0 4508 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1565
timestamp 1623621585
transform 1 0 6348 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_162_49
timestamp 1623621585
transform 1 0 5612 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_162_58
timestamp 1623621585
transform 1 0 6440 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_70
timestamp 1623621585
transform 1 0 7544 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_82
timestamp 1623621585
transform 1 0 8648 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_94
timestamp 1623621585
transform 1 0 9752 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1566
timestamp 1623621585
transform 1 0 11592 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_162_106
timestamp 1623621585
transform 1 0 10856 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_162_115
timestamp 1623621585
transform 1 0 11684 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_127
timestamp 1623621585
transform 1 0 12788 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_139
timestamp 1623621585
transform 1 0 13892 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_151
timestamp 1623621585
transform 1 0 14996 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_162_163
timestamp 1623621585
transform 1 0 16100 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1567
timestamp 1623621585
transform 1 0 16836 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_172
timestamp 1623621585
transform 1 0 16928 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_184
timestamp 1623621585
transform 1 0 18032 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_196
timestamp 1623621585
transform 1 0 19136 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_208
timestamp 1623621585
transform 1 0 20240 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1568
timestamp 1623621585
transform 1 0 22080 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_162_220
timestamp 1623621585
transform 1 0 21344 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_162_229
timestamp 1623621585
transform 1 0 22172 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_241
timestamp 1623621585
transform 1 0 23276 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_253
timestamp 1623621585
transform 1 0 24380 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_265
timestamp 1623621585
transform 1 0 25484 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1569
timestamp 1623621585
transform 1 0 27324 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_162_277
timestamp 1623621585
transform 1 0 26588 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_162_286
timestamp 1623621585
transform 1 0 27416 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_298
timestamp 1623621585
transform 1 0 28520 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_310
timestamp 1623621585
transform 1 0 29624 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_322
timestamp 1623621585
transform 1 0 30728 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1570
timestamp 1623621585
transform 1 0 32568 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_162_334
timestamp 1623621585
transform 1 0 31832 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_162_343
timestamp 1623621585
transform 1 0 32660 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_355
timestamp 1623621585
transform 1 0 33764 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_367
timestamp 1623621585
transform 1 0 34868 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_379
timestamp 1623621585
transform 1 0 35972 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_162_391
timestamp 1623621585
transform 1 0 37076 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_325
timestamp 1623621585
transform -1 0 38824 0 -1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1571
timestamp 1623621585
transform 1 0 37812 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_162_400
timestamp 1623621585
transform 1 0 37904 0 -1 90848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_406
timestamp 1623621585
transform 1 0 38456 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _710_
timestamp 1623621585
transform 1 0 1380 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_326
timestamp 1623621585
transform 1 0 1104 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_163_6
timestamp 1623621585
transform 1 0 1656 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_163_18
timestamp 1623621585
transform 1 0 2760 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1572
timestamp 1623621585
transform 1 0 3772 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_163_26
timestamp 1623621585
transform 1 0 3496 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_163_30
timestamp 1623621585
transform 1 0 3864 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_42
timestamp 1623621585
transform 1 0 4968 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_54
timestamp 1623621585
transform 1 0 6072 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_66
timestamp 1623621585
transform 1 0 7176 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_163_78
timestamp 1623621585
transform 1 0 8280 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1573
timestamp 1623621585
transform 1 0 9016 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_87
timestamp 1623621585
transform 1 0 9108 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_99
timestamp 1623621585
transform 1 0 10212 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_111
timestamp 1623621585
transform 1 0 11316 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_123
timestamp 1623621585
transform 1 0 12420 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1574
timestamp 1623621585
transform 1 0 14260 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_163_135
timestamp 1623621585
transform 1 0 13524 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_163_144
timestamp 1623621585
transform 1 0 14352 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_156
timestamp 1623621585
transform 1 0 15456 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_168
timestamp 1623621585
transform 1 0 16560 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_180
timestamp 1623621585
transform 1 0 17664 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1575
timestamp 1623621585
transform 1 0 19504 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_163_192
timestamp 1623621585
transform 1 0 18768 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_163_201
timestamp 1623621585
transform 1 0 19596 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_213
timestamp 1623621585
transform 1 0 20700 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_225
timestamp 1623621585
transform 1 0 21804 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_237
timestamp 1623621585
transform 1 0 22908 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_163_249
timestamp 1623621585
transform 1 0 24012 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1576
timestamp 1623621585
transform 1 0 24748 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_258
timestamp 1623621585
transform 1 0 24840 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_270
timestamp 1623621585
transform 1 0 25944 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_282
timestamp 1623621585
transform 1 0 27048 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_294
timestamp 1623621585
transform 1 0 28152 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_163_306
timestamp 1623621585
transform 1 0 29256 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1577
timestamp 1623621585
transform 1 0 29992 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_315
timestamp 1623621585
transform 1 0 30084 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_327
timestamp 1623621585
transform 1 0 31188 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_339
timestamp 1623621585
transform 1 0 32292 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_351
timestamp 1623621585
transform 1 0 33396 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1578
timestamp 1623621585
transform 1 0 35236 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_163_363
timestamp 1623621585
transform 1 0 34500 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_163_372
timestamp 1623621585
transform 1 0 35328 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input257
timestamp 1623621585
transform 1 0 37260 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_163_384
timestamp 1623621585
transform 1 0 36432 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_163_392
timestamp 1623621585
transform 1 0 37168 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_327
timestamp 1623621585
transform -1 0 38824 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input256
timestamp 1623621585
transform 1 0 37904 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_163_396
timestamp 1623621585
transform 1 0 37536 0 1 90848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_163_403
timestamp 1623621585
transform 1 0 38180 0 1 90848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_328
timestamp 1623621585
transform 1 0 1104 0 -1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input424
timestamp 1623621585
transform 1 0 1380 0 -1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_164_6
timestamp 1623621585
transform 1 0 1656 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_18
timestamp 1623621585
transform 1 0 2760 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_30
timestamp 1623621585
transform 1 0 3864 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1579
timestamp 1623621585
transform 1 0 6348 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_42
timestamp 1623621585
transform 1 0 4968 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_164_54
timestamp 1623621585
transform 1 0 6072 0 -1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_164_58
timestamp 1623621585
transform 1 0 6440 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_70
timestamp 1623621585
transform 1 0 7544 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_82
timestamp 1623621585
transform 1 0 8648 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_94
timestamp 1623621585
transform 1 0 9752 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1580
timestamp 1623621585
transform 1 0 11592 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_164_106
timestamp 1623621585
transform 1 0 10856 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_164_115
timestamp 1623621585
transform 1 0 11684 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_127
timestamp 1623621585
transform 1 0 12788 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_139
timestamp 1623621585
transform 1 0 13892 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_151
timestamp 1623621585
transform 1 0 14996 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_164_163
timestamp 1623621585
transform 1 0 16100 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1581
timestamp 1623621585
transform 1 0 16836 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_172
timestamp 1623621585
transform 1 0 16928 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_184
timestamp 1623621585
transform 1 0 18032 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_196
timestamp 1623621585
transform 1 0 19136 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_208
timestamp 1623621585
transform 1 0 20240 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1582
timestamp 1623621585
transform 1 0 22080 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_164_220
timestamp 1623621585
transform 1 0 21344 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_164_229
timestamp 1623621585
transform 1 0 22172 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_241
timestamp 1623621585
transform 1 0 23276 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_253
timestamp 1623621585
transform 1 0 24380 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_265
timestamp 1623621585
transform 1 0 25484 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1583
timestamp 1623621585
transform 1 0 27324 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_164_277
timestamp 1623621585
transform 1 0 26588 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_164_286
timestamp 1623621585
transform 1 0 27416 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_298
timestamp 1623621585
transform 1 0 28520 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_310
timestamp 1623621585
transform 1 0 29624 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_322
timestamp 1623621585
transform 1 0 30728 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1584
timestamp 1623621585
transform 1 0 32568 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_164_334
timestamp 1623621585
transform 1 0 31832 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_164_343
timestamp 1623621585
transform 1 0 32660 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_355
timestamp 1623621585
transform 1 0 33764 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_367
timestamp 1623621585
transform 1 0 34868 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input259
timestamp 1623621585
transform 1 0 37168 0 -1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_164_379
timestamp 1623621585
transform 1 0 35972 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_164_391
timestamp 1623621585
transform 1 0 37076 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_164_395
timestamp 1623621585
transform 1 0 37444 0 -1 91936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_329
timestamp 1623621585
transform -1 0 38824 0 -1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1585
timestamp 1623621585
transform 1 0 37812 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_164_400
timestamp 1623621585
transform 1 0 37904 0 -1 91936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_406
timestamp 1623621585
transform 1 0 38456 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _723_
timestamp 1623621585
transform 1 0 2116 0 -1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_330
timestamp 1623621585
transform 1 0 1104 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_332
timestamp 1623621585
transform 1 0 1104 0 -1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input425
timestamp 1623621585
transform 1 0 1380 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_165_6
timestamp 1623621585
transform 1 0 1656 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_18
timestamp 1623621585
transform 1 0 2760 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_166_3
timestamp 1623621585
transform 1 0 1380 0 -1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_14
timestamp 1623621585
transform 1 0 2392 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1586
timestamp 1623621585
transform 1 0 3772 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_165_26
timestamp 1623621585
transform 1 0 3496 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_165_30
timestamp 1623621585
transform 1 0 3864 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_26
timestamp 1623621585
transform 1 0 3496 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_38
timestamp 1623621585
transform 1 0 4600 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1593
timestamp 1623621585
transform 1 0 6348 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_42
timestamp 1623621585
transform 1 0 4968 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_54
timestamp 1623621585
transform 1 0 6072 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_50
timestamp 1623621585
transform 1 0 5704 0 -1 93024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_56
timestamp 1623621585
transform 1 0 6256 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_58
timestamp 1623621585
transform 1 0 6440 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_66
timestamp 1623621585
transform 1 0 7176 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_78
timestamp 1623621585
transform 1 0 8280 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_70
timestamp 1623621585
transform 1 0 7544 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_82
timestamp 1623621585
transform 1 0 8648 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1587
timestamp 1623621585
transform 1 0 9016 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_87
timestamp 1623621585
transform 1 0 9108 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_99
timestamp 1623621585
transform 1 0 10212 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_94
timestamp 1623621585
transform 1 0 9752 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1594
timestamp 1623621585
transform 1 0 11592 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_111
timestamp 1623621585
transform 1 0 11316 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_123
timestamp 1623621585
transform 1 0 12420 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_106
timestamp 1623621585
transform 1 0 10856 0 -1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_115
timestamp 1623621585
transform 1 0 11684 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1588
timestamp 1623621585
transform 1 0 14260 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_165_135
timestamp 1623621585
transform 1 0 13524 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_165_144
timestamp 1623621585
transform 1 0 14352 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_127
timestamp 1623621585
transform 1 0 12788 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_139
timestamp 1623621585
transform 1 0 13892 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_156
timestamp 1623621585
transform 1 0 15456 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_151
timestamp 1623621585
transform 1 0 14996 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_163
timestamp 1623621585
transform 1 0 16100 0 -1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1595
timestamp 1623621585
transform 1 0 16836 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_168
timestamp 1623621585
transform 1 0 16560 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_180
timestamp 1623621585
transform 1 0 17664 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_172
timestamp 1623621585
transform 1 0 16928 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_184
timestamp 1623621585
transform 1 0 18032 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1589
timestamp 1623621585
transform 1 0 19504 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_165_192
timestamp 1623621585
transform 1 0 18768 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_165_201
timestamp 1623621585
transform 1 0 19596 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_196
timestamp 1623621585
transform 1 0 19136 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_208
timestamp 1623621585
transform 1 0 20240 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1596
timestamp 1623621585
transform 1 0 22080 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_213
timestamp 1623621585
transform 1 0 20700 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_225
timestamp 1623621585
transform 1 0 21804 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_220
timestamp 1623621585
transform 1 0 21344 0 -1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_229
timestamp 1623621585
transform 1 0 22172 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_237
timestamp 1623621585
transform 1 0 22908 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_249
timestamp 1623621585
transform 1 0 24012 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_241
timestamp 1623621585
transform 1 0 23276 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1590
timestamp 1623621585
transform 1 0 24748 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_258
timestamp 1623621585
transform 1 0 24840 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_270
timestamp 1623621585
transform 1 0 25944 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_253
timestamp 1623621585
transform 1 0 24380 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_265
timestamp 1623621585
transform 1 0 25484 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1597
timestamp 1623621585
transform 1 0 27324 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_282
timestamp 1623621585
transform 1 0 27048 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_277
timestamp 1623621585
transform 1 0 26588 0 -1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_286
timestamp 1623621585
transform 1 0 27416 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_294
timestamp 1623621585
transform 1 0 28152 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_306
timestamp 1623621585
transform 1 0 29256 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_298
timestamp 1623621585
transform 1 0 28520 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_310
timestamp 1623621585
transform 1 0 29624 0 -1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _739_
timestamp 1623621585
transform 1 0 30452 0 -1 93024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1591
timestamp 1623621585
transform 1 0 29992 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_315
timestamp 1623621585
transform 1 0 30084 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_327
timestamp 1623621585
transform 1 0 31188 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_166_318
timestamp 1623621585
transform 1 0 30360 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_323
timestamp 1623621585
transform 1 0 30820 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1598
timestamp 1623621585
transform 1 0 32568 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_339
timestamp 1623621585
transform 1 0 32292 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_351
timestamp 1623621585
transform 1 0 33396 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_335
timestamp 1623621585
transform 1 0 31924 0 -1 93024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_341
timestamp 1623621585
transform 1 0 32476 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_343
timestamp 1623621585
transform 1 0 32660 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1592
timestamp 1623621585
transform 1 0 35236 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_165_363
timestamp 1623621585
transform 1 0 34500 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_165_372
timestamp 1623621585
transform 1 0 35328 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_355
timestamp 1623621585
transform 1 0 33764 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_367
timestamp 1623621585
transform 1 0 34868 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input260
timestamp 1623621585
transform 1 0 37260 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_165_384
timestamp 1623621585
transform 1 0 36432 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_165_392
timestamp 1623621585
transform 1 0 37168 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_379
timestamp 1623621585
transform 1 0 35972 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_391
timestamp 1623621585
transform 1 0 37076 0 -1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_331
timestamp 1623621585
transform -1 0 38824 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_333
timestamp 1623621585
transform -1 0 38824 0 -1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1599
timestamp 1623621585
transform 1 0 37812 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input258
timestamp 1623621585
transform 1 0 37904 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_165_396
timestamp 1623621585
transform 1 0 37536 0 1 91936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_165_403
timestamp 1623621585
transform 1 0 38180 0 1 91936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_166_400
timestamp 1623621585
transform 1 0 37904 0 -1 93024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_406
timestamp 1623621585
transform 1 0 38456 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_334
timestamp 1623621585
transform 1 0 1104 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input427
timestamp 1623621585
transform 1 0 1380 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_167_6
timestamp 1623621585
transform 1 0 1656 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_167_18
timestamp 1623621585
transform 1 0 2760 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1600
timestamp 1623621585
transform 1 0 3772 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_167_26
timestamp 1623621585
transform 1 0 3496 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_167_30
timestamp 1623621585
transform 1 0 3864 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_42
timestamp 1623621585
transform 1 0 4968 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_54
timestamp 1623621585
transform 1 0 6072 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_66
timestamp 1623621585
transform 1 0 7176 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_167_78
timestamp 1623621585
transform 1 0 8280 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1601
timestamp 1623621585
transform 1 0 9016 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_87
timestamp 1623621585
transform 1 0 9108 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_99
timestamp 1623621585
transform 1 0 10212 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_111
timestamp 1623621585
transform 1 0 11316 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_123
timestamp 1623621585
transform 1 0 12420 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1602
timestamp 1623621585
transform 1 0 14260 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_167_135
timestamp 1623621585
transform 1 0 13524 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_167_144
timestamp 1623621585
transform 1 0 14352 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_156
timestamp 1623621585
transform 1 0 15456 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_168
timestamp 1623621585
transform 1 0 16560 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_180
timestamp 1623621585
transform 1 0 17664 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1603
timestamp 1623621585
transform 1 0 19504 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_167_192
timestamp 1623621585
transform 1 0 18768 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_167_201
timestamp 1623621585
transform 1 0 19596 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_213
timestamp 1623621585
transform 1 0 20700 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_225
timestamp 1623621585
transform 1 0 21804 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_237
timestamp 1623621585
transform 1 0 22908 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_167_249
timestamp 1623621585
transform 1 0 24012 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1604
timestamp 1623621585
transform 1 0 24748 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_258
timestamp 1623621585
transform 1 0 24840 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_270
timestamp 1623621585
transform 1 0 25944 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_282
timestamp 1623621585
transform 1 0 27048 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_294
timestamp 1623621585
transform 1 0 28152 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_167_306
timestamp 1623621585
transform 1 0 29256 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1605
timestamp 1623621585
transform 1 0 29992 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_315
timestamp 1623621585
transform 1 0 30084 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_327
timestamp 1623621585
transform 1 0 31188 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_339
timestamp 1623621585
transform 1 0 32292 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_351
timestamp 1623621585
transform 1 0 33396 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1606
timestamp 1623621585
transform 1 0 35236 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_167_363
timestamp 1623621585
transform 1 0 34500 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_167_372
timestamp 1623621585
transform 1 0 35328 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input262
timestamp 1623621585
transform 1 0 37260 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_167_384
timestamp 1623621585
transform 1 0 36432 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_167_392
timestamp 1623621585
transform 1 0 37168 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_335
timestamp 1623621585
transform -1 0 38824 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input261
timestamp 1623621585
transform 1 0 37904 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_167_396
timestamp 1623621585
transform 1 0 37536 0 1 93024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_167_403
timestamp 1623621585
transform 1 0 38180 0 1 93024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_336
timestamp 1623621585
transform 1 0 1104 0 -1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input428
timestamp 1623621585
transform 1 0 1380 0 -1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_168_6
timestamp 1623621585
transform 1 0 1656 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_18
timestamp 1623621585
transform 1 0 2760 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_30
timestamp 1623621585
transform 1 0 3864 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1607
timestamp 1623621585
transform 1 0 6348 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_42
timestamp 1623621585
transform 1 0 4968 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_168_54
timestamp 1623621585
transform 1 0 6072 0 -1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_168_58
timestamp 1623621585
transform 1 0 6440 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_70
timestamp 1623621585
transform 1 0 7544 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_82
timestamp 1623621585
transform 1 0 8648 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_94
timestamp 1623621585
transform 1 0 9752 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1608
timestamp 1623621585
transform 1 0 11592 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_168_106
timestamp 1623621585
transform 1 0 10856 0 -1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_168_115
timestamp 1623621585
transform 1 0 11684 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_127
timestamp 1623621585
transform 1 0 12788 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_139
timestamp 1623621585
transform 1 0 13892 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_151
timestamp 1623621585
transform 1 0 14996 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_168_163
timestamp 1623621585
transform 1 0 16100 0 -1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1609
timestamp 1623621585
transform 1 0 16836 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_172
timestamp 1623621585
transform 1 0 16928 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_184
timestamp 1623621585
transform 1 0 18032 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_196
timestamp 1623621585
transform 1 0 19136 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_208
timestamp 1623621585
transform 1 0 20240 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1610
timestamp 1623621585
transform 1 0 22080 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_168_220
timestamp 1623621585
transform 1 0 21344 0 -1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_168_229
timestamp 1623621585
transform 1 0 22172 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_241
timestamp 1623621585
transform 1 0 23276 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_253
timestamp 1623621585
transform 1 0 24380 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_265
timestamp 1623621585
transform 1 0 25484 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1611
timestamp 1623621585
transform 1 0 27324 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_168_277
timestamp 1623621585
transform 1 0 26588 0 -1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_168_286
timestamp 1623621585
transform 1 0 27416 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_298
timestamp 1623621585
transform 1 0 28520 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_310
timestamp 1623621585
transform 1 0 29624 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_322
timestamp 1623621585
transform 1 0 30728 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1612
timestamp 1623621585
transform 1 0 32568 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_168_334
timestamp 1623621585
transform 1 0 31832 0 -1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_168_343
timestamp 1623621585
transform 1 0 32660 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_355
timestamp 1623621585
transform 1 0 33764 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_367
timestamp 1623621585
transform 1 0 34868 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input263
timestamp 1623621585
transform 1 0 37168 0 -1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_168_379
timestamp 1623621585
transform 1 0 35972 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_168_391
timestamp 1623621585
transform 1 0 37076 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_168_395
timestamp 1623621585
transform 1 0 37444 0 -1 94112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_337
timestamp 1623621585
transform -1 0 38824 0 -1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1613
timestamp 1623621585
transform 1 0 37812 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_168_400
timestamp 1623621585
transform 1 0 37904 0 -1 94112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_406
timestamp 1623621585
transform 1 0 38456 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _712_
timestamp 1623621585
transform 1 0 2668 0 1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_338
timestamp 1623621585
transform 1 0 1104 0 1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input429
timestamp 1623621585
transform 1 0 1380 0 1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_169_6
timestamp 1623621585
transform 1 0 1656 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_169_14
timestamp 1623621585
transform 1 0 2392 0 1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_169_20
timestamp 1623621585
transform 1 0 2944 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1614
timestamp 1623621585
transform 1 0 3772 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_169_28
timestamp 1623621585
transform 1 0 3680 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_30
timestamp 1623621585
transform 1 0 3864 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_42
timestamp 1623621585
transform 1 0 4968 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_54
timestamp 1623621585
transform 1 0 6072 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_66
timestamp 1623621585
transform 1 0 7176 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_169_78
timestamp 1623621585
transform 1 0 8280 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1615
timestamp 1623621585
transform 1 0 9016 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_87
timestamp 1623621585
transform 1 0 9108 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_99
timestamp 1623621585
transform 1 0 10212 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_111
timestamp 1623621585
transform 1 0 11316 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_123
timestamp 1623621585
transform 1 0 12420 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1616
timestamp 1623621585
transform 1 0 14260 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_169_135
timestamp 1623621585
transform 1 0 13524 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_169_144
timestamp 1623621585
transform 1 0 14352 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_156
timestamp 1623621585
transform 1 0 15456 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_168
timestamp 1623621585
transform 1 0 16560 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_180
timestamp 1623621585
transform 1 0 17664 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1617
timestamp 1623621585
transform 1 0 19504 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_169_192
timestamp 1623621585
transform 1 0 18768 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_169_201
timestamp 1623621585
transform 1 0 19596 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_213
timestamp 1623621585
transform 1 0 20700 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_225
timestamp 1623621585
transform 1 0 21804 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_237
timestamp 1623621585
transform 1 0 22908 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_169_249
timestamp 1623621585
transform 1 0 24012 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1618
timestamp 1623621585
transform 1 0 24748 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_258
timestamp 1623621585
transform 1 0 24840 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_270
timestamp 1623621585
transform 1 0 25944 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_282
timestamp 1623621585
transform 1 0 27048 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_294
timestamp 1623621585
transform 1 0 28152 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_169_306
timestamp 1623621585
transform 1 0 29256 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1619
timestamp 1623621585
transform 1 0 29992 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_315
timestamp 1623621585
transform 1 0 30084 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_327
timestamp 1623621585
transform 1 0 31188 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_339
timestamp 1623621585
transform 1 0 32292 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_351
timestamp 1623621585
transform 1 0 33396 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1620
timestamp 1623621585
transform 1 0 35236 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_169_363
timestamp 1623621585
transform 1 0 34500 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_169_372
timestamp 1623621585
transform 1 0 35328 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input265
timestamp 1623621585
transform 1 0 37076 0 1 94112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_169_384
timestamp 1623621585
transform 1 0 36432 0 1 94112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_390
timestamp 1623621585
transform 1 0 36984 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_169_395
timestamp 1623621585
transform 1 0 37444 0 1 94112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_339
timestamp 1623621585
transform -1 0 38824 0 1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input264
timestamp 1623621585
transform 1 0 37812 0 1 94112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_169_403
timestamp 1623621585
transform 1 0 38180 0 1 94112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_340
timestamp 1623621585
transform 1 0 1104 0 -1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_170_3
timestamp 1623621585
transform 1 0 1380 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_15
timestamp 1623621585
transform 1 0 2484 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_27
timestamp 1623621585
transform 1 0 3588 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_39
timestamp 1623621585
transform 1 0 4692 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1621
timestamp 1623621585
transform 1 0 6348 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_170_51
timestamp 1623621585
transform 1 0 5796 0 -1 95200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_170_58
timestamp 1623621585
transform 1 0 6440 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_70
timestamp 1623621585
transform 1 0 7544 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_82
timestamp 1623621585
transform 1 0 8648 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_94
timestamp 1623621585
transform 1 0 9752 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1622
timestamp 1623621585
transform 1 0 11592 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_170_106
timestamp 1623621585
transform 1 0 10856 0 -1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_170_115
timestamp 1623621585
transform 1 0 11684 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_127
timestamp 1623621585
transform 1 0 12788 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_139
timestamp 1623621585
transform 1 0 13892 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_151
timestamp 1623621585
transform 1 0 14996 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_170_163
timestamp 1623621585
transform 1 0 16100 0 -1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1623
timestamp 1623621585
transform 1 0 16836 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_172
timestamp 1623621585
transform 1 0 16928 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_184
timestamp 1623621585
transform 1 0 18032 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_196
timestamp 1623621585
transform 1 0 19136 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_208
timestamp 1623621585
transform 1 0 20240 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1624
timestamp 1623621585
transform 1 0 22080 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_170_220
timestamp 1623621585
transform 1 0 21344 0 -1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_170_229
timestamp 1623621585
transform 1 0 22172 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_241
timestamp 1623621585
transform 1 0 23276 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_253
timestamp 1623621585
transform 1 0 24380 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_265
timestamp 1623621585
transform 1 0 25484 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1625
timestamp 1623621585
transform 1 0 27324 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_170_277
timestamp 1623621585
transform 1 0 26588 0 -1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_170_286
timestamp 1623621585
transform 1 0 27416 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_298
timestamp 1623621585
transform 1 0 28520 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_310
timestamp 1623621585
transform 1 0 29624 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_322
timestamp 1623621585
transform 1 0 30728 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1626
timestamp 1623621585
transform 1 0 32568 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_170_334
timestamp 1623621585
transform 1 0 31832 0 -1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_170_343
timestamp 1623621585
transform 1 0 32660 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_355
timestamp 1623621585
transform 1 0 33764 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_367
timestamp 1623621585
transform 1 0 34868 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input267
timestamp 1623621585
transform 1 0 37076 0 -1 95200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_170_379
timestamp 1623621585
transform 1 0 35972 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_170_395
timestamp 1623621585
transform 1 0 37444 0 -1 95200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_341
timestamp 1623621585
transform -1 0 38824 0 -1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1627
timestamp 1623621585
transform 1 0 37812 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_170_400
timestamp 1623621585
transform 1 0 37904 0 -1 95200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_406
timestamp 1623621585
transform 1 0 38456 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _724_
timestamp 1623621585
transform 1 0 2760 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_342
timestamp 1623621585
transform 1 0 1104 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_344
timestamp 1623621585
transform 1 0 1104 0 -1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input430
timestamp 1623621585
transform 1 0 1380 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input431
timestamp 1623621585
transform 1 0 1380 0 -1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_171_6
timestamp 1623621585
transform 1 0 1656 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_6
timestamp 1623621585
transform 1 0 1656 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_18
timestamp 1623621585
transform 1 0 2760 0 -1 96288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _713_
timestamp 1623621585
transform 1 0 3312 0 -1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1628
timestamp 1623621585
transform 1 0 3772 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_21
timestamp 1623621585
transform 1 0 3036 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_171_30
timestamp 1623621585
transform 1 0 3864 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_27
timestamp 1623621585
transform 1 0 3588 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_39
timestamp 1623621585
transform 1 0 4692 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1635
timestamp 1623621585
transform 1 0 6348 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_42
timestamp 1623621585
transform 1 0 4968 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_54
timestamp 1623621585
transform 1 0 6072 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_51
timestamp 1623621585
transform 1 0 5796 0 -1 96288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_172_58
timestamp 1623621585
transform 1 0 6440 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_66
timestamp 1623621585
transform 1 0 7176 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_171_78
timestamp 1623621585
transform 1 0 8280 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_70
timestamp 1623621585
transform 1 0 7544 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_82
timestamp 1623621585
transform 1 0 8648 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1629
timestamp 1623621585
transform 1 0 9016 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_87
timestamp 1623621585
transform 1 0 9108 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_99
timestamp 1623621585
transform 1 0 10212 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_94
timestamp 1623621585
transform 1 0 9752 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1636
timestamp 1623621585
transform 1 0 11592 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_111
timestamp 1623621585
transform 1 0 11316 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_123
timestamp 1623621585
transform 1 0 12420 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_106
timestamp 1623621585
transform 1 0 10856 0 -1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_115
timestamp 1623621585
transform 1 0 11684 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1630
timestamp 1623621585
transform 1 0 14260 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_135
timestamp 1623621585
transform 1 0 13524 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_171_144
timestamp 1623621585
transform 1 0 14352 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_127
timestamp 1623621585
transform 1 0 12788 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_139
timestamp 1623621585
transform 1 0 13892 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_156
timestamp 1623621585
transform 1 0 15456 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_151
timestamp 1623621585
transform 1 0 14996 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_163
timestamp 1623621585
transform 1 0 16100 0 -1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1637
timestamp 1623621585
transform 1 0 16836 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_168
timestamp 1623621585
transform 1 0 16560 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_180
timestamp 1623621585
transform 1 0 17664 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_172
timestamp 1623621585
transform 1 0 16928 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_184
timestamp 1623621585
transform 1 0 18032 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1631
timestamp 1623621585
transform 1 0 19504 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_192
timestamp 1623621585
transform 1 0 18768 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_171_201
timestamp 1623621585
transform 1 0 19596 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_196
timestamp 1623621585
transform 1 0 19136 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_208
timestamp 1623621585
transform 1 0 20240 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1638
timestamp 1623621585
transform 1 0 22080 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_213
timestamp 1623621585
transform 1 0 20700 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_225
timestamp 1623621585
transform 1 0 21804 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_220
timestamp 1623621585
transform 1 0 21344 0 -1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_229
timestamp 1623621585
transform 1 0 22172 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_237
timestamp 1623621585
transform 1 0 22908 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_171_249
timestamp 1623621585
transform 1 0 24012 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_241
timestamp 1623621585
transform 1 0 23276 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1632
timestamp 1623621585
transform 1 0 24748 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_258
timestamp 1623621585
transform 1 0 24840 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_270
timestamp 1623621585
transform 1 0 25944 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_253
timestamp 1623621585
transform 1 0 24380 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_265
timestamp 1623621585
transform 1 0 25484 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1639
timestamp 1623621585
transform 1 0 27324 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_282
timestamp 1623621585
transform 1 0 27048 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_277
timestamp 1623621585
transform 1 0 26588 0 -1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_286
timestamp 1623621585
transform 1 0 27416 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_294
timestamp 1623621585
transform 1 0 28152 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_171_306
timestamp 1623621585
transform 1 0 29256 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_298
timestamp 1623621585
transform 1 0 28520 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_310
timestamp 1623621585
transform 1 0 29624 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1633
timestamp 1623621585
transform 1 0 29992 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_315
timestamp 1623621585
transform 1 0 30084 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_327
timestamp 1623621585
transform 1 0 31188 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_322
timestamp 1623621585
transform 1 0 30728 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1640
timestamp 1623621585
transform 1 0 32568 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_339
timestamp 1623621585
transform 1 0 32292 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_351
timestamp 1623621585
transform 1 0 33396 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_334
timestamp 1623621585
transform 1 0 31832 0 -1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_343
timestamp 1623621585
transform 1 0 32660 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1634
timestamp 1623621585
transform 1 0 35236 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_363
timestamp 1623621585
transform 1 0 34500 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_171_372
timestamp 1623621585
transform 1 0 35328 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_355
timestamp 1623621585
transform 1 0 33764 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_367
timestamp 1623621585
transform 1 0 34868 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input269
timestamp 1623621585
transform 1 0 37076 0 -1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_171_384
timestamp 1623621585
transform 1 0 36432 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_379
timestamp 1623621585
transform 1 0 35972 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_172_395
timestamp 1623621585
transform 1 0 37444 0 -1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_343
timestamp 1623621585
transform -1 0 38824 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_345
timestamp 1623621585
transform -1 0 38824 0 -1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1641
timestamp 1623621585
transform 1 0 37812 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input268
timestamp 1623621585
transform 1 0 37812 0 1 95200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_171_396
timestamp 1623621585
transform 1 0 37536 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_171_403
timestamp 1623621585
transform 1 0 38180 0 1 95200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_172_400
timestamp 1623621585
transform 1 0 37904 0 -1 96288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_406
timestamp 1623621585
transform 1 0 38456 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_346
timestamp 1623621585
transform 1 0 1104 0 1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_173_3
timestamp 1623621585
transform 1 0 1380 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_15
timestamp 1623621585
transform 1 0 2484 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1642
timestamp 1623621585
transform 1 0 3772 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_173_27
timestamp 1623621585
transform 1 0 3588 0 1 96288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_173_30
timestamp 1623621585
transform 1 0 3864 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_42
timestamp 1623621585
transform 1 0 4968 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_54
timestamp 1623621585
transform 1 0 6072 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_66
timestamp 1623621585
transform 1 0 7176 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_173_78
timestamp 1623621585
transform 1 0 8280 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1643
timestamp 1623621585
transform 1 0 9016 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_87
timestamp 1623621585
transform 1 0 9108 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_99
timestamp 1623621585
transform 1 0 10212 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_111
timestamp 1623621585
transform 1 0 11316 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_123
timestamp 1623621585
transform 1 0 12420 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1644
timestamp 1623621585
transform 1 0 14260 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_173_135
timestamp 1623621585
transform 1 0 13524 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_173_144
timestamp 1623621585
transform 1 0 14352 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_156
timestamp 1623621585
transform 1 0 15456 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_168
timestamp 1623621585
transform 1 0 16560 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_180
timestamp 1623621585
transform 1 0 17664 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1645
timestamp 1623621585
transform 1 0 19504 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_173_192
timestamp 1623621585
transform 1 0 18768 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_173_201
timestamp 1623621585
transform 1 0 19596 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_213
timestamp 1623621585
transform 1 0 20700 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_225
timestamp 1623621585
transform 1 0 21804 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_237
timestamp 1623621585
transform 1 0 22908 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_173_249
timestamp 1623621585
transform 1 0 24012 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1646
timestamp 1623621585
transform 1 0 24748 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_258
timestamp 1623621585
transform 1 0 24840 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_270
timestamp 1623621585
transform 1 0 25944 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_282
timestamp 1623621585
transform 1 0 27048 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_294
timestamp 1623621585
transform 1 0 28152 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_173_306
timestamp 1623621585
transform 1 0 29256 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1647
timestamp 1623621585
transform 1 0 29992 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_315
timestamp 1623621585
transform 1 0 30084 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_327
timestamp 1623621585
transform 1 0 31188 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_339
timestamp 1623621585
transform 1 0 32292 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_351
timestamp 1623621585
transform 1 0 33396 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1648
timestamp 1623621585
transform 1 0 35236 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_173_363
timestamp 1623621585
transform 1 0 34500 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_173_372
timestamp 1623621585
transform 1 0 35328 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  input271
timestamp 1623621585
transform 1 0 37076 0 1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_173_384
timestamp 1623621585
transform 1 0 36432 0 1 96288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_390
timestamp 1623621585
transform 1 0 36984 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_173_395
timestamp 1623621585
transform 1 0 37444 0 1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_347
timestamp 1623621585
transform -1 0 38824 0 1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input270
timestamp 1623621585
transform 1 0 37812 0 1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_173_403
timestamp 1623621585
transform 1 0 38180 0 1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_348
timestamp 1623621585
transform 1 0 1104 0 -1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input432
timestamp 1623621585
transform 1 0 1380 0 -1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_174_6
timestamp 1623621585
transform 1 0 1656 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_18
timestamp 1623621585
transform 1 0 2760 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_30
timestamp 1623621585
transform 1 0 3864 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1649
timestamp 1623621585
transform 1 0 6348 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_42
timestamp 1623621585
transform 1 0 4968 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_54
timestamp 1623621585
transform 1 0 6072 0 -1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_174_58
timestamp 1623621585
transform 1 0 6440 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_70
timestamp 1623621585
transform 1 0 7544 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_82
timestamp 1623621585
transform 1 0 8648 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_94
timestamp 1623621585
transform 1 0 9752 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1650
timestamp 1623621585
transform 1 0 11592 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_174_106
timestamp 1623621585
transform 1 0 10856 0 -1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_174_115
timestamp 1623621585
transform 1 0 11684 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_127
timestamp 1623621585
transform 1 0 12788 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_139
timestamp 1623621585
transform 1 0 13892 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_151
timestamp 1623621585
transform 1 0 14996 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_174_163
timestamp 1623621585
transform 1 0 16100 0 -1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1651
timestamp 1623621585
transform 1 0 16836 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_172
timestamp 1623621585
transform 1 0 16928 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_184
timestamp 1623621585
transform 1 0 18032 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_196
timestamp 1623621585
transform 1 0 19136 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_208
timestamp 1623621585
transform 1 0 20240 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1652
timestamp 1623621585
transform 1 0 22080 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_174_220
timestamp 1623621585
transform 1 0 21344 0 -1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_174_229
timestamp 1623621585
transform 1 0 22172 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_241
timestamp 1623621585
transform 1 0 23276 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_253
timestamp 1623621585
transform 1 0 24380 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_265
timestamp 1623621585
transform 1 0 25484 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1653
timestamp 1623621585
transform 1 0 27324 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_174_277
timestamp 1623621585
transform 1 0 26588 0 -1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_174_286
timestamp 1623621585
transform 1 0 27416 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_298
timestamp 1623621585
transform 1 0 28520 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_310
timestamp 1623621585
transform 1 0 29624 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_322
timestamp 1623621585
transform 1 0 30728 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1654
timestamp 1623621585
transform 1 0 32568 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_174_334
timestamp 1623621585
transform 1 0 31832 0 -1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_174_343
timestamp 1623621585
transform 1 0 32660 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_355
timestamp 1623621585
transform 1 0 33764 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_367
timestamp 1623621585
transform 1 0 34868 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  input272
timestamp 1623621585
transform 1 0 37076 0 -1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_174_379
timestamp 1623621585
transform 1 0 35972 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_174_395
timestamp 1623621585
transform 1 0 37444 0 -1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_349
timestamp 1623621585
transform -1 0 38824 0 -1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1655
timestamp 1623621585
transform 1 0 37812 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_174_400
timestamp 1623621585
transform 1 0 37904 0 -1 97376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_406
timestamp 1623621585
transform 1 0 38456 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_350
timestamp 1623621585
transform 1 0 1104 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input433
timestamp 1623621585
transform 1 0 1380 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_175_6
timestamp 1623621585
transform 1 0 1656 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_175_18
timestamp 1623621585
transform 1 0 2760 0 1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _714_
timestamp 1623621585
transform 1 0 4232 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1656
timestamp 1623621585
transform 1 0 3772 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_175_26
timestamp 1623621585
transform 1 0 3496 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_175_30
timestamp 1623621585
transform 1 0 3864 0 1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_175_37
timestamp 1623621585
transform 1 0 4508 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_49
timestamp 1623621585
transform 1 0 5612 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_61
timestamp 1623621585
transform 1 0 6716 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_73
timestamp 1623621585
transform 1 0 7820 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1657
timestamp 1623621585
transform 1 0 9016 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_175_85
timestamp 1623621585
transform 1 0 8924 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_87
timestamp 1623621585
transform 1 0 9108 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_99
timestamp 1623621585
transform 1 0 10212 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_111
timestamp 1623621585
transform 1 0 11316 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_123
timestamp 1623621585
transform 1 0 12420 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1658
timestamp 1623621585
transform 1 0 14260 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_175_135
timestamp 1623621585
transform 1 0 13524 0 1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_175_144
timestamp 1623621585
transform 1 0 14352 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_156
timestamp 1623621585
transform 1 0 15456 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_168
timestamp 1623621585
transform 1 0 16560 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_180
timestamp 1623621585
transform 1 0 17664 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1659
timestamp 1623621585
transform 1 0 19504 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_175_192
timestamp 1623621585
transform 1 0 18768 0 1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_175_201
timestamp 1623621585
transform 1 0 19596 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_213
timestamp 1623621585
transform 1 0 20700 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_225
timestamp 1623621585
transform 1 0 21804 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_237
timestamp 1623621585
transform 1 0 22908 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_175_249
timestamp 1623621585
transform 1 0 24012 0 1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1660
timestamp 1623621585
transform 1 0 24748 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_258
timestamp 1623621585
transform 1 0 24840 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_270
timestamp 1623621585
transform 1 0 25944 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_282
timestamp 1623621585
transform 1 0 27048 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_294
timestamp 1623621585
transform 1 0 28152 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_175_306
timestamp 1623621585
transform 1 0 29256 0 1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1661
timestamp 1623621585
transform 1 0 29992 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_315
timestamp 1623621585
transform 1 0 30084 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_327
timestamp 1623621585
transform 1 0 31188 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_339
timestamp 1623621585
transform 1 0 32292 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_351
timestamp 1623621585
transform 1 0 33396 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1662
timestamp 1623621585
transform 1 0 35236 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_175_363
timestamp 1623621585
transform 1 0 34500 0 1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_175_372
timestamp 1623621585
transform 1 0 35328 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_384
timestamp 1623621585
transform 1 0 36432 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_351
timestamp 1623621585
transform -1 0 38824 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input273
timestamp 1623621585
transform 1 0 37812 0 1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_175_396
timestamp 1623621585
transform 1 0 37536 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_175_403
timestamp 1623621585
transform 1 0 38180 0 1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_352
timestamp 1623621585
transform 1 0 1104 0 -1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_176_3
timestamp 1623621585
transform 1 0 1380 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_15
timestamp 1623621585
transform 1 0 2484 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _716_
timestamp 1623621585
transform 1 0 4876 0 -1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_176_27
timestamp 1623621585
transform 1 0 3588 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_176_39
timestamp 1623621585
transform 1 0 4692 0 -1 98464
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1663
timestamp 1623621585
transform 1 0 6348 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_44
timestamp 1623621585
transform 1 0 5152 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_176_56
timestamp 1623621585
transform 1 0 6256 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_58
timestamp 1623621585
transform 1 0 6440 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_70
timestamp 1623621585
transform 1 0 7544 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_82
timestamp 1623621585
transform 1 0 8648 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_94
timestamp 1623621585
transform 1 0 9752 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1664
timestamp 1623621585
transform 1 0 11592 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_176_106
timestamp 1623621585
transform 1 0 10856 0 -1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_176_115
timestamp 1623621585
transform 1 0 11684 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_127
timestamp 1623621585
transform 1 0 12788 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_139
timestamp 1623621585
transform 1 0 13892 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_151
timestamp 1623621585
transform 1 0 14996 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_176_163
timestamp 1623621585
transform 1 0 16100 0 -1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1665
timestamp 1623621585
transform 1 0 16836 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_172
timestamp 1623621585
transform 1 0 16928 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_184
timestamp 1623621585
transform 1 0 18032 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_196
timestamp 1623621585
transform 1 0 19136 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_208
timestamp 1623621585
transform 1 0 20240 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1666
timestamp 1623621585
transform 1 0 22080 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_176_220
timestamp 1623621585
transform 1 0 21344 0 -1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_176_229
timestamp 1623621585
transform 1 0 22172 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_241
timestamp 1623621585
transform 1 0 23276 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_253
timestamp 1623621585
transform 1 0 24380 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_265
timestamp 1623621585
transform 1 0 25484 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1667
timestamp 1623621585
transform 1 0 27324 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_176_277
timestamp 1623621585
transform 1 0 26588 0 -1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_176_286
timestamp 1623621585
transform 1 0 27416 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_298
timestamp 1623621585
transform 1 0 28520 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_310
timestamp 1623621585
transform 1 0 29624 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_322
timestamp 1623621585
transform 1 0 30728 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1668
timestamp 1623621585
transform 1 0 32568 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_176_334
timestamp 1623621585
transform 1 0 31832 0 -1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_176_343
timestamp 1623621585
transform 1 0 32660 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_355
timestamp 1623621585
transform 1 0 33764 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_367
timestamp 1623621585
transform 1 0 34868 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  input274
timestamp 1623621585
transform 1 0 37076 0 -1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_176_379
timestamp 1623621585
transform 1 0 35972 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_176_395
timestamp 1623621585
transform 1 0 37444 0 -1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_353
timestamp 1623621585
transform -1 0 38824 0 -1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1669
timestamp 1623621585
transform 1 0 37812 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_176_400
timestamp 1623621585
transform 1 0 37904 0 -1 98464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_406
timestamp 1623621585
transform 1 0 38456 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_354
timestamp 1623621585
transform 1 0 1104 0 1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input434
timestamp 1623621585
transform 1 0 1380 0 1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_177_6
timestamp 1623621585
transform 1 0 1656 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_177_18
timestamp 1623621585
transform 1 0 2760 0 1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1670
timestamp 1623621585
transform 1 0 3772 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_177_26
timestamp 1623621585
transform 1 0 3496 0 1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_177_30
timestamp 1623621585
transform 1 0 3864 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_42
timestamp 1623621585
transform 1 0 4968 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_54
timestamp 1623621585
transform 1 0 6072 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_66
timestamp 1623621585
transform 1 0 7176 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_177_78
timestamp 1623621585
transform 1 0 8280 0 1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1671
timestamp 1623621585
transform 1 0 9016 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_87
timestamp 1623621585
transform 1 0 9108 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_99
timestamp 1623621585
transform 1 0 10212 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_111
timestamp 1623621585
transform 1 0 11316 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_123
timestamp 1623621585
transform 1 0 12420 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1672
timestamp 1623621585
transform 1 0 14260 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_177_135
timestamp 1623621585
transform 1 0 13524 0 1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_177_144
timestamp 1623621585
transform 1 0 14352 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_156
timestamp 1623621585
transform 1 0 15456 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_168
timestamp 1623621585
transform 1 0 16560 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_180
timestamp 1623621585
transform 1 0 17664 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1673
timestamp 1623621585
transform 1 0 19504 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_177_192
timestamp 1623621585
transform 1 0 18768 0 1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_177_201
timestamp 1623621585
transform 1 0 19596 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_213
timestamp 1623621585
transform 1 0 20700 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_225
timestamp 1623621585
transform 1 0 21804 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_237
timestamp 1623621585
transform 1 0 22908 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_177_249
timestamp 1623621585
transform 1 0 24012 0 1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1674
timestamp 1623621585
transform 1 0 24748 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_258
timestamp 1623621585
transform 1 0 24840 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_270
timestamp 1623621585
transform 1 0 25944 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_282
timestamp 1623621585
transform 1 0 27048 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_294
timestamp 1623621585
transform 1 0 28152 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_177_306
timestamp 1623621585
transform 1 0 29256 0 1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1675
timestamp 1623621585
transform 1 0 29992 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_315
timestamp 1623621585
transform 1 0 30084 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_327
timestamp 1623621585
transform 1 0 31188 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_339
timestamp 1623621585
transform 1 0 32292 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_351
timestamp 1623621585
transform 1 0 33396 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1676
timestamp 1623621585
transform 1 0 35236 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_177_363
timestamp 1623621585
transform 1 0 34500 0 1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_177_372
timestamp 1623621585
transform 1 0 35328 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_384
timestamp 1623621585
transform 1 0 36432 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_355
timestamp 1623621585
transform -1 0 38824 0 1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input275
timestamp 1623621585
transform 1 0 37904 0 1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_177_396
timestamp 1623621585
transform 1 0 37536 0 1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_177_403
timestamp 1623621585
transform 1 0 38180 0 1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_356
timestamp 1623621585
transform 1 0 1104 0 -1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_358
timestamp 1623621585
transform 1 0 1104 0 1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input435
timestamp 1623621585
transform 1 0 1380 0 -1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_178_6
timestamp 1623621585
transform 1 0 1656 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_18
timestamp 1623621585
transform 1 0 2760 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_3
timestamp 1623621585
transform 1 0 1380 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_15
timestamp 1623621585
transform 1 0 2484 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1684
timestamp 1623621585
transform 1 0 3772 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_30
timestamp 1623621585
transform 1 0 3864 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_179_27
timestamp 1623621585
transform 1 0 3588 0 1 99552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_179_30
timestamp 1623621585
transform 1 0 3864 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _728_
timestamp 1623621585
transform 1 0 5060 0 -1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _730_
timestamp 1623621585
transform 1 0 6072 0 1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1677
timestamp 1623621585
transform 1 0 6348 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_178_42
timestamp 1623621585
transform 1 0 4968 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_178_46
timestamp 1623621585
transform 1 0 5336 0 -1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_178_54
timestamp 1623621585
transform 1 0 6072 0 -1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_178_58
timestamp 1623621585
transform 1 0 6440 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_42
timestamp 1623621585
transform 1 0 4968 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_57
timestamp 1623621585
transform 1 0 6348 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_70
timestamp 1623621585
transform 1 0 7544 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_82
timestamp 1623621585
transform 1 0 8648 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_69
timestamp 1623621585
transform 1 0 7452 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_179_81
timestamp 1623621585
transform 1 0 8556 0 1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1685
timestamp 1623621585
transform 1 0 9016 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_94
timestamp 1623621585
transform 1 0 9752 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_179_85
timestamp 1623621585
transform 1 0 8924 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_87
timestamp 1623621585
transform 1 0 9108 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_99
timestamp 1623621585
transform 1 0 10212 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1678
timestamp 1623621585
transform 1 0 11592 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_178_106
timestamp 1623621585
transform 1 0 10856 0 -1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_178_115
timestamp 1623621585
transform 1 0 11684 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_111
timestamp 1623621585
transform 1 0 11316 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_123
timestamp 1623621585
transform 1 0 12420 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1686
timestamp 1623621585
transform 1 0 14260 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_127
timestamp 1623621585
transform 1 0 12788 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_139
timestamp 1623621585
transform 1 0 13892 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_179_135
timestamp 1623621585
transform 1 0 13524 0 1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_179_144
timestamp 1623621585
transform 1 0 14352 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_151
timestamp 1623621585
transform 1 0 14996 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_178_163
timestamp 1623621585
transform 1 0 16100 0 -1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_179_156
timestamp 1623621585
transform 1 0 15456 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1679
timestamp 1623621585
transform 1 0 16836 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_172
timestamp 1623621585
transform 1 0 16928 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_184
timestamp 1623621585
transform 1 0 18032 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_168
timestamp 1623621585
transform 1 0 16560 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_180
timestamp 1623621585
transform 1 0 17664 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1687
timestamp 1623621585
transform 1 0 19504 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_196
timestamp 1623621585
transform 1 0 19136 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_208
timestamp 1623621585
transform 1 0 20240 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_179_192
timestamp 1623621585
transform 1 0 18768 0 1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_179_201
timestamp 1623621585
transform 1 0 19596 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1680
timestamp 1623621585
transform 1 0 22080 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_178_220
timestamp 1623621585
transform 1 0 21344 0 -1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_178_229
timestamp 1623621585
transform 1 0 22172 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_213
timestamp 1623621585
transform 1 0 20700 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_225
timestamp 1623621585
transform 1 0 21804 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_241
timestamp 1623621585
transform 1 0 23276 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_237
timestamp 1623621585
transform 1 0 22908 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_179_249
timestamp 1623621585
transform 1 0 24012 0 1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1688
timestamp 1623621585
transform 1 0 24748 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_253
timestamp 1623621585
transform 1 0 24380 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_265
timestamp 1623621585
transform 1 0 25484 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_258
timestamp 1623621585
transform 1 0 24840 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_270
timestamp 1623621585
transform 1 0 25944 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1681
timestamp 1623621585
transform 1 0 27324 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_178_277
timestamp 1623621585
transform 1 0 26588 0 -1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_178_286
timestamp 1623621585
transform 1 0 27416 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_282
timestamp 1623621585
transform 1 0 27048 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_298
timestamp 1623621585
transform 1 0 28520 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_310
timestamp 1623621585
transform 1 0 29624 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_294
timestamp 1623621585
transform 1 0 28152 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_179_306
timestamp 1623621585
transform 1 0 29256 0 1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1689
timestamp 1623621585
transform 1 0 29992 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_322
timestamp 1623621585
transform 1 0 30728 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_315
timestamp 1623621585
transform 1 0 30084 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_327
timestamp 1623621585
transform 1 0 31188 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1682
timestamp 1623621585
transform 1 0 32568 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_178_334
timestamp 1623621585
transform 1 0 31832 0 -1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_178_343
timestamp 1623621585
transform 1 0 32660 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_339
timestamp 1623621585
transform 1 0 32292 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_351
timestamp 1623621585
transform 1 0 33396 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1690
timestamp 1623621585
transform 1 0 35236 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_355
timestamp 1623621585
transform 1 0 33764 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_367
timestamp 1623621585
transform 1 0 34868 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_179_363
timestamp 1623621585
transform 1 0 34500 0 1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_179_372
timestamp 1623621585
transform 1 0 35328 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input278
timestamp 1623621585
transform 1 0 37168 0 -1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input279
timestamp 1623621585
transform 1 0 37260 0 1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_178_379
timestamp 1623621585
transform 1 0 35972 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_178_391
timestamp 1623621585
transform 1 0 37076 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_178_395
timestamp 1623621585
transform 1 0 37444 0 -1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_179_384
timestamp 1623621585
transform 1 0 36432 0 1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_179_392
timestamp 1623621585
transform 1 0 37168 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_357
timestamp 1623621585
transform -1 0 38824 0 -1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_359
timestamp 1623621585
transform -1 0 38824 0 1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1683
timestamp 1623621585
transform 1 0 37812 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input276
timestamp 1623621585
transform 1 0 37904 0 1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_178_400
timestamp 1623621585
transform 1 0 37904 0 -1 99552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_406
timestamp 1623621585
transform 1 0 38456 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_179_396
timestamp 1623621585
transform 1 0 37536 0 1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_179_403
timestamp 1623621585
transform 1 0 38180 0 1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_360
timestamp 1623621585
transform 1 0 1104 0 -1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input436
timestamp 1623621585
transform 1 0 1380 0 -1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_180_6
timestamp 1623621585
transform 1 0 1656 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_18
timestamp 1623621585
transform 1 0 2760 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_30
timestamp 1623621585
transform 1 0 3864 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1691
timestamp 1623621585
transform 1 0 6348 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_42
timestamp 1623621585
transform 1 0 4968 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_180_54
timestamp 1623621585
transform 1 0 6072 0 -1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_180_58
timestamp 1623621585
transform 1 0 6440 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_70
timestamp 1623621585
transform 1 0 7544 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_82
timestamp 1623621585
transform 1 0 8648 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_94
timestamp 1623621585
transform 1 0 9752 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1692
timestamp 1623621585
transform 1 0 11592 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_180_106
timestamp 1623621585
transform 1 0 10856 0 -1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_180_115
timestamp 1623621585
transform 1 0 11684 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_127
timestamp 1623621585
transform 1 0 12788 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_139
timestamp 1623621585
transform 1 0 13892 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_151
timestamp 1623621585
transform 1 0 14996 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_180_163
timestamp 1623621585
transform 1 0 16100 0 -1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1693
timestamp 1623621585
transform 1 0 16836 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_172
timestamp 1623621585
transform 1 0 16928 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_184
timestamp 1623621585
transform 1 0 18032 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_196
timestamp 1623621585
transform 1 0 19136 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_208
timestamp 1623621585
transform 1 0 20240 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1694
timestamp 1623621585
transform 1 0 22080 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_180_220
timestamp 1623621585
transform 1 0 21344 0 -1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_180_229
timestamp 1623621585
transform 1 0 22172 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_241
timestamp 1623621585
transform 1 0 23276 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_253
timestamp 1623621585
transform 1 0 24380 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_265
timestamp 1623621585
transform 1 0 25484 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1695
timestamp 1623621585
transform 1 0 27324 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_180_277
timestamp 1623621585
transform 1 0 26588 0 -1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_180_286
timestamp 1623621585
transform 1 0 27416 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_298
timestamp 1623621585
transform 1 0 28520 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_310
timestamp 1623621585
transform 1 0 29624 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_322
timestamp 1623621585
transform 1 0 30728 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1696
timestamp 1623621585
transform 1 0 32568 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_180_334
timestamp 1623621585
transform 1 0 31832 0 -1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_180_343
timestamp 1623621585
transform 1 0 32660 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_355
timestamp 1623621585
transform 1 0 33764 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_367
timestamp 1623621585
transform 1 0 34868 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input287
timestamp 1623621585
transform 1 0 37076 0 -1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_180_379
timestamp 1623621585
transform 1 0 35972 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_180_395
timestamp 1623621585
transform 1 0 37444 0 -1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_361
timestamp 1623621585
transform -1 0 38824 0 -1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1697
timestamp 1623621585
transform 1 0 37812 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_180_400
timestamp 1623621585
transform 1 0 37904 0 -1 100640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_406
timestamp 1623621585
transform 1 0 38456 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_362
timestamp 1623621585
transform 1 0 1104 0 1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input438
timestamp 1623621585
transform 1 0 1380 0 1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_181_6
timestamp 1623621585
transform 1 0 1656 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_181_18
timestamp 1623621585
transform 1 0 2760 0 1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1698
timestamp 1623621585
transform 1 0 3772 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_181_26
timestamp 1623621585
transform 1 0 3496 0 1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_181_30
timestamp 1623621585
transform 1 0 3864 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _719_
timestamp 1623621585
transform 1 0 6348 0 1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_181_42
timestamp 1623621585
transform 1 0 4968 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_181_54
timestamp 1623621585
transform 1 0 6072 0 1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_181_60
timestamp 1623621585
transform 1 0 6624 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_72
timestamp 1623621585
transform 1 0 7728 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1699
timestamp 1623621585
transform 1 0 9016 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_181_84
timestamp 1623621585
transform 1 0 8832 0 1 100640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_181_87
timestamp 1623621585
transform 1 0 9108 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_99
timestamp 1623621585
transform 1 0 10212 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_111
timestamp 1623621585
transform 1 0 11316 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_123
timestamp 1623621585
transform 1 0 12420 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1700
timestamp 1623621585
transform 1 0 14260 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_181_135
timestamp 1623621585
transform 1 0 13524 0 1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_181_144
timestamp 1623621585
transform 1 0 14352 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_156
timestamp 1623621585
transform 1 0 15456 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_168
timestamp 1623621585
transform 1 0 16560 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_180
timestamp 1623621585
transform 1 0 17664 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1701
timestamp 1623621585
transform 1 0 19504 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_181_192
timestamp 1623621585
transform 1 0 18768 0 1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_181_201
timestamp 1623621585
transform 1 0 19596 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_213
timestamp 1623621585
transform 1 0 20700 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_225
timestamp 1623621585
transform 1 0 21804 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_237
timestamp 1623621585
transform 1 0 22908 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_181_249
timestamp 1623621585
transform 1 0 24012 0 1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1702
timestamp 1623621585
transform 1 0 24748 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_258
timestamp 1623621585
transform 1 0 24840 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_270
timestamp 1623621585
transform 1 0 25944 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_282
timestamp 1623621585
transform 1 0 27048 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_294
timestamp 1623621585
transform 1 0 28152 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_181_306
timestamp 1623621585
transform 1 0 29256 0 1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1703
timestamp 1623621585
transform 1 0 29992 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_315
timestamp 1623621585
transform 1 0 30084 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_327
timestamp 1623621585
transform 1 0 31188 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_339
timestamp 1623621585
transform 1 0 32292 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_351
timestamp 1623621585
transform 1 0 33396 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1704
timestamp 1623621585
transform 1 0 35236 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_181_363
timestamp 1623621585
transform 1 0 34500 0 1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_181_372
timestamp 1623621585
transform 1 0 35328 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_384
timestamp 1623621585
transform 1 0 36432 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_363
timestamp 1623621585
transform -1 0 38824 0 1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input298
timestamp 1623621585
transform 1 0 37812 0 1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_181_396
timestamp 1623621585
transform 1 0 37536 0 1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_181_403
timestamp 1623621585
transform 1 0 38180 0 1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_364
timestamp 1623621585
transform 1 0 1104 0 -1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_182_3
timestamp 1623621585
transform 1 0 1380 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_15
timestamp 1623621585
transform 1 0 2484 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_27
timestamp 1623621585
transform 1 0 3588 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_39
timestamp 1623621585
transform 1 0 4692 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1705
timestamp 1623621585
transform 1 0 6348 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_182_51
timestamp 1623621585
transform 1 0 5796 0 -1 101728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_182_58
timestamp 1623621585
transform 1 0 6440 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_70
timestamp 1623621585
transform 1 0 7544 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_82
timestamp 1623621585
transform 1 0 8648 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_94
timestamp 1623621585
transform 1 0 9752 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1706
timestamp 1623621585
transform 1 0 11592 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_182_106
timestamp 1623621585
transform 1 0 10856 0 -1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_182_115
timestamp 1623621585
transform 1 0 11684 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_127
timestamp 1623621585
transform 1 0 12788 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_139
timestamp 1623621585
transform 1 0 13892 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_151
timestamp 1623621585
transform 1 0 14996 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_182_163
timestamp 1623621585
transform 1 0 16100 0 -1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1707
timestamp 1623621585
transform 1 0 16836 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_172
timestamp 1623621585
transform 1 0 16928 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_184
timestamp 1623621585
transform 1 0 18032 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_196
timestamp 1623621585
transform 1 0 19136 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_208
timestamp 1623621585
transform 1 0 20240 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1708
timestamp 1623621585
transform 1 0 22080 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_182_220
timestamp 1623621585
transform 1 0 21344 0 -1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_182_229
timestamp 1623621585
transform 1 0 22172 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_241
timestamp 1623621585
transform 1 0 23276 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_253
timestamp 1623621585
transform 1 0 24380 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_265
timestamp 1623621585
transform 1 0 25484 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1709
timestamp 1623621585
transform 1 0 27324 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_182_277
timestamp 1623621585
transform 1 0 26588 0 -1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_182_286
timestamp 1623621585
transform 1 0 27416 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_298
timestamp 1623621585
transform 1 0 28520 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_310
timestamp 1623621585
transform 1 0 29624 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_322
timestamp 1623621585
transform 1 0 30728 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1710
timestamp 1623621585
transform 1 0 32568 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_182_334
timestamp 1623621585
transform 1 0 31832 0 -1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_182_343
timestamp 1623621585
transform 1 0 32660 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_355
timestamp 1623621585
transform 1 0 33764 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_367
timestamp 1623621585
transform 1 0 34868 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input309
timestamp 1623621585
transform 1 0 37076 0 -1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_182_379
timestamp 1623621585
transform 1 0 35972 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_182_395
timestamp 1623621585
transform 1 0 37444 0 -1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_365
timestamp 1623621585
transform -1 0 38824 0 -1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1711
timestamp 1623621585
transform 1 0 37812 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_182_400
timestamp 1623621585
transform 1 0 37904 0 -1 101728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_406
timestamp 1623621585
transform 1 0 38456 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_366
timestamp 1623621585
transform 1 0 1104 0 1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input439
timestamp 1623621585
transform 1 0 1380 0 1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_183_6
timestamp 1623621585
transform 1 0 1656 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_183_18
timestamp 1623621585
transform 1 0 2760 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1712
timestamp 1623621585
transform 1 0 3772 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_183_26
timestamp 1623621585
transform 1 0 3496 0 1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_183_30
timestamp 1623621585
transform 1 0 3864 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_42
timestamp 1623621585
transform 1 0 4968 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_54
timestamp 1623621585
transform 1 0 6072 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_66
timestamp 1623621585
transform 1 0 7176 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_183_78
timestamp 1623621585
transform 1 0 8280 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _736_
timestamp 1623621585
transform 1 0 9476 0 1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1713
timestamp 1623621585
transform 1 0 9016 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_183_87
timestamp 1623621585
transform 1 0 9108 0 1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_183_94
timestamp 1623621585
transform 1 0 9752 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_106
timestamp 1623621585
transform 1 0 10856 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_118
timestamp 1623621585
transform 1 0 11960 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1714
timestamp 1623621585
transform 1 0 14260 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_130
timestamp 1623621585
transform 1 0 13064 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_183_142
timestamp 1623621585
transform 1 0 14168 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_144
timestamp 1623621585
transform 1 0 14352 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_156
timestamp 1623621585
transform 1 0 15456 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_168
timestamp 1623621585
transform 1 0 16560 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_180
timestamp 1623621585
transform 1 0 17664 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1715
timestamp 1623621585
transform 1 0 19504 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_183_192
timestamp 1623621585
transform 1 0 18768 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_183_201
timestamp 1623621585
transform 1 0 19596 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_213
timestamp 1623621585
transform 1 0 20700 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_225
timestamp 1623621585
transform 1 0 21804 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_237
timestamp 1623621585
transform 1 0 22908 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_183_249
timestamp 1623621585
transform 1 0 24012 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _729_
timestamp 1623621585
transform 1 0 25576 0 1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1716
timestamp 1623621585
transform 1 0 24748 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_183_258
timestamp 1623621585
transform 1 0 24840 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_183_270
timestamp 1623621585
transform 1 0 25944 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_282
timestamp 1623621585
transform 1 0 27048 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_294
timestamp 1623621585
transform 1 0 28152 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_183_306
timestamp 1623621585
transform 1 0 29256 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1717
timestamp 1623621585
transform 1 0 29992 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_315
timestamp 1623621585
transform 1 0 30084 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_327
timestamp 1623621585
transform 1 0 31188 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_339
timestamp 1623621585
transform 1 0 32292 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_351
timestamp 1623621585
transform 1 0 33396 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1718
timestamp 1623621585
transform 1 0 35236 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_183_363
timestamp 1623621585
transform 1 0 34500 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_183_372
timestamp 1623621585
transform 1 0 35328 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input313
timestamp 1623621585
transform 1 0 37076 0 1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_183_384
timestamp 1623621585
transform 1 0 36432 0 1 101728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_390
timestamp 1623621585
transform 1 0 36984 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_183_395
timestamp 1623621585
transform 1 0 37444 0 1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_367
timestamp 1623621585
transform -1 0 38824 0 1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input312
timestamp 1623621585
transform 1 0 37812 0 1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_183_403
timestamp 1623621585
transform 1 0 38180 0 1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_368
timestamp 1623621585
transform 1 0 1104 0 -1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output672
timestamp 1623621585
transform 1 0 1748 0 -1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_184_3
timestamp 1623621585
transform 1 0 1380 0 -1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_184_11
timestamp 1623621585
transform 1 0 2116 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_23
timestamp 1623621585
transform 1 0 3220 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_35
timestamp 1623621585
transform 1 0 4324 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1719
timestamp 1623621585
transform 1 0 6348 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_184_47
timestamp 1623621585
transform 1 0 5428 0 -1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_184_55
timestamp 1623621585
transform 1 0 6164 0 -1 102816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_184_58
timestamp 1623621585
transform 1 0 6440 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _733_
timestamp 1623621585
transform 1 0 7544 0 -1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_184_73
timestamp 1623621585
transform 1 0 7820 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_85
timestamp 1623621585
transform 1 0 8924 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_97
timestamp 1623621585
transform 1 0 10028 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1720
timestamp 1623621585
transform 1 0 11592 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_184_109
timestamp 1623621585
transform 1 0 11132 0 -1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_184_113
timestamp 1623621585
transform 1 0 11500 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_115
timestamp 1623621585
transform 1 0 11684 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_127
timestamp 1623621585
transform 1 0 12788 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_139
timestamp 1623621585
transform 1 0 13892 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_151
timestamp 1623621585
transform 1 0 14996 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_184_163
timestamp 1623621585
transform 1 0 16100 0 -1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1721
timestamp 1623621585
transform 1 0 16836 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_172
timestamp 1623621585
transform 1 0 16928 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_184
timestamp 1623621585
transform 1 0 18032 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_196
timestamp 1623621585
transform 1 0 19136 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_208
timestamp 1623621585
transform 1 0 20240 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1722
timestamp 1623621585
transform 1 0 22080 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_184_220
timestamp 1623621585
transform 1 0 21344 0 -1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_184_229
timestamp 1623621585
transform 1 0 22172 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_241
timestamp 1623621585
transform 1 0 23276 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_253
timestamp 1623621585
transform 1 0 24380 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_265
timestamp 1623621585
transform 1 0 25484 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1723
timestamp 1623621585
transform 1 0 27324 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_184_277
timestamp 1623621585
transform 1 0 26588 0 -1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_184_286
timestamp 1623621585
transform 1 0 27416 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_298
timestamp 1623621585
transform 1 0 28520 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_310
timestamp 1623621585
transform 1 0 29624 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_322
timestamp 1623621585
transform 1 0 30728 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1724
timestamp 1623621585
transform 1 0 32568 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_184_334
timestamp 1623621585
transform 1 0 31832 0 -1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_184_343
timestamp 1623621585
transform 1 0 32660 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_355
timestamp 1623621585
transform 1 0 33764 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_367
timestamp 1623621585
transform 1 0 34868 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input314
timestamp 1623621585
transform 1 0 37076 0 -1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_184_379
timestamp 1623621585
transform 1 0 35972 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_184_395
timestamp 1623621585
transform 1 0 37444 0 -1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_369
timestamp 1623621585
transform -1 0 38824 0 -1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1725
timestamp 1623621585
transform 1 0 37812 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_184_400
timestamp 1623621585
transform 1 0 37904 0 -1 102816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_406
timestamp 1623621585
transform 1 0 38456 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_370
timestamp 1623621585
transform 1 0 1104 0 1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_372
timestamp 1623621585
transform 1 0 1104 0 -1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output616
timestamp 1623621585
transform 1 0 1748 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_185_3
timestamp 1623621585
transform 1 0 1380 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_15
timestamp 1623621585
transform 1 0 2484 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_186_3
timestamp 1623621585
transform 1 0 1380 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_186_11
timestamp 1623621585
transform 1 0 2116 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1726
timestamp 1623621585
transform 1 0 3772 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_185_27
timestamp 1623621585
transform 1 0 3588 0 1 102816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_185_30
timestamp 1623621585
transform 1 0 3864 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_23
timestamp 1623621585
transform 1 0 3220 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_35
timestamp 1623621585
transform 1 0 4324 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1733
timestamp 1623621585
transform 1 0 6348 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_42
timestamp 1623621585
transform 1 0 4968 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_185_54
timestamp 1623621585
transform 1 0 6072 0 1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_185_62
timestamp 1623621585
transform 1 0 6808 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_186_47
timestamp 1623621585
transform 1 0 5428 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_186_55
timestamp 1623621585
transform 1 0 6164 0 -1 103904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_186_58
timestamp 1623621585
transform 1 0 6440 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _720_
timestamp 1623621585
transform 1 0 6900 0 1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_185_66
timestamp 1623621585
transform 1 0 7176 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_185_78
timestamp 1623621585
transform 1 0 8280 0 1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_186_70
timestamp 1623621585
transform 1 0 7544 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_82
timestamp 1623621585
transform 1 0 8648 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1727
timestamp 1623621585
transform 1 0 9016 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_87
timestamp 1623621585
transform 1 0 9108 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_99
timestamp 1623621585
transform 1 0 10212 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_94
timestamp 1623621585
transform 1 0 9752 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1734
timestamp 1623621585
transform 1 0 11592 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_111
timestamp 1623621585
transform 1 0 11316 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_123
timestamp 1623621585
transform 1 0 12420 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_186_106
timestamp 1623621585
transform 1 0 10856 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_186_115
timestamp 1623621585
transform 1 0 11684 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1728
timestamp 1623621585
transform 1 0 14260 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_185_135
timestamp 1623621585
transform 1 0 13524 0 1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_185_144
timestamp 1623621585
transform 1 0 14352 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_127
timestamp 1623621585
transform 1 0 12788 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_139
timestamp 1623621585
transform 1 0 13892 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_156
timestamp 1623621585
transform 1 0 15456 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_151
timestamp 1623621585
transform 1 0 14996 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_186_163
timestamp 1623621585
transform 1 0 16100 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1735
timestamp 1623621585
transform 1 0 16836 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_168
timestamp 1623621585
transform 1 0 16560 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_180
timestamp 1623621585
transform 1 0 17664 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_172
timestamp 1623621585
transform 1 0 16928 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_184
timestamp 1623621585
transform 1 0 18032 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1729
timestamp 1623621585
transform 1 0 19504 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_185_192
timestamp 1623621585
transform 1 0 18768 0 1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_185_201
timestamp 1623621585
transform 1 0 19596 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_196
timestamp 1623621585
transform 1 0 19136 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_208
timestamp 1623621585
transform 1 0 20240 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1736
timestamp 1623621585
transform 1 0 22080 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_213
timestamp 1623621585
transform 1 0 20700 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_225
timestamp 1623621585
transform 1 0 21804 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_186_220
timestamp 1623621585
transform 1 0 21344 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_186_229
timestamp 1623621585
transform 1 0 22172 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_237
timestamp 1623621585
transform 1 0 22908 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_185_249
timestamp 1623621585
transform 1 0 24012 0 1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_186_241
timestamp 1623621585
transform 1 0 23276 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _717_
timestamp 1623621585
transform 1 0 25392 0 1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1730
timestamp 1623621585
transform 1 0 24748 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_185_258
timestamp 1623621585
transform 1 0 24840 0 1 102816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_185_268
timestamp 1623621585
transform 1 0 25760 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_253
timestamp 1623621585
transform 1 0 24380 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_265
timestamp 1623621585
transform 1 0 25484 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1737
timestamp 1623621585
transform 1 0 27324 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_280
timestamp 1623621585
transform 1 0 26864 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_186_277
timestamp 1623621585
transform 1 0 26588 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_186_286
timestamp 1623621585
transform 1 0 27416 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_292
timestamp 1623621585
transform 1 0 27968 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_185_304
timestamp 1623621585
transform 1 0 29072 0 1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_185_312
timestamp 1623621585
transform 1 0 29808 0 1 102816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_186_298
timestamp 1623621585
transform 1 0 28520 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_186_310
timestamp 1623621585
transform 1 0 29624 0 -1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _588_
timestamp 1623621585
transform 1 0 30820 0 -1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _592_
timestamp 1623621585
transform 1 0 30452 0 1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _597_
timestamp 1623621585
transform 1 0 29900 0 -1 103904
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1731
timestamp 1623621585
transform 1 0 29992 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_185_315
timestamp 1623621585
transform 1 0 30084 0 1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_185_322
timestamp 1623621585
transform 1 0 30728 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_186_319
timestamp 1623621585
transform 1 0 30452 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_186_326
timestamp 1623621585
transform 1 0 31096 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1738
timestamp 1623621585
transform 1 0 32568 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_334
timestamp 1623621585
transform 1 0 31832 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_346
timestamp 1623621585
transform 1 0 32936 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_186_338
timestamp 1623621585
transform 1 0 32200 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_186_343
timestamp 1623621585
transform 1 0 32660 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1732
timestamp 1623621585
transform 1 0 35236 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_358
timestamp 1623621585
transform 1 0 34040 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_185_370
timestamp 1623621585
transform 1 0 35144 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_372
timestamp 1623621585
transform 1 0 35328 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_355
timestamp 1623621585
transform 1 0 33764 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_367
timestamp 1623621585
transform 1 0 34868 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input316
timestamp 1623621585
transform 1 0 37076 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_185_384
timestamp 1623621585
transform 1 0 36432 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_379
timestamp 1623621585
transform 1 0 35972 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_186_395
timestamp 1623621585
transform 1 0 37444 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_371
timestamp 1623621585
transform -1 0 38824 0 1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_373
timestamp 1623621585
transform -1 0 38824 0 -1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1739
timestamp 1623621585
transform 1 0 37812 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input315
timestamp 1623621585
transform 1 0 37812 0 1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_185_396
timestamp 1623621585
transform 1 0 37536 0 1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_185_403
timestamp 1623621585
transform 1 0 38180 0 1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_186_400
timestamp 1623621585
transform 1 0 37904 0 -1 103904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_406
timestamp 1623621585
transform 1 0 38456 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_374
timestamp 1623621585
transform 1 0 1104 0 1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input54
timestamp 1623621585
transform 1 0 1380 0 1 103904
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_187_12
timestamp 1623621585
transform 1 0 2208 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1740
timestamp 1623621585
transform 1 0 3772 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_187_24
timestamp 1623621585
transform 1 0 3312 0 1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_187_28
timestamp 1623621585
transform 1 0 3680 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_30
timestamp 1623621585
transform 1 0 3864 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_42
timestamp 1623621585
transform 1 0 4968 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_54
timestamp 1623621585
transform 1 0 6072 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_66
timestamp 1623621585
transform 1 0 7176 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_187_78
timestamp 1623621585
transform 1 0 8280 0 1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1741
timestamp 1623621585
transform 1 0 9016 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_87
timestamp 1623621585
transform 1 0 9108 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_99
timestamp 1623621585
transform 1 0 10212 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_111
timestamp 1623621585
transform 1 0 11316 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_123
timestamp 1623621585
transform 1 0 12420 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1742
timestamp 1623621585
transform 1 0 14260 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_187_135
timestamp 1623621585
transform 1 0 13524 0 1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_187_144
timestamp 1623621585
transform 1 0 14352 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_156
timestamp 1623621585
transform 1 0 15456 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_168
timestamp 1623621585
transform 1 0 16560 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_180
timestamp 1623621585
transform 1 0 17664 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1743
timestamp 1623621585
transform 1 0 19504 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_187_192
timestamp 1623621585
transform 1 0 18768 0 1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_187_201
timestamp 1623621585
transform 1 0 19596 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_213
timestamp 1623621585
transform 1 0 20700 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_225
timestamp 1623621585
transform 1 0 21804 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_237
timestamp 1623621585
transform 1 0 22908 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_187_249
timestamp 1623621585
transform 1 0 24012 0 1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1744
timestamp 1623621585
transform 1 0 24748 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_258
timestamp 1623621585
transform 1 0 24840 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_270
timestamp 1623621585
transform 1 0 25944 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_282
timestamp 1623621585
transform 1 0 27048 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_294
timestamp 1623621585
transform 1 0 28152 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_187_306
timestamp 1623621585
transform 1 0 29256 0 1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _595_
timestamp 1623621585
transform 1 0 30452 0 1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1745
timestamp 1623621585
transform 1 0 29992 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_187_315
timestamp 1623621585
transform 1 0 30084 0 1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_187_323
timestamp 1623621585
transform 1 0 30820 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_335
timestamp 1623621585
transform 1 0 31924 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_347
timestamp 1623621585
transform 1 0 33028 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1746
timestamp 1623621585
transform 1 0 35236 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_359
timestamp 1623621585
transform 1 0 34132 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_372
timestamp 1623621585
transform 1 0 35328 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input318
timestamp 1623621585
transform 1 0 37076 0 1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_187_384
timestamp 1623621585
transform 1 0 36432 0 1 103904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_390
timestamp 1623621585
transform 1 0 36984 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_187_395
timestamp 1623621585
transform 1 0 37444 0 1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_375
timestamp 1623621585
transform -1 0 38824 0 1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input317
timestamp 1623621585
transform 1 0 37812 0 1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_187_403
timestamp 1623621585
transform 1 0 38180 0 1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_376
timestamp 1623621585
transform 1 0 1104 0 -1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_188_3
timestamp 1623621585
transform 1 0 1380 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_15
timestamp 1623621585
transform 1 0 2484 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_27
timestamp 1623621585
transform 1 0 3588 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_39
timestamp 1623621585
transform 1 0 4692 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1747
timestamp 1623621585
transform 1 0 6348 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_188_51
timestamp 1623621585
transform 1 0 5796 0 -1 104992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_188_58
timestamp 1623621585
transform 1 0 6440 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_70
timestamp 1623621585
transform 1 0 7544 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_82
timestamp 1623621585
transform 1 0 8648 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_94
timestamp 1623621585
transform 1 0 9752 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1748
timestamp 1623621585
transform 1 0 11592 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_188_106
timestamp 1623621585
transform 1 0 10856 0 -1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_188_115
timestamp 1623621585
transform 1 0 11684 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_127
timestamp 1623621585
transform 1 0 12788 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_139
timestamp 1623621585
transform 1 0 13892 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_151
timestamp 1623621585
transform 1 0 14996 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_188_163
timestamp 1623621585
transform 1 0 16100 0 -1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1749
timestamp 1623621585
transform 1 0 16836 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_172
timestamp 1623621585
transform 1 0 16928 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_184
timestamp 1623621585
transform 1 0 18032 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_196
timestamp 1623621585
transform 1 0 19136 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_208
timestamp 1623621585
transform 1 0 20240 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1750
timestamp 1623621585
transform 1 0 22080 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_188_220
timestamp 1623621585
transform 1 0 21344 0 -1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_188_229
timestamp 1623621585
transform 1 0 22172 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_241
timestamp 1623621585
transform 1 0 23276 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_253
timestamp 1623621585
transform 1 0 24380 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_265
timestamp 1623621585
transform 1 0 25484 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1751
timestamp 1623621585
transform 1 0 27324 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_188_277
timestamp 1623621585
transform 1 0 26588 0 -1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_188_286
timestamp 1623621585
transform 1 0 27416 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_298
timestamp 1623621585
transform 1 0 28520 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_310
timestamp 1623621585
transform 1 0 29624 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_322
timestamp 1623621585
transform 1 0 30728 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1752
timestamp 1623621585
transform 1 0 32568 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_188_334
timestamp 1623621585
transform 1 0 31832 0 -1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_188_343
timestamp 1623621585
transform 1 0 32660 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_355
timestamp 1623621585
transform 1 0 33764 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_367
timestamp 1623621585
transform 1 0 34868 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input288
timestamp 1623621585
transform 1 0 37076 0 -1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_188_379
timestamp 1623621585
transform 1 0 35972 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_188_395
timestamp 1623621585
transform 1 0 37444 0 -1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_377
timestamp 1623621585
transform -1 0 38824 0 -1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1753
timestamp 1623621585
transform 1 0 37812 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_188_400
timestamp 1623621585
transform 1 0 37904 0 -1 104992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_406
timestamp 1623621585
transform 1 0 38456 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_378
timestamp 1623621585
transform 1 0 1104 0 1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output651
timestamp 1623621585
transform 1 0 1748 0 1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_189_3
timestamp 1623621585
transform 1 0 1380 0 1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_189_11
timestamp 1623621585
transform 1 0 2116 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1754
timestamp 1623621585
transform 1 0 3772 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_189_23
timestamp 1623621585
transform 1 0 3220 0 1 104992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_189_30
timestamp 1623621585
transform 1 0 3864 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_42
timestamp 1623621585
transform 1 0 4968 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_54
timestamp 1623621585
transform 1 0 6072 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_66
timestamp 1623621585
transform 1 0 7176 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_189_78
timestamp 1623621585
transform 1 0 8280 0 1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1755
timestamp 1623621585
transform 1 0 9016 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_87
timestamp 1623621585
transform 1 0 9108 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_99
timestamp 1623621585
transform 1 0 10212 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_111
timestamp 1623621585
transform 1 0 11316 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_123
timestamp 1623621585
transform 1 0 12420 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1756
timestamp 1623621585
transform 1 0 14260 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_189_135
timestamp 1623621585
transform 1 0 13524 0 1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_189_144
timestamp 1623621585
transform 1 0 14352 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_156
timestamp 1623621585
transform 1 0 15456 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_168
timestamp 1623621585
transform 1 0 16560 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_180
timestamp 1623621585
transform 1 0 17664 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1757
timestamp 1623621585
transform 1 0 19504 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_189_192
timestamp 1623621585
transform 1 0 18768 0 1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_189_201
timestamp 1623621585
transform 1 0 19596 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_213
timestamp 1623621585
transform 1 0 20700 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_225
timestamp 1623621585
transform 1 0 21804 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_237
timestamp 1623621585
transform 1 0 22908 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_189_249
timestamp 1623621585
transform 1 0 24012 0 1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1758
timestamp 1623621585
transform 1 0 24748 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_258
timestamp 1623621585
transform 1 0 24840 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_270
timestamp 1623621585
transform 1 0 25944 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_282
timestamp 1623621585
transform 1 0 27048 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_294
timestamp 1623621585
transform 1 0 28152 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_189_306
timestamp 1623621585
transform 1 0 29256 0 1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1759
timestamp 1623621585
transform 1 0 29992 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_315
timestamp 1623621585
transform 1 0 30084 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_327
timestamp 1623621585
transform 1 0 31188 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_339
timestamp 1623621585
transform 1 0 32292 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_351
timestamp 1623621585
transform 1 0 33396 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1760
timestamp 1623621585
transform 1 0 35236 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_189_363
timestamp 1623621585
transform 1 0 34500 0 1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_189_372
timestamp 1623621585
transform 1 0 35328 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_384
timestamp 1623621585
transform 1 0 36432 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_379
timestamp 1623621585
transform -1 0 38824 0 1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input289
timestamp 1623621585
transform 1 0 37812 0 1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_189_396
timestamp 1623621585
transform 1 0 37536 0 1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_189_403
timestamp 1623621585
transform 1 0 38180 0 1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_380
timestamp 1623621585
transform 1 0 1104 0 -1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input55
timestamp 1623621585
transform 1 0 1380 0 -1 106080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_190_9
timestamp 1623621585
transform 1 0 1932 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_21
timestamp 1623621585
transform 1 0 3036 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_33
timestamp 1623621585
transform 1 0 4140 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1761
timestamp 1623621585
transform 1 0 6348 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_45
timestamp 1623621585
transform 1 0 5244 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_58
timestamp 1623621585
transform 1 0 6440 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_70
timestamp 1623621585
transform 1 0 7544 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_82
timestamp 1623621585
transform 1 0 8648 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _738_
timestamp 1623621585
transform 1 0 9936 0 -1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_190_94
timestamp 1623621585
transform 1 0 9752 0 -1 106080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_190_99
timestamp 1623621585
transform 1 0 10212 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1762
timestamp 1623621585
transform 1 0 11592 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_190_111
timestamp 1623621585
transform 1 0 11316 0 -1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_190_115
timestamp 1623621585
transform 1 0 11684 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_127
timestamp 1623621585
transform 1 0 12788 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_139
timestamp 1623621585
transform 1 0 13892 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_151
timestamp 1623621585
transform 1 0 14996 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_190_163
timestamp 1623621585
transform 1 0 16100 0 -1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1763
timestamp 1623621585
transform 1 0 16836 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_172
timestamp 1623621585
transform 1 0 16928 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_184
timestamp 1623621585
transform 1 0 18032 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_196
timestamp 1623621585
transform 1 0 19136 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_208
timestamp 1623621585
transform 1 0 20240 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1764
timestamp 1623621585
transform 1 0 22080 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_190_220
timestamp 1623621585
transform 1 0 21344 0 -1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_190_229
timestamp 1623621585
transform 1 0 22172 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_241
timestamp 1623621585
transform 1 0 23276 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_253
timestamp 1623621585
transform 1 0 24380 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_265
timestamp 1623621585
transform 1 0 25484 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1765
timestamp 1623621585
transform 1 0 27324 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_190_277
timestamp 1623621585
transform 1 0 26588 0 -1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_190_286
timestamp 1623621585
transform 1 0 27416 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_298
timestamp 1623621585
transform 1 0 28520 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_310
timestamp 1623621585
transform 1 0 29624 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_322
timestamp 1623621585
transform 1 0 30728 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1766
timestamp 1623621585
transform 1 0 32568 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  repeater714
timestamp 1623621585
transform 1 0 33028 0 -1 106080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_190_334
timestamp 1623621585
transform 1 0 31832 0 -1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_190_343
timestamp 1623621585
transform 1 0 32660 0 -1 106080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_190_353
timestamp 1623621585
transform 1 0 33580 0 -1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_4  _594_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 34500 0 -1 106080
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_190_361
timestamp 1623621585
transform 1 0 34316 0 -1 106080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_190_374
timestamp 1623621585
transform 1 0 35512 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input290
timestamp 1623621585
transform 1 0 37076 0 -1 106080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_190_386
timestamp 1623621585
transform 1 0 36616 0 -1 106080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_190_390
timestamp 1623621585
transform 1 0 36984 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_190_395
timestamp 1623621585
transform 1 0 37444 0 -1 106080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_381
timestamp 1623621585
transform -1 0 38824 0 -1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1767
timestamp 1623621585
transform 1 0 37812 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_190_400
timestamp 1623621585
transform 1 0 37904 0 -1 106080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_406
timestamp 1623621585
transform 1 0 38456 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_382
timestamp 1623621585
transform 1 0 1104 0 1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_384
timestamp 1623621585
transform 1 0 1104 0 -1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output620
timestamp 1623621585
transform 1 0 1748 0 -1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_191_3
timestamp 1623621585
transform 1 0 1380 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_15
timestamp 1623621585
transform 1 0 2484 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_192_3
timestamp 1623621585
transform 1 0 1380 0 -1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_192_11
timestamp 1623621585
transform 1 0 2116 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1768
timestamp 1623621585
transform 1 0 3772 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_191_27
timestamp 1623621585
transform 1 0 3588 0 1 106080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_191_30
timestamp 1623621585
transform 1 0 3864 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_23
timestamp 1623621585
transform 1 0 3220 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_35
timestamp 1623621585
transform 1 0 4324 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1775
timestamp 1623621585
transform 1 0 6348 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_42
timestamp 1623621585
transform 1 0 4968 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_54
timestamp 1623621585
transform 1 0 6072 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_47
timestamp 1623621585
transform 1 0 5428 0 -1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_192_55
timestamp 1623621585
transform 1 0 6164 0 -1 107168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_192_58
timestamp 1623621585
transform 1 0 6440 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_66
timestamp 1623621585
transform 1 0 7176 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_191_78
timestamp 1623621585
transform 1 0 8280 0 1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_70
timestamp 1623621585
transform 1 0 7544 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_82
timestamp 1623621585
transform 1 0 8648 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1769
timestamp 1623621585
transform 1 0 9016 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_87
timestamp 1623621585
transform 1 0 9108 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_99
timestamp 1623621585
transform 1 0 10212 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_94
timestamp 1623621585
transform 1 0 9752 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1776
timestamp 1623621585
transform 1 0 11592 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_111
timestamp 1623621585
transform 1 0 11316 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_123
timestamp 1623621585
transform 1 0 12420 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_106
timestamp 1623621585
transform 1 0 10856 0 -1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_115
timestamp 1623621585
transform 1 0 11684 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1770
timestamp 1623621585
transform 1 0 14260 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_191_135
timestamp 1623621585
transform 1 0 13524 0 1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_191_144
timestamp 1623621585
transform 1 0 14352 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_127
timestamp 1623621585
transform 1 0 12788 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_139
timestamp 1623621585
transform 1 0 13892 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_156
timestamp 1623621585
transform 1 0 15456 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_151
timestamp 1623621585
transform 1 0 14996 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_163
timestamp 1623621585
transform 1 0 16100 0 -1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1777
timestamp 1623621585
transform 1 0 16836 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_168
timestamp 1623621585
transform 1 0 16560 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_180
timestamp 1623621585
transform 1 0 17664 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_172
timestamp 1623621585
transform 1 0 16928 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_184
timestamp 1623621585
transform 1 0 18032 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1771
timestamp 1623621585
transform 1 0 19504 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_191_192
timestamp 1623621585
transform 1 0 18768 0 1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_191_201
timestamp 1623621585
transform 1 0 19596 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_196
timestamp 1623621585
transform 1 0 19136 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_208
timestamp 1623621585
transform 1 0 20240 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1778
timestamp 1623621585
transform 1 0 22080 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_213
timestamp 1623621585
transform 1 0 20700 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_225
timestamp 1623621585
transform 1 0 21804 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_220
timestamp 1623621585
transform 1 0 21344 0 -1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_229
timestamp 1623621585
transform 1 0 22172 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_237
timestamp 1623621585
transform 1 0 22908 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_191_249
timestamp 1623621585
transform 1 0 24012 0 1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_241
timestamp 1623621585
transform 1 0 23276 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1772
timestamp 1623621585
transform 1 0 24748 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_258
timestamp 1623621585
transform 1 0 24840 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_270
timestamp 1623621585
transform 1 0 25944 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_253
timestamp 1623621585
transform 1 0 24380 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_265
timestamp 1623621585
transform 1 0 25484 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1779
timestamp 1623621585
transform 1 0 27324 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_282
timestamp 1623621585
transform 1 0 27048 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_277
timestamp 1623621585
transform 1 0 26588 0 -1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_286
timestamp 1623621585
transform 1 0 27416 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_294
timestamp 1623621585
transform 1 0 28152 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_191_306
timestamp 1623621585
transform 1 0 29256 0 1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_298
timestamp 1623621585
transform 1 0 28520 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_310
timestamp 1623621585
transform 1 0 29624 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1773
timestamp 1623621585
transform 1 0 29992 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_315
timestamp 1623621585
transform 1 0 30084 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_327
timestamp 1623621585
transform 1 0 31188 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_322
timestamp 1623621585
transform 1 0 30728 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1780
timestamp 1623621585
transform 1 0 32568 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_339
timestamp 1623621585
transform 1 0 32292 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_351
timestamp 1623621585
transform 1 0 33396 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_334
timestamp 1623621585
transform 1 0 31832 0 -1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_343
timestamp 1623621585
transform 1 0 32660 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1774
timestamp 1623621585
transform 1 0 35236 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_191_363
timestamp 1623621585
transform 1 0 34500 0 1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_191_372
timestamp 1623621585
transform 1 0 35328 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_355
timestamp 1623621585
transform 1 0 33764 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_367
timestamp 1623621585
transform 1 0 34868 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input292
timestamp 1623621585
transform 1 0 37076 0 -1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_191_384
timestamp 1623621585
transform 1 0 36432 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_379
timestamp 1623621585
transform 1 0 35972 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_192_395
timestamp 1623621585
transform 1 0 37444 0 -1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_383
timestamp 1623621585
transform -1 0 38824 0 1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_385
timestamp 1623621585
transform -1 0 38824 0 -1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1781
timestamp 1623621585
transform 1 0 37812 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input291
timestamp 1623621585
transform 1 0 37812 0 1 106080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_191_396
timestamp 1623621585
transform 1 0 37536 0 1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_191_403
timestamp 1623621585
transform 1 0 38180 0 1 106080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_192_400
timestamp 1623621585
transform 1 0 37904 0 -1 107168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_406
timestamp 1623621585
transform 1 0 38456 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_386
timestamp 1623621585
transform 1 0 1104 0 1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output662
timestamp 1623621585
transform 1 0 1748 0 1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_193_3
timestamp 1623621585
transform 1 0 1380 0 1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_193_11
timestamp 1623621585
transform 1 0 2116 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1782
timestamp 1623621585
transform 1 0 3772 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_193_23
timestamp 1623621585
transform 1 0 3220 0 1 107168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_193_30
timestamp 1623621585
transform 1 0 3864 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_42
timestamp 1623621585
transform 1 0 4968 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_54
timestamp 1623621585
transform 1 0 6072 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_66
timestamp 1623621585
transform 1 0 7176 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_193_78
timestamp 1623621585
transform 1 0 8280 0 1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1783
timestamp 1623621585
transform 1 0 9016 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_87
timestamp 1623621585
transform 1 0 9108 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_99
timestamp 1623621585
transform 1 0 10212 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_111
timestamp 1623621585
transform 1 0 11316 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_123
timestamp 1623621585
transform 1 0 12420 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1784
timestamp 1623621585
transform 1 0 14260 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_193_135
timestamp 1623621585
transform 1 0 13524 0 1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_193_144
timestamp 1623621585
transform 1 0 14352 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_156
timestamp 1623621585
transform 1 0 15456 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_168
timestamp 1623621585
transform 1 0 16560 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_180
timestamp 1623621585
transform 1 0 17664 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1785
timestamp 1623621585
transform 1 0 19504 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_193_192
timestamp 1623621585
transform 1 0 18768 0 1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_193_201
timestamp 1623621585
transform 1 0 19596 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_213
timestamp 1623621585
transform 1 0 20700 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_225
timestamp 1623621585
transform 1 0 21804 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_237
timestamp 1623621585
transform 1 0 22908 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_193_249
timestamp 1623621585
transform 1 0 24012 0 1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1786
timestamp 1623621585
transform 1 0 24748 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_258
timestamp 1623621585
transform 1 0 24840 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_270
timestamp 1623621585
transform 1 0 25944 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_282
timestamp 1623621585
transform 1 0 27048 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_294
timestamp 1623621585
transform 1 0 28152 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_193_306
timestamp 1623621585
transform 1 0 29256 0 1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1787
timestamp 1623621585
transform 1 0 29992 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_315
timestamp 1623621585
transform 1 0 30084 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_327
timestamp 1623621585
transform 1 0 31188 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _591_
timestamp 1623621585
transform 1 0 32936 0 1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_193_339
timestamp 1623621585
transform 1 0 32292 0 1 107168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_345
timestamp 1623621585
transform 1 0 32844 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_349
timestamp 1623621585
transform 1 0 33212 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1788
timestamp 1623621585
transform 1 0 35236 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_193_361
timestamp 1623621585
transform 1 0 34316 0 1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_193_369
timestamp 1623621585
transform 1 0 35052 0 1 107168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_193_372
timestamp 1623621585
transform 1 0 35328 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input294
timestamp 1623621585
transform 1 0 37076 0 1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_193_384
timestamp 1623621585
transform 1 0 36432 0 1 107168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_390
timestamp 1623621585
transform 1 0 36984 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_193_395
timestamp 1623621585
transform 1 0 37444 0 1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_387
timestamp 1623621585
transform -1 0 38824 0 1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input293
timestamp 1623621585
transform 1 0 37812 0 1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_193_403
timestamp 1623621585
transform 1 0 38180 0 1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_388
timestamp 1623621585
transform 1 0 1104 0 -1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output621
timestamp 1623621585
transform 1 0 1748 0 -1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_194_3
timestamp 1623621585
transform 1 0 1380 0 -1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_194_11
timestamp 1623621585
transform 1 0 2116 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_23
timestamp 1623621585
transform 1 0 3220 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_35
timestamp 1623621585
transform 1 0 4324 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1789
timestamp 1623621585
transform 1 0 6348 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_194_47
timestamp 1623621585
transform 1 0 5428 0 -1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_194_55
timestamp 1623621585
transform 1 0 6164 0 -1 108256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_194_58
timestamp 1623621585
transform 1 0 6440 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_70
timestamp 1623621585
transform 1 0 7544 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_82
timestamp 1623621585
transform 1 0 8648 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_94
timestamp 1623621585
transform 1 0 9752 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1790
timestamp 1623621585
transform 1 0 11592 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_194_106
timestamp 1623621585
transform 1 0 10856 0 -1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_194_115
timestamp 1623621585
transform 1 0 11684 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_127
timestamp 1623621585
transform 1 0 12788 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_139
timestamp 1623621585
transform 1 0 13892 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_151
timestamp 1623621585
transform 1 0 14996 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_194_163
timestamp 1623621585
transform 1 0 16100 0 -1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1791
timestamp 1623621585
transform 1 0 16836 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_172
timestamp 1623621585
transform 1 0 16928 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_184
timestamp 1623621585
transform 1 0 18032 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_196
timestamp 1623621585
transform 1 0 19136 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_208
timestamp 1623621585
transform 1 0 20240 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1792
timestamp 1623621585
transform 1 0 22080 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_194_220
timestamp 1623621585
transform 1 0 21344 0 -1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_194_229
timestamp 1623621585
transform 1 0 22172 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_241
timestamp 1623621585
transform 1 0 23276 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_253
timestamp 1623621585
transform 1 0 24380 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_265
timestamp 1623621585
transform 1 0 25484 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1793
timestamp 1623621585
transform 1 0 27324 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_194_277
timestamp 1623621585
transform 1 0 26588 0 -1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_194_286
timestamp 1623621585
transform 1 0 27416 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_298
timestamp 1623621585
transform 1 0 28520 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_310
timestamp 1623621585
transform 1 0 29624 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_322
timestamp 1623621585
transform 1 0 30728 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _589_
timestamp 1623621585
transform 1 0 33304 0 -1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1794
timestamp 1623621585
transform 1 0 32568 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_194_334
timestamp 1623621585
transform 1 0 31832 0 -1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_194_343
timestamp 1623621585
transform 1 0 32660 0 -1 108256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_349
timestamp 1623621585
transform 1 0 33212 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_354
timestamp 1623621585
transform 1 0 33672 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_366
timestamp 1623621585
transform 1 0 34776 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input295
timestamp 1623621585
transform 1 0 37076 0 -1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_194_378
timestamp 1623621585
transform 1 0 35880 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_194_390
timestamp 1623621585
transform 1 0 36984 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_194_395
timestamp 1623621585
transform 1 0 37444 0 -1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_389
timestamp 1623621585
transform -1 0 38824 0 -1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1795
timestamp 1623621585
transform 1 0 37812 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_194_400
timestamp 1623621585
transform 1 0 37904 0 -1 108256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_406
timestamp 1623621585
transform 1 0 38456 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_390
timestamp 1623621585
transform 1 0 1104 0 1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_195_3
timestamp 1623621585
transform 1 0 1380 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_15
timestamp 1623621585
transform 1 0 2484 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1796
timestamp 1623621585
transform 1 0 3772 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_195_27
timestamp 1623621585
transform 1 0 3588 0 1 108256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_195_30
timestamp 1623621585
transform 1 0 3864 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_42
timestamp 1623621585
transform 1 0 4968 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_54
timestamp 1623621585
transform 1 0 6072 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_66
timestamp 1623621585
transform 1 0 7176 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_195_78
timestamp 1623621585
transform 1 0 8280 0 1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1797
timestamp 1623621585
transform 1 0 9016 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_87
timestamp 1623621585
transform 1 0 9108 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_99
timestamp 1623621585
transform 1 0 10212 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_111
timestamp 1623621585
transform 1 0 11316 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_195_123
timestamp 1623621585
transform 1 0 12420 0 1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _744_
timestamp 1623621585
transform 1 0 12880 0 1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1798
timestamp 1623621585
transform 1 0 14260 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_195_127
timestamp 1623621585
transform 1 0 12788 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_131
timestamp 1623621585
transform 1 0 13156 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_144
timestamp 1623621585
transform 1 0 14352 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_156
timestamp 1623621585
transform 1 0 15456 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_168
timestamp 1623621585
transform 1 0 16560 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_180
timestamp 1623621585
transform 1 0 17664 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1799
timestamp 1623621585
transform 1 0 19504 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_195_192
timestamp 1623621585
transform 1 0 18768 0 1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_195_201
timestamp 1623621585
transform 1 0 19596 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_213
timestamp 1623621585
transform 1 0 20700 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_225
timestamp 1623621585
transform 1 0 21804 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_237
timestamp 1623621585
transform 1 0 22908 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_195_249
timestamp 1623621585
transform 1 0 24012 0 1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1800
timestamp 1623621585
transform 1 0 24748 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_258
timestamp 1623621585
transform 1 0 24840 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_270
timestamp 1623621585
transform 1 0 25944 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_282
timestamp 1623621585
transform 1 0 27048 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _735_
timestamp 1623621585
transform 1 0 28520 0 1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_195_294
timestamp 1623621585
transform 1 0 28152 0 1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_195_301
timestamp 1623621585
transform 1 0 28796 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1801
timestamp 1623621585
transform 1 0 29992 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_195_313
timestamp 1623621585
transform 1 0 29900 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_315
timestamp 1623621585
transform 1 0 30084 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_327
timestamp 1623621585
transform 1 0 31188 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 33120 0 1 108256
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_195_339
timestamp 1623621585
transform 1 0 32292 0 1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_195_347
timestamp 1623621585
transform 1 0 33028 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _593_
timestamp 1623621585
transform 1 0 34132 0 1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1802
timestamp 1623621585
transform 1 0 35236 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_195_355
timestamp 1623621585
transform 1 0 33764 0 1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_195_363
timestamp 1623621585
transform 1 0 34500 0 1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_195_372
timestamp 1623621585
transform 1 0 35328 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_384
timestamp 1623621585
transform 1 0 36432 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_391
timestamp 1623621585
transform -1 0 38824 0 1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input296
timestamp 1623621585
transform 1 0 37812 0 1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_195_396
timestamp 1623621585
transform 1 0 37536 0 1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_195_403
timestamp 1623621585
transform 1 0 38180 0 1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_392
timestamp 1623621585
transform 1 0 1104 0 -1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input57
timestamp 1623621585
transform 1 0 1748 0 -1 109344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_196_3
timestamp 1623621585
transform 1 0 1380 0 -1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_196_13
timestamp 1623621585
transform 1 0 2300 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_25
timestamp 1623621585
transform 1 0 3404 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_37
timestamp 1623621585
transform 1 0 4508 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1803
timestamp 1623621585
transform 1 0 6348 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_196_49
timestamp 1623621585
transform 1 0 5612 0 -1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_196_58
timestamp 1623621585
transform 1 0 6440 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_70
timestamp 1623621585
transform 1 0 7544 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_82
timestamp 1623621585
transform 1 0 8648 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_94
timestamp 1623621585
transform 1 0 9752 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1804
timestamp 1623621585
transform 1 0 11592 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_196_106
timestamp 1623621585
transform 1 0 10856 0 -1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_196_115
timestamp 1623621585
transform 1 0 11684 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_127
timestamp 1623621585
transform 1 0 12788 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_139
timestamp 1623621585
transform 1 0 13892 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_151
timestamp 1623621585
transform 1 0 14996 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_196_163
timestamp 1623621585
transform 1 0 16100 0 -1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1805
timestamp 1623621585
transform 1 0 16836 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_172
timestamp 1623621585
transform 1 0 16928 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_184
timestamp 1623621585
transform 1 0 18032 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_196
timestamp 1623621585
transform 1 0 19136 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_208
timestamp 1623621585
transform 1 0 20240 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1806
timestamp 1623621585
transform 1 0 22080 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_196_220
timestamp 1623621585
transform 1 0 21344 0 -1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_196_229
timestamp 1623621585
transform 1 0 22172 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_241
timestamp 1623621585
transform 1 0 23276 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_253
timestamp 1623621585
transform 1 0 24380 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_265
timestamp 1623621585
transform 1 0 25484 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1807
timestamp 1623621585
transform 1 0 27324 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_196_277
timestamp 1623621585
transform 1 0 26588 0 -1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_196_286
timestamp 1623621585
transform 1 0 27416 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_298
timestamp 1623621585
transform 1 0 28520 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_310
timestamp 1623621585
transform 1 0 29624 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_322
timestamp 1623621585
transform 1 0 30728 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1808
timestamp 1623621585
transform 1 0 32568 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_196_334
timestamp 1623621585
transform 1 0 31832 0 -1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_196_343
timestamp 1623621585
transform 1 0 32660 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_1  _607_
timestamp 1623621585
transform 1 0 33764 0 -1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_196_363
timestamp 1623621585
transform 1 0 34500 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_375
timestamp 1623621585
transform 1 0 35604 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  input297
timestamp 1623621585
transform 1 0 37076 0 -1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_196_387
timestamp 1623621585
transform 1 0 36708 0 -1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_196_395
timestamp 1623621585
transform 1 0 37444 0 -1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_393
timestamp 1623621585
transform -1 0 38824 0 -1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1809
timestamp 1623621585
transform 1 0 37812 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_196_400
timestamp 1623621585
transform 1 0 37904 0 -1 109344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_406
timestamp 1623621585
transform 1 0 38456 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_394
timestamp 1623621585
transform 1 0 1104 0 1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output622
timestamp 1623621585
transform 1 0 1748 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_197_3
timestamp 1623621585
transform 1 0 1380 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_197_11
timestamp 1623621585
transform 1 0 2116 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1810
timestamp 1623621585
transform 1 0 3772 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_197_23
timestamp 1623621585
transform 1 0 3220 0 1 109344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_197_30
timestamp 1623621585
transform 1 0 3864 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_42
timestamp 1623621585
transform 1 0 4968 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_54
timestamp 1623621585
transform 1 0 6072 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_66
timestamp 1623621585
transform 1 0 7176 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_197_78
timestamp 1623621585
transform 1 0 8280 0 1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1811
timestamp 1623621585
transform 1 0 9016 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_87
timestamp 1623621585
transform 1 0 9108 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_99
timestamp 1623621585
transform 1 0 10212 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_111
timestamp 1623621585
transform 1 0 11316 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_123
timestamp 1623621585
transform 1 0 12420 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1812
timestamp 1623621585
transform 1 0 14260 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_197_135
timestamp 1623621585
transform 1 0 13524 0 1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_197_144
timestamp 1623621585
transform 1 0 14352 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_156
timestamp 1623621585
transform 1 0 15456 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_168
timestamp 1623621585
transform 1 0 16560 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_180
timestamp 1623621585
transform 1 0 17664 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1813
timestamp 1623621585
transform 1 0 19504 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_197_192
timestamp 1623621585
transform 1 0 18768 0 1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_197_201
timestamp 1623621585
transform 1 0 19596 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_213
timestamp 1623621585
transform 1 0 20700 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_225
timestamp 1623621585
transform 1 0 21804 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_237
timestamp 1623621585
transform 1 0 22908 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_197_249
timestamp 1623621585
transform 1 0 24012 0 1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1814
timestamp 1623621585
transform 1 0 24748 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_258
timestamp 1623621585
transform 1 0 24840 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_270
timestamp 1623621585
transform 1 0 25944 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_282
timestamp 1623621585
transform 1 0 27048 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_294
timestamp 1623621585
transform 1 0 28152 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_197_306
timestamp 1623621585
transform 1 0 29256 0 1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1815
timestamp 1623621585
transform 1 0 29992 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_315
timestamp 1623621585
transform 1 0 30084 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_327
timestamp 1623621585
transform 1 0 31188 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__nor4_2  _585_
timestamp 1623621585
transform 1 0 32660 0 1 109344
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_197_339
timestamp 1623621585
transform 1 0 32292 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_197_353
timestamp 1623621585
transform 1 0 33580 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _608_
timestamp 1623621585
transform 1 0 33948 0 1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1816
timestamp 1623621585
transform 1 0 35236 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_197_365
timestamp 1623621585
transform 1 0 34684 0 1 109344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_197_372
timestamp 1623621585
transform 1 0 35328 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  input300
timestamp 1623621585
transform 1 0 37076 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_197_384
timestamp 1623621585
transform 1 0 36432 0 1 109344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_390
timestamp 1623621585
transform 1 0 36984 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_197_395
timestamp 1623621585
transform 1 0 37444 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_395
timestamp 1623621585
transform -1 0 38824 0 1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input299
timestamp 1623621585
transform 1 0 37812 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_197_403
timestamp 1623621585
transform 1 0 38180 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_396
timestamp 1623621585
transform 1 0 1104 0 -1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_398
timestamp 1623621585
transform 1 0 1104 0 1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output624
timestamp 1623621585
transform 1 0 1748 0 1 110432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_198_3
timestamp 1623621585
transform 1 0 1380 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_15
timestamp 1623621585
transform 1 0 2484 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_199_3
timestamp 1623621585
transform 1 0 1380 0 1 110432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_199_11
timestamp 1623621585
transform 1 0 2116 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1824
timestamp 1623621585
transform 1 0 3772 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_27
timestamp 1623621585
transform 1 0 3588 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_39
timestamp 1623621585
transform 1 0 4692 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_23
timestamp 1623621585
transform 1 0 3220 0 1 110432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_199_30
timestamp 1623621585
transform 1 0 3864 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1817
timestamp 1623621585
transform 1 0 6348 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_198_51
timestamp 1623621585
transform 1 0 5796 0 -1 110432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_198_58
timestamp 1623621585
transform 1 0 6440 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_42
timestamp 1623621585
transform 1 0 4968 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_54
timestamp 1623621585
transform 1 0 6072 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_70
timestamp 1623621585
transform 1 0 7544 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_82
timestamp 1623621585
transform 1 0 8648 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_66
timestamp 1623621585
transform 1 0 7176 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_78
timestamp 1623621585
transform 1 0 8280 0 1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1825
timestamp 1623621585
transform 1 0 9016 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_94
timestamp 1623621585
transform 1 0 9752 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_87
timestamp 1623621585
transform 1 0 9108 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_99
timestamp 1623621585
transform 1 0 10212 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1818
timestamp 1623621585
transform 1 0 11592 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_198_106
timestamp 1623621585
transform 1 0 10856 0 -1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_198_115
timestamp 1623621585
transform 1 0 11684 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_111
timestamp 1623621585
transform 1 0 11316 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_123
timestamp 1623621585
transform 1 0 12420 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1826
timestamp 1623621585
transform 1 0 14260 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_127
timestamp 1623621585
transform 1 0 12788 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_139
timestamp 1623621585
transform 1 0 13892 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_135
timestamp 1623621585
transform 1 0 13524 0 1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_199_144
timestamp 1623621585
transform 1 0 14352 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_151
timestamp 1623621585
transform 1 0 14996 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_198_163
timestamp 1623621585
transform 1 0 16100 0 -1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_199_156
timestamp 1623621585
transform 1 0 15456 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1819
timestamp 1623621585
transform 1 0 16836 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_172
timestamp 1623621585
transform 1 0 16928 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_184
timestamp 1623621585
transform 1 0 18032 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_168
timestamp 1623621585
transform 1 0 16560 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_180
timestamp 1623621585
transform 1 0 17664 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1827
timestamp 1623621585
transform 1 0 19504 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_196
timestamp 1623621585
transform 1 0 19136 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_208
timestamp 1623621585
transform 1 0 20240 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_192
timestamp 1623621585
transform 1 0 18768 0 1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_199_201
timestamp 1623621585
transform 1 0 19596 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1820
timestamp 1623621585
transform 1 0 22080 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_198_220
timestamp 1623621585
transform 1 0 21344 0 -1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_198_229
timestamp 1623621585
transform 1 0 22172 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_213
timestamp 1623621585
transform 1 0 20700 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_225
timestamp 1623621585
transform 1 0 21804 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_241
timestamp 1623621585
transform 1 0 23276 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_237
timestamp 1623621585
transform 1 0 22908 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_249
timestamp 1623621585
transform 1 0 24012 0 1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1828
timestamp 1623621585
transform 1 0 24748 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_253
timestamp 1623621585
transform 1 0 24380 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_265
timestamp 1623621585
transform 1 0 25484 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_258
timestamp 1623621585
transform 1 0 24840 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_270
timestamp 1623621585
transform 1 0 25944 0 1 110432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _731_
timestamp 1623621585
transform 1 0 26588 0 1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1821
timestamp 1623621585
transform 1 0 27324 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_198_277
timestamp 1623621585
transform 1 0 26588 0 -1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_198_286
timestamp 1623621585
transform 1 0 27416 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_199_276
timestamp 1623621585
transform 1 0 26496 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_280
timestamp 1623621585
transform 1 0 26864 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_298
timestamp 1623621585
transform 1 0 28520 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_310
timestamp 1623621585
transform 1 0 29624 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_292
timestamp 1623621585
transform 1 0 27968 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_304
timestamp 1623621585
transform 1 0 29072 0 1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_199_312
timestamp 1623621585
transform 1 0 29808 0 1 110432
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1829
timestamp 1623621585
transform 1 0 29992 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_322
timestamp 1623621585
transform 1 0 30728 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_315
timestamp 1623621585
transform 1 0 30084 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_327
timestamp 1623621585
transform 1 0 31188 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1822
timestamp 1623621585
transform 1 0 32568 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_198_334
timestamp 1623621585
transform 1 0 31832 0 -1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_198_343
timestamp 1623621585
transform 1 0 32660 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_339
timestamp 1623621585
transform 1 0 32292 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_351
timestamp 1623621585
transform 1 0 33396 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1830
timestamp 1623621585
transform 1 0 35236 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_355
timestamp 1623621585
transform 1 0 33764 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_367
timestamp 1623621585
transform 1 0 34868 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_363
timestamp 1623621585
transform 1 0 34500 0 1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_199_372
timestamp 1623621585
transform 1 0 35328 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  input301
timestamp 1623621585
transform 1 0 37076 0 -1 110432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_198_379
timestamp 1623621585
transform 1 0 35972 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_198_395
timestamp 1623621585
transform 1 0 37444 0 -1 110432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_199_384
timestamp 1623621585
transform 1 0 36432 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_397
timestamp 1623621585
transform -1 0 38824 0 -1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_399
timestamp 1623621585
transform -1 0 38824 0 1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1823
timestamp 1623621585
transform 1 0 37812 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input302
timestamp 1623621585
transform 1 0 37812 0 1 110432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_198_400
timestamp 1623621585
transform 1 0 37904 0 -1 110432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_406
timestamp 1623621585
transform 1 0 38456 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_199_396
timestamp 1623621585
transform 1 0 37536 0 1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_199_403
timestamp 1623621585
transform 1 0 38180 0 1 110432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_400
timestamp 1623621585
transform 1 0 1104 0 -1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output668
timestamp 1623621585
transform 1 0 1748 0 -1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_200_3
timestamp 1623621585
transform 1 0 1380 0 -1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_200_11
timestamp 1623621585
transform 1 0 2116 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_23
timestamp 1623621585
transform 1 0 3220 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_35
timestamp 1623621585
transform 1 0 4324 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1831
timestamp 1623621585
transform 1 0 6348 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_200_47
timestamp 1623621585
transform 1 0 5428 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_200_55
timestamp 1623621585
transform 1 0 6164 0 -1 111520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_200_58
timestamp 1623621585
transform 1 0 6440 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_70
timestamp 1623621585
transform 1 0 7544 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_82
timestamp 1623621585
transform 1 0 8648 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_94
timestamp 1623621585
transform 1 0 9752 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1832
timestamp 1623621585
transform 1 0 11592 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_200_106
timestamp 1623621585
transform 1 0 10856 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_200_115
timestamp 1623621585
transform 1 0 11684 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_127
timestamp 1623621585
transform 1 0 12788 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_139
timestamp 1623621585
transform 1 0 13892 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_151
timestamp 1623621585
transform 1 0 14996 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_200_163
timestamp 1623621585
transform 1 0 16100 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1833
timestamp 1623621585
transform 1 0 16836 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_172
timestamp 1623621585
transform 1 0 16928 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_184
timestamp 1623621585
transform 1 0 18032 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_196
timestamp 1623621585
transform 1 0 19136 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_208
timestamp 1623621585
transform 1 0 20240 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1834
timestamp 1623621585
transform 1 0 22080 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_200_220
timestamp 1623621585
transform 1 0 21344 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_200_229
timestamp 1623621585
transform 1 0 22172 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_241
timestamp 1623621585
transform 1 0 23276 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_253
timestamp 1623621585
transform 1 0 24380 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_265
timestamp 1623621585
transform 1 0 25484 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1835
timestamp 1623621585
transform 1 0 27324 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_200_277
timestamp 1623621585
transform 1 0 26588 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_200_286
timestamp 1623621585
transform 1 0 27416 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_298
timestamp 1623621585
transform 1 0 28520 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_310
timestamp 1623621585
transform 1 0 29624 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_322
timestamp 1623621585
transform 1 0 30728 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1836
timestamp 1623621585
transform 1 0 32568 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_200_334
timestamp 1623621585
transform 1 0 31832 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_200_343
timestamp 1623621585
transform 1 0 32660 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_1  _598_
timestamp 1623621585
transform 1 0 35328 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_200_355
timestamp 1623621585
transform 1 0 33764 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_200_367
timestamp 1623621585
transform 1 0 34868 0 -1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_200_371
timestamp 1623621585
transform 1 0 35236 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input303
timestamp 1623621585
transform 1 0 37076 0 -1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_200_380
timestamp 1623621585
transform 1 0 36064 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_200_388
timestamp 1623621585
transform 1 0 36800 0 -1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_200_395
timestamp 1623621585
transform 1 0 37444 0 -1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_401
timestamp 1623621585
transform -1 0 38824 0 -1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1837
timestamp 1623621585
transform 1 0 37812 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_200_400
timestamp 1623621585
transform 1 0 37904 0 -1 111520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_406
timestamp 1623621585
transform 1 0 38456 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_402
timestamp 1623621585
transform 1 0 1104 0 1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_201_3
timestamp 1623621585
transform 1 0 1380 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_15
timestamp 1623621585
transform 1 0 2484 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1838
timestamp 1623621585
transform 1 0 3772 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_201_27
timestamp 1623621585
transform 1 0 3588 0 1 111520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_201_30
timestamp 1623621585
transform 1 0 3864 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_42
timestamp 1623621585
transform 1 0 4968 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_54
timestamp 1623621585
transform 1 0 6072 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_66
timestamp 1623621585
transform 1 0 7176 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_201_78
timestamp 1623621585
transform 1 0 8280 0 1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1839
timestamp 1623621585
transform 1 0 9016 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_87
timestamp 1623621585
transform 1 0 9108 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_99
timestamp 1623621585
transform 1 0 10212 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_111
timestamp 1623621585
transform 1 0 11316 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_123
timestamp 1623621585
transform 1 0 12420 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1840
timestamp 1623621585
transform 1 0 14260 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_201_135
timestamp 1623621585
transform 1 0 13524 0 1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_201_144
timestamp 1623621585
transform 1 0 14352 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_156
timestamp 1623621585
transform 1 0 15456 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_168
timestamp 1623621585
transform 1 0 16560 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_180
timestamp 1623621585
transform 1 0 17664 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1841
timestamp 1623621585
transform 1 0 19504 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_201_192
timestamp 1623621585
transform 1 0 18768 0 1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_201_201
timestamp 1623621585
transform 1 0 19596 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_213
timestamp 1623621585
transform 1 0 20700 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_225
timestamp 1623621585
transform 1 0 21804 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_237
timestamp 1623621585
transform 1 0 22908 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_201_249
timestamp 1623621585
transform 1 0 24012 0 1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1842
timestamp 1623621585
transform 1 0 24748 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_258
timestamp 1623621585
transform 1 0 24840 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_270
timestamp 1623621585
transform 1 0 25944 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_282
timestamp 1623621585
transform 1 0 27048 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_294
timestamp 1623621585
transform 1 0 28152 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_201_306
timestamp 1623621585
transform 1 0 29256 0 1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1843
timestamp 1623621585
transform 1 0 29992 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_315
timestamp 1623621585
transform 1 0 30084 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_327
timestamp 1623621585
transform 1 0 31188 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_339
timestamp 1623621585
transform 1 0 32292 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_351
timestamp 1623621585
transform 1 0 33396 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1844
timestamp 1623621585
transform 1 0 35236 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_201_363
timestamp 1623621585
transform 1 0 34500 0 1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_201_372
timestamp 1623621585
transform 1 0 35328 0 1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _606_
timestamp 1623621585
transform 1 0 35696 0 1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input305
timestamp 1623621585
transform 1 0 37076 0 1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_201_384
timestamp 1623621585
transform 1 0 36432 0 1 111520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_390
timestamp 1623621585
transform 1 0 36984 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_201_395
timestamp 1623621585
transform 1 0 37444 0 1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_403
timestamp 1623621585
transform -1 0 38824 0 1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input304
timestamp 1623621585
transform 1 0 37812 0 1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_201_403
timestamp 1623621585
transform 1 0 38180 0 1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_404
timestamp 1623621585
transform 1 0 1104 0 -1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output670
timestamp 1623621585
transform 1 0 1748 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_202_3
timestamp 1623621585
transform 1 0 1380 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_202_11
timestamp 1623621585
transform 1 0 2116 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_23
timestamp 1623621585
transform 1 0 3220 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_35
timestamp 1623621585
transform 1 0 4324 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1845
timestamp 1623621585
transform 1 0 6348 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_202_47
timestamp 1623621585
transform 1 0 5428 0 -1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_202_55
timestamp 1623621585
transform 1 0 6164 0 -1 112608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_202_58
timestamp 1623621585
transform 1 0 6440 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_70
timestamp 1623621585
transform 1 0 7544 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_82
timestamp 1623621585
transform 1 0 8648 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_94
timestamp 1623621585
transform 1 0 9752 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1846
timestamp 1623621585
transform 1 0 11592 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_202_106
timestamp 1623621585
transform 1 0 10856 0 -1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_202_115
timestamp 1623621585
transform 1 0 11684 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_127
timestamp 1623621585
transform 1 0 12788 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_139
timestamp 1623621585
transform 1 0 13892 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_151
timestamp 1623621585
transform 1 0 14996 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_202_163
timestamp 1623621585
transform 1 0 16100 0 -1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1847
timestamp 1623621585
transform 1 0 16836 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_172
timestamp 1623621585
transform 1 0 16928 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_184
timestamp 1623621585
transform 1 0 18032 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_196
timestamp 1623621585
transform 1 0 19136 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_208
timestamp 1623621585
transform 1 0 20240 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1848
timestamp 1623621585
transform 1 0 22080 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_202_220
timestamp 1623621585
transform 1 0 21344 0 -1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_202_229
timestamp 1623621585
transform 1 0 22172 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_241
timestamp 1623621585
transform 1 0 23276 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_253
timestamp 1623621585
transform 1 0 24380 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_265
timestamp 1623621585
transform 1 0 25484 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1849
timestamp 1623621585
transform 1 0 27324 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_202_277
timestamp 1623621585
transform 1 0 26588 0 -1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_202_286
timestamp 1623621585
transform 1 0 27416 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_298
timestamp 1623621585
transform 1 0 28520 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_310
timestamp 1623621585
transform 1 0 29624 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_322
timestamp 1623621585
transform 1 0 30728 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1850
timestamp 1623621585
transform 1 0 32568 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_202_334
timestamp 1623621585
transform 1 0 31832 0 -1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_202_343
timestamp 1623621585
transform 1 0 32660 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1623621585
transform 1 0 34040 0 -1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_202_355
timestamp 1623621585
transform 1 0 33764 0 -1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_202_361
timestamp 1623621585
transform 1 0 34316 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_202_373
timestamp 1623621585
transform 1 0 35420 0 -1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1623621585
transform 1 0 35696 0 -1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input306
timestamp 1623621585
transform 1 0 37076 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output671
timestamp 1623621585
transform 1 0 36340 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_202_379
timestamp 1623621585
transform 1 0 35972 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_202_387
timestamp 1623621585
transform 1 0 36708 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_202_395
timestamp 1623621585
transform 1 0 37444 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_405
timestamp 1623621585
transform -1 0 38824 0 -1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1851
timestamp 1623621585
transform 1 0 37812 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_202_400
timestamp 1623621585
transform 1 0 37904 0 -1 112608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_406
timestamp 1623621585
transform 1 0 38456 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_406
timestamp 1623621585
transform 1 0 1104 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output627
timestamp 1623621585
transform 1 0 1748 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_203_3
timestamp 1623621585
transform 1 0 1380 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_203_11
timestamp 1623621585
transform 1 0 2116 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1852
timestamp 1623621585
transform 1 0 3772 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_203_23
timestamp 1623621585
transform 1 0 3220 0 1 112608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_203_30
timestamp 1623621585
transform 1 0 3864 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_42
timestamp 1623621585
transform 1 0 4968 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_54
timestamp 1623621585
transform 1 0 6072 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_66
timestamp 1623621585
transform 1 0 7176 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_203_78
timestamp 1623621585
transform 1 0 8280 0 1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1853
timestamp 1623621585
transform 1 0 9016 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_87
timestamp 1623621585
transform 1 0 9108 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_99
timestamp 1623621585
transform 1 0 10212 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_111
timestamp 1623621585
transform 1 0 11316 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_123
timestamp 1623621585
transform 1 0 12420 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1854
timestamp 1623621585
transform 1 0 14260 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_203_135
timestamp 1623621585
transform 1 0 13524 0 1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_203_144
timestamp 1623621585
transform 1 0 14352 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_156
timestamp 1623621585
transform 1 0 15456 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_168
timestamp 1623621585
transform 1 0 16560 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_180
timestamp 1623621585
transform 1 0 17664 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1855
timestamp 1623621585
transform 1 0 19504 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_203_192
timestamp 1623621585
transform 1 0 18768 0 1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_203_201
timestamp 1623621585
transform 1 0 19596 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_213
timestamp 1623621585
transform 1 0 20700 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_225
timestamp 1623621585
transform 1 0 21804 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_237
timestamp 1623621585
transform 1 0 22908 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_203_249
timestamp 1623621585
transform 1 0 24012 0 1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1856
timestamp 1623621585
transform 1 0 24748 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_258
timestamp 1623621585
transform 1 0 24840 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_270
timestamp 1623621585
transform 1 0 25944 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_282
timestamp 1623621585
transform 1 0 27048 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_4  _613_
timestamp 1623621585
transform 1 0 28796 0 1 112608
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_203_294
timestamp 1623621585
transform 1 0 28152 0 1 112608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_300
timestamp 1623621585
transform 1 0 28704 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_203_310
timestamp 1623621585
transform 1 0 29624 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1857
timestamp 1623621585
transform 1 0 29992 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input452
timestamp 1623621585
transform 1 0 31280 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_203_315
timestamp 1623621585
transform 1 0 30084 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_203_327
timestamp 1623621585
transform 1 0 31188 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_203_331
timestamp 1623621585
transform 1 0 31556 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1623621585
transform 1 0 33396 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input453
timestamp 1623621585
transform 1 0 31924 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input454
timestamp 1623621585
transform 1 0 32568 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_203_338
timestamp 1623621585
transform 1 0 32200 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_203_345
timestamp 1623621585
transform 1 0 32844 0 1 112608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_203_354
timestamp 1623621585
transform 1 0 33672 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _596_
timestamp 1623621585
transform 1 0 34040 0 1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1858
timestamp 1623621585
transform 1 0 35236 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_203_366
timestamp 1623621585
transform 1 0 34776 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_203_370
timestamp 1623621585
transform 1 0 35144 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_203_372
timestamp 1623621585
transform 1 0 35328 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1623621585
transform 1 0 35696 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output646
timestamp 1623621585
transform 1 0 37076 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output653
timestamp 1623621585
transform 1 0 36340 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_203_379
timestamp 1623621585
transform 1 0 35972 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_203_387
timestamp 1623621585
transform 1 0 36708 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_203_395
timestamp 1623621585
transform 1 0 37444 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_407
timestamp 1623621585
transform -1 0 38824 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input307
timestamp 1623621585
transform 1 0 37812 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_203_403
timestamp 1623621585
transform 1 0 38180 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_3
timestamp 1623621585
transform 1 0 1380 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_204_3
timestamp 1623621585
transform 1 0 1380 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1623621585
transform 1 0 1748 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_410
timestamp 1623621585
transform 1 0 1104 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_408
timestamp 1623621585
transform 1 0 1104 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_205_11
timestamp 1623621585
transform 1 0 2116 0 1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_204_14
timestamp 1623621585
transform 1 0 2392 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1623621585
transform 1 0 2116 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1623621585
transform 1 0 2760 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _662_
timestamp 1623621585
transform 1 0 2852 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_205_22
timestamp 1623621585
transform 1 0 3128 0 1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_204_21
timestamp 1623621585
transform 1 0 3036 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1623621585
transform 1 0 3404 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_30
timestamp 1623621585
transform 1 0 3864 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_205_28
timestamp 1623621585
transform 1 0 3680 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_204_28
timestamp 1623621585
transform 1 0 3680 0 -1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1623621585
transform 1 0 4232 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1866
timestamp 1623621585
transform 1 0 3772 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _665_
timestamp 1623621585
transform 1 0 4232 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_205_41
timestamp 1623621585
transform 1 0 4876 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_205_37
timestamp 1623621585
transform 1 0 4508 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_37
timestamp 1623621585
transform 1 0 4508 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1623621585
transform 1 0 4876 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_45
timestamp 1623621585
transform 1 0 5244 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_44
timestamp 1623621585
transform 1 0 5152 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1623621585
transform 1 0 5520 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _693_
timestamp 1623621585
transform 1 0 4968 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_52
timestamp 1623621585
transform 1 0 5888 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_204_51
timestamp 1623621585
transform 1 0 5796 0 -1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _667_
timestamp 1623621585
transform 1 0 5612 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_59
timestamp 1623621585
transform 1 0 6532 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_58
timestamp 1623621585
transform 1 0 6440 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1623621585
transform 1 0 6808 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1859
timestamp 1623621585
transform 1 0 6348 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _694_
timestamp 1623621585
transform 1 0 6256 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_66
timestamp 1623621585
transform 1 0 7176 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_65
timestamp 1623621585
transform 1 0 7084 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1623621585
transform 1 0 7452 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _695_
timestamp 1623621585
transform 1 0 6900 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_73
timestamp 1623621585
transform 1 0 7820 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_204_72
timestamp 1623621585
transform 1 0 7728 0 -1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _696_
timestamp 1623621585
transform 1 0 7544 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_205_80
timestamp 1623621585
transform 1 0 8464 0 1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_204_82
timestamp 1623621585
transform 1 0 8648 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_204_78
timestamp 1623621585
transform 1 0 8280 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1623621585
transform 1 0 8372 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _699_
timestamp 1623621585
transform 1 0 8188 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1867
timestamp 1623621585
transform 1 0 9016 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1623621585
transform 1 0 9016 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_204_89
timestamp 1623621585
transform 1 0 9292 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_101
timestamp 1623621585
transform 1 0 10396 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_87
timestamp 1623621585
transform 1 0 9108 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_99
timestamp 1623621585
transform 1 0 10212 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1860
timestamp 1623621585
transform 1 0 11592 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_204_113
timestamp 1623621585
transform 1 0 11500 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_115
timestamp 1623621585
transform 1 0 11684 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_111
timestamp 1623621585
transform 1 0 11316 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_123
timestamp 1623621585
transform 1 0 12420 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1868
timestamp 1623621585
transform 1 0 14260 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_127
timestamp 1623621585
transform 1 0 12788 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_139
timestamp 1623621585
transform 1 0 13892 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_205_135
timestamp 1623621585
transform 1 0 13524 0 1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_205_144
timestamp 1623621585
transform 1 0 14352 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_151
timestamp 1623621585
transform 1 0 14996 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_204_163
timestamp 1623621585
transform 1 0 16100 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_205_156
timestamp 1623621585
transform 1 0 15456 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1861
timestamp 1623621585
transform 1 0 16836 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_172
timestamp 1623621585
transform 1 0 16928 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_184
timestamp 1623621585
transform 1 0 18032 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_168
timestamp 1623621585
transform 1 0 16560 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_180
timestamp 1623621585
transform 1 0 17664 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1869
timestamp 1623621585
transform 1 0 19504 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_196
timestamp 1623621585
transform 1 0 19136 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_208
timestamp 1623621585
transform 1 0 20240 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_205_192
timestamp 1623621585
transform 1 0 18768 0 1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_205_201
timestamp 1623621585
transform 1 0 19596 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1862
timestamp 1623621585
transform 1 0 22080 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1623621585
transform 1 0 21988 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_204_220
timestamp 1623621585
transform 1 0 21344 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_204_229
timestamp 1623621585
transform 1 0 22172 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_213
timestamp 1623621585
transform 1 0 20700 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_205_225
timestamp 1623621585
transform 1 0 21804 0 1 113696
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1623621585
transform 1 0 23368 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_204_241
timestamp 1623621585
transform 1 0 23276 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_230
timestamp 1623621585
transform 1 0 22264 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_245
timestamp 1623621585
transform 1 0 23644 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1870
timestamp 1623621585
transform 1 0 24748 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_253
timestamp 1623621585
transform 1 0 24380 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_265
timestamp 1623621585
transform 1 0 25484 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_258
timestamp 1623621585
transform 1 0 24840 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_205_270
timestamp 1623621585
transform 1 0 25944 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_276
timestamp 1623621585
transform 1 0 26496 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_204_277
timestamp 1623621585
transform 1 0 26588 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1623621585
transform 1 0 26864 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1623621585
transform 1 0 26220 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_205_287
timestamp 1623621585
transform 1 0 27508 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_205_283
timestamp 1623621585
transform 1 0 27140 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1623621585
transform 1 0 27600 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1863
timestamp 1623621585
transform 1 0 27324 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_291
timestamp 1623621585
transform 1 0 27876 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_286
timestamp 1623621585
transform 1 0 27416 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_298
timestamp 1623621585
transform 1 0 28520 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_310
timestamp 1623621585
transform 1 0 29624 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_205_303
timestamp 1623621585
transform 1 0 28980 0 1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_205_311
timestamp 1623621585
transform 1 0 29716 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_315
timestamp 1623621585
transform 1 0 30084 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input448
timestamp 1623621585
transform 1 0 30452 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1871
timestamp 1623621585
transform 1 0 29992 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_205_329
timestamp 1623621585
transform 1 0 31372 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_322
timestamp 1623621585
transform 1 0 30728 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_326
timestamp 1623621585
transform 1 0 31096 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_204_322
timestamp 1623621585
transform 1 0 30728 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input451
timestamp 1623621585
transform 1 0 31464 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input450
timestamp 1623621585
transform 1 0 30820 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input449
timestamp 1623621585
transform 1 0 31096 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_205_333
timestamp 1623621585
transform 1 0 31740 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_204_333
timestamp 1623621585
transform 1 0 31740 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_205_337
timestamp 1623621585
transform 1 0 32108 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1623621585
transform 1 0 31832 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_344
timestamp 1623621585
transform 1 0 32752 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_204_347
timestamp 1623621585
transform 1 0 33028 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_204_343
timestamp 1623621585
transform 1 0 32660 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_204_341
timestamp 1623621585
transform 1 0 32476 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1623621585
transform 1 0 32476 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1864
timestamp 1623621585
transform 1 0 32568 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_205_351
timestamp 1623621585
transform 1 0 33396 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_204_351
timestamp 1623621585
transform 1 0 33396 0 -1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1623621585
transform 1 0 33120 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1623621585
transform 1 0 33120 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_359
timestamp 1623621585
transform 1 0 34132 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_205_355
timestamp 1623621585
transform 1 0 33764 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output663
timestamp 1623621585
transform 1 0 34500 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1623621585
transform 1 0 33856 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _599_
timestamp 1623621585
transform 1 0 33948 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_205_367
timestamp 1623621585
transform 1 0 34868 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_204_365
timestamp 1623621585
transform 1 0 34684 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1872
timestamp 1623621585
transform 1 0 35236 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_205_372
timestamp 1623621585
transform 1 0 35328 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_204_373
timestamp 1623621585
transform 1 0 35420 0 -1 113696
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output661
timestamp 1623621585
transform 1 0 35604 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _604_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 35696 0 1 113696
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  input308
timestamp 1623621585
transform 1 0 37076 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output644
timestamp 1623621585
transform 1 0 36340 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_379
timestamp 1623621585
transform 1 0 35972 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_387
timestamp 1623621585
transform 1 0 36708 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_395
timestamp 1623621585
transform 1 0 37444 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_205_389
timestamp 1623621585
transform 1 0 36892 0 1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_409
timestamp 1623621585
transform -1 0 38824 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_411
timestamp 1623621585
transform -1 0 38824 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1865
timestamp 1623621585
transform 1 0 37812 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input310
timestamp 1623621585
transform 1 0 37812 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_204_400
timestamp 1623621585
transform 1 0 37904 0 -1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_406
timestamp 1623621585
transform 1 0 38456 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_205_397
timestamp 1623621585
transform 1 0 37628 0 1 113696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_205_403
timestamp 1623621585
transform 1 0 38180 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_412
timestamp 1623621585
transform 1 0 1104 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output617
timestamp 1623621585
transform 1 0 1748 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output658
timestamp 1623621585
transform 1 0 2484 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_3
timestamp 1623621585
transform 1 0 1380 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_11
timestamp 1623621585
transform 1 0 2116 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_19
timestamp 1623621585
transform 1 0 2852 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _663_
timestamp 1623621585
transform 1 0 3956 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _664_
timestamp 1623621585
transform 1 0 4600 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output659
timestamp 1623621585
transform 1 0 3220 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_27
timestamp 1623621585
transform 1 0 3588 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_34
timestamp 1623621585
transform 1 0 4232 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_41
timestamp 1623621585
transform 1 0 4876 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _666_
timestamp 1623621585
transform 1 0 5244 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _668_
timestamp 1623621585
transform 1 0 6808 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1873
timestamp 1623621585
transform 1 0 6348 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_206_48
timestamp 1623621585
transform 1 0 5520 0 -1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_206_56
timestamp 1623621585
transform 1 0 6256 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_206_58
timestamp 1623621585
transform 1 0 6440 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _697_
timestamp 1623621585
transform 1 0 7452 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _698_
timestamp 1623621585
transform 1 0 8096 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _700_
timestamp 1623621585
transform 1 0 8740 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_65
timestamp 1623621585
transform 1 0 7084 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_72
timestamp 1623621585
transform 1 0 7728 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_79
timestamp 1623621585
transform 1 0 8372 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1623621585
transform 1 0 9384 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1623621585
transform 1 0 10028 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1623621585
transform 1 0 10672 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_86
timestamp 1623621585
transform 1 0 9016 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_93
timestamp 1623621585
transform 1 0 9660 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_100
timestamp 1623621585
transform 1 0 10304 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1874
timestamp 1623621585
transform 1 0 11592 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1623621585
transform 1 0 12052 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_206_107
timestamp 1623621585
transform 1 0 10948 0 -1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_113
timestamp 1623621585
transform 1 0 11500 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_206_115
timestamp 1623621585
transform 1 0 11684 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_122
timestamp 1623621585
transform 1 0 12328 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1623621585
transform 1 0 12696 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1623621585
transform 1 0 13340 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1623621585
transform 1 0 13984 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_129
timestamp 1623621585
transform 1 0 12972 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_136
timestamp 1623621585
transform 1 0 13616 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_143
timestamp 1623621585
transform 1 0 14260 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1623621585
transform 1 0 14628 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1623621585
transform 1 0 15272 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1623621585
transform 1 0 15916 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_150
timestamp 1623621585
transform 1 0 14904 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_157
timestamp 1623621585
transform 1 0 15548 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_206_164
timestamp 1623621585
transform 1 0 16192 0 -1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1875
timestamp 1623621585
transform 1 0 16836 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1623621585
transform 1 0 17848 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_206_170
timestamp 1623621585
transform 1 0 16744 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_206_172
timestamp 1623621585
transform 1 0 16928 0 -1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_206_180
timestamp 1623621585
transform 1 0 17664 0 -1 114784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_206_185
timestamp 1623621585
transform 1 0 18124 0 -1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1623621585
transform 1 0 19228 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1623621585
transform 1 0 19964 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_200
timestamp 1623621585
transform 1 0 19504 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_206_204
timestamp 1623621585
transform 1 0 19872 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_208
timestamp 1623621585
transform 1 0 20240 0 -1 114784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1876
timestamp 1623621585
transform 1 0 22080 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_206_220
timestamp 1623621585
transform 1 0 21344 0 -1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_206_229
timestamp 1623621585
transform 1 0 22172 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _759_
timestamp 1623621585
transform 1 0 22632 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1623621585
transform 1 0 23276 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_206_233
timestamp 1623621585
transform 1 0 22540 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_206_237
timestamp 1623621585
transform 1 0 22908 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_206_244
timestamp 1623621585
transform 1 0 23552 0 -1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _761_
timestamp 1623621585
transform 1 0 24288 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1623621585
transform 1 0 24932 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1623621585
transform 1 0 25576 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_255
timestamp 1623621585
transform 1 0 24564 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_262
timestamp 1623621585
transform 1 0 25208 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_269
timestamp 1623621585
transform 1 0 25852 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _703_
timestamp 1623621585
transform 1 0 27784 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1877
timestamp 1623621585
transform 1 0 27324 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1623621585
transform 1 0 26220 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_206_276
timestamp 1623621585
transform 1 0 26496 0 -1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_206_284
timestamp 1623621585
transform 1 0 27232 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_206_286
timestamp 1623621585
transform 1 0 27416 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _705_
timestamp 1623621585
transform 1 0 28428 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _707_
timestamp 1623621585
transform 1 0 29072 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_293
timestamp 1623621585
transform 1 0 28060 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_300
timestamp 1623621585
transform 1 0 28704 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_206_307
timestamp 1623621585
transform 1 0 29348 0 -1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1623621585
transform 1 0 31280 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input447
timestamp 1623621585
transform 1 0 30636 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output680
timestamp 1623621585
transform 1 0 29900 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_317
timestamp 1623621585
transform 1 0 30268 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_324
timestamp 1623621585
transform 1 0 30912 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_331
timestamp 1623621585
transform 1 0 31556 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1878
timestamp 1623621585
transform 1 0 32568 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1623621585
transform 1 0 31924 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output665
timestamp 1623621585
transform 1 0 33120 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_338
timestamp 1623621585
transform 1 0 32200 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_343
timestamp 1623621585
transform 1 0 32660 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_206_347
timestamp 1623621585
transform 1 0 33028 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_206_352
timestamp 1623621585
transform 1 0 33488 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _601_
timestamp 1623621585
transform 1 0 34592 0 -1 114784
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  output655
timestamp 1623621585
transform 1 0 33856 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_360
timestamp 1623621585
transform 1 0 34224 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _602_
timestamp 1623621585
transform 1 0 36156 0 -1 114784
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_206_377
timestamp 1623621585
transform 1 0 35788 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_394
timestamp 1623621585
transform 1 0 37352 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_413
timestamp 1623621585
transform -1 0 38824 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1879
timestamp 1623621585
transform 1 0 37812 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_206_398
timestamp 1623621585
transform 1 0 37720 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_206_400
timestamp 1623621585
transform 1 0 37904 0 -1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_406
timestamp 1623621585
transform 1 0 38456 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_414
timestamp 1623621585
transform 1 0 1104 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output647
timestamp 1623621585
transform 1 0 2484 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output654
timestamp 1623621585
transform 1 0 1748 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_3
timestamp 1623621585
transform 1 0 1380 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_11
timestamp 1623621585
transform 1 0 2116 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_207_19
timestamp 1623621585
transform 1 0 2852 0 1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _635_
timestamp 1623621585
transform 1 0 4232 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _637_
timestamp 1623621585
transform 1 0 4876 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1880
timestamp 1623621585
transform 1 0 3772 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_207_27
timestamp 1623621585
transform 1 0 3588 0 1 114784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_207_30
timestamp 1623621585
transform 1 0 3864 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_37
timestamp 1623621585
transform 1 0 4508 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _638_
timestamp 1623621585
transform 1 0 5520 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _640_
timestamp 1623621585
transform 1 0 6164 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _641_
timestamp 1623621585
transform 1 0 6808 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_44
timestamp 1623621585
transform 1 0 5152 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_51
timestamp 1623621585
transform 1 0 5796 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_58
timestamp 1623621585
transform 1 0 6440 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _669_
timestamp 1623621585
transform 1 0 7452 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _670_
timestamp 1623621585
transform 1 0 8096 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_65
timestamp 1623621585
transform 1 0 7084 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_72
timestamp 1623621585
transform 1 0 7728 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_207_79
timestamp 1623621585
transform 1 0 8372 0 1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _671_
timestamp 1623621585
transform 1 0 9476 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _672_
timestamp 1623621585
transform 1 0 10120 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1881
timestamp 1623621585
transform 1 0 9016 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_207_85
timestamp 1623621585
transform 1 0 8924 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_87
timestamp 1623621585
transform 1 0 9108 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_94
timestamp 1623621585
transform 1 0 9752 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_101
timestamp 1623621585
transform 1 0 10396 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _673_
timestamp 1623621585
transform 1 0 10764 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _676_
timestamp 1623621585
transform 1 0 12604 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1623621585
transform 1 0 11408 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_108
timestamp 1623621585
transform 1 0 11040 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_207_115
timestamp 1623621585
transform 1 0 11684 0 1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_207_123
timestamp 1623621585
transform 1 0 12420 0 1 114784
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _677_
timestamp 1623621585
transform 1 0 13248 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1882
timestamp 1623621585
transform 1 0 14260 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_128
timestamp 1623621585
transform 1 0 12880 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_207_135
timestamp 1623621585
transform 1 0 13524 0 1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_207_144
timestamp 1623621585
transform 1 0 14352 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _679_
timestamp 1623621585
transform 1 0 14720 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _680_
timestamp 1623621585
transform 1 0 15364 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _681_
timestamp 1623621585
transform 1 0 16100 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_151
timestamp 1623621585
transform 1 0 14996 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_158
timestamp 1623621585
transform 1 0 15640 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_207_162
timestamp 1623621585
transform 1 0 16008 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_166
timestamp 1623621585
transform 1 0 16376 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _684_
timestamp 1623621585
transform 1 0 18124 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1623621585
transform 1 0 16744 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1623621585
transform 1 0 17388 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_173
timestamp 1623621585
transform 1 0 17020 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_180
timestamp 1623621585
transform 1 0 17664 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_207_184
timestamp 1623621585
transform 1 0 18032 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _686_
timestamp 1623621585
transform 1 0 19964 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1883
timestamp 1623621585
transform 1 0 19504 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1623621585
transform 1 0 18768 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_188
timestamp 1623621585
transform 1 0 18400 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_195
timestamp 1623621585
transform 1 0 19044 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_207_199
timestamp 1623621585
transform 1 0 19412 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_201
timestamp 1623621585
transform 1 0 19596 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_208
timestamp 1623621585
transform 1 0 20240 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _687_
timestamp 1623621585
transform 1 0 20608 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1623621585
transform 1 0 21252 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1623621585
transform 1 0 21896 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_215
timestamp 1623621585
transform 1 0 20884 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_222
timestamp 1623621585
transform 1 0 21528 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_207_229
timestamp 1623621585
transform 1 0 22172 0 1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _756_
timestamp 1623621585
transform 1 0 22724 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _757_
timestamp 1623621585
transform 1 0 23460 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _760_
timestamp 1623621585
transform 1 0 24104 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_238
timestamp 1623621585
transform 1 0 23000 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_207_242
timestamp 1623621585
transform 1 0 23368 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_246
timestamp 1623621585
transform 1 0 23736 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _762_
timestamp 1623621585
transform 1 0 25208 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1884
timestamp 1623621585
transform 1 0 24748 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_253
timestamp 1623621585
transform 1 0 24380 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_258
timestamp 1623621585
transform 1 0 24840 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_207_265
timestamp 1623621585
transform 1 0 25484 0 1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _689_
timestamp 1623621585
transform 1 0 27140 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _690_
timestamp 1623621585
transform 1 0 27876 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _701_
timestamp 1623621585
transform 1 0 26220 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_207_276
timestamp 1623621585
transform 1 0 26496 0 1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_282
timestamp 1623621585
transform 1 0 27048 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_286
timestamp 1623621585
transform 1 0 27416 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_207_290
timestamp 1623621585
transform 1 0 27784 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _704_
timestamp 1623621585
transform 1 0 28520 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _706_
timestamp 1623621585
transform 1 0 29164 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_294
timestamp 1623621585
transform 1 0 28152 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_301
timestamp 1623621585
transform 1 0 28796 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_207_308
timestamp 1623621585
transform 1 0 29440 0 1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1885
timestamp 1623621585
transform 1 0 29992 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1623621585
transform 1 0 31280 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output679
timestamp 1623621585
transform 1 0 30452 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_315
timestamp 1623621585
transform 1 0 30084 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_323
timestamp 1623621585
transform 1 0 30820 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_207_327
timestamp 1623621585
transform 1 0 31188 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_331
timestamp 1623621585
transform 1 0 31556 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1623621585
transform 1 0 31924 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output664
timestamp 1623621585
transform 1 0 33028 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_207_338
timestamp 1623621585
transform 1 0 32200 0 1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_207_346
timestamp 1623621585
transform 1 0 32936 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_351
timestamp 1623621585
transform 1 0 33396 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1886
timestamp 1623621585
transform 1 0 35236 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output639
timestamp 1623621585
transform 1 0 34500 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output648
timestamp 1623621585
transform 1 0 33764 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_359
timestamp 1623621585
transform 1 0 34132 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_367
timestamp 1623621585
transform 1 0 34868 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_372
timestamp 1623621585
transform 1 0 35328 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _603_
timestamp 1623621585
transform 1 0 35696 0 1 114784
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_207_389
timestamp 1623621585
transform 1 0 36892 0 1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_415
timestamp 1623621585
transform -1 0 38824 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input311
timestamp 1623621585
transform 1 0 37812 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_207_397
timestamp 1623621585
transform 1 0 37628 0 1 114784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_207_403
timestamp 1623621585
transform 1 0 38180 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_416
timestamp 1623621585
transform 1 0 1104 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output642
timestamp 1623621585
transform 1 0 1748 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_3
timestamp 1623621585
transform 1 0 1380 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_208_11
timestamp 1623621585
transform 1 0 2116 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_208_19
timestamp 1623621585
transform 1 0 2852 0 -1 115872
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _634_
timestamp 1623621585
transform 1 0 3772 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output584
timestamp 1623621585
transform 1 0 3036 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output604
timestamp 1623621585
transform 1 0 4416 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_25
timestamp 1623621585
transform 1 0 3404 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_32
timestamp 1623621585
transform 1 0 4048 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_40
timestamp 1623621585
transform 1 0 4784 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1887
timestamp 1623621585
transform 1 0 6348 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output605
timestamp 1623621585
transform 1 0 5152 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_208_48
timestamp 1623621585
transform 1 0 5520 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_208_56
timestamp 1623621585
transform 1 0 6256 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_208_58
timestamp 1623621585
transform 1 0 6440 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _624_
timestamp 1623621585
transform 1 0 7268 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _625_
timestamp 1623621585
transform 1 0 8648 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output609
timestamp 1623621585
transform 1 0 7912 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_208_66
timestamp 1623621585
transform 1 0 7176 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_208_70
timestamp 1623621585
transform 1 0 7544 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_78
timestamp 1623621585
transform 1 0 8280 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _642_
timestamp 1623621585
transform 1 0 9292 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _643_
timestamp 1623621585
transform 1 0 9936 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _644_
timestamp 1623621585
transform 1 0 10580 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_208_85
timestamp 1623621585
transform 1 0 8924 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_92
timestamp 1623621585
transform 1 0 9568 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_99
timestamp 1623621585
transform 1 0 10212 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _674_
timestamp 1623621585
transform 1 0 12052 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1888
timestamp 1623621585
transform 1 0 11592 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_208_106
timestamp 1623621585
transform 1 0 10856 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_208_115
timestamp 1623621585
transform 1 0 11684 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_122
timestamp 1623621585
transform 1 0 12328 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _649_
timestamp 1623621585
transform 1 0 13708 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _650_
timestamp 1623621585
transform 1 0 14444 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _675_
timestamp 1623621585
transform 1 0 12696 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_208_129
timestamp 1623621585
transform 1 0 12972 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_208_140
timestamp 1623621585
transform 1 0 13984 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_208_144
timestamp 1623621585
transform 1 0 14352 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _652_
timestamp 1623621585
transform 1 0 15824 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _678_
timestamp 1623621585
transform 1 0 15088 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_208_148
timestamp 1623621585
transform 1 0 14720 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_155
timestamp 1623621585
transform 1 0 15364 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_208_159
timestamp 1623621585
transform 1 0 15732 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_208_163
timestamp 1623621585
transform 1 0 16100 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _682_
timestamp 1623621585
transform 1 0 17296 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _683_
timestamp 1623621585
transform 1 0 17940 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1889
timestamp 1623621585
transform 1 0 16836 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_208_172
timestamp 1623621585
transform 1 0 16928 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_179
timestamp 1623621585
transform 1 0 17572 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_186
timestamp 1623621585
transform 1 0 18216 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _656_
timestamp 1623621585
transform 1 0 18584 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _658_
timestamp 1623621585
transform 1 0 19964 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _685_
timestamp 1623621585
transform 1 0 19228 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_208_193
timestamp 1623621585
transform 1 0 18860 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_200
timestamp 1623621585
transform 1 0 19504 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_208_204
timestamp 1623621585
transform 1 0 19872 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_208_208
timestamp 1623621585
transform 1 0 20240 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _659_
timestamp 1623621585
transform 1 0 20700 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _688_
timestamp 1623621585
transform 1 0 21344 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1890
timestamp 1623621585
transform 1 0 22080 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_208_212
timestamp 1623621585
transform 1 0 20608 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_208_216
timestamp 1623621585
transform 1 0 20976 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_223
timestamp 1623621585
transform 1 0 21620 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_208_227
timestamp 1623621585
transform 1 0 21988 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_208_229
timestamp 1623621585
transform 1 0 22172 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _629_
timestamp 1623621585
transform 1 0 23552 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _755_
timestamp 1623621585
transform 1 0 22540 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_208_236
timestamp 1623621585
transform 1 0 22816 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_208_247
timestamp 1623621585
transform 1 0 23828 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _630_
timestamp 1623621585
transform 1 0 24288 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _702_
timestamp 1623621585
transform 1 0 25668 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _758_
timestamp 1623621585
transform 1 0 24932 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_208_251
timestamp 1623621585
transform 1 0 24196 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_208_255
timestamp 1623621585
transform 1 0 24564 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_262
timestamp 1623621585
transform 1 0 25208 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_208_266
timestamp 1623621585
transform 1 0 25576 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_208_270
timestamp 1623621585
transform 1 0 25944 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _633_
timestamp 1623621585
transform 1 0 26312 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _661_
timestamp 1623621585
transform 1 0 27784 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1891
timestamp 1623621585
transform 1 0 27324 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_208_277
timestamp 1623621585
transform 1 0 26588 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_208_286
timestamp 1623621585
transform 1 0 27416 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output676
timestamp 1623621585
transform 1 0 28980 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output677
timestamp 1623621585
transform 1 0 29716 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_208_293
timestamp 1623621585
transform 1 0 28060 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_208_301
timestamp 1623621585
transform 1 0 28796 0 -1 115872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_208_307
timestamp 1623621585
transform 1 0 29348 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _708_
timestamp 1623621585
transform 1 0 31188 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output678
timestamp 1623621585
transform 1 0 30452 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_315
timestamp 1623621585
transform 1 0 30084 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_323
timestamp 1623621585
transform 1 0 30820 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_330
timestamp 1623621585
transform 1 0 31464 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1892
timestamp 1623621585
transform 1 0 32568 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output640
timestamp 1623621585
transform 1 0 33396 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output669
timestamp 1623621585
transform 1 0 31832 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_338
timestamp 1623621585
transform 1 0 32200 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_208_343
timestamp 1623621585
transform 1 0 32660 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output634
timestamp 1623621585
transform 1 0 35604 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output636
timestamp 1623621585
transform 1 0 34868 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output638
timestamp 1623621585
transform 1 0 34132 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_355
timestamp 1623621585
transform 1 0 33764 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_363
timestamp 1623621585
transform 1 0 34500 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_371
timestamp 1623621585
transform 1 0 35236 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output625
timestamp 1623621585
transform 1 0 37076 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output632
timestamp 1623621585
transform 1 0 36340 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_379
timestamp 1623621585
transform 1 0 35972 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_387
timestamp 1623621585
transform 1 0 36708 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_395
timestamp 1623621585
transform 1 0 37444 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_417
timestamp 1623621585
transform -1 0 38824 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1893
timestamp 1623621585
transform 1 0 37812 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_208_400
timestamp 1623621585
transform 1 0 37904 0 -1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_406
timestamp 1623621585
transform 1 0 38456 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_418
timestamp 1623621585
transform 1 0 1104 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output645
timestamp 1623621585
transform 1 0 1748 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_3
timestamp 1623621585
transform 1 0 1380 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_11
timestamp 1623621585
transform 1 0 2116 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_209_19
timestamp 1623621585
transform 1 0 2852 0 1 115872
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1894
timestamp 1623621585
transform 1 0 3772 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output573
timestamp 1623621585
transform 1 0 3036 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output595
timestamp 1623621585
transform 1 0 4232 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_25
timestamp 1623621585
transform 1 0 3404 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_30
timestamp 1623621585
transform 1 0 3864 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_38
timestamp 1623621585
transform 1 0 4600 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _636_
timestamp 1623621585
transform 1 0 4968 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output568
timestamp 1623621585
transform 1 0 5612 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output606
timestamp 1623621585
transform 1 0 6348 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_45
timestamp 1623621585
transform 1 0 5244 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_53
timestamp 1623621585
transform 1 0 5980 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_61
timestamp 1623621585
transform 1 0 6716 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output607
timestamp 1623621585
transform 1 0 7084 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output608
timestamp 1623621585
transform 1 0 7820 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_69
timestamp 1623621585
transform 1 0 7452 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_77
timestamp 1623621585
transform 1 0 8188 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1895
timestamp 1623621585
transform 1 0 9016 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output576
timestamp 1623621585
transform 1 0 10672 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output610
timestamp 1623621585
transform 1 0 9476 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_209_85
timestamp 1623621585
transform 1 0 8924 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_209_87
timestamp 1623621585
transform 1 0 9108 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_95
timestamp 1623621585
transform 1 0 9844 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_209_103
timestamp 1623621585
transform 1 0 10580 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _645_
timestamp 1623621585
transform 1 0 11408 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _646_
timestamp 1623621585
transform 1 0 12052 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_209_108
timestamp 1623621585
transform 1 0 11040 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_115
timestamp 1623621585
transform 1 0 11684 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_122
timestamp 1623621585
transform 1 0 12328 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _647_
timestamp 1623621585
transform 1 0 12696 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _648_
timestamp 1623621585
transform 1 0 13340 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1896
timestamp 1623621585
transform 1 0 14260 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_209_129
timestamp 1623621585
transform 1 0 12972 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_209_136
timestamp 1623621585
transform 1 0 13616 0 1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_142
timestamp 1623621585
transform 1 0 14168 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_209_144
timestamp 1623621585
transform 1 0 14352 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _651_
timestamp 1623621585
transform 1 0 15548 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output582
timestamp 1623621585
transform 1 0 14812 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output585
timestamp 1623621585
transform 1 0 16284 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_209_148
timestamp 1623621585
transform 1 0 14720 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_209_153
timestamp 1623621585
transform 1 0 15180 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_160
timestamp 1623621585
transform 1 0 15824 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_209_164
timestamp 1623621585
transform 1 0 16192 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _653_
timestamp 1623621585
transform 1 0 17020 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _654_
timestamp 1623621585
transform 1 0 17664 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _655_
timestamp 1623621585
transform 1 0 18308 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_209_169
timestamp 1623621585
transform 1 0 16652 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_176
timestamp 1623621585
transform 1 0 17296 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_183
timestamp 1623621585
transform 1 0 17940 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _657_
timestamp 1623621585
transform 1 0 19964 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1897
timestamp 1623621585
transform 1 0 19504 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_209_190
timestamp 1623621585
transform 1 0 18584 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_209_198
timestamp 1623621585
transform 1 0 19320 0 1 115872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_209_201
timestamp 1623621585
transform 1 0 19596 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_208
timestamp 1623621585
transform 1 0 20240 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _626_
timestamp 1623621585
transform 1 0 21804 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output592
timestamp 1623621585
transform 1 0 21068 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_209_216
timestamp 1623621585
transform 1 0 20976 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_209_221
timestamp 1623621585
transform 1 0 21436 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_228
timestamp 1623621585
transform 1 0 22080 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _627_
timestamp 1623621585
transform 1 0 22448 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _628_
timestamp 1623621585
transform 1 0 23092 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output597
timestamp 1623621585
transform 1 0 23828 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_235
timestamp 1623621585
transform 1 0 22724 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_242
timestamp 1623621585
transform 1 0 23368 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_209_246
timestamp 1623621585
transform 1 0 23736 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _631_
timestamp 1623621585
transform 1 0 25208 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _632_
timestamp 1623621585
transform 1 0 25852 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1898
timestamp 1623621585
transform 1 0 24748 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_209_251
timestamp 1623621585
transform 1 0 24196 0 1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_209_258
timestamp 1623621585
transform 1 0 24840 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_265
timestamp 1623621585
transform 1 0 25484 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _660_
timestamp 1623621585
transform 1 0 27416 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output601
timestamp 1623621585
transform 1 0 26680 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_209_272
timestamp 1623621585
transform 1 0 26128 0 1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_209_282
timestamp 1623621585
transform 1 0 27048 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_209_289
timestamp 1623621585
transform 1 0 27692 0 1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output673
timestamp 1623621585
transform 1 0 28244 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output675
timestamp 1623621585
transform 1 0 28980 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_299
timestamp 1623621585
transform 1 0 28612 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_209_307
timestamp 1623621585
transform 1 0 29348 0 1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _611_
timestamp 1623621585
transform 1 0 31004 0 1 115872
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1899
timestamp 1623621585
transform 1 0 29992 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_209_313
timestamp 1623621585
transform 1 0 29900 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_209_315
timestamp 1623621585
transform 1 0 30084 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_209_323
timestamp 1623621585
transform 1 0 30820 0 1 115872
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _610_
timestamp 1623621585
transform 1 0 32200 0 1 115872
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _612_
timestamp 1623621585
transform 1 0 33396 0 1 115872
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_209_334
timestamp 1623621585
transform 1 0 31832 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_347
timestamp 1623621585
transform 1 0 33028 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1900
timestamp 1623621585
transform 1 0 35236 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1623621585
transform 1 0 34592 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_209_360
timestamp 1623621585
transform 1 0 34224 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_367
timestamp 1623621585
transform 1 0 34868 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_372
timestamp 1623621585
transform 1 0 35328 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output626
timestamp 1623621585
transform 1 0 36800 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output633
timestamp 1623621585
transform 1 0 35696 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_380
timestamp 1623621585
transform 1 0 36064 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_209_392
timestamp 1623621585
transform 1 0 37168 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_419
timestamp 1623621585
transform -1 0 38824 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input60
timestamp 1623621585
transform 1 0 37536 0 1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_209_402
timestamp 1623621585
transform 1 0 38088 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_209_406
timestamp 1623621585
transform 1 0 38456 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_420
timestamp 1623621585
transform 1 0 1104 0 -1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output534
timestamp 1623621585
transform 1 0 1748 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output535
timestamp 1623621585
transform 1 0 2484 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_3
timestamp 1623621585
transform 1 0 1380 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_11
timestamp 1623621585
transform 1 0 2116 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_19
timestamp 1623621585
transform 1 0 2852 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output529
timestamp 1623621585
transform 1 0 3220 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output566
timestamp 1623621585
transform 1 0 4232 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_210_27
timestamp 1623621585
transform 1 0 3588 0 -1 116960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_33
timestamp 1623621585
transform 1 0 4140 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_210_38
timestamp 1623621585
transform 1 0 4600 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _639_
timestamp 1623621585
transform 1 0 5704 0 -1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1901
timestamp 1623621585
transform 1 0 6348 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output567
timestamp 1623621585
transform 1 0 4968 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output569
timestamp 1623621585
transform 1 0 6808 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_46
timestamp 1623621585
transform 1 0 5336 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_53
timestamp 1623621585
transform 1 0 5980 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_58
timestamp 1623621585
transform 1 0 6440 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output570
timestamp 1623621585
transform 1 0 7544 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output571
timestamp 1623621585
transform 1 0 8280 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_66
timestamp 1623621585
transform 1 0 7176 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_74
timestamp 1623621585
transform 1 0 7912 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_82
timestamp 1623621585
transform 1 0 8648 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output572
timestamp 1623621585
transform 1 0 9016 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output574
timestamp 1623621585
transform 1 0 9752 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output575
timestamp 1623621585
transform 1 0 10488 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_90
timestamp 1623621585
transform 1 0 9384 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_98
timestamp 1623621585
transform 1 0 10120 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1902
timestamp 1623621585
transform 1 0 11592 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output577
timestamp 1623621585
transform 1 0 12052 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_210_106
timestamp 1623621585
transform 1 0 10856 0 -1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_210_115
timestamp 1623621585
transform 1 0 11684 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_123
timestamp 1623621585
transform 1 0 12420 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output578
timestamp 1623621585
transform 1 0 12788 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output579
timestamp 1623621585
transform 1 0 13524 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output580
timestamp 1623621585
transform 1 0 14260 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_131
timestamp 1623621585
transform 1 0 13156 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_139
timestamp 1623621585
transform 1 0 13892 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output581
timestamp 1623621585
transform 1 0 14996 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output583
timestamp 1623621585
transform 1 0 15732 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_147
timestamp 1623621585
transform 1 0 14628 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_155
timestamp 1623621585
transform 1 0 15364 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_210_163
timestamp 1623621585
transform 1 0 16100 0 -1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1903
timestamp 1623621585
transform 1 0 16836 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output586
timestamp 1623621585
transform 1 0 17296 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output587
timestamp 1623621585
transform 1 0 18032 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_172
timestamp 1623621585
transform 1 0 16928 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_180
timestamp 1623621585
transform 1 0 17664 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output588
timestamp 1623621585
transform 1 0 18768 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output589
timestamp 1623621585
transform 1 0 19504 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output590
timestamp 1623621585
transform 1 0 20240 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_188
timestamp 1623621585
transform 1 0 18400 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_196
timestamp 1623621585
transform 1 0 19136 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_204
timestamp 1623621585
transform 1 0 19872 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1904
timestamp 1623621585
transform 1 0 22080 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output591
timestamp 1623621585
transform 1 0 20976 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_212
timestamp 1623621585
transform 1 0 20608 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_210_220
timestamp 1623621585
transform 1 0 21344 0 -1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_210_229
timestamp 1623621585
transform 1 0 22172 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output593
timestamp 1623621585
transform 1 0 22540 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output594
timestamp 1623621585
transform 1 0 23276 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output596
timestamp 1623621585
transform 1 0 24012 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_237
timestamp 1623621585
transform 1 0 22908 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_245
timestamp 1623621585
transform 1 0 23644 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output598
timestamp 1623621585
transform 1 0 24748 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output599
timestamp 1623621585
transform 1 0 25484 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_253
timestamp 1623621585
transform 1 0 24380 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_261
timestamp 1623621585
transform 1 0 25116 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_269
timestamp 1623621585
transform 1 0 25852 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1905
timestamp 1623621585
transform 1 0 27324 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output565
timestamp 1623621585
transform 1 0 27784 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output600
timestamp 1623621585
transform 1 0 26220 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_210_277
timestamp 1623621585
transform 1 0 26588 0 -1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_210_286
timestamp 1623621585
transform 1 0 27416 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output603
timestamp 1623621585
transform 1 0 28520 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output674
timestamp 1623621585
transform 1 0 29256 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_294
timestamp 1623621585
transform 1 0 28152 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_302
timestamp 1623621585
transform 1 0 28888 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_210_310
timestamp 1623621585
transform 1 0 29624 0 -1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output649
timestamp 1623621585
transform 1 0 31096 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output656
timestamp 1623621585
transform 1 0 30360 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_322
timestamp 1623621585
transform 1 0 30728 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_330
timestamp 1623621585
transform 1 0 31464 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1906
timestamp 1623621585
transform 1 0 32568 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output637
timestamp 1623621585
transform 1 0 33396 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output643
timestamp 1623621585
transform 1 0 31832 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_338
timestamp 1623621585
transform 1 0 32200 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_210_343
timestamp 1623621585
transform 1 0 32660 0 -1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output629
timestamp 1623621585
transform 1 0 35604 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output631
timestamp 1623621585
transform 1 0 34868 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output635
timestamp 1623621585
transform 1 0 34132 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_355
timestamp 1623621585
transform 1 0 33764 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_363
timestamp 1623621585
transform 1 0 34500 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_371
timestamp 1623621585
transform 1 0 35236 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1623621585
transform 1 0 36340 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output623
timestamp 1623621585
transform 1 0 37076 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_379
timestamp 1623621585
transform 1 0 35972 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_387
timestamp 1623621585
transform 1 0 36708 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_395
timestamp 1623621585
transform 1 0 37444 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_421
timestamp 1623621585
transform -1 0 38824 0 -1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1907
timestamp 1623621585
transform 1 0 37812 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_210_400
timestamp 1623621585
transform 1 0 37904 0 -1 116960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_406
timestamp 1623621585
transform 1 0 38456 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_422
timestamp 1623621585
transform 1 0 1104 0 1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output527
timestamp 1623621585
transform 1 0 1748 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output528
timestamp 1623621585
transform 1 0 2484 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_3
timestamp 1623621585
transform 1 0 1380 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_11
timestamp 1623621585
transform 1 0 2116 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_211_19
timestamp 1623621585
transform 1 0 2852 0 1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1908
timestamp 1623621585
transform 1 0 3772 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output530
timestamp 1623621585
transform 1 0 4232 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_211_27
timestamp 1623621585
transform 1 0 3588 0 1 116960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_211_30
timestamp 1623621585
transform 1 0 3864 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_38
timestamp 1623621585
transform 1 0 4600 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1909
timestamp 1623621585
transform 1 0 6440 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output531
timestamp 1623621585
transform 1 0 4968 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output532
timestamp 1623621585
transform 1 0 5704 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_46
timestamp 1623621585
transform 1 0 5336 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_54
timestamp 1623621585
transform 1 0 6072 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_59
timestamp 1623621585
transform 1 0 6532 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output533
timestamp 1623621585
transform 1 0 6900 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output546
timestamp 1623621585
transform 1 0 7636 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output557
timestamp 1623621585
transform 1 0 8372 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_67
timestamp 1623621585
transform 1 0 7268 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_75
timestamp 1623621585
transform 1 0 8004 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_83
timestamp 1623621585
transform 1 0 8740 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1910
timestamp 1623621585
transform 1 0 9108 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output536
timestamp 1623621585
transform 1 0 9568 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output537
timestamp 1623621585
transform 1 0 10304 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_88
timestamp 1623621585
transform 1 0 9200 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_96
timestamp 1623621585
transform 1 0 9936 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_104
timestamp 1623621585
transform 1 0 10672 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1911
timestamp 1623621585
transform 1 0 11776 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output538
timestamp 1623621585
transform 1 0 11040 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output539
timestamp 1623621585
transform 1 0 12236 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_112
timestamp 1623621585
transform 1 0 11408 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_117
timestamp 1623621585
transform 1 0 11868 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_125
timestamp 1623621585
transform 1 0 12604 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1912
timestamp 1623621585
transform 1 0 14444 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output540
timestamp 1623621585
transform 1 0 12972 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output541
timestamp 1623621585
transform 1 0 13708 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_133
timestamp 1623621585
transform 1 0 13340 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_141
timestamp 1623621585
transform 1 0 14076 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output542
timestamp 1623621585
transform 1 0 14904 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output543
timestamp 1623621585
transform 1 0 15640 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output544
timestamp 1623621585
transform 1 0 16376 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_146
timestamp 1623621585
transform 1 0 14536 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_154
timestamp 1623621585
transform 1 0 15272 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_162
timestamp 1623621585
transform 1 0 16008 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1913
timestamp 1623621585
transform 1 0 17112 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output545
timestamp 1623621585
transform 1 0 17572 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output547
timestamp 1623621585
transform 1 0 18308 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_170
timestamp 1623621585
transform 1 0 16744 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_175
timestamp 1623621585
transform 1 0 17204 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_183
timestamp 1623621585
transform 1 0 17940 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1914
timestamp 1623621585
transform 1 0 19780 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output548
timestamp 1623621585
transform 1 0 19044 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output549
timestamp 1623621585
transform 1 0 20240 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_191
timestamp 1623621585
transform 1 0 18676 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_199
timestamp 1623621585
transform 1 0 19412 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_204
timestamp 1623621585
transform 1 0 19872 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output550
timestamp 1623621585
transform 1 0 20976 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output551
timestamp 1623621585
transform 1 0 21712 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_212
timestamp 1623621585
transform 1 0 20608 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_220
timestamp 1623621585
transform 1 0 21344 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_228
timestamp 1623621585
transform 1 0 22080 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1915
timestamp 1623621585
transform 1 0 22448 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output552
timestamp 1623621585
transform 1 0 22908 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output553
timestamp 1623621585
transform 1 0 23644 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_233
timestamp 1623621585
transform 1 0 22540 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_241
timestamp 1623621585
transform 1 0 23276 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_249
timestamp 1623621585
transform 1 0 24012 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1916
timestamp 1623621585
transform 1 0 25116 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output554
timestamp 1623621585
transform 1 0 24380 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output555
timestamp 1623621585
transform 1 0 25576 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_257
timestamp 1623621585
transform 1 0 24748 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_262
timestamp 1623621585
transform 1 0 25208 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_270
timestamp 1623621585
transform 1 0 25944 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1917
timestamp 1623621585
transform 1 0 27784 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output556
timestamp 1623621585
transform 1 0 26312 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output558
timestamp 1623621585
transform 1 0 27048 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_278
timestamp 1623621585
transform 1 0 26680 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_286
timestamp 1623621585
transform 1 0 27416 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_291
timestamp 1623621585
transform 1 0 27876 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output559
timestamp 1623621585
transform 1 0 28244 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output560
timestamp 1623621585
transform 1 0 28980 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output561
timestamp 1623621585
transform 1 0 29716 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_299
timestamp 1623621585
transform 1 0 28612 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_307
timestamp 1623621585
transform 1 0 29348 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1918
timestamp 1623621585
transform 1 0 30452 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output562
timestamp 1623621585
transform 1 0 30912 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output563
timestamp 1623621585
transform 1 0 31648 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_315
timestamp 1623621585
transform 1 0 30084 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_320
timestamp 1623621585
transform 1 0 30544 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_328
timestamp 1623621585
transform 1 0 31280 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1919
timestamp 1623621585
transform 1 0 33120 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output564
timestamp 1623621585
transform 1 0 32384 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output602
timestamp 1623621585
transform 1 0 33580 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_336
timestamp 1623621585
transform 1 0 32016 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_344
timestamp 1623621585
transform 1 0 32752 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_349
timestamp 1623621585
transform 1 0 33212 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output615
timestamp 1623621585
transform 1 0 34776 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_211_357
timestamp 1623621585
transform 1 0 33948 0 1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_211_365
timestamp 1623621585
transform 1 0 34684 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_211_370
timestamp 1623621585
transform 1 0 35144 0 1 116960
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1920
timestamp 1623621585
transform 1 0 35788 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1623621585
transform 1 0 36248 0 1 116960
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input59
timestamp 1623621585
transform 1 0 37168 0 1 116960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_211_376
timestamp 1623621585
transform 1 0 35696 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_211_378
timestamp 1623621585
transform 1 0 35880 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_388
timestamp 1623621585
transform 1 0 36800 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_423
timestamp 1623621585
transform -1 0 38824 0 1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1921
timestamp 1623621585
transform 1 0 38456 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_211_398
timestamp 1623621585
transform 1 0 37720 0 1 116960
box -38 -48 774 592
<< labels >>
rlabel metal2 s 110 119200 166 120800 6 dsi[0]
port 0 nsew signal tristate
rlabel metal2 s 294 119200 350 120800 6 dsi[1]
port 1 nsew signal tristate
rlabel metal2 s 570 119200 626 120800 6 dsi[2]
port 2 nsew signal tristate
rlabel metal2 s 754 119200 810 120800 6 dsi[3]
port 3 nsew signal tristate
rlabel metal2 s 1030 119200 1086 120800 6 dsi[4]
port 4 nsew signal tristate
rlabel metal2 s 1214 119200 1270 120800 6 dsi[5]
port 5 nsew signal tristate
rlabel metal2 s 1490 119200 1546 120800 6 dsi[6]
port 6 nsew signal tristate
rlabel metal2 s 1674 119200 1730 120800 6 dsi[7]
port 7 nsew signal tristate
rlabel metal2 s 1950 119200 2006 120800 6 io_in[0]
port 8 nsew signal input
rlabel metal2 s 8850 119200 8906 120800 6 io_in[10]
port 9 nsew signal input
rlabel metal2 s 9586 119200 9642 120800 6 io_in[11]
port 10 nsew signal input
rlabel metal2 s 10230 119200 10286 120800 6 io_in[12]
port 11 nsew signal input
rlabel metal2 s 10966 119200 11022 120800 6 io_in[13]
port 12 nsew signal input
rlabel metal2 s 11610 119200 11666 120800 6 io_in[14]
port 13 nsew signal input
rlabel metal2 s 12346 119200 12402 120800 6 io_in[15]
port 14 nsew signal input
rlabel metal2 s 12990 119200 13046 120800 6 io_in[16]
port 15 nsew signal input
rlabel metal2 s 13726 119200 13782 120800 6 io_in[17]
port 16 nsew signal input
rlabel metal2 s 14370 119200 14426 120800 6 io_in[18]
port 17 nsew signal input
rlabel metal2 s 15106 119200 15162 120800 6 io_in[19]
port 18 nsew signal input
rlabel metal2 s 2594 119200 2650 120800 6 io_in[1]
port 19 nsew signal input
rlabel metal2 s 15750 119200 15806 120800 6 io_in[20]
port 20 nsew signal input
rlabel metal2 s 16486 119200 16542 120800 6 io_in[21]
port 21 nsew signal input
rlabel metal2 s 17222 119200 17278 120800 6 io_in[22]
port 22 nsew signal input
rlabel metal2 s 17866 119200 17922 120800 6 io_in[23]
port 23 nsew signal input
rlabel metal2 s 18602 119200 18658 120800 6 io_in[24]
port 24 nsew signal input
rlabel metal2 s 19246 119200 19302 120800 6 io_in[25]
port 25 nsew signal input
rlabel metal2 s 19982 119200 20038 120800 6 io_in[26]
port 26 nsew signal input
rlabel metal2 s 20626 119200 20682 120800 6 io_in[27]
port 27 nsew signal input
rlabel metal2 s 21362 119200 21418 120800 6 io_in[28]
port 28 nsew signal input
rlabel metal2 s 22006 119200 22062 120800 6 io_in[29]
port 29 nsew signal input
rlabel metal2 s 3330 119200 3386 120800 6 io_in[2]
port 30 nsew signal input
rlabel metal2 s 22742 119200 22798 120800 6 io_in[30]
port 31 nsew signal input
rlabel metal2 s 23386 119200 23442 120800 6 io_in[31]
port 32 nsew signal input
rlabel metal2 s 24122 119200 24178 120800 6 io_in[32]
port 33 nsew signal input
rlabel metal2 s 24858 119200 24914 120800 6 io_in[33]
port 34 nsew signal input
rlabel metal2 s 25502 119200 25558 120800 6 io_in[34]
port 35 nsew signal input
rlabel metal2 s 26238 119200 26294 120800 6 io_in[35]
port 36 nsew signal input
rlabel metal2 s 26882 119200 26938 120800 6 io_in[36]
port 37 nsew signal input
rlabel metal2 s 27618 119200 27674 120800 6 io_in[37]
port 38 nsew signal input
rlabel metal2 s 3974 119200 4030 120800 6 io_in[3]
port 39 nsew signal input
rlabel metal2 s 4710 119200 4766 120800 6 io_in[4]
port 40 nsew signal input
rlabel metal2 s 5354 119200 5410 120800 6 io_in[5]
port 41 nsew signal input
rlabel metal2 s 6090 119200 6146 120800 6 io_in[6]
port 42 nsew signal input
rlabel metal2 s 6734 119200 6790 120800 6 io_in[7]
port 43 nsew signal input
rlabel metal2 s 7470 119200 7526 120800 6 io_in[8]
port 44 nsew signal input
rlabel metal2 s 8206 119200 8262 120800 6 io_in[9]
port 45 nsew signal input
rlabel metal2 s 2134 119200 2190 120800 6 io_oeb[0]
port 46 nsew signal tristate
rlabel metal2 s 9126 119200 9182 120800 6 io_oeb[10]
port 47 nsew signal tristate
rlabel metal2 s 9770 119200 9826 120800 6 io_oeb[11]
port 48 nsew signal tristate
rlabel metal2 s 10506 119200 10562 120800 6 io_oeb[12]
port 49 nsew signal tristate
rlabel metal2 s 11150 119200 11206 120800 6 io_oeb[13]
port 50 nsew signal tristate
rlabel metal2 s 11886 119200 11942 120800 6 io_oeb[14]
port 51 nsew signal tristate
rlabel metal2 s 12530 119200 12586 120800 6 io_oeb[15]
port 52 nsew signal tristate
rlabel metal2 s 13266 119200 13322 120800 6 io_oeb[16]
port 53 nsew signal tristate
rlabel metal2 s 13910 119200 13966 120800 6 io_oeb[17]
port 54 nsew signal tristate
rlabel metal2 s 14646 119200 14702 120800 6 io_oeb[18]
port 55 nsew signal tristate
rlabel metal2 s 15290 119200 15346 120800 6 io_oeb[19]
port 56 nsew signal tristate
rlabel metal2 s 2870 119200 2926 120800 6 io_oeb[1]
port 57 nsew signal tristate
rlabel metal2 s 16026 119200 16082 120800 6 io_oeb[20]
port 58 nsew signal tristate
rlabel metal2 s 16762 119200 16818 120800 6 io_oeb[21]
port 59 nsew signal tristate
rlabel metal2 s 17406 119200 17462 120800 6 io_oeb[22]
port 60 nsew signal tristate
rlabel metal2 s 18142 119200 18198 120800 6 io_oeb[23]
port 61 nsew signal tristate
rlabel metal2 s 18786 119200 18842 120800 6 io_oeb[24]
port 62 nsew signal tristate
rlabel metal2 s 19522 119200 19578 120800 6 io_oeb[25]
port 63 nsew signal tristate
rlabel metal2 s 20166 119200 20222 120800 6 io_oeb[26]
port 64 nsew signal tristate
rlabel metal2 s 20902 119200 20958 120800 6 io_oeb[27]
port 65 nsew signal tristate
rlabel metal2 s 21546 119200 21602 120800 6 io_oeb[28]
port 66 nsew signal tristate
rlabel metal2 s 22282 119200 22338 120800 6 io_oeb[29]
port 67 nsew signal tristate
rlabel metal2 s 3514 119200 3570 120800 6 io_oeb[2]
port 68 nsew signal tristate
rlabel metal2 s 22926 119200 22982 120800 6 io_oeb[30]
port 69 nsew signal tristate
rlabel metal2 s 23662 119200 23718 120800 6 io_oeb[31]
port 70 nsew signal tristate
rlabel metal2 s 24398 119200 24454 120800 6 io_oeb[32]
port 71 nsew signal tristate
rlabel metal2 s 25042 119200 25098 120800 6 io_oeb[33]
port 72 nsew signal tristate
rlabel metal2 s 25778 119200 25834 120800 6 io_oeb[34]
port 73 nsew signal tristate
rlabel metal2 s 26422 119200 26478 120800 6 io_oeb[35]
port 74 nsew signal tristate
rlabel metal2 s 27158 119200 27214 120800 6 io_oeb[36]
port 75 nsew signal tristate
rlabel metal2 s 27802 119200 27858 120800 6 io_oeb[37]
port 76 nsew signal tristate
rlabel metal2 s 4250 119200 4306 120800 6 io_oeb[3]
port 77 nsew signal tristate
rlabel metal2 s 4894 119200 4950 120800 6 io_oeb[4]
port 78 nsew signal tristate
rlabel metal2 s 5630 119200 5686 120800 6 io_oeb[5]
port 79 nsew signal tristate
rlabel metal2 s 6274 119200 6330 120800 6 io_oeb[6]
port 80 nsew signal tristate
rlabel metal2 s 7010 119200 7066 120800 6 io_oeb[7]
port 81 nsew signal tristate
rlabel metal2 s 7654 119200 7710 120800 6 io_oeb[8]
port 82 nsew signal tristate
rlabel metal2 s 8390 119200 8446 120800 6 io_oeb[9]
port 83 nsew signal tristate
rlabel metal2 s 2410 119200 2466 120800 6 io_out[0]
port 84 nsew signal tristate
rlabel metal2 s 9310 119200 9366 120800 6 io_out[10]
port 85 nsew signal tristate
rlabel metal2 s 10046 119200 10102 120800 6 io_out[11]
port 86 nsew signal tristate
rlabel metal2 s 10690 119200 10746 120800 6 io_out[12]
port 87 nsew signal tristate
rlabel metal2 s 11426 119200 11482 120800 6 io_out[13]
port 88 nsew signal tristate
rlabel metal2 s 12070 119200 12126 120800 6 io_out[14]
port 89 nsew signal tristate
rlabel metal2 s 12806 119200 12862 120800 6 io_out[15]
port 90 nsew signal tristate
rlabel metal2 s 13450 119200 13506 120800 6 io_out[16]
port 91 nsew signal tristate
rlabel metal2 s 14186 119200 14242 120800 6 io_out[17]
port 92 nsew signal tristate
rlabel metal2 s 14830 119200 14886 120800 6 io_out[18]
port 93 nsew signal tristate
rlabel metal2 s 15566 119200 15622 120800 6 io_out[19]
port 94 nsew signal tristate
rlabel metal2 s 3054 119200 3110 120800 6 io_out[1]
port 95 nsew signal tristate
rlabel metal2 s 16302 119200 16358 120800 6 io_out[20]
port 96 nsew signal tristate
rlabel metal2 s 16946 119200 17002 120800 6 io_out[21]
port 97 nsew signal tristate
rlabel metal2 s 17682 119200 17738 120800 6 io_out[22]
port 98 nsew signal tristate
rlabel metal2 s 18326 119200 18382 120800 6 io_out[23]
port 99 nsew signal tristate
rlabel metal2 s 19062 119200 19118 120800 6 io_out[24]
port 100 nsew signal tristate
rlabel metal2 s 19706 119200 19762 120800 6 io_out[25]
port 101 nsew signal tristate
rlabel metal2 s 20442 119200 20498 120800 6 io_out[26]
port 102 nsew signal tristate
rlabel metal2 s 21086 119200 21142 120800 6 io_out[27]
port 103 nsew signal tristate
rlabel metal2 s 21822 119200 21878 120800 6 io_out[28]
port 104 nsew signal tristate
rlabel metal2 s 22466 119200 22522 120800 6 io_out[29]
port 105 nsew signal tristate
rlabel metal2 s 3790 119200 3846 120800 6 io_out[2]
port 106 nsew signal tristate
rlabel metal2 s 23202 119200 23258 120800 6 io_out[30]
port 107 nsew signal tristate
rlabel metal2 s 23846 119200 23902 120800 6 io_out[31]
port 108 nsew signal tristate
rlabel metal2 s 24582 119200 24638 120800 6 io_out[32]
port 109 nsew signal tristate
rlabel metal2 s 25318 119200 25374 120800 6 io_out[33]
port 110 nsew signal tristate
rlabel metal2 s 25962 119200 26018 120800 6 io_out[34]
port 111 nsew signal tristate
rlabel metal2 s 26698 119200 26754 120800 6 io_out[35]
port 112 nsew signal tristate
rlabel metal2 s 27342 119200 27398 120800 6 io_out[36]
port 113 nsew signal tristate
rlabel metal2 s 28078 119200 28134 120800 6 io_out[37]
port 114 nsew signal tristate
rlabel metal2 s 4434 119200 4490 120800 6 io_out[3]
port 115 nsew signal tristate
rlabel metal2 s 5170 119200 5226 120800 6 io_out[4]
port 116 nsew signal tristate
rlabel metal2 s 5814 119200 5870 120800 6 io_out[5]
port 117 nsew signal tristate
rlabel metal2 s 6550 119200 6606 120800 6 io_out[6]
port 118 nsew signal tristate
rlabel metal2 s 7194 119200 7250 120800 6 io_out[7]
port 119 nsew signal tristate
rlabel metal2 s 7930 119200 7986 120800 6 io_out[8]
port 120 nsew signal tristate
rlabel metal2 s 8666 119200 8722 120800 6 io_out[9]
port 121 nsew signal tristate
rlabel metal2 s 754 -800 810 800 8 irq[0]
port 122 nsew signal tristate
rlabel metal2 s 1030 -800 1086 800 8 irq[1]
port 123 nsew signal tristate
rlabel metal2 s 1398 -800 1454 800 8 irq[2]
port 124 nsew signal tristate
rlabel metal2 s 31942 119200 31998 120800 6 m_irqs[0]
port 125 nsew signal input
rlabel metal2 s 34334 119200 34390 120800 6 m_irqs[10]
port 126 nsew signal input
rlabel metal2 s 34518 119200 34574 120800 6 m_irqs[11]
port 127 nsew signal input
rlabel metal2 s 32218 119200 32274 120800 6 m_irqs[1]
port 128 nsew signal input
rlabel metal2 s 32494 119200 32550 120800 6 m_irqs[2]
port 129 nsew signal input
rlabel metal2 s 32678 119200 32734 120800 6 m_irqs[3]
port 130 nsew signal input
rlabel metal2 s 32954 119200 33010 120800 6 m_irqs[4]
port 131 nsew signal input
rlabel metal2 s 33138 119200 33194 120800 6 m_irqs[5]
port 132 nsew signal input
rlabel metal2 s 33414 119200 33470 120800 6 m_irqs[6]
port 133 nsew signal input
rlabel metal2 s 33598 119200 33654 120800 6 m_irqs[7]
port 134 nsew signal input
rlabel metal2 s 33874 119200 33930 120800 6 m_irqs[8]
port 135 nsew signal input
rlabel metal2 s 34058 119200 34114 120800 6 m_irqs[9]
port 136 nsew signal input
rlabel metal2 s 35530 -800 35586 800 8 m_wb_clk_i
port 137 nsew signal tristate
rlabel metal2 s 34794 119200 34850 120800 6 m_wb_rst_i
port 138 nsew signal tristate
rlabel metal2 s 35898 -800 35954 800 8 m_wbs_ack_o[0]
port 139 nsew signal input
rlabel metal3 s -800 113704 800 113824 4 m_wbs_ack_o[10]
port 140 nsew signal input
rlabel metal2 s 38474 119200 38530 120800 6 m_wbs_ack_o[11]
port 141 nsew signal input
rlabel metal3 s -800 104184 800 104304 4 m_wbs_ack_o[1]
port 142 nsew signal input
rlabel metal3 s -800 105816 800 105936 4 m_wbs_ack_o[2]
port 143 nsew signal input
rlabel metal2 s 35438 119200 35494 120800 6 m_wbs_ack_o[3]
port 144 nsew signal input
rlabel metal3 s -800 108944 800 109064 4 m_wbs_ack_o[4]
port 145 nsew signal input
rlabel metal2 s 36358 119200 36414 120800 6 m_wbs_ack_o[5]
port 146 nsew signal input
rlabel metal2 s 37094 119200 37150 120800 6 m_wbs_ack_o[6]
port 147 nsew signal input
rlabel metal2 s 37554 119200 37610 120800 6 m_wbs_ack_o[7]
port 148 nsew signal input
rlabel metal3 s 39200 116016 40800 116136 6 m_wbs_ack_o[8]
port 149 nsew signal input
rlabel metal2 s 37462 -800 37518 800 8 m_wbs_ack_o[9]
port 150 nsew signal input
rlabel metal3 s -800 103368 800 103488 4 m_wbs_adr_i[0]
port 151 nsew signal tristate
rlabel metal3 s -800 114520 800 114640 4 m_wbs_adr_i[10]
port 152 nsew signal tristate
rlabel metal2 s 38106 -800 38162 800 8 m_wbs_adr_i[11]
port 153 nsew signal tristate
rlabel metal2 s 36542 -800 36598 800 8 m_wbs_adr_i[1]
port 154 nsew signal tristate
rlabel metal3 s -800 106632 800 106752 4 m_wbs_adr_i[2]
port 155 nsew signal tristate
rlabel metal3 s -800 108128 800 108248 4 m_wbs_adr_i[3]
port 156 nsew signal tristate
rlabel metal3 s -800 109760 800 109880 4 m_wbs_adr_i[4]
port 157 nsew signal tristate
rlabel metal2 s 36634 119200 36690 120800 6 m_wbs_adr_i[5]
port 158 nsew signal tristate
rlabel metal3 s -800 110576 800 110696 4 m_wbs_adr_i[6]
port 159 nsew signal tristate
rlabel metal3 s 39200 115064 40800 115184 6 m_wbs_adr_i[7]
port 160 nsew signal tristate
rlabel metal2 s 38014 119200 38070 120800 6 m_wbs_adr_i[8]
port 161 nsew signal tristate
rlabel metal3 s -800 113024 800 113144 4 m_wbs_adr_i[9]
port 162 nsew signal tristate
rlabel metal2 s 36174 -800 36230 800 8 m_wbs_cs_i[0]
port 163 nsew signal tristate
rlabel metal2 s 38198 119200 38254 120800 6 m_wbs_cs_i[10]
port 164 nsew signal tristate
rlabel metal2 s 38474 -800 38530 800 8 m_wbs_cs_i[11]
port 165 nsew signal tristate
rlabel metal2 s 35254 119200 35310 120800 6 m_wbs_cs_i[1]
port 166 nsew signal tristate
rlabel metal3 s 39200 114656 40800 114776 6 m_wbs_cs_i[2]
port 167 nsew signal tristate
rlabel metal2 s 35714 119200 35770 120800 6 m_wbs_cs_i[3]
port 168 nsew signal tristate
rlabel metal2 s 36174 119200 36230 120800 6 m_wbs_cs_i[4]
port 169 nsew signal tristate
rlabel metal2 s 36818 119200 36874 120800 6 m_wbs_cs_i[5]
port 170 nsew signal tristate
rlabel metal2 s 37278 119200 37334 120800 6 m_wbs_cs_i[6]
port 171 nsew signal tristate
rlabel metal2 s 37738 119200 37794 120800 6 m_wbs_cs_i[7]
port 172 nsew signal tristate
rlabel metal3 s 39200 116424 40800 116544 6 m_wbs_cs_i[8]
port 173 nsew signal tristate
rlabel metal3 s 39200 116832 40800 116952 6 m_wbs_cs_i[9]
port 174 nsew signal tristate
rlabel metal2 s 34978 119200 35034 120800 6 m_wbs_dat_i[0]
port 175 nsew signal tristate
rlabel metal2 s 37830 -800 37886 800 8 m_wbs_dat_i[10]
port 176 nsew signal tristate
rlabel metal3 s -800 115336 800 115456 4 m_wbs_dat_i[11]
port 177 nsew signal tristate
rlabel metal2 s 38658 119200 38714 120800 6 m_wbs_dat_i[12]
port 178 nsew signal tristate
rlabel metal3 s 39200 117784 40800 117904 6 m_wbs_dat_i[13]
port 179 nsew signal tristate
rlabel metal3 s -800 116152 800 116272 4 m_wbs_dat_i[14]
port 180 nsew signal tristate
rlabel metal2 s 38934 119200 38990 120800 6 m_wbs_dat_i[15]
port 181 nsew signal tristate
rlabel metal3 s -800 116968 800 117088 4 m_wbs_dat_i[16]
port 182 nsew signal tristate
rlabel metal3 s 39200 118192 40800 118312 6 m_wbs_dat_i[17]
port 183 nsew signal tristate
rlabel metal3 s 39200 118736 40800 118856 6 m_wbs_dat_i[18]
port 184 nsew signal tristate
rlabel metal2 s 38750 -800 38806 800 8 m_wbs_dat_i[19]
port 185 nsew signal tristate
rlabel metal3 s -800 105000 800 105120 4 m_wbs_dat_i[1]
port 186 nsew signal tristate
rlabel metal2 s 39118 -800 39174 800 8 m_wbs_dat_i[20]
port 187 nsew signal tristate
rlabel metal2 s 39118 119200 39174 120800 6 m_wbs_dat_i[21]
port 188 nsew signal tristate
rlabel metal3 s -800 117784 800 117904 4 m_wbs_dat_i[22]
port 189 nsew signal tristate
rlabel metal2 s 39394 119200 39450 120800 6 m_wbs_dat_i[23]
port 190 nsew signal tristate
rlabel metal2 s 39578 119200 39634 120800 6 m_wbs_dat_i[24]
port 191 nsew signal tristate
rlabel metal2 s 39394 -800 39450 800 8 m_wbs_dat_i[25]
port 192 nsew signal tristate
rlabel metal3 s -800 118600 800 118720 4 m_wbs_dat_i[26]
port 193 nsew signal tristate
rlabel metal3 s -800 119416 800 119536 4 m_wbs_dat_i[27]
port 194 nsew signal tristate
rlabel metal2 s 39762 -800 39818 800 8 m_wbs_dat_i[28]
port 195 nsew signal tristate
rlabel metal3 s 39200 119144 40800 119264 6 m_wbs_dat_i[29]
port 196 nsew signal tristate
rlabel metal3 s -800 107312 800 107432 4 m_wbs_dat_i[2]
port 197 nsew signal tristate
rlabel metal3 s 39200 119552 40800 119672 6 m_wbs_dat_i[30]
port 198 nsew signal tristate
rlabel metal2 s 39854 119200 39910 120800 6 m_wbs_dat_i[31]
port 199 nsew signal tristate
rlabel metal2 s 35898 119200 35954 120800 6 m_wbs_dat_i[3]
port 200 nsew signal tristate
rlabel metal2 s 36818 -800 36874 800 8 m_wbs_dat_i[4]
port 201 nsew signal tristate
rlabel metal2 s 37186 -800 37242 800 8 m_wbs_dat_i[5]
port 202 nsew signal tristate
rlabel metal3 s -800 111392 800 111512 4 m_wbs_dat_i[6]
port 203 nsew signal tristate
rlabel metal3 s 39200 115608 40800 115728 6 m_wbs_dat_i[7]
port 204 nsew signal tristate
rlabel metal3 s -800 112208 800 112328 4 m_wbs_dat_i[8]
port 205 nsew signal tristate
rlabel metal3 s 39200 117376 40800 117496 6 m_wbs_dat_i[9]
port 206 nsew signal tristate
rlabel metal3 s 39200 144 40800 264 6 m_wbs_dat_o_0[0]
port 207 nsew signal input
rlabel metal3 s 39200 4496 40800 4616 6 m_wbs_dat_o_0[10]
port 208 nsew signal input
rlabel metal3 s 39200 5040 40800 5160 6 m_wbs_dat_o_0[11]
port 209 nsew signal input
rlabel metal3 s 39200 5448 40800 5568 6 m_wbs_dat_o_0[12]
port 210 nsew signal input
rlabel metal3 s 39200 5856 40800 5976 6 m_wbs_dat_o_0[13]
port 211 nsew signal input
rlabel metal3 s 39200 6400 40800 6520 6 m_wbs_dat_o_0[14]
port 212 nsew signal input
rlabel metal3 s 39200 6808 40800 6928 6 m_wbs_dat_o_0[15]
port 213 nsew signal input
rlabel metal3 s 39200 7216 40800 7336 6 m_wbs_dat_o_0[16]
port 214 nsew signal input
rlabel metal3 s 39200 7624 40800 7744 6 m_wbs_dat_o_0[17]
port 215 nsew signal input
rlabel metal3 s 39200 8168 40800 8288 6 m_wbs_dat_o_0[18]
port 216 nsew signal input
rlabel metal3 s 39200 8576 40800 8696 6 m_wbs_dat_o_0[19]
port 217 nsew signal input
rlabel metal3 s 39200 552 40800 672 6 m_wbs_dat_o_0[1]
port 218 nsew signal input
rlabel metal3 s 39200 8984 40800 9104 6 m_wbs_dat_o_0[20]
port 219 nsew signal input
rlabel metal3 s 39200 9528 40800 9648 6 m_wbs_dat_o_0[21]
port 220 nsew signal input
rlabel metal3 s 39200 9936 40800 10056 6 m_wbs_dat_o_0[22]
port 221 nsew signal input
rlabel metal3 s 39200 10344 40800 10464 6 m_wbs_dat_o_0[23]
port 222 nsew signal input
rlabel metal3 s 39200 10752 40800 10872 6 m_wbs_dat_o_0[24]
port 223 nsew signal input
rlabel metal3 s 39200 11296 40800 11416 6 m_wbs_dat_o_0[25]
port 224 nsew signal input
rlabel metal3 s 39200 11704 40800 11824 6 m_wbs_dat_o_0[26]
port 225 nsew signal input
rlabel metal3 s 39200 12112 40800 12232 6 m_wbs_dat_o_0[27]
port 226 nsew signal input
rlabel metal3 s 39200 12656 40800 12776 6 m_wbs_dat_o_0[28]
port 227 nsew signal input
rlabel metal3 s 39200 13064 40800 13184 6 m_wbs_dat_o_0[29]
port 228 nsew signal input
rlabel metal3 s 39200 960 40800 1080 6 m_wbs_dat_o_0[2]
port 229 nsew signal input
rlabel metal3 s 39200 13472 40800 13592 6 m_wbs_dat_o_0[30]
port 230 nsew signal input
rlabel metal3 s 39200 14016 40800 14136 6 m_wbs_dat_o_0[31]
port 231 nsew signal input
rlabel metal3 s 39200 1368 40800 1488 6 m_wbs_dat_o_0[3]
port 232 nsew signal input
rlabel metal3 s 39200 1912 40800 2032 6 m_wbs_dat_o_0[4]
port 233 nsew signal input
rlabel metal3 s 39200 2320 40800 2440 6 m_wbs_dat_o_0[5]
port 234 nsew signal input
rlabel metal3 s 39200 2728 40800 2848 6 m_wbs_dat_o_0[6]
port 235 nsew signal input
rlabel metal3 s 39200 3272 40800 3392 6 m_wbs_dat_o_0[7]
port 236 nsew signal input
rlabel metal3 s 39200 3680 40800 3800 6 m_wbs_dat_o_0[8]
port 237 nsew signal input
rlabel metal3 s 39200 4088 40800 4208 6 m_wbs_dat_o_0[9]
port 238 nsew signal input
rlabel metal3 s 39200 14832 40800 14952 6 m_wbs_dat_o_10[0]
port 239 nsew signal input
rlabel metal3 s 39200 28296 40800 28416 6 m_wbs_dat_o_10[10]
port 240 nsew signal input
rlabel metal3 s 39200 29656 40800 29776 6 m_wbs_dat_o_10[11]
port 241 nsew signal input
rlabel metal3 s 39200 31016 40800 31136 6 m_wbs_dat_o_10[12]
port 242 nsew signal input
rlabel metal3 s 39200 32240 40800 32360 6 m_wbs_dat_o_10[13]
port 243 nsew signal input
rlabel metal3 s 39200 33600 40800 33720 6 m_wbs_dat_o_10[14]
port 244 nsew signal input
rlabel metal3 s 39200 34960 40800 35080 6 m_wbs_dat_o_10[15]
port 245 nsew signal input
rlabel metal3 s 39200 36320 40800 36440 6 m_wbs_dat_o_10[16]
port 246 nsew signal input
rlabel metal3 s 39200 37680 40800 37800 6 m_wbs_dat_o_10[17]
port 247 nsew signal input
rlabel metal3 s 39200 39040 40800 39160 6 m_wbs_dat_o_10[18]
port 248 nsew signal input
rlabel metal3 s 39200 40400 40800 40520 6 m_wbs_dat_o_10[19]
port 249 nsew signal input
rlabel metal3 s 39200 16192 40800 16312 6 m_wbs_dat_o_10[1]
port 250 nsew signal input
rlabel metal3 s 39200 41760 40800 41880 6 m_wbs_dat_o_10[20]
port 251 nsew signal input
rlabel metal3 s 39200 42984 40800 43104 6 m_wbs_dat_o_10[21]
port 252 nsew signal input
rlabel metal3 s 39200 44344 40800 44464 6 m_wbs_dat_o_10[22]
port 253 nsew signal input
rlabel metal3 s 39200 45704 40800 45824 6 m_wbs_dat_o_10[23]
port 254 nsew signal input
rlabel metal3 s 39200 47064 40800 47184 6 m_wbs_dat_o_10[24]
port 255 nsew signal input
rlabel metal3 s 39200 48424 40800 48544 6 m_wbs_dat_o_10[25]
port 256 nsew signal input
rlabel metal3 s 39200 49784 40800 49904 6 m_wbs_dat_o_10[26]
port 257 nsew signal input
rlabel metal3 s 39200 51144 40800 51264 6 m_wbs_dat_o_10[27]
port 258 nsew signal input
rlabel metal3 s 39200 52504 40800 52624 6 m_wbs_dat_o_10[28]
port 259 nsew signal input
rlabel metal3 s 39200 53728 40800 53848 6 m_wbs_dat_o_10[29]
port 260 nsew signal input
rlabel metal3 s 39200 17552 40800 17672 6 m_wbs_dat_o_10[2]
port 261 nsew signal input
rlabel metal3 s 39200 55088 40800 55208 6 m_wbs_dat_o_10[30]
port 262 nsew signal input
rlabel metal3 s 39200 56448 40800 56568 6 m_wbs_dat_o_10[31]
port 263 nsew signal input
rlabel metal3 s 39200 18912 40800 19032 6 m_wbs_dat_o_10[3]
port 264 nsew signal input
rlabel metal3 s 39200 20272 40800 20392 6 m_wbs_dat_o_10[4]
port 265 nsew signal input
rlabel metal3 s 39200 21496 40800 21616 6 m_wbs_dat_o_10[5]
port 266 nsew signal input
rlabel metal3 s 39200 22856 40800 22976 6 m_wbs_dat_o_10[6]
port 267 nsew signal input
rlabel metal3 s 39200 24216 40800 24336 6 m_wbs_dat_o_10[7]
port 268 nsew signal input
rlabel metal3 s 39200 25576 40800 25696 6 m_wbs_dat_o_10[8]
port 269 nsew signal input
rlabel metal3 s 39200 26936 40800 27056 6 m_wbs_dat_o_10[9]
port 270 nsew signal input
rlabel metal3 s 39200 15240 40800 15360 6 m_wbs_dat_o_11[0]
port 271 nsew signal input
rlabel metal3 s 39200 28704 40800 28824 6 m_wbs_dat_o_11[10]
port 272 nsew signal input
rlabel metal3 s 39200 30064 40800 30184 6 m_wbs_dat_o_11[11]
port 273 nsew signal input
rlabel metal3 s 39200 31424 40800 31544 6 m_wbs_dat_o_11[12]
port 274 nsew signal input
rlabel metal3 s 39200 32784 40800 32904 6 m_wbs_dat_o_11[13]
port 275 nsew signal input
rlabel metal3 s 39200 34144 40800 34264 6 m_wbs_dat_o_11[14]
port 276 nsew signal input
rlabel metal3 s 39200 35368 40800 35488 6 m_wbs_dat_o_11[15]
port 277 nsew signal input
rlabel metal3 s 39200 36728 40800 36848 6 m_wbs_dat_o_11[16]
port 278 nsew signal input
rlabel metal3 s 39200 38088 40800 38208 6 m_wbs_dat_o_11[17]
port 279 nsew signal input
rlabel metal3 s 39200 39448 40800 39568 6 m_wbs_dat_o_11[18]
port 280 nsew signal input
rlabel metal3 s 39200 40808 40800 40928 6 m_wbs_dat_o_11[19]
port 281 nsew signal input
rlabel metal3 s 39200 16600 40800 16720 6 m_wbs_dat_o_11[1]
port 282 nsew signal input
rlabel metal3 s 39200 42168 40800 42288 6 m_wbs_dat_o_11[20]
port 283 nsew signal input
rlabel metal3 s 39200 43528 40800 43648 6 m_wbs_dat_o_11[21]
port 284 nsew signal input
rlabel metal3 s 39200 44888 40800 45008 6 m_wbs_dat_o_11[22]
port 285 nsew signal input
rlabel metal3 s 39200 46112 40800 46232 6 m_wbs_dat_o_11[23]
port 286 nsew signal input
rlabel metal3 s 39200 47472 40800 47592 6 m_wbs_dat_o_11[24]
port 287 nsew signal input
rlabel metal3 s 39200 48832 40800 48952 6 m_wbs_dat_o_11[25]
port 288 nsew signal input
rlabel metal3 s 39200 50192 40800 50312 6 m_wbs_dat_o_11[26]
port 289 nsew signal input
rlabel metal3 s 39200 51552 40800 51672 6 m_wbs_dat_o_11[27]
port 290 nsew signal input
rlabel metal3 s 39200 52912 40800 53032 6 m_wbs_dat_o_11[28]
port 291 nsew signal input
rlabel metal3 s 39200 54272 40800 54392 6 m_wbs_dat_o_11[29]
port 292 nsew signal input
rlabel metal3 s 39200 17960 40800 18080 6 m_wbs_dat_o_11[2]
port 293 nsew signal input
rlabel metal3 s 39200 55632 40800 55752 6 m_wbs_dat_o_11[30]
port 294 nsew signal input
rlabel metal3 s 39200 56856 40800 56976 6 m_wbs_dat_o_11[31]
port 295 nsew signal input
rlabel metal3 s 39200 19320 40800 19440 6 m_wbs_dat_o_11[3]
port 296 nsew signal input
rlabel metal3 s 39200 20680 40800 20800 6 m_wbs_dat_o_11[4]
port 297 nsew signal input
rlabel metal3 s 39200 22040 40800 22160 6 m_wbs_dat_o_11[5]
port 298 nsew signal input
rlabel metal3 s 39200 23400 40800 23520 6 m_wbs_dat_o_11[6]
port 299 nsew signal input
rlabel metal3 s 39200 24760 40800 24880 6 m_wbs_dat_o_11[7]
port 300 nsew signal input
rlabel metal3 s 39200 25984 40800 26104 6 m_wbs_dat_o_11[8]
port 301 nsew signal input
rlabel metal3 s 39200 27344 40800 27464 6 m_wbs_dat_o_11[9]
port 302 nsew signal input
rlabel metal3 s 39200 14424 40800 14544 6 m_wbs_dat_o_1[0]
port 303 nsew signal input
rlabel metal3 s 39200 27888 40800 28008 6 m_wbs_dat_o_1[10]
port 304 nsew signal input
rlabel metal3 s 39200 29112 40800 29232 6 m_wbs_dat_o_1[11]
port 305 nsew signal input
rlabel metal3 s 39200 30472 40800 30592 6 m_wbs_dat_o_1[12]
port 306 nsew signal input
rlabel metal3 s 39200 31832 40800 31952 6 m_wbs_dat_o_1[13]
port 307 nsew signal input
rlabel metal3 s 39200 33192 40800 33312 6 m_wbs_dat_o_1[14]
port 308 nsew signal input
rlabel metal3 s 39200 34552 40800 34672 6 m_wbs_dat_o_1[15]
port 309 nsew signal input
rlabel metal3 s 39200 35912 40800 36032 6 m_wbs_dat_o_1[16]
port 310 nsew signal input
rlabel metal3 s 39200 37272 40800 37392 6 m_wbs_dat_o_1[17]
port 311 nsew signal input
rlabel metal3 s 39200 38632 40800 38752 6 m_wbs_dat_o_1[18]
port 312 nsew signal input
rlabel metal3 s 39200 39856 40800 39976 6 m_wbs_dat_o_1[19]
port 313 nsew signal input
rlabel metal3 s 39200 15784 40800 15904 6 m_wbs_dat_o_1[1]
port 314 nsew signal input
rlabel metal3 s 39200 41216 40800 41336 6 m_wbs_dat_o_1[20]
port 315 nsew signal input
rlabel metal3 s 39200 42576 40800 42696 6 m_wbs_dat_o_1[21]
port 316 nsew signal input
rlabel metal3 s 39200 43936 40800 44056 6 m_wbs_dat_o_1[22]
port 317 nsew signal input
rlabel metal3 s 39200 45296 40800 45416 6 m_wbs_dat_o_1[23]
port 318 nsew signal input
rlabel metal3 s 39200 46656 40800 46776 6 m_wbs_dat_o_1[24]
port 319 nsew signal input
rlabel metal3 s 39200 48016 40800 48136 6 m_wbs_dat_o_1[25]
port 320 nsew signal input
rlabel metal3 s 39200 49376 40800 49496 6 m_wbs_dat_o_1[26]
port 321 nsew signal input
rlabel metal3 s 39200 50600 40800 50720 6 m_wbs_dat_o_1[27]
port 322 nsew signal input
rlabel metal3 s 39200 51960 40800 52080 6 m_wbs_dat_o_1[28]
port 323 nsew signal input
rlabel metal3 s 39200 53320 40800 53440 6 m_wbs_dat_o_1[29]
port 324 nsew signal input
rlabel metal3 s 39200 17144 40800 17264 6 m_wbs_dat_o_1[2]
port 325 nsew signal input
rlabel metal3 s 39200 54680 40800 54800 6 m_wbs_dat_o_1[30]
port 326 nsew signal input
rlabel metal3 s 39200 56040 40800 56160 6 m_wbs_dat_o_1[31]
port 327 nsew signal input
rlabel metal3 s 39200 18368 40800 18488 6 m_wbs_dat_o_1[3]
port 328 nsew signal input
rlabel metal3 s 39200 19728 40800 19848 6 m_wbs_dat_o_1[4]
port 329 nsew signal input
rlabel metal3 s 39200 21088 40800 21208 6 m_wbs_dat_o_1[5]
port 330 nsew signal input
rlabel metal3 s 39200 22448 40800 22568 6 m_wbs_dat_o_1[6]
port 331 nsew signal input
rlabel metal3 s 39200 23808 40800 23928 6 m_wbs_dat_o_1[7]
port 332 nsew signal input
rlabel metal3 s 39200 25168 40800 25288 6 m_wbs_dat_o_1[8]
port 333 nsew signal input
rlabel metal3 s 39200 26528 40800 26648 6 m_wbs_dat_o_1[9]
port 334 nsew signal input
rlabel metal3 s 39200 57400 40800 57520 6 m_wbs_dat_o_2[0]
port 335 nsew signal input
rlabel metal3 s 39200 61888 40800 62008 6 m_wbs_dat_o_2[10]
port 336 nsew signal input
rlabel metal3 s 39200 62296 40800 62416 6 m_wbs_dat_o_2[11]
port 337 nsew signal input
rlabel metal3 s 39200 62704 40800 62824 6 m_wbs_dat_o_2[12]
port 338 nsew signal input
rlabel metal3 s 39200 63248 40800 63368 6 m_wbs_dat_o_2[13]
port 339 nsew signal input
rlabel metal3 s 39200 63656 40800 63776 6 m_wbs_dat_o_2[14]
port 340 nsew signal input
rlabel metal3 s 39200 64064 40800 64184 6 m_wbs_dat_o_2[15]
port 341 nsew signal input
rlabel metal3 s 39200 64472 40800 64592 6 m_wbs_dat_o_2[16]
port 342 nsew signal input
rlabel metal3 s 39200 65016 40800 65136 6 m_wbs_dat_o_2[17]
port 343 nsew signal input
rlabel metal3 s 39200 65424 40800 65544 6 m_wbs_dat_o_2[18]
port 344 nsew signal input
rlabel metal3 s 39200 65832 40800 65952 6 m_wbs_dat_o_2[19]
port 345 nsew signal input
rlabel metal3 s 39200 57808 40800 57928 6 m_wbs_dat_o_2[1]
port 346 nsew signal input
rlabel metal3 s 39200 66376 40800 66496 6 m_wbs_dat_o_2[20]
port 347 nsew signal input
rlabel metal3 s 39200 66784 40800 66904 6 m_wbs_dat_o_2[21]
port 348 nsew signal input
rlabel metal3 s 39200 67192 40800 67312 6 m_wbs_dat_o_2[22]
port 349 nsew signal input
rlabel metal3 s 39200 67600 40800 67720 6 m_wbs_dat_o_2[23]
port 350 nsew signal input
rlabel metal3 s 39200 68144 40800 68264 6 m_wbs_dat_o_2[24]
port 351 nsew signal input
rlabel metal3 s 39200 68552 40800 68672 6 m_wbs_dat_o_2[25]
port 352 nsew signal input
rlabel metal3 s 39200 68960 40800 69080 6 m_wbs_dat_o_2[26]
port 353 nsew signal input
rlabel metal3 s 39200 69504 40800 69624 6 m_wbs_dat_o_2[27]
port 354 nsew signal input
rlabel metal3 s 39200 69912 40800 70032 6 m_wbs_dat_o_2[28]
port 355 nsew signal input
rlabel metal3 s 39200 70320 40800 70440 6 m_wbs_dat_o_2[29]
port 356 nsew signal input
rlabel metal3 s 39200 58216 40800 58336 6 m_wbs_dat_o_2[2]
port 357 nsew signal input
rlabel metal3 s 39200 70728 40800 70848 6 m_wbs_dat_o_2[30]
port 358 nsew signal input
rlabel metal3 s 39200 71272 40800 71392 6 m_wbs_dat_o_2[31]
port 359 nsew signal input
rlabel metal3 s 39200 58760 40800 58880 6 m_wbs_dat_o_2[3]
port 360 nsew signal input
rlabel metal3 s 39200 59168 40800 59288 6 m_wbs_dat_o_2[4]
port 361 nsew signal input
rlabel metal3 s 39200 59576 40800 59696 6 m_wbs_dat_o_2[5]
port 362 nsew signal input
rlabel metal3 s 39200 60120 40800 60240 6 m_wbs_dat_o_2[6]
port 363 nsew signal input
rlabel metal3 s 39200 60528 40800 60648 6 m_wbs_dat_o_2[7]
port 364 nsew signal input
rlabel metal3 s 39200 60936 40800 61056 6 m_wbs_dat_o_2[8]
port 365 nsew signal input
rlabel metal3 s 39200 61344 40800 61464 6 m_wbs_dat_o_2[9]
port 366 nsew signal input
rlabel metal3 s 39200 71680 40800 71800 6 m_wbs_dat_o_3[0]
port 367 nsew signal input
rlabel metal3 s 39200 76168 40800 76288 6 m_wbs_dat_o_3[10]
port 368 nsew signal input
rlabel metal3 s 39200 76576 40800 76696 6 m_wbs_dat_o_3[11]
port 369 nsew signal input
rlabel metal3 s 39200 77120 40800 77240 6 m_wbs_dat_o_3[12]
port 370 nsew signal input
rlabel metal3 s 39200 77528 40800 77648 6 m_wbs_dat_o_3[13]
port 371 nsew signal input
rlabel metal3 s 39200 77936 40800 78056 6 m_wbs_dat_o_3[14]
port 372 nsew signal input
rlabel metal3 s 39200 78344 40800 78464 6 m_wbs_dat_o_3[15]
port 373 nsew signal input
rlabel metal3 s 39200 78888 40800 79008 6 m_wbs_dat_o_3[16]
port 374 nsew signal input
rlabel metal3 s 39200 79296 40800 79416 6 m_wbs_dat_o_3[17]
port 375 nsew signal input
rlabel metal3 s 39200 79704 40800 79824 6 m_wbs_dat_o_3[18]
port 376 nsew signal input
rlabel metal3 s 39200 80248 40800 80368 6 m_wbs_dat_o_3[19]
port 377 nsew signal input
rlabel metal3 s 39200 72088 40800 72208 6 m_wbs_dat_o_3[1]
port 378 nsew signal input
rlabel metal3 s 39200 80656 40800 80776 6 m_wbs_dat_o_3[20]
port 379 nsew signal input
rlabel metal3 s 39200 81064 40800 81184 6 m_wbs_dat_o_3[21]
port 380 nsew signal input
rlabel metal3 s 39200 81472 40800 81592 6 m_wbs_dat_o_3[22]
port 381 nsew signal input
rlabel metal3 s 39200 82016 40800 82136 6 m_wbs_dat_o_3[23]
port 382 nsew signal input
rlabel metal3 s 39200 82424 40800 82544 6 m_wbs_dat_o_3[24]
port 383 nsew signal input
rlabel metal3 s 39200 82832 40800 82952 6 m_wbs_dat_o_3[25]
port 384 nsew signal input
rlabel metal3 s 39200 83376 40800 83496 6 m_wbs_dat_o_3[26]
port 385 nsew signal input
rlabel metal3 s 39200 83784 40800 83904 6 m_wbs_dat_o_3[27]
port 386 nsew signal input
rlabel metal3 s 39200 84192 40800 84312 6 m_wbs_dat_o_3[28]
port 387 nsew signal input
rlabel metal3 s 39200 84736 40800 84856 6 m_wbs_dat_o_3[29]
port 388 nsew signal input
rlabel metal3 s 39200 72632 40800 72752 6 m_wbs_dat_o_3[2]
port 389 nsew signal input
rlabel metal3 s 39200 85144 40800 85264 6 m_wbs_dat_o_3[30]
port 390 nsew signal input
rlabel metal3 s 39200 85552 40800 85672 6 m_wbs_dat_o_3[31]
port 391 nsew signal input
rlabel metal3 s 39200 73040 40800 73160 6 m_wbs_dat_o_3[3]
port 392 nsew signal input
rlabel metal3 s 39200 73448 40800 73568 6 m_wbs_dat_o_3[4]
port 393 nsew signal input
rlabel metal3 s 39200 73992 40800 74112 6 m_wbs_dat_o_3[5]
port 394 nsew signal input
rlabel metal3 s 39200 74400 40800 74520 6 m_wbs_dat_o_3[6]
port 395 nsew signal input
rlabel metal3 s 39200 74808 40800 74928 6 m_wbs_dat_o_3[7]
port 396 nsew signal input
rlabel metal3 s 39200 75216 40800 75336 6 m_wbs_dat_o_3[8]
port 397 nsew signal input
rlabel metal3 s 39200 75760 40800 75880 6 m_wbs_dat_o_3[9]
port 398 nsew signal input
rlabel metal3 s 39200 85960 40800 86080 6 m_wbs_dat_o_4[0]
port 399 nsew signal input
rlabel metal3 s 39200 90448 40800 90568 6 m_wbs_dat_o_4[10]
port 400 nsew signal input
rlabel metal3 s 39200 90992 40800 91112 6 m_wbs_dat_o_4[11]
port 401 nsew signal input
rlabel metal3 s 39200 91400 40800 91520 6 m_wbs_dat_o_4[12]
port 402 nsew signal input
rlabel metal3 s 39200 91808 40800 91928 6 m_wbs_dat_o_4[13]
port 403 nsew signal input
rlabel metal3 s 39200 92216 40800 92336 6 m_wbs_dat_o_4[14]
port 404 nsew signal input
rlabel metal3 s 39200 92760 40800 92880 6 m_wbs_dat_o_4[15]
port 405 nsew signal input
rlabel metal3 s 39200 93168 40800 93288 6 m_wbs_dat_o_4[16]
port 406 nsew signal input
rlabel metal3 s 39200 93576 40800 93696 6 m_wbs_dat_o_4[17]
port 407 nsew signal input
rlabel metal3 s 39200 94120 40800 94240 6 m_wbs_dat_o_4[18]
port 408 nsew signal input
rlabel metal3 s 39200 94528 40800 94648 6 m_wbs_dat_o_4[19]
port 409 nsew signal input
rlabel metal3 s 39200 86504 40800 86624 6 m_wbs_dat_o_4[1]
port 410 nsew signal input
rlabel metal3 s 39200 94936 40800 95056 6 m_wbs_dat_o_4[20]
port 411 nsew signal input
rlabel metal3 s 39200 95344 40800 95464 6 m_wbs_dat_o_4[21]
port 412 nsew signal input
rlabel metal3 s 39200 95888 40800 96008 6 m_wbs_dat_o_4[22]
port 413 nsew signal input
rlabel metal3 s 39200 96296 40800 96416 6 m_wbs_dat_o_4[23]
port 414 nsew signal input
rlabel metal3 s 39200 96704 40800 96824 6 m_wbs_dat_o_4[24]
port 415 nsew signal input
rlabel metal3 s 39200 97248 40800 97368 6 m_wbs_dat_o_4[25]
port 416 nsew signal input
rlabel metal3 s 39200 97656 40800 97776 6 m_wbs_dat_o_4[26]
port 417 nsew signal input
rlabel metal3 s 39200 98064 40800 98184 6 m_wbs_dat_o_4[27]
port 418 nsew signal input
rlabel metal3 s 39200 98608 40800 98728 6 m_wbs_dat_o_4[28]
port 419 nsew signal input
rlabel metal3 s 39200 99016 40800 99136 6 m_wbs_dat_o_4[29]
port 420 nsew signal input
rlabel metal3 s 39200 86912 40800 87032 6 m_wbs_dat_o_4[2]
port 421 nsew signal input
rlabel metal3 s 39200 99424 40800 99544 6 m_wbs_dat_o_4[30]
port 422 nsew signal input
rlabel metal3 s 39200 99832 40800 99952 6 m_wbs_dat_o_4[31]
port 423 nsew signal input
rlabel metal3 s 39200 87320 40800 87440 6 m_wbs_dat_o_4[3]
port 424 nsew signal input
rlabel metal3 s 39200 87864 40800 87984 6 m_wbs_dat_o_4[4]
port 425 nsew signal input
rlabel metal3 s 39200 88272 40800 88392 6 m_wbs_dat_o_4[5]
port 426 nsew signal input
rlabel metal3 s 39200 88680 40800 88800 6 m_wbs_dat_o_4[6]
port 427 nsew signal input
rlabel metal3 s 39200 89088 40800 89208 6 m_wbs_dat_o_4[7]
port 428 nsew signal input
rlabel metal3 s 39200 89632 40800 89752 6 m_wbs_dat_o_4[8]
port 429 nsew signal input
rlabel metal3 s 39200 90040 40800 90160 6 m_wbs_dat_o_4[9]
port 430 nsew signal input
rlabel metal3 s 39200 100376 40800 100496 6 m_wbs_dat_o_5[0]
port 431 nsew signal input
rlabel metal3 s 39200 104864 40800 104984 6 m_wbs_dat_o_5[10]
port 432 nsew signal input
rlabel metal3 s 39200 105272 40800 105392 6 m_wbs_dat_o_5[11]
port 433 nsew signal input
rlabel metal3 s 39200 105680 40800 105800 6 m_wbs_dat_o_5[12]
port 434 nsew signal input
rlabel metal3 s 39200 106088 40800 106208 6 m_wbs_dat_o_5[13]
port 435 nsew signal input
rlabel metal3 s 39200 106632 40800 106752 6 m_wbs_dat_o_5[14]
port 436 nsew signal input
rlabel metal3 s 39200 107040 40800 107160 6 m_wbs_dat_o_5[15]
port 437 nsew signal input
rlabel metal3 s 39200 107448 40800 107568 6 m_wbs_dat_o_5[16]
port 438 nsew signal input
rlabel metal3 s 39200 107992 40800 108112 6 m_wbs_dat_o_5[17]
port 439 nsew signal input
rlabel metal3 s 39200 108400 40800 108520 6 m_wbs_dat_o_5[18]
port 440 nsew signal input
rlabel metal3 s 39200 108808 40800 108928 6 m_wbs_dat_o_5[19]
port 441 nsew signal input
rlabel metal3 s 39200 100784 40800 100904 6 m_wbs_dat_o_5[1]
port 442 nsew signal input
rlabel metal3 s 39200 109352 40800 109472 6 m_wbs_dat_o_5[20]
port 443 nsew signal input
rlabel metal3 s 39200 109760 40800 109880 6 m_wbs_dat_o_5[21]
port 444 nsew signal input
rlabel metal3 s 39200 110168 40800 110288 6 m_wbs_dat_o_5[22]
port 445 nsew signal input
rlabel metal3 s 39200 110576 40800 110696 6 m_wbs_dat_o_5[23]
port 446 nsew signal input
rlabel metal3 s 39200 111120 40800 111240 6 m_wbs_dat_o_5[24]
port 447 nsew signal input
rlabel metal3 s 39200 111528 40800 111648 6 m_wbs_dat_o_5[25]
port 448 nsew signal input
rlabel metal3 s 39200 111936 40800 112056 6 m_wbs_dat_o_5[26]
port 449 nsew signal input
rlabel metal3 s 39200 112480 40800 112600 6 m_wbs_dat_o_5[27]
port 450 nsew signal input
rlabel metal3 s 39200 112888 40800 113008 6 m_wbs_dat_o_5[28]
port 451 nsew signal input
rlabel metal3 s 39200 113296 40800 113416 6 m_wbs_dat_o_5[29]
port 452 nsew signal input
rlabel metal3 s 39200 101192 40800 101312 6 m_wbs_dat_o_5[2]
port 453 nsew signal input
rlabel metal3 s 39200 113704 40800 113824 6 m_wbs_dat_o_5[30]
port 454 nsew signal input
rlabel metal3 s 39200 114248 40800 114368 6 m_wbs_dat_o_5[31]
port 455 nsew signal input
rlabel metal3 s 39200 101736 40800 101856 6 m_wbs_dat_o_5[3]
port 456 nsew signal input
rlabel metal3 s 39200 102144 40800 102264 6 m_wbs_dat_o_5[4]
port 457 nsew signal input
rlabel metal3 s 39200 102552 40800 102672 6 m_wbs_dat_o_5[5]
port 458 nsew signal input
rlabel metal3 s 39200 102960 40800 103080 6 m_wbs_dat_o_5[6]
port 459 nsew signal input
rlabel metal3 s 39200 103504 40800 103624 6 m_wbs_dat_o_5[7]
port 460 nsew signal input
rlabel metal3 s 39200 103912 40800 104032 6 m_wbs_dat_o_5[8]
port 461 nsew signal input
rlabel metal3 s 39200 104320 40800 104440 6 m_wbs_dat_o_5[9]
port 462 nsew signal input
rlabel metal3 s -800 280 800 400 4 m_wbs_dat_o_6[0]
port 463 nsew signal input
rlabel metal3 s -800 8168 800 8288 4 m_wbs_dat_o_6[10]
port 464 nsew signal input
rlabel metal3 s -800 8984 800 9104 4 m_wbs_dat_o_6[11]
port 465 nsew signal input
rlabel metal3 s -800 9800 800 9920 4 m_wbs_dat_o_6[12]
port 466 nsew signal input
rlabel metal3 s -800 10616 800 10736 4 m_wbs_dat_o_6[13]
port 467 nsew signal input
rlabel metal3 s -800 11432 800 11552 4 m_wbs_dat_o_6[14]
port 468 nsew signal input
rlabel metal3 s -800 12248 800 12368 4 m_wbs_dat_o_6[15]
port 469 nsew signal input
rlabel metal3 s -800 13064 800 13184 4 m_wbs_dat_o_6[16]
port 470 nsew signal input
rlabel metal3 s -800 13744 800 13864 4 m_wbs_dat_o_6[17]
port 471 nsew signal input
rlabel metal3 s -800 14560 800 14680 4 m_wbs_dat_o_6[18]
port 472 nsew signal input
rlabel metal3 s -800 15376 800 15496 4 m_wbs_dat_o_6[19]
port 473 nsew signal input
rlabel metal3 s -800 960 800 1080 4 m_wbs_dat_o_6[1]
port 474 nsew signal input
rlabel metal3 s -800 16192 800 16312 4 m_wbs_dat_o_6[20]
port 475 nsew signal input
rlabel metal3 s -800 17008 800 17128 4 m_wbs_dat_o_6[21]
port 476 nsew signal input
rlabel metal3 s -800 17824 800 17944 4 m_wbs_dat_o_6[22]
port 477 nsew signal input
rlabel metal3 s -800 18640 800 18760 4 m_wbs_dat_o_6[23]
port 478 nsew signal input
rlabel metal3 s -800 19456 800 19576 4 m_wbs_dat_o_6[24]
port 479 nsew signal input
rlabel metal3 s -800 20272 800 20392 4 m_wbs_dat_o_6[25]
port 480 nsew signal input
rlabel metal3 s -800 20952 800 21072 4 m_wbs_dat_o_6[26]
port 481 nsew signal input
rlabel metal3 s -800 21768 800 21888 4 m_wbs_dat_o_6[27]
port 482 nsew signal input
rlabel metal3 s -800 22584 800 22704 4 m_wbs_dat_o_6[28]
port 483 nsew signal input
rlabel metal3 s -800 23400 800 23520 4 m_wbs_dat_o_6[29]
port 484 nsew signal input
rlabel metal3 s -800 1776 800 1896 4 m_wbs_dat_o_6[2]
port 485 nsew signal input
rlabel metal3 s -800 24216 800 24336 4 m_wbs_dat_o_6[30]
port 486 nsew signal input
rlabel metal3 s -800 25032 800 25152 4 m_wbs_dat_o_6[31]
port 487 nsew signal input
rlabel metal3 s -800 2592 800 2712 4 m_wbs_dat_o_6[3]
port 488 nsew signal input
rlabel metal3 s -800 3408 800 3528 4 m_wbs_dat_o_6[4]
port 489 nsew signal input
rlabel metal3 s -800 4224 800 4344 4 m_wbs_dat_o_6[5]
port 490 nsew signal input
rlabel metal3 s -800 5040 800 5160 4 m_wbs_dat_o_6[6]
port 491 nsew signal input
rlabel metal3 s -800 5856 800 5976 4 m_wbs_dat_o_6[7]
port 492 nsew signal input
rlabel metal3 s -800 6672 800 6792 4 m_wbs_dat_o_6[8]
port 493 nsew signal input
rlabel metal3 s -800 7352 800 7472 4 m_wbs_dat_o_6[9]
port 494 nsew signal input
rlabel metal3 s -800 25848 800 25968 4 m_wbs_dat_o_7[0]
port 495 nsew signal input
rlabel metal3 s -800 33736 800 33856 4 m_wbs_dat_o_7[10]
port 496 nsew signal input
rlabel metal3 s -800 34552 800 34672 4 m_wbs_dat_o_7[11]
port 497 nsew signal input
rlabel metal3 s -800 35368 800 35488 4 m_wbs_dat_o_7[12]
port 498 nsew signal input
rlabel metal3 s -800 36184 800 36304 4 m_wbs_dat_o_7[13]
port 499 nsew signal input
rlabel metal3 s -800 37000 800 37120 4 m_wbs_dat_o_7[14]
port 500 nsew signal input
rlabel metal3 s -800 37816 800 37936 4 m_wbs_dat_o_7[15]
port 501 nsew signal input
rlabel metal3 s -800 38632 800 38752 4 m_wbs_dat_o_7[16]
port 502 nsew signal input
rlabel metal3 s -800 39448 800 39568 4 m_wbs_dat_o_7[17]
port 503 nsew signal input
rlabel metal3 s -800 40264 800 40384 4 m_wbs_dat_o_7[18]
port 504 nsew signal input
rlabel metal3 s -800 40944 800 41064 4 m_wbs_dat_o_7[19]
port 505 nsew signal input
rlabel metal3 s -800 26664 800 26784 4 m_wbs_dat_o_7[1]
port 506 nsew signal input
rlabel metal3 s -800 41760 800 41880 4 m_wbs_dat_o_7[20]
port 507 nsew signal input
rlabel metal3 s -800 42576 800 42696 4 m_wbs_dat_o_7[21]
port 508 nsew signal input
rlabel metal3 s -800 43392 800 43512 4 m_wbs_dat_o_7[22]
port 509 nsew signal input
rlabel metal3 s -800 44208 800 44328 4 m_wbs_dat_o_7[23]
port 510 nsew signal input
rlabel metal3 s -800 45024 800 45144 4 m_wbs_dat_o_7[24]
port 511 nsew signal input
rlabel metal3 s -800 45840 800 45960 4 m_wbs_dat_o_7[25]
port 512 nsew signal input
rlabel metal3 s -800 46656 800 46776 4 m_wbs_dat_o_7[26]
port 513 nsew signal input
rlabel metal3 s -800 47336 800 47456 4 m_wbs_dat_o_7[27]
port 514 nsew signal input
rlabel metal3 s -800 48152 800 48272 4 m_wbs_dat_o_7[28]
port 515 nsew signal input
rlabel metal3 s -800 48968 800 49088 4 m_wbs_dat_o_7[29]
port 516 nsew signal input
rlabel metal3 s -800 27344 800 27464 4 m_wbs_dat_o_7[2]
port 517 nsew signal input
rlabel metal3 s -800 49784 800 49904 4 m_wbs_dat_o_7[30]
port 518 nsew signal input
rlabel metal3 s -800 50600 800 50720 4 m_wbs_dat_o_7[31]
port 519 nsew signal input
rlabel metal3 s -800 28160 800 28280 4 m_wbs_dat_o_7[3]
port 520 nsew signal input
rlabel metal3 s -800 28976 800 29096 4 m_wbs_dat_o_7[4]
port 521 nsew signal input
rlabel metal3 s -800 29792 800 29912 4 m_wbs_dat_o_7[5]
port 522 nsew signal input
rlabel metal3 s -800 30608 800 30728 4 m_wbs_dat_o_7[6]
port 523 nsew signal input
rlabel metal3 s -800 31424 800 31544 4 m_wbs_dat_o_7[7]
port 524 nsew signal input
rlabel metal3 s -800 32240 800 32360 4 m_wbs_dat_o_7[8]
port 525 nsew signal input
rlabel metal3 s -800 33056 800 33176 4 m_wbs_dat_o_7[9]
port 526 nsew signal input
rlabel metal3 s -800 51416 800 51536 4 m_wbs_dat_o_8[0]
port 527 nsew signal input
rlabel metal3 s -800 59440 800 59560 4 m_wbs_dat_o_8[10]
port 528 nsew signal input
rlabel metal3 s -800 60256 800 60376 4 m_wbs_dat_o_8[11]
port 529 nsew signal input
rlabel metal3 s -800 60936 800 61056 4 m_wbs_dat_o_8[12]
port 530 nsew signal input
rlabel metal3 s -800 61752 800 61872 4 m_wbs_dat_o_8[13]
port 531 nsew signal input
rlabel metal3 s -800 62568 800 62688 4 m_wbs_dat_o_8[14]
port 532 nsew signal input
rlabel metal3 s -800 63384 800 63504 4 m_wbs_dat_o_8[15]
port 533 nsew signal input
rlabel metal3 s -800 64200 800 64320 4 m_wbs_dat_o_8[16]
port 534 nsew signal input
rlabel metal3 s -800 65016 800 65136 4 m_wbs_dat_o_8[17]
port 535 nsew signal input
rlabel metal3 s -800 65832 800 65952 4 m_wbs_dat_o_8[18]
port 536 nsew signal input
rlabel metal3 s -800 66648 800 66768 4 m_wbs_dat_o_8[19]
port 537 nsew signal input
rlabel metal3 s -800 52232 800 52352 4 m_wbs_dat_o_8[1]
port 538 nsew signal input
rlabel metal3 s -800 67328 800 67448 4 m_wbs_dat_o_8[20]
port 539 nsew signal input
rlabel metal3 s -800 68144 800 68264 4 m_wbs_dat_o_8[21]
port 540 nsew signal input
rlabel metal3 s -800 68960 800 69080 4 m_wbs_dat_o_8[22]
port 541 nsew signal input
rlabel metal3 s -800 69776 800 69896 4 m_wbs_dat_o_8[23]
port 542 nsew signal input
rlabel metal3 s -800 70592 800 70712 4 m_wbs_dat_o_8[24]
port 543 nsew signal input
rlabel metal3 s -800 71408 800 71528 4 m_wbs_dat_o_8[25]
port 544 nsew signal input
rlabel metal3 s -800 72224 800 72344 4 m_wbs_dat_o_8[26]
port 545 nsew signal input
rlabel metal3 s -800 73040 800 73160 4 m_wbs_dat_o_8[27]
port 546 nsew signal input
rlabel metal3 s -800 73720 800 73840 4 m_wbs_dat_o_8[28]
port 547 nsew signal input
rlabel metal3 s -800 74536 800 74656 4 m_wbs_dat_o_8[29]
port 548 nsew signal input
rlabel metal3 s -800 53048 800 53168 4 m_wbs_dat_o_8[2]
port 549 nsew signal input
rlabel metal3 s -800 75352 800 75472 4 m_wbs_dat_o_8[30]
port 550 nsew signal input
rlabel metal3 s -800 76168 800 76288 4 m_wbs_dat_o_8[31]
port 551 nsew signal input
rlabel metal3 s -800 53728 800 53848 4 m_wbs_dat_o_8[3]
port 552 nsew signal input
rlabel metal3 s -800 54544 800 54664 4 m_wbs_dat_o_8[4]
port 553 nsew signal input
rlabel metal3 s -800 55360 800 55480 4 m_wbs_dat_o_8[5]
port 554 nsew signal input
rlabel metal3 s -800 56176 800 56296 4 m_wbs_dat_o_8[6]
port 555 nsew signal input
rlabel metal3 s -800 56992 800 57112 4 m_wbs_dat_o_8[7]
port 556 nsew signal input
rlabel metal3 s -800 57808 800 57928 4 m_wbs_dat_o_8[8]
port 557 nsew signal input
rlabel metal3 s -800 58624 800 58744 4 m_wbs_dat_o_8[9]
port 558 nsew signal input
rlabel metal3 s -800 76984 800 77104 4 m_wbs_dat_o_9[0]
port 559 nsew signal input
rlabel metal3 s -800 85008 800 85128 4 m_wbs_dat_o_9[10]
port 560 nsew signal input
rlabel metal3 s -800 85824 800 85944 4 m_wbs_dat_o_9[11]
port 561 nsew signal input
rlabel metal3 s -800 86640 800 86760 4 m_wbs_dat_o_9[12]
port 562 nsew signal input
rlabel metal3 s -800 87320 800 87440 4 m_wbs_dat_o_9[13]
port 563 nsew signal input
rlabel metal3 s -800 88136 800 88256 4 m_wbs_dat_o_9[14]
port 564 nsew signal input
rlabel metal3 s -800 88952 800 89072 4 m_wbs_dat_o_9[15]
port 565 nsew signal input
rlabel metal3 s -800 89768 800 89888 4 m_wbs_dat_o_9[16]
port 566 nsew signal input
rlabel metal3 s -800 90584 800 90704 4 m_wbs_dat_o_9[17]
port 567 nsew signal input
rlabel metal3 s -800 91400 800 91520 4 m_wbs_dat_o_9[18]
port 568 nsew signal input
rlabel metal3 s -800 92216 800 92336 4 m_wbs_dat_o_9[19]
port 569 nsew signal input
rlabel metal3 s -800 77800 800 77920 4 m_wbs_dat_o_9[1]
port 570 nsew signal input
rlabel metal3 s -800 93032 800 93152 4 m_wbs_dat_o_9[20]
port 571 nsew signal input
rlabel metal3 s -800 93712 800 93832 4 m_wbs_dat_o_9[21]
port 572 nsew signal input
rlabel metal3 s -800 94528 800 94648 4 m_wbs_dat_o_9[22]
port 573 nsew signal input
rlabel metal3 s -800 95344 800 95464 4 m_wbs_dat_o_9[23]
port 574 nsew signal input
rlabel metal3 s -800 96160 800 96280 4 m_wbs_dat_o_9[24]
port 575 nsew signal input
rlabel metal3 s -800 96976 800 97096 4 m_wbs_dat_o_9[25]
port 576 nsew signal input
rlabel metal3 s -800 97792 800 97912 4 m_wbs_dat_o_9[26]
port 577 nsew signal input
rlabel metal3 s -800 98608 800 98728 4 m_wbs_dat_o_9[27]
port 578 nsew signal input
rlabel metal3 s -800 99424 800 99544 4 m_wbs_dat_o_9[28]
port 579 nsew signal input
rlabel metal3 s -800 100240 800 100360 4 m_wbs_dat_o_9[29]
port 580 nsew signal input
rlabel metal3 s -800 78616 800 78736 4 m_wbs_dat_o_9[2]
port 581 nsew signal input
rlabel metal3 s -800 100920 800 101040 4 m_wbs_dat_o_9[30]
port 582 nsew signal input
rlabel metal3 s -800 101736 800 101856 4 m_wbs_dat_o_9[31]
port 583 nsew signal input
rlabel metal3 s -800 79432 800 79552 4 m_wbs_dat_o_9[3]
port 584 nsew signal input
rlabel metal3 s -800 80248 800 80368 4 m_wbs_dat_o_9[4]
port 585 nsew signal input
rlabel metal3 s -800 80928 800 81048 4 m_wbs_dat_o_9[5]
port 586 nsew signal input
rlabel metal3 s -800 81744 800 81864 4 m_wbs_dat_o_9[6]
port 587 nsew signal input
rlabel metal3 s -800 82560 800 82680 4 m_wbs_dat_o_9[7]
port 588 nsew signal input
rlabel metal3 s -800 83376 800 83496 4 m_wbs_dat_o_9[8]
port 589 nsew signal input
rlabel metal3 s -800 84192 800 84312 4 m_wbs_dat_o_9[9]
port 590 nsew signal input
rlabel metal3 s -800 102552 800 102672 4 m_wbs_we_i
port 591 nsew signal tristate
rlabel metal2 s 28262 119200 28318 120800 6 mt_QEI_ChA_0
port 592 nsew signal tristate
rlabel metal2 s 28538 119200 28594 120800 6 mt_QEI_ChA_1
port 593 nsew signal tristate
rlabel metal2 s 28722 119200 28778 120800 6 mt_QEI_ChA_2
port 594 nsew signal tristate
rlabel metal2 s 28998 119200 29054 120800 6 mt_QEI_ChA_3
port 595 nsew signal tristate
rlabel metal2 s 29182 119200 29238 120800 6 mt_QEI_ChB_0
port 596 nsew signal tristate
rlabel metal2 s 29458 119200 29514 120800 6 mt_QEI_ChB_1
port 597 nsew signal tristate
rlabel metal2 s 29642 119200 29698 120800 6 mt_QEI_ChB_2
port 598 nsew signal tristate
rlabel metal2 s 29918 119200 29974 120800 6 mt_QEI_ChB_3
port 599 nsew signal tristate
rlabel metal2 s 30102 119200 30158 120800 6 mt_pwm_h_0
port 600 nsew signal input
rlabel metal2 s 30378 119200 30434 120800 6 mt_pwm_h_1
port 601 nsew signal input
rlabel metal2 s 30562 119200 30618 120800 6 mt_pwm_h_2
port 602 nsew signal input
rlabel metal2 s 30838 119200 30894 120800 6 mt_pwm_h_3
port 603 nsew signal input
rlabel metal2 s 31022 119200 31078 120800 6 mt_pwm_l_0
port 604 nsew signal input
rlabel metal2 s 31298 119200 31354 120800 6 mt_pwm_l_1
port 605 nsew signal input
rlabel metal2 s 31482 119200 31538 120800 6 mt_pwm_l_2
port 606 nsew signal input
rlabel metal2 s 31758 119200 31814 120800 6 mt_pwm_l_3
port 607 nsew signal input
rlabel metal2 s 110 -800 166 800 8 wb_clk_i
port 608 nsew signal input
rlabel metal2 s 386 -800 442 800 8 wb_rst_i
port 609 nsew signal input
rlabel metal2 s 1674 -800 1730 800 8 wbs_ack_o
port 610 nsew signal tristate
rlabel metal2 s 2962 -800 3018 800 8 wbs_adr_i[0]
port 611 nsew signal input
rlabel metal2 s 14094 -800 14150 800 8 wbs_adr_i[10]
port 612 nsew signal input
rlabel metal2 s 15014 -800 15070 800 8 wbs_adr_i[11]
port 613 nsew signal input
rlabel metal2 s 16026 -800 16082 800 8 wbs_adr_i[12]
port 614 nsew signal input
rlabel metal2 s 16946 -800 17002 800 8 wbs_adr_i[13]
port 615 nsew signal input
rlabel metal2 s 17958 -800 18014 800 8 wbs_adr_i[14]
port 616 nsew signal input
rlabel metal2 s 18970 -800 19026 800 8 wbs_adr_i[15]
port 617 nsew signal input
rlabel metal2 s 19890 -800 19946 800 8 wbs_adr_i[16]
port 618 nsew signal input
rlabel metal2 s 20902 -800 20958 800 8 wbs_adr_i[17]
port 619 nsew signal input
rlabel metal2 s 21822 -800 21878 800 8 wbs_adr_i[18]
port 620 nsew signal input
rlabel metal2 s 22834 -800 22890 800 8 wbs_adr_i[19]
port 621 nsew signal input
rlabel metal2 s 4250 -800 4306 800 8 wbs_adr_i[1]
port 622 nsew signal input
rlabel metal2 s 23846 -800 23902 800 8 wbs_adr_i[20]
port 623 nsew signal input
rlabel metal2 s 24766 -800 24822 800 8 wbs_adr_i[21]
port 624 nsew signal input
rlabel metal2 s 25778 -800 25834 800 8 wbs_adr_i[22]
port 625 nsew signal input
rlabel metal2 s 26790 -800 26846 800 8 wbs_adr_i[23]
port 626 nsew signal input
rlabel metal2 s 27710 -800 27766 800 8 wbs_adr_i[24]
port 627 nsew signal input
rlabel metal2 s 28722 -800 28778 800 8 wbs_adr_i[25]
port 628 nsew signal input
rlabel metal2 s 29642 -800 29698 800 8 wbs_adr_i[26]
port 629 nsew signal input
rlabel metal2 s 30654 -800 30710 800 8 wbs_adr_i[27]
port 630 nsew signal input
rlabel metal2 s 31666 -800 31722 800 8 wbs_adr_i[28]
port 631 nsew signal input
rlabel metal2 s 32586 -800 32642 800 8 wbs_adr_i[29]
port 632 nsew signal input
rlabel metal2 s 5630 -800 5686 800 8 wbs_adr_i[2]
port 633 nsew signal input
rlabel metal2 s 33598 -800 33654 800 8 wbs_adr_i[30]
port 634 nsew signal input
rlabel metal2 s 34518 -800 34574 800 8 wbs_adr_i[31]
port 635 nsew signal input
rlabel metal2 s 6918 -800 6974 800 8 wbs_adr_i[3]
port 636 nsew signal input
rlabel metal2 s 8206 -800 8262 800 8 wbs_adr_i[4]
port 637 nsew signal input
rlabel metal2 s 9218 -800 9274 800 8 wbs_adr_i[5]
port 638 nsew signal input
rlabel metal2 s 10138 -800 10194 800 8 wbs_adr_i[6]
port 639 nsew signal input
rlabel metal2 s 11150 -800 11206 800 8 wbs_adr_i[7]
port 640 nsew signal input
rlabel metal2 s 12070 -800 12126 800 8 wbs_adr_i[8]
port 641 nsew signal input
rlabel metal2 s 13082 -800 13138 800 8 wbs_adr_i[9]
port 642 nsew signal input
rlabel metal2 s 2042 -800 2098 800 8 wbs_cyc_i
port 643 nsew signal input
rlabel metal2 s 3330 -800 3386 800 8 wbs_dat_i[0]
port 644 nsew signal input
rlabel metal2 s 14370 -800 14426 800 8 wbs_dat_i[10]
port 645 nsew signal input
rlabel metal2 s 15382 -800 15438 800 8 wbs_dat_i[11]
port 646 nsew signal input
rlabel metal2 s 16302 -800 16358 800 8 wbs_dat_i[12]
port 647 nsew signal input
rlabel metal2 s 17314 -800 17370 800 8 wbs_dat_i[13]
port 648 nsew signal input
rlabel metal2 s 18326 -800 18382 800 8 wbs_dat_i[14]
port 649 nsew signal input
rlabel metal2 s 19246 -800 19302 800 8 wbs_dat_i[15]
port 650 nsew signal input
rlabel metal2 s 20258 -800 20314 800 8 wbs_dat_i[16]
port 651 nsew signal input
rlabel metal2 s 21178 -800 21234 800 8 wbs_dat_i[17]
port 652 nsew signal input
rlabel metal2 s 22190 -800 22246 800 8 wbs_dat_i[18]
port 653 nsew signal input
rlabel metal2 s 23202 -800 23258 800 8 wbs_dat_i[19]
port 654 nsew signal input
rlabel metal2 s 4618 -800 4674 800 8 wbs_dat_i[1]
port 655 nsew signal input
rlabel metal2 s 24122 -800 24178 800 8 wbs_dat_i[20]
port 656 nsew signal input
rlabel metal2 s 25134 -800 25190 800 8 wbs_dat_i[21]
port 657 nsew signal input
rlabel metal2 s 26054 -800 26110 800 8 wbs_dat_i[22]
port 658 nsew signal input
rlabel metal2 s 27066 -800 27122 800 8 wbs_dat_i[23]
port 659 nsew signal input
rlabel metal2 s 28078 -800 28134 800 8 wbs_dat_i[24]
port 660 nsew signal input
rlabel metal2 s 28998 -800 29054 800 8 wbs_dat_i[25]
port 661 nsew signal input
rlabel metal2 s 30010 -800 30066 800 8 wbs_dat_i[26]
port 662 nsew signal input
rlabel metal2 s 30930 -800 30986 800 8 wbs_dat_i[27]
port 663 nsew signal input
rlabel metal2 s 31942 -800 31998 800 8 wbs_dat_i[28]
port 664 nsew signal input
rlabel metal2 s 32954 -800 33010 800 8 wbs_dat_i[29]
port 665 nsew signal input
rlabel metal2 s 5906 -800 5962 800 8 wbs_dat_i[2]
port 666 nsew signal input
rlabel metal2 s 33874 -800 33930 800 8 wbs_dat_i[30]
port 667 nsew signal input
rlabel metal2 s 34886 -800 34942 800 8 wbs_dat_i[31]
port 668 nsew signal input
rlabel metal2 s 7194 -800 7250 800 8 wbs_dat_i[3]
port 669 nsew signal input
rlabel metal2 s 8482 -800 8538 800 8 wbs_dat_i[4]
port 670 nsew signal input
rlabel metal2 s 9494 -800 9550 800 8 wbs_dat_i[5]
port 671 nsew signal input
rlabel metal2 s 10506 -800 10562 800 8 wbs_dat_i[6]
port 672 nsew signal input
rlabel metal2 s 11426 -800 11482 800 8 wbs_dat_i[7]
port 673 nsew signal input
rlabel metal2 s 12438 -800 12494 800 8 wbs_dat_i[8]
port 674 nsew signal input
rlabel metal2 s 13450 -800 13506 800 8 wbs_dat_i[9]
port 675 nsew signal input
rlabel metal2 s 3606 -800 3662 800 8 wbs_dat_o[0]
port 676 nsew signal tristate
rlabel metal2 s 14738 -800 14794 800 8 wbs_dat_o[10]
port 677 nsew signal tristate
rlabel metal2 s 15658 -800 15714 800 8 wbs_dat_o[11]
port 678 nsew signal tristate
rlabel metal2 s 16670 -800 16726 800 8 wbs_dat_o[12]
port 679 nsew signal tristate
rlabel metal2 s 17590 -800 17646 800 8 wbs_dat_o[13]
port 680 nsew signal tristate
rlabel metal2 s 18602 -800 18658 800 8 wbs_dat_o[14]
port 681 nsew signal tristate
rlabel metal2 s 19614 -800 19670 800 8 wbs_dat_o[15]
port 682 nsew signal tristate
rlabel metal2 s 20534 -800 20590 800 8 wbs_dat_o[16]
port 683 nsew signal tristate
rlabel metal2 s 21546 -800 21602 800 8 wbs_dat_o[17]
port 684 nsew signal tristate
rlabel metal2 s 22558 -800 22614 800 8 wbs_dat_o[18]
port 685 nsew signal tristate
rlabel metal2 s 23478 -800 23534 800 8 wbs_dat_o[19]
port 686 nsew signal tristate
rlabel metal2 s 4986 -800 5042 800 8 wbs_dat_o[1]
port 687 nsew signal tristate
rlabel metal2 s 24490 -800 24546 800 8 wbs_dat_o[20]
port 688 nsew signal tristate
rlabel metal2 s 25410 -800 25466 800 8 wbs_dat_o[21]
port 689 nsew signal tristate
rlabel metal2 s 26422 -800 26478 800 8 wbs_dat_o[22]
port 690 nsew signal tristate
rlabel metal2 s 27434 -800 27490 800 8 wbs_dat_o[23]
port 691 nsew signal tristate
rlabel metal2 s 28354 -800 28410 800 8 wbs_dat_o[24]
port 692 nsew signal tristate
rlabel metal2 s 29366 -800 29422 800 8 wbs_dat_o[25]
port 693 nsew signal tristate
rlabel metal2 s 30286 -800 30342 800 8 wbs_dat_o[26]
port 694 nsew signal tristate
rlabel metal2 s 31298 -800 31354 800 8 wbs_dat_o[27]
port 695 nsew signal tristate
rlabel metal2 s 32310 -800 32366 800 8 wbs_dat_o[28]
port 696 nsew signal tristate
rlabel metal2 s 33230 -800 33286 800 8 wbs_dat_o[29]
port 697 nsew signal tristate
rlabel metal2 s 6274 -800 6330 800 8 wbs_dat_o[2]
port 698 nsew signal tristate
rlabel metal2 s 34242 -800 34298 800 8 wbs_dat_o[30]
port 699 nsew signal tristate
rlabel metal2 s 35162 -800 35218 800 8 wbs_dat_o[31]
port 700 nsew signal tristate
rlabel metal2 s 7562 -800 7618 800 8 wbs_dat_o[3]
port 701 nsew signal tristate
rlabel metal2 s 8850 -800 8906 800 8 wbs_dat_o[4]
port 702 nsew signal tristate
rlabel metal2 s 9862 -800 9918 800 8 wbs_dat_o[5]
port 703 nsew signal tristate
rlabel metal2 s 10782 -800 10838 800 8 wbs_dat_o[6]
port 704 nsew signal tristate
rlabel metal2 s 11794 -800 11850 800 8 wbs_dat_o[7]
port 705 nsew signal tristate
rlabel metal2 s 12714 -800 12770 800 8 wbs_dat_o[8]
port 706 nsew signal tristate
rlabel metal2 s 13726 -800 13782 800 8 wbs_dat_o[9]
port 707 nsew signal tristate
rlabel metal2 s 3974 -800 4030 800 8 wbs_sel_i[0]
port 708 nsew signal input
rlabel metal2 s 5262 -800 5318 800 8 wbs_sel_i[1]
port 709 nsew signal input
rlabel metal2 s 6550 -800 6606 800 8 wbs_sel_i[2]
port 710 nsew signal input
rlabel metal2 s 7838 -800 7894 800 8 wbs_sel_i[3]
port 711 nsew signal input
rlabel metal2 s 2318 -800 2374 800 8 wbs_stb_i
port 712 nsew signal input
rlabel metal2 s 2686 -800 2742 800 8 wbs_we_i
port 713 nsew signal input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 714 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 715 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 716 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 120000
<< end >>
